VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_128x16m4w8
    CLASS BLOCK  ;
    FOREIGN sram22_128x16m4w8   ;
    SIZE 250.840 BY 224.320 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 139.830 0.000 139.970 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 145.930 0.000 146.070 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 152.030 0.000 152.170 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 158.130 0.000 158.270 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 164.230 0.000 164.370 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 170.330 0.000 170.470 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 176.430 0.000 176.570 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 182.530 0.000 182.670 0.140 ; 
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 188.630 0.000 188.770 0.140 ; 
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 194.730 0.000 194.870 0.140 ; 
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 200.830 0.000 200.970 0.140 ; 
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 206.930 0.000 207.070 0.140 ; 
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 213.030 0.000 213.170 0.140 ; 
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 219.130 0.000 219.270 0.140 ; 
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 225.230 0.000 225.370 0.140 ; 
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 231.330 0.000 231.470 0.140 ; 
        END 
    END dout[15] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 139.410 0.000 139.550 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 145.510 0.000 145.650 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 151.610 0.000 151.750 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 157.710 0.000 157.850 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 163.810 0.000 163.950 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 169.910 0.000 170.050 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 176.010 0.000 176.150 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 182.110 0.000 182.250 0.140 ; 
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 188.210 0.000 188.350 0.140 ; 
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 194.310 0.000 194.450 0.140 ; 
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 200.410 0.000 200.550 0.140 ; 
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 206.510 0.000 206.650 0.140 ; 
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 212.610 0.000 212.750 0.140 ; 
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 218.710 0.000 218.850 0.140 ; 
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 224.810 0.000 224.950 0.140 ; 
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 230.910 0.000 231.050 0.140 ; 
        END 
    END din[15] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.831200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 139.060 0.000 139.200 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.831200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 187.860 0.000 188.000 0.140 ; 
        END 
    END wmask[1] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 97.720 0.000 98.040 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 91.600 0.000 91.920 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 85.480 0.000 85.800 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 79.360 0.000 79.680 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 73.240 0.000 73.560 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 67.120 0.000 67.440 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 61.000 0.000 61.320 0.320 ; 
        END 
    END addr[6] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 109.960 0.000 110.280 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 103.840 0.000 104.160 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 12.555000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 112.680 0.000 113.000 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 16.461000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 113.360 0.000 113.680 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 138.840 6.240 ; 
                RECT 140.560 5.920 144.960 6.240 ; 
                RECT 146.680 5.920 151.080 6.240 ; 
                RECT 152.800 5.920 157.200 6.240 ; 
                RECT 158.920 5.920 163.320 6.240 ; 
                RECT 165.040 5.920 169.440 6.240 ; 
                RECT 171.160 5.920 175.560 6.240 ; 
                RECT 177.280 5.920 181.680 6.240 ; 
                RECT 183.400 5.920 187.800 6.240 ; 
                RECT 189.520 5.920 193.920 6.240 ; 
                RECT 195.640 5.920 200.040 6.240 ; 
                RECT 201.760 5.920 206.160 6.240 ; 
                RECT 207.880 5.920 212.280 6.240 ; 
                RECT 214.000 5.920 218.400 6.240 ; 
                RECT 220.120 5.920 224.520 6.240 ; 
                RECT 226.240 5.920 230.640 6.240 ; 
                RECT 232.360 5.920 250.680 6.240 ; 
                RECT 0.160 7.280 250.680 7.600 ; 
                RECT 0.160 8.640 250.680 8.960 ; 
                RECT 0.160 10.000 112.320 10.320 ; 
                RECT 135.120 10.000 250.680 10.320 ; 
                RECT 0.160 11.360 250.680 11.680 ; 
                RECT 0.160 12.720 250.680 13.040 ; 
                RECT 0.160 14.080 57.240 14.400 ; 
                RECT 114.040 14.080 250.680 14.400 ; 
                RECT 0.160 15.440 250.680 15.760 ; 
                RECT 0.160 16.800 250.680 17.120 ; 
                RECT 0.160 18.160 57.240 18.480 ; 
                RECT 113.360 18.160 138.160 18.480 ; 
                RECT 188.840 18.160 250.680 18.480 ; 
                RECT 0.160 19.520 128.640 19.840 ; 
                RECT 240.520 19.520 250.680 19.840 ; 
                RECT 0.160 20.880 128.640 21.200 ; 
                RECT 240.520 20.880 250.680 21.200 ; 
                RECT 0.160 22.240 128.640 22.560 ; 
                RECT 240.520 22.240 250.680 22.560 ; 
                RECT 0.160 23.600 128.640 23.920 ; 
                RECT 240.520 23.600 250.680 23.920 ; 
                RECT 0.160 24.960 128.640 25.280 ; 
                RECT 240.520 24.960 250.680 25.280 ; 
                RECT 0.160 26.320 128.640 26.640 ; 
                RECT 240.520 26.320 250.680 26.640 ; 
                RECT 0.160 27.680 128.640 28.000 ; 
                RECT 240.520 27.680 250.680 28.000 ; 
                RECT 0.160 29.040 128.640 29.360 ; 
                RECT 240.520 29.040 250.680 29.360 ; 
                RECT 0.160 30.400 128.640 30.720 ; 
                RECT 240.520 30.400 250.680 30.720 ; 
                RECT 0.160 31.760 128.640 32.080 ; 
                RECT 240.520 31.760 250.680 32.080 ; 
                RECT 0.160 33.120 79.680 33.440 ; 
                RECT 90.920 33.120 128.640 33.440 ; 
                RECT 240.520 33.120 250.680 33.440 ; 
                RECT 0.160 34.480 78.320 34.800 ; 
                RECT 97.040 34.480 128.640 34.800 ; 
                RECT 240.520 34.480 250.680 34.800 ; 
                RECT 0.160 35.840 59.280 36.160 ; 
                RECT 114.040 35.840 128.640 36.160 ; 
                RECT 240.520 35.840 250.680 36.160 ; 
                RECT 0.160 37.200 57.920 37.520 ; 
                RECT 109.960 37.200 127.960 37.520 ; 
                RECT 240.520 37.200 250.680 37.520 ; 
                RECT 0.160 38.560 128.640 38.880 ; 
                RECT 240.520 38.560 250.680 38.880 ; 
                RECT 0.160 39.920 128.640 40.240 ; 
                RECT 240.520 39.920 250.680 40.240 ; 
                RECT 0.160 41.280 128.640 41.600 ; 
                RECT 240.520 41.280 250.680 41.600 ; 
                RECT 0.160 42.640 128.640 42.960 ; 
                RECT 240.520 42.640 250.680 42.960 ; 
                RECT 0.160 44.000 54.520 44.320 ; 
                RECT 65.760 44.000 128.640 44.320 ; 
                RECT 240.520 44.000 250.680 44.320 ; 
                RECT 0.160 45.360 55.880 45.680 ; 
                RECT 61.680 45.360 69.480 45.680 ; 
                RECT 71.880 45.360 128.640 45.680 ; 
                RECT 240.520 45.360 250.680 45.680 ; 
                RECT 0.160 46.720 57.240 47.040 ; 
                RECT 61.000 46.720 128.640 47.040 ; 
                RECT 240.520 46.720 250.680 47.040 ; 
                RECT 0.160 48.080 128.640 48.400 ; 
                RECT 240.520 48.080 250.680 48.400 ; 
                RECT 0.160 49.440 64.040 49.760 ; 
                RECT 72.560 49.440 128.640 49.760 ; 
                RECT 240.520 49.440 250.680 49.760 ; 
                RECT 0.160 50.800 56.560 51.120 ; 
                RECT 65.760 50.800 128.640 51.120 ; 
                RECT 240.520 50.800 250.680 51.120 ; 
                RECT 0.160 52.160 59.960 52.480 ; 
                RECT 65.080 52.160 128.640 52.480 ; 
                RECT 240.520 52.160 250.680 52.480 ; 
                RECT 0.160 53.520 128.640 53.840 ; 
                RECT 240.520 53.520 250.680 53.840 ; 
                RECT 0.160 54.880 55.880 55.200 ; 
                RECT 65.760 54.880 106.200 55.200 ; 
                RECT 112.000 54.880 128.640 55.200 ; 
                RECT 240.520 54.880 250.680 55.200 ; 
                RECT 0.160 56.240 62.680 56.560 ; 
                RECT 71.200 56.240 106.200 56.560 ; 
                RECT 112.000 56.240 128.640 56.560 ; 
                RECT 240.520 56.240 250.680 56.560 ; 
                RECT 0.160 57.600 106.200 57.920 ; 
                RECT 240.520 57.600 250.680 57.920 ; 
                RECT 0.160 58.960 64.040 59.280 ; 
                RECT 69.840 58.960 106.200 59.280 ; 
                RECT 112.000 58.960 128.640 59.280 ; 
                RECT 240.520 58.960 250.680 59.280 ; 
                RECT 0.160 60.320 66.760 60.640 ; 
                RECT 71.880 60.320 128.640 60.640 ; 
                RECT 240.520 60.320 250.680 60.640 ; 
                RECT 0.160 61.680 60.640 62.000 ; 
                RECT 65.760 61.680 128.640 62.000 ; 
                RECT 240.520 61.680 250.680 62.000 ; 
                RECT 0.160 63.040 128.640 63.360 ; 
                RECT 240.520 63.040 250.680 63.360 ; 
                RECT 0.160 64.400 53.840 64.720 ; 
                RECT 76.640 64.400 89.880 64.720 ; 
                RECT 111.320 64.400 128.640 64.720 ; 
                RECT 240.520 64.400 250.680 64.720 ; 
                RECT 0.160 65.760 64.040 66.080 ; 
                RECT 71.880 65.760 79.000 66.080 ; 
                RECT 84.120 65.760 89.880 66.080 ; 
                RECT 111.320 65.760 128.640 66.080 ; 
                RECT 240.520 65.760 250.680 66.080 ; 
                RECT 0.160 67.120 62.680 67.440 ; 
                RECT 65.760 67.120 72.200 67.440 ; 
                RECT 78.680 67.120 80.360 67.440 ; 
                RECT 82.760 67.120 89.880 67.440 ; 
                RECT 120.840 67.120 128.640 67.440 ; 
                RECT 240.520 67.120 250.680 67.440 ; 
                RECT 0.160 68.480 54.520 68.800 ; 
                RECT 68.480 68.480 89.880 68.800 ; 
                RECT 120.840 68.480 128.640 68.800 ; 
                RECT 240.520 68.480 250.680 68.800 ; 
                RECT 0.160 69.840 63.360 70.160 ; 
                RECT 71.880 69.840 89.880 70.160 ; 
                RECT 119.480 69.840 128.640 70.160 ; 
                RECT 240.520 69.840 250.680 70.160 ; 
                RECT 0.160 71.200 60.640 71.520 ; 
                RECT 65.080 71.200 89.880 71.520 ; 
                RECT 120.840 71.200 128.640 71.520 ; 
                RECT 240.520 71.200 250.680 71.520 ; 
                RECT 0.160 72.560 56.560 72.880 ; 
                RECT 61.000 72.560 64.040 72.880 ; 
                RECT 72.560 72.560 89.880 72.880 ; 
                RECT 123.560 72.560 128.640 72.880 ; 
                RECT 240.520 72.560 250.680 72.880 ; 
                RECT 0.160 73.920 59.280 74.240 ; 
                RECT 62.360 73.920 89.880 74.240 ; 
                RECT 111.320 73.920 128.640 74.240 ; 
                RECT 240.520 73.920 250.680 74.240 ; 
                RECT 0.160 75.280 55.880 75.600 ; 
                RECT 59.640 75.280 89.880 75.600 ; 
                RECT 123.560 75.280 128.640 75.600 ; 
                RECT 240.520 75.280 250.680 75.600 ; 
                RECT 0.160 76.640 59.960 76.960 ; 
                RECT 65.760 76.640 89.880 76.960 ; 
                RECT 122.200 76.640 128.640 76.960 ; 
                RECT 240.520 76.640 250.680 76.960 ; 
                RECT 0.160 78.000 55.880 78.320 ; 
                RECT 71.200 78.000 89.880 78.320 ; 
                RECT 123.560 78.000 128.640 78.320 ; 
                RECT 240.520 78.000 250.680 78.320 ; 
                RECT 0.160 79.360 89.880 79.680 ; 
                RECT 126.280 79.360 128.640 79.680 ; 
                RECT 240.520 79.360 250.680 79.680 ; 
                RECT 0.160 80.720 62.680 81.040 ; 
                RECT 65.080 80.720 89.880 81.040 ; 
                RECT 126.280 80.720 128.640 81.040 ; 
                RECT 240.520 80.720 250.680 81.040 ; 
                RECT 0.160 82.080 64.040 82.400 ; 
                RECT 65.760 82.080 89.880 82.400 ; 
                RECT 124.920 82.080 128.640 82.400 ; 
                RECT 240.520 82.080 250.680 82.400 ; 
                RECT 0.160 83.440 54.520 83.760 ; 
                RECT 65.080 83.440 89.880 83.760 ; 
                RECT 111.320 83.440 128.640 83.760 ; 
                RECT 240.520 83.440 250.680 83.760 ; 
                RECT 0.160 84.800 59.960 85.120 ; 
                RECT 71.880 84.800 89.880 85.120 ; 
                RECT 124.920 84.800 128.640 85.120 ; 
                RECT 240.520 84.800 250.680 85.120 ; 
                RECT 0.160 86.160 54.520 86.480 ; 
                RECT 65.760 86.160 89.880 86.480 ; 
                RECT 240.520 86.160 250.680 86.480 ; 
                RECT 0.160 87.520 63.360 87.840 ; 
                RECT 65.760 87.520 89.880 87.840 ; 
                RECT 240.520 87.520 250.680 87.840 ; 
                RECT 0.160 88.880 89.880 89.200 ; 
                RECT 240.520 88.880 250.680 89.200 ; 
                RECT 0.160 90.240 89.880 90.560 ; 
                RECT 240.520 90.240 250.680 90.560 ; 
                RECT 0.160 91.600 51.120 91.920 ; 
                RECT 68.480 91.600 89.880 91.920 ; 
                RECT 111.320 91.600 128.640 91.920 ; 
                RECT 240.520 91.600 250.680 91.920 ; 
                RECT 0.160 92.960 128.640 93.280 ; 
                RECT 240.520 92.960 250.680 93.280 ; 
                RECT 0.160 94.320 128.640 94.640 ; 
                RECT 240.520 94.320 250.680 94.640 ; 
                RECT 0.160 95.680 59.280 96.000 ; 
                RECT 71.880 95.680 128.640 96.000 ; 
                RECT 240.520 95.680 250.680 96.000 ; 
                RECT 0.160 97.040 66.760 97.360 ; 
                RECT 73.920 97.040 128.640 97.360 ; 
                RECT 240.520 97.040 250.680 97.360 ; 
                RECT 0.160 98.400 77.640 98.720 ; 
                RECT 88.880 98.400 91.920 98.720 ; 
                RECT 112.000 98.400 128.640 98.720 ; 
                RECT 240.520 98.400 250.680 98.720 ; 
                RECT 0.160 99.760 91.920 100.080 ; 
                RECT 112.000 99.760 128.640 100.080 ; 
                RECT 240.520 99.760 250.680 100.080 ; 
                RECT 0.160 101.120 53.840 101.440 ; 
                RECT 59.640 101.120 91.920 101.440 ; 
                RECT 112.000 101.120 128.640 101.440 ; 
                RECT 240.520 101.120 250.680 101.440 ; 
                RECT 0.160 102.480 91.920 102.800 ; 
                RECT 112.000 102.480 128.640 102.800 ; 
                RECT 240.520 102.480 250.680 102.800 ; 
                RECT 0.160 103.840 91.920 104.160 ; 
                RECT 112.000 103.840 128.640 104.160 ; 
                RECT 240.520 103.840 250.680 104.160 ; 
                RECT 0.160 105.200 69.480 105.520 ; 
                RECT 72.560 105.200 91.920 105.520 ; 
                RECT 112.000 105.200 128.640 105.520 ; 
                RECT 240.520 105.200 250.680 105.520 ; 
                RECT 0.160 106.560 91.920 106.880 ; 
                RECT 112.000 106.560 128.640 106.880 ; 
                RECT 240.520 106.560 250.680 106.880 ; 
                RECT 0.160 107.920 91.920 108.240 ; 
                RECT 112.000 107.920 128.640 108.240 ; 
                RECT 240.520 107.920 250.680 108.240 ; 
                RECT 0.160 109.280 91.920 109.600 ; 
                RECT 240.520 109.280 250.680 109.600 ; 
                RECT 0.160 110.640 56.560 110.960 ; 
                RECT 61.000 110.640 91.920 110.960 ; 
                RECT 112.000 110.640 125.920 110.960 ; 
                RECT 240.520 110.640 250.680 110.960 ; 
                RECT 0.160 112.000 91.920 112.320 ; 
                RECT 112.000 112.000 123.200 112.320 ; 
                RECT 240.520 112.000 250.680 112.320 ; 
                RECT 0.160 113.360 32.760 113.680 ; 
                RECT 51.480 113.360 62.680 113.680 ; 
                RECT 71.200 113.360 91.920 113.680 ; 
                RECT 112.000 113.360 120.480 113.680 ; 
                RECT 240.520 113.360 250.680 113.680 ; 
                RECT 0.160 114.720 32.760 115.040 ; 
                RECT 51.480 114.720 117.760 115.040 ; 
                RECT 240.520 114.720 250.680 115.040 ; 
                RECT 0.160 116.080 32.760 116.400 ; 
                RECT 51.480 116.080 59.280 116.400 ; 
                RECT 61.680 116.080 128.640 116.400 ; 
                RECT 240.520 116.080 250.680 116.400 ; 
                RECT 0.160 117.440 32.760 117.760 ; 
                RECT 51.480 117.440 55.880 117.760 ; 
                RECT 58.960 117.440 128.640 117.760 ; 
                RECT 240.520 117.440 250.680 117.760 ; 
                RECT 0.160 118.800 32.760 119.120 ; 
                RECT 52.160 118.800 128.640 119.120 ; 
                RECT 240.520 118.800 250.680 119.120 ; 
                RECT 0.160 120.160 32.760 120.480 ; 
                RECT 51.480 120.160 91.920 120.480 ; 
                RECT 112.000 120.160 128.640 120.480 ; 
                RECT 240.520 120.160 250.680 120.480 ; 
                RECT 0.160 121.520 32.760 121.840 ; 
                RECT 51.480 121.520 91.920 121.840 ; 
                RECT 112.000 121.520 128.640 121.840 ; 
                RECT 240.520 121.520 250.680 121.840 ; 
                RECT 0.160 122.880 32.760 123.200 ; 
                RECT 51.480 122.880 91.920 123.200 ; 
                RECT 112.000 122.880 128.640 123.200 ; 
                RECT 240.520 122.880 250.680 123.200 ; 
                RECT 0.160 124.240 32.760 124.560 ; 
                RECT 51.480 124.240 91.920 124.560 ; 
                RECT 112.000 124.240 119.120 124.560 ; 
                RECT 240.520 124.240 250.680 124.560 ; 
                RECT 0.160 125.600 32.760 125.920 ; 
                RECT 51.480 125.600 91.920 125.920 ; 
                RECT 112.000 125.600 121.840 125.920 ; 
                RECT 240.520 125.600 250.680 125.920 ; 
                RECT 0.160 126.960 32.760 127.280 ; 
                RECT 51.480 126.960 57.920 127.280 ; 
                RECT 61.680 126.960 91.920 127.280 ; 
                RECT 112.000 126.960 124.560 127.280 ; 
                RECT 240.520 126.960 250.680 127.280 ; 
                RECT 0.160 128.320 91.920 128.640 ; 
                RECT 112.000 128.320 127.280 128.640 ; 
                RECT 240.520 128.320 250.680 128.640 ; 
                RECT 0.160 129.680 91.920 130.000 ; 
                RECT 240.520 129.680 250.680 130.000 ; 
                RECT 0.160 131.040 16.440 131.360 ; 
                RECT 32.440 131.040 59.960 131.360 ; 
                RECT 65.760 131.040 91.920 131.360 ; 
                RECT 112.000 131.040 128.640 131.360 ; 
                RECT 240.520 131.040 250.680 131.360 ; 
                RECT 0.160 132.400 16.440 132.720 ; 
                RECT 32.440 132.400 38.880 132.720 ; 
                RECT 46.040 132.400 91.920 132.720 ; 
                RECT 112.000 132.400 128.640 132.720 ; 
                RECT 240.520 132.400 250.680 132.720 ; 
                RECT 0.160 133.760 16.440 134.080 ; 
                RECT 32.440 133.760 33.440 134.080 ; 
                RECT 50.800 133.760 91.920 134.080 ; 
                RECT 112.000 133.760 128.640 134.080 ; 
                RECT 240.520 133.760 250.680 134.080 ; 
                RECT 0.160 135.120 16.440 135.440 ; 
                RECT 32.440 135.120 33.440 135.440 ; 
                RECT 50.800 135.120 91.920 135.440 ; 
                RECT 240.520 135.120 250.680 135.440 ; 
                RECT 0.160 136.480 16.440 136.800 ; 
                RECT 32.440 136.480 38.880 136.800 ; 
                RECT 46.040 136.480 54.520 136.800 ; 
                RECT 64.400 136.480 91.920 136.800 ; 
                RECT 112.000 136.480 115.040 136.800 ; 
                RECT 240.520 136.480 250.680 136.800 ; 
                RECT 0.160 137.840 17.120 138.160 ; 
                RECT 45.360 137.840 91.920 138.160 ; 
                RECT 112.000 137.840 250.680 138.160 ; 
                RECT 0.160 139.200 45.000 139.520 ; 
                RECT 89.560 139.200 250.680 139.520 ; 
                RECT 0.160 140.560 125.920 140.880 ; 
                RECT 243.240 140.560 250.680 140.880 ; 
                RECT 0.160 141.920 125.920 142.240 ; 
                RECT 243.240 141.920 250.680 142.240 ; 
                RECT 0.160 143.280 125.920 143.600 ; 
                RECT 243.240 143.280 250.680 143.600 ; 
                RECT 0.160 144.640 34.800 144.960 ; 
                RECT 41.280 144.640 42.960 144.960 ; 
                RECT 54.200 144.640 84.440 144.960 ; 
                RECT 243.240 144.640 250.680 144.960 ; 
                RECT 0.160 146.000 32.760 146.320 ; 
                RECT 53.520 146.000 67.440 146.320 ; 
                RECT 73.240 146.000 84.440 146.320 ; 
                RECT 243.240 146.000 250.680 146.320 ; 
                RECT 0.160 147.360 32.760 147.680 ; 
                RECT 52.840 147.360 65.400 147.680 ; 
                RECT 73.240 147.360 84.440 147.680 ; 
                RECT 243.240 147.360 250.680 147.680 ; 
                RECT 0.160 148.720 32.760 149.040 ; 
                RECT 43.320 148.720 65.400 149.040 ; 
                RECT 69.160 148.720 84.440 149.040 ; 
                RECT 243.240 148.720 250.680 149.040 ; 
                RECT 0.160 150.080 65.400 150.400 ; 
                RECT 73.240 150.080 84.440 150.400 ; 
                RECT 243.240 150.080 250.680 150.400 ; 
                RECT 0.160 151.440 32.760 151.760 ; 
                RECT 43.320 151.440 65.400 151.760 ; 
                RECT 73.240 151.440 84.440 151.760 ; 
                RECT 243.240 151.440 250.680 151.760 ; 
                RECT 0.160 152.800 32.760 153.120 ; 
                RECT 43.320 152.800 84.440 153.120 ; 
                RECT 243.240 152.800 250.680 153.120 ; 
                RECT 0.160 154.160 69.480 154.480 ; 
                RECT 73.240 154.160 84.440 154.480 ; 
                RECT 243.240 154.160 250.680 154.480 ; 
                RECT 0.160 155.520 65.400 155.840 ; 
                RECT 73.240 155.520 84.440 155.840 ; 
                RECT 243.240 155.520 250.680 155.840 ; 
                RECT 0.160 156.880 15.760 157.200 ; 
                RECT 28.360 156.880 65.400 157.200 ; 
                RECT 73.240 156.880 84.440 157.200 ; 
                RECT 243.240 156.880 250.680 157.200 ; 
                RECT 0.160 158.240 65.400 158.560 ; 
                RECT 67.120 158.240 84.440 158.560 ; 
                RECT 243.240 158.240 250.680 158.560 ; 
                RECT 0.160 159.600 15.080 159.920 ; 
                RECT 28.360 159.600 41.600 159.920 ; 
                RECT 44.680 159.600 65.400 159.920 ; 
                RECT 73.240 159.600 84.440 159.920 ; 
                RECT 243.240 159.600 250.680 159.920 ; 
                RECT 0.160 160.960 14.400 161.280 ; 
                RECT 28.360 160.960 41.600 161.280 ; 
                RECT 45.360 160.960 84.440 161.280 ; 
                RECT 243.240 160.960 250.680 161.280 ; 
                RECT 0.160 162.320 13.720 162.640 ; 
                RECT 28.360 162.320 41.600 162.640 ; 
                RECT 46.040 162.320 67.440 162.640 ; 
                RECT 73.240 162.320 84.440 162.640 ; 
                RECT 243.240 162.320 250.680 162.640 ; 
                RECT 0.160 163.680 65.400 164.000 ; 
                RECT 73.240 163.680 84.440 164.000 ; 
                RECT 243.240 163.680 250.680 164.000 ; 
                RECT 0.160 165.040 13.040 165.360 ; 
                RECT 28.360 165.040 41.600 165.360 ; 
                RECT 46.720 165.040 65.400 165.360 ; 
                RECT 73.240 165.040 84.440 165.360 ; 
                RECT 243.240 165.040 250.680 165.360 ; 
                RECT 0.160 166.400 12.360 166.720 ; 
                RECT 28.360 166.400 65.400 166.720 ; 
                RECT 73.240 166.400 84.440 166.720 ; 
                RECT 243.240 166.400 250.680 166.720 ; 
                RECT 0.160 167.760 11.680 168.080 ; 
                RECT 28.360 167.760 65.400 168.080 ; 
                RECT 71.880 167.760 84.440 168.080 ; 
                RECT 243.240 167.760 250.680 168.080 ; 
                RECT 0.160 169.120 11.000 169.440 ; 
                RECT 28.360 169.120 84.440 169.440 ; 
                RECT 243.240 169.120 250.680 169.440 ; 
                RECT 0.160 170.480 65.400 170.800 ; 
                RECT 73.240 170.480 84.440 170.800 ; 
                RECT 243.240 170.480 250.680 170.800 ; 
                RECT 0.160 171.840 10.320 172.160 ; 
                RECT 28.360 171.840 65.400 172.160 ; 
                RECT 73.240 171.840 84.440 172.160 ; 
                RECT 243.240 171.840 250.680 172.160 ; 
                RECT 0.160 173.200 9.640 173.520 ; 
                RECT 28.360 173.200 65.400 173.520 ; 
                RECT 73.240 173.200 84.440 173.520 ; 
                RECT 243.240 173.200 250.680 173.520 ; 
                RECT 0.160 174.560 65.400 174.880 ; 
                RECT 73.240 174.560 84.440 174.880 ; 
                RECT 243.240 174.560 250.680 174.880 ; 
                RECT 0.160 175.920 65.400 176.240 ; 
                RECT 72.560 175.920 84.440 176.240 ; 
                RECT 243.240 175.920 250.680 176.240 ; 
                RECT 0.160 177.280 67.440 177.600 ; 
                RECT 73.240 177.280 84.440 177.600 ; 
                RECT 243.240 177.280 250.680 177.600 ; 
                RECT 0.160 178.640 84.440 178.960 ; 
                RECT 243.240 178.640 250.680 178.960 ; 
                RECT 0.160 180.000 68.120 180.320 ; 
                RECT 73.240 180.000 84.440 180.320 ; 
                RECT 243.240 180.000 250.680 180.320 ; 
                RECT 0.160 181.360 68.800 181.680 ; 
                RECT 73.240 181.360 84.440 181.680 ; 
                RECT 243.240 181.360 250.680 181.680 ; 
                RECT 0.160 182.720 68.800 183.040 ; 
                RECT 73.240 182.720 84.440 183.040 ; 
                RECT 243.240 182.720 250.680 183.040 ; 
                RECT 0.160 184.080 45.000 184.400 ; 
                RECT 53.520 184.080 84.440 184.400 ; 
                RECT 243.240 184.080 250.680 184.400 ; 
                RECT 0.160 185.440 43.640 185.760 ; 
                RECT 52.840 185.440 65.400 185.760 ; 
                RECT 73.240 185.440 84.440 185.760 ; 
                RECT 243.240 185.440 250.680 185.760 ; 
                RECT 0.160 186.800 65.400 187.120 ; 
                RECT 73.240 186.800 84.440 187.120 ; 
                RECT 243.240 186.800 250.680 187.120 ; 
                RECT 0.160 188.160 65.400 188.480 ; 
                RECT 67.800 188.160 84.440 188.480 ; 
                RECT 243.240 188.160 250.680 188.480 ; 
                RECT 0.160 189.520 65.400 189.840 ; 
                RECT 73.240 189.520 84.440 189.840 ; 
                RECT 243.240 189.520 250.680 189.840 ; 
                RECT 0.160 190.880 65.400 191.200 ; 
                RECT 73.240 190.880 84.440 191.200 ; 
                RECT 243.240 190.880 250.680 191.200 ; 
                RECT 0.160 192.240 65.400 192.560 ; 
                RECT 68.480 192.240 84.440 192.560 ; 
                RECT 243.240 192.240 250.680 192.560 ; 
                RECT 0.160 193.600 67.440 193.920 ; 
                RECT 73.240 193.600 84.440 193.920 ; 
                RECT 243.240 193.600 250.680 193.920 ; 
                RECT 0.160 194.960 68.120 195.280 ; 
                RECT 73.240 194.960 84.440 195.280 ; 
                RECT 243.240 194.960 250.680 195.280 ; 
                RECT 0.160 196.320 68.800 196.640 ; 
                RECT 73.240 196.320 84.440 196.640 ; 
                RECT 243.240 196.320 250.680 196.640 ; 
                RECT 0.160 197.680 84.440 198.000 ; 
                RECT 243.240 197.680 250.680 198.000 ; 
                RECT 0.160 199.040 68.800 199.360 ; 
                RECT 73.240 199.040 84.440 199.360 ; 
                RECT 243.240 199.040 250.680 199.360 ; 
                RECT 0.160 200.400 84.440 200.720 ; 
                RECT 243.240 200.400 250.680 200.720 ; 
                RECT 0.160 201.760 69.480 202.080 ; 
                RECT 73.240 201.760 84.440 202.080 ; 
                RECT 243.240 201.760 250.680 202.080 ; 
                RECT 0.160 203.120 70.160 203.440 ; 
                RECT 73.240 203.120 84.440 203.440 ; 
                RECT 243.240 203.120 250.680 203.440 ; 
                RECT 0.160 204.480 70.160 204.800 ; 
                RECT 73.240 204.480 84.440 204.800 ; 
                RECT 243.240 204.480 250.680 204.800 ; 
                RECT 0.160 205.840 70.840 206.160 ; 
                RECT 73.240 205.840 84.440 206.160 ; 
                RECT 243.240 205.840 250.680 206.160 ; 
                RECT 0.160 207.200 84.440 207.520 ; 
                RECT 243.240 207.200 250.680 207.520 ; 
                RECT 0.160 208.560 84.440 208.880 ; 
                RECT 243.240 208.560 250.680 208.880 ; 
                RECT 0.160 209.920 125.920 210.240 ; 
                RECT 243.240 209.920 250.680 210.240 ; 
                RECT 0.160 211.280 125.920 211.600 ; 
                RECT 243.240 211.280 250.680 211.600 ; 
                RECT 0.160 212.640 125.920 212.960 ; 
                RECT 243.240 212.640 250.680 212.960 ; 
                RECT 0.160 214.000 250.680 214.320 ; 
                RECT 0.160 215.360 250.680 215.680 ; 
                RECT 0.160 216.720 250.680 217.040 ; 
                RECT 0.160 218.080 250.680 218.400 ; 
                RECT 0.160 0.160 250.680 1.520 ; 
                RECT 0.160 222.800 250.680 224.160 ; 
                RECT 130.060 40.720 135.860 42.090 ; 
                RECT 233.160 40.720 238.960 42.090 ; 
                RECT 130.060 45.835 135.860 47.255 ; 
                RECT 233.160 45.835 238.960 47.255 ; 
                RECT 130.060 51.155 135.860 52.675 ; 
                RECT 233.160 51.155 238.960 52.675 ; 
                RECT 130.060 56.625 135.860 58.145 ; 
                RECT 233.160 56.625 238.960 58.145 ; 
                RECT 130.060 132.560 238.960 133.910 ; 
                RECT 130.060 84.400 238.960 85.200 ; 
                RECT 130.060 65.030 238.960 66.830 ; 
                RECT 130.060 90.715 238.960 91.785 ; 
                RECT 130.060 95.005 238.960 95.295 ; 
                RECT 130.060 79.510 238.960 80.310 ; 
                RECT 130.060 117.310 238.960 118.280 ; 
                RECT 130.060 76.500 238.960 77.300 ; 
                RECT 130.060 24.965 238.960 26.765 ; 
                RECT 89.830 144.355 91.750 209.135 ; 
                RECT 93.670 144.355 95.590 209.135 ; 
                RECT 106.955 144.355 108.875 209.135 ; 
                RECT 110.795 144.355 112.715 209.135 ; 
                RECT 114.635 144.355 116.555 209.135 ; 
                RECT 118.475 144.355 120.395 209.135 ; 
                RECT 122.315 144.355 124.235 209.135 ; 
                RECT 93.275 65.060 95.195 91.860 ; 
                RECT 100.035 65.060 101.955 91.860 ; 
                RECT 108.515 65.060 110.435 91.860 ; 
                RECT 96.050 119.500 97.970 137.720 ; 
                RECT 103.025 119.500 104.945 137.720 ; 
                RECT 109.655 119.500 111.405 137.720 ; 
                RECT 95.620 97.860 97.540 113.500 ; 
                RECT 102.595 97.860 104.515 113.500 ; 
                RECT 109.355 97.860 111.275 113.500 ; 
                RECT 109.675 55.480 111.425 59.060 ; 
                RECT 33.450 146.625 42.610 147.375 ; 
                RECT 33.450 151.250 42.610 153.000 ; 
                RECT 34.020 134.410 50.060 135.210 ; 
                RECT 17.220 135.070 32.060 136.760 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 138.840 5.560 ; 
                RECT 140.560 5.240 144.960 5.560 ; 
                RECT 146.680 5.240 151.080 5.560 ; 
                RECT 152.800 5.240 157.200 5.560 ; 
                RECT 158.920 5.240 163.320 5.560 ; 
                RECT 165.040 5.240 169.440 5.560 ; 
                RECT 171.160 5.240 175.560 5.560 ; 
                RECT 177.280 5.240 181.680 5.560 ; 
                RECT 183.400 5.240 187.800 5.560 ; 
                RECT 189.520 5.240 193.920 5.560 ; 
                RECT 195.640 5.240 200.040 5.560 ; 
                RECT 201.760 5.240 206.160 5.560 ; 
                RECT 207.880 5.240 212.280 5.560 ; 
                RECT 214.000 5.240 218.400 5.560 ; 
                RECT 220.120 5.240 224.520 5.560 ; 
                RECT 226.240 5.240 230.640 5.560 ; 
                RECT 232.360 5.240 247.960 5.560 ; 
                RECT 2.880 6.600 247.960 6.920 ; 
                RECT 2.880 7.960 247.960 8.280 ; 
                RECT 2.880 9.320 113.000 9.640 ; 
                RECT 134.440 9.320 247.960 9.640 ; 
                RECT 2.880 10.680 247.960 11.000 ; 
                RECT 2.880 12.040 247.960 12.360 ; 
                RECT 2.880 13.400 57.240 13.720 ; 
                RECT 114.040 13.400 247.960 13.720 ; 
                RECT 2.880 14.760 247.960 15.080 ; 
                RECT 2.880 16.120 247.960 16.440 ; 
                RECT 2.880 17.480 57.240 17.800 ; 
                RECT 113.360 17.480 247.960 17.800 ; 
                RECT 2.880 18.840 128.640 19.160 ; 
                RECT 240.520 18.840 247.960 19.160 ; 
                RECT 2.880 20.200 128.640 20.520 ; 
                RECT 240.520 20.200 247.960 20.520 ; 
                RECT 2.880 21.560 128.640 21.880 ; 
                RECT 240.520 21.560 247.960 21.880 ; 
                RECT 2.880 22.920 128.640 23.240 ; 
                RECT 240.520 22.920 247.960 23.240 ; 
                RECT 2.880 24.280 128.640 24.600 ; 
                RECT 240.520 24.280 247.960 24.600 ; 
                RECT 2.880 25.640 128.640 25.960 ; 
                RECT 240.520 25.640 247.960 25.960 ; 
                RECT 2.880 27.000 128.640 27.320 ; 
                RECT 240.520 27.000 247.960 27.320 ; 
                RECT 2.880 28.360 128.640 28.680 ; 
                RECT 240.520 28.360 247.960 28.680 ; 
                RECT 2.880 29.720 128.640 30.040 ; 
                RECT 240.520 29.720 247.960 30.040 ; 
                RECT 2.880 31.080 128.640 31.400 ; 
                RECT 240.520 31.080 247.960 31.400 ; 
                RECT 2.880 32.440 80.360 32.760 ; 
                RECT 92.280 32.440 128.640 32.760 ; 
                RECT 240.520 32.440 247.960 32.760 ; 
                RECT 2.880 33.800 79.000 34.120 ; 
                RECT 98.400 33.800 128.640 34.120 ; 
                RECT 240.520 33.800 247.960 34.120 ; 
                RECT 2.880 35.160 56.560 35.480 ; 
                RECT 113.360 35.160 128.640 35.480 ; 
                RECT 240.520 35.160 247.960 35.480 ; 
                RECT 2.880 36.520 57.240 36.840 ; 
                RECT 103.840 36.520 127.960 36.840 ; 
                RECT 240.520 36.520 247.960 36.840 ; 
                RECT 2.880 37.880 128.640 38.200 ; 
                RECT 240.520 37.880 247.960 38.200 ; 
                RECT 2.880 39.240 128.640 39.560 ; 
                RECT 240.520 39.240 247.960 39.560 ; 
                RECT 2.880 40.600 128.640 40.920 ; 
                RECT 240.520 40.600 247.960 40.920 ; 
                RECT 2.880 41.960 128.640 42.280 ; 
                RECT 240.520 41.960 247.960 42.280 ; 
                RECT 2.880 43.320 54.520 43.640 ; 
                RECT 65.760 43.320 128.640 43.640 ; 
                RECT 240.520 43.320 247.960 43.640 ; 
                RECT 2.880 44.680 55.880 45.000 ; 
                RECT 58.280 44.680 128.640 45.000 ; 
                RECT 240.520 44.680 247.960 45.000 ; 
                RECT 2.880 46.040 57.240 46.360 ; 
                RECT 61.680 46.040 69.480 46.360 ; 
                RECT 71.880 46.040 128.640 46.360 ; 
                RECT 240.520 46.040 247.960 46.360 ; 
                RECT 2.880 47.400 57.240 47.720 ; 
                RECT 61.000 47.400 128.640 47.720 ; 
                RECT 240.520 47.400 247.960 47.720 ; 
                RECT 2.880 48.760 64.040 49.080 ; 
                RECT 72.560 48.760 128.640 49.080 ; 
                RECT 240.520 48.760 247.960 49.080 ; 
                RECT 2.880 50.120 59.280 50.440 ; 
                RECT 65.760 50.120 128.640 50.440 ; 
                RECT 240.520 50.120 247.960 50.440 ; 
                RECT 2.880 51.480 56.560 51.800 ; 
                RECT 65.760 51.480 128.640 51.800 ; 
                RECT 240.520 51.480 247.960 51.800 ; 
                RECT 2.880 52.840 128.640 53.160 ; 
                RECT 240.520 52.840 247.960 53.160 ; 
                RECT 2.880 54.200 55.880 54.520 ; 
                RECT 65.760 54.200 128.640 54.520 ; 
                RECT 240.520 54.200 247.960 54.520 ; 
                RECT 2.880 55.560 64.040 55.880 ; 
                RECT 71.200 55.560 106.200 55.880 ; 
                RECT 112.000 55.560 128.640 55.880 ; 
                RECT 240.520 55.560 247.960 55.880 ; 
                RECT 2.880 56.920 62.680 57.240 ; 
                RECT 65.760 56.920 106.200 57.240 ; 
                RECT 240.520 56.920 247.960 57.240 ; 
                RECT 2.880 58.280 76.960 58.600 ; 
                RECT 103.840 58.280 106.200 58.600 ; 
                RECT 112.000 58.280 128.640 58.600 ; 
                RECT 240.520 58.280 247.960 58.600 ; 
                RECT 2.880 59.640 64.040 59.960 ; 
                RECT 71.880 59.640 128.640 59.960 ; 
                RECT 240.520 59.640 247.960 59.960 ; 
                RECT 2.880 61.000 60.640 61.320 ; 
                RECT 65.760 61.000 128.640 61.320 ; 
                RECT 240.520 61.000 247.960 61.320 ; 
                RECT 2.880 62.360 62.680 62.680 ; 
                RECT 65.760 62.360 128.640 62.680 ; 
                RECT 240.520 62.360 247.960 62.680 ; 
                RECT 2.880 63.720 128.640 64.040 ; 
                RECT 240.520 63.720 247.960 64.040 ; 
                RECT 2.880 65.080 53.840 65.400 ; 
                RECT 84.800 65.080 89.880 65.400 ; 
                RECT 111.320 65.080 128.640 65.400 ; 
                RECT 240.520 65.080 247.960 65.400 ; 
                RECT 2.880 66.440 72.200 66.760 ; 
                RECT 78.000 66.440 79.680 66.760 ; 
                RECT 83.440 66.440 89.880 66.760 ; 
                RECT 120.840 66.440 128.640 66.760 ; 
                RECT 240.520 66.440 247.960 66.760 ; 
                RECT 2.880 67.800 62.680 68.120 ; 
                RECT 65.760 67.800 74.920 68.120 ; 
                RECT 78.680 67.800 89.880 68.120 ; 
                RECT 119.480 67.800 128.640 68.120 ; 
                RECT 240.520 67.800 247.960 68.120 ; 
                RECT 2.880 69.160 54.520 69.480 ; 
                RECT 68.480 69.160 89.880 69.480 ; 
                RECT 120.840 69.160 128.640 69.480 ; 
                RECT 240.520 69.160 247.960 69.480 ; 
                RECT 2.880 70.520 63.360 70.840 ; 
                RECT 71.880 70.520 89.880 70.840 ; 
                RECT 120.840 70.520 128.640 70.840 ; 
                RECT 240.520 70.520 247.960 70.840 ; 
                RECT 2.880 71.880 60.640 72.200 ; 
                RECT 72.560 71.880 89.880 72.200 ; 
                RECT 111.320 71.880 128.640 72.200 ; 
                RECT 240.520 71.880 247.960 72.200 ; 
                RECT 2.880 73.240 56.560 73.560 ; 
                RECT 62.360 73.240 89.880 73.560 ; 
                RECT 122.200 73.240 128.640 73.560 ; 
                RECT 240.520 73.240 247.960 73.560 ; 
                RECT 2.880 74.600 89.880 74.920 ; 
                RECT 111.320 74.600 128.640 74.920 ; 
                RECT 240.520 74.600 247.960 74.920 ; 
                RECT 2.880 75.960 55.880 76.280 ; 
                RECT 59.640 75.960 89.880 76.280 ; 
                RECT 123.560 75.960 128.640 76.280 ; 
                RECT 240.520 75.960 247.960 76.280 ; 
                RECT 2.880 77.320 55.880 77.640 ; 
                RECT 65.760 77.320 89.880 77.640 ; 
                RECT 123.560 77.320 128.640 77.640 ; 
                RECT 240.520 77.320 247.960 77.640 ; 
                RECT 2.880 78.680 59.960 79.000 ; 
                RECT 71.200 78.680 89.880 79.000 ; 
                RECT 126.280 78.680 128.640 79.000 ; 
                RECT 240.520 78.680 247.960 79.000 ; 
                RECT 2.880 80.040 62.680 80.360 ; 
                RECT 65.080 80.040 89.880 80.360 ; 
                RECT 124.920 80.040 128.640 80.360 ; 
                RECT 240.520 80.040 247.960 80.360 ; 
                RECT 2.880 81.400 64.040 81.720 ; 
                RECT 65.760 81.400 89.880 81.720 ; 
                RECT 126.280 81.400 128.640 81.720 ; 
                RECT 240.520 81.400 247.960 81.720 ; 
                RECT 2.880 82.760 89.880 83.080 ; 
                RECT 111.320 82.760 128.640 83.080 ; 
                RECT 240.520 82.760 247.960 83.080 ; 
                RECT 2.880 84.120 54.520 84.440 ; 
                RECT 71.880 84.120 89.880 84.440 ; 
                RECT 126.280 84.120 128.640 84.440 ; 
                RECT 240.520 84.120 247.960 84.440 ; 
                RECT 2.880 85.480 54.520 85.800 ; 
                RECT 65.760 85.480 69.480 85.800 ; 
                RECT 71.880 85.480 89.880 85.800 ; 
                RECT 240.520 85.480 247.960 85.800 ; 
                RECT 2.880 86.840 63.360 87.160 ; 
                RECT 65.760 86.840 89.880 87.160 ; 
                RECT 240.520 86.840 247.960 87.160 ; 
                RECT 2.880 88.200 89.880 88.520 ; 
                RECT 240.520 88.200 247.960 88.520 ; 
                RECT 2.880 89.560 89.880 89.880 ; 
                RECT 240.520 89.560 247.960 89.880 ; 
                RECT 2.880 90.920 51.120 91.240 ; 
                RECT 64.400 90.920 89.880 91.240 ; 
                RECT 240.520 90.920 247.960 91.240 ; 
                RECT 2.880 92.280 60.640 92.600 ; 
                RECT 68.480 92.280 128.640 92.600 ; 
                RECT 240.520 92.280 247.960 92.600 ; 
                RECT 2.880 93.640 128.640 93.960 ; 
                RECT 240.520 93.640 247.960 93.960 ; 
                RECT 2.880 95.000 128.640 95.320 ; 
                RECT 240.520 95.000 247.960 95.320 ; 
                RECT 2.880 96.360 59.280 96.680 ; 
                RECT 73.920 96.360 128.640 96.680 ; 
                RECT 240.520 96.360 247.960 96.680 ; 
                RECT 2.880 97.720 91.920 98.040 ; 
                RECT 112.000 97.720 128.640 98.040 ; 
                RECT 240.520 97.720 247.960 98.040 ; 
                RECT 2.880 99.080 91.920 99.400 ; 
                RECT 112.000 99.080 128.640 99.400 ; 
                RECT 240.520 99.080 247.960 99.400 ; 
                RECT 2.880 100.440 56.560 100.760 ; 
                RECT 59.640 100.440 91.920 100.760 ; 
                RECT 112.000 100.440 128.640 100.760 ; 
                RECT 240.520 100.440 247.960 100.760 ; 
                RECT 2.880 101.800 53.840 102.120 ; 
                RECT 58.280 101.800 91.920 102.120 ; 
                RECT 112.000 101.800 128.640 102.120 ; 
                RECT 240.520 101.800 247.960 102.120 ; 
                RECT 2.880 103.160 91.920 103.480 ; 
                RECT 112.000 103.160 128.640 103.480 ; 
                RECT 240.520 103.160 247.960 103.480 ; 
                RECT 2.880 104.520 69.480 104.840 ; 
                RECT 72.560 104.520 91.920 104.840 ; 
                RECT 112.000 104.520 128.640 104.840 ; 
                RECT 240.520 104.520 247.960 104.840 ; 
                RECT 2.880 105.880 91.920 106.200 ; 
                RECT 112.000 105.880 128.640 106.200 ; 
                RECT 240.520 105.880 247.960 106.200 ; 
                RECT 2.880 107.240 91.920 107.560 ; 
                RECT 112.000 107.240 128.640 107.560 ; 
                RECT 240.520 107.240 247.960 107.560 ; 
                RECT 2.880 108.600 91.920 108.920 ; 
                RECT 240.520 108.600 247.960 108.920 ; 
                RECT 2.880 109.960 56.560 110.280 ; 
                RECT 61.000 109.960 91.920 110.280 ; 
                RECT 112.000 109.960 125.920 110.280 ; 
                RECT 240.520 109.960 247.960 110.280 ; 
                RECT 2.880 111.320 91.920 111.640 ; 
                RECT 112.000 111.320 123.200 111.640 ; 
                RECT 240.520 111.320 247.960 111.640 ; 
                RECT 2.880 112.680 32.760 113.000 ; 
                RECT 51.480 112.680 62.680 113.000 ; 
                RECT 71.200 112.680 91.920 113.000 ; 
                RECT 112.000 112.680 120.480 113.000 ; 
                RECT 240.520 112.680 247.960 113.000 ; 
                RECT 2.880 114.040 32.760 114.360 ; 
                RECT 51.480 114.040 117.760 114.360 ; 
                RECT 240.520 114.040 247.960 114.360 ; 
                RECT 2.880 115.400 32.760 115.720 ; 
                RECT 51.480 115.400 59.280 115.720 ; 
                RECT 61.680 115.400 117.760 115.720 ; 
                RECT 240.520 115.400 247.960 115.720 ; 
                RECT 2.880 116.760 32.760 117.080 ; 
                RECT 51.480 116.760 55.880 117.080 ; 
                RECT 58.960 116.760 128.640 117.080 ; 
                RECT 240.520 116.760 247.960 117.080 ; 
                RECT 2.880 118.120 32.760 118.440 ; 
                RECT 51.480 118.120 128.640 118.440 ; 
                RECT 240.520 118.120 247.960 118.440 ; 
                RECT 2.880 119.480 32.760 119.800 ; 
                RECT 51.480 119.480 91.920 119.800 ; 
                RECT 112.000 119.480 128.640 119.800 ; 
                RECT 240.520 119.480 247.960 119.800 ; 
                RECT 2.880 120.840 32.760 121.160 ; 
                RECT 51.480 120.840 91.920 121.160 ; 
                RECT 112.000 120.840 128.640 121.160 ; 
                RECT 240.520 120.840 247.960 121.160 ; 
                RECT 2.880 122.200 32.760 122.520 ; 
                RECT 51.480 122.200 91.920 122.520 ; 
                RECT 112.000 122.200 128.640 122.520 ; 
                RECT 240.520 122.200 247.960 122.520 ; 
                RECT 2.880 123.560 32.760 123.880 ; 
                RECT 51.480 123.560 91.920 123.880 ; 
                RECT 112.000 123.560 119.120 123.880 ; 
                RECT 240.520 123.560 247.960 123.880 ; 
                RECT 2.880 124.920 32.760 125.240 ; 
                RECT 51.480 124.920 91.920 125.240 ; 
                RECT 112.000 124.920 119.120 125.240 ; 
                RECT 240.520 124.920 247.960 125.240 ; 
                RECT 2.880 126.280 32.760 126.600 ; 
                RECT 51.480 126.280 57.920 126.600 ; 
                RECT 61.680 126.280 91.920 126.600 ; 
                RECT 112.000 126.280 121.840 126.600 ; 
                RECT 240.520 126.280 247.960 126.600 ; 
                RECT 2.880 127.640 91.920 127.960 ; 
                RECT 112.000 127.640 124.560 127.960 ; 
                RECT 240.520 127.640 247.960 127.960 ; 
                RECT 2.880 129.000 91.920 129.320 ; 
                RECT 240.520 129.000 247.960 129.320 ; 
                RECT 2.880 130.360 91.920 130.680 ; 
                RECT 240.520 130.360 247.960 130.680 ; 
                RECT 2.880 131.720 16.440 132.040 ; 
                RECT 32.440 131.720 59.960 132.040 ; 
                RECT 65.760 131.720 91.920 132.040 ; 
                RECT 112.000 131.720 128.640 132.040 ; 
                RECT 240.520 131.720 247.960 132.040 ; 
                RECT 2.880 133.080 16.440 133.400 ; 
                RECT 32.440 133.080 38.880 133.400 ; 
                RECT 46.040 133.080 91.920 133.400 ; 
                RECT 112.000 133.080 128.640 133.400 ; 
                RECT 240.520 133.080 247.960 133.400 ; 
                RECT 2.880 134.440 16.440 134.760 ; 
                RECT 32.440 134.440 33.440 134.760 ; 
                RECT 50.800 134.440 91.920 134.760 ; 
                RECT 112.000 134.440 128.640 134.760 ; 
                RECT 240.520 134.440 247.960 134.760 ; 
                RECT 2.880 135.800 16.440 136.120 ; 
                RECT 32.440 135.800 91.920 136.120 ; 
                RECT 240.520 135.800 247.960 136.120 ; 
                RECT 2.880 137.160 17.120 137.480 ; 
                RECT 46.040 137.160 54.520 137.480 ; 
                RECT 64.400 137.160 91.920 137.480 ; 
                RECT 112.000 137.160 128.640 137.480 ; 
                RECT 240.520 137.160 247.960 137.480 ; 
                RECT 2.880 138.520 38.880 138.840 ; 
                RECT 58.960 138.520 247.960 138.840 ; 
                RECT 2.880 139.880 39.560 140.200 ; 
                RECT 58.280 139.880 247.960 140.200 ; 
                RECT 2.880 141.240 125.920 141.560 ; 
                RECT 243.240 141.240 247.960 141.560 ; 
                RECT 2.880 142.600 125.920 142.920 ; 
                RECT 243.240 142.600 247.960 142.920 ; 
                RECT 2.880 143.960 34.800 144.280 ; 
                RECT 41.280 143.960 84.440 144.280 ; 
                RECT 243.240 143.960 247.960 144.280 ; 
                RECT 2.880 145.320 32.760 145.640 ; 
                RECT 54.200 145.320 84.440 145.640 ; 
                RECT 243.240 145.320 247.960 145.640 ; 
                RECT 2.880 146.680 32.760 147.000 ; 
                RECT 52.840 146.680 65.400 147.000 ; 
                RECT 73.240 146.680 84.440 147.000 ; 
                RECT 243.240 146.680 247.960 147.000 ; 
                RECT 2.880 148.040 46.360 148.360 ; 
                RECT 52.160 148.040 65.400 148.360 ; 
                RECT 73.240 148.040 84.440 148.360 ; 
                RECT 243.240 148.040 247.960 148.360 ; 
                RECT 2.880 149.400 32.760 149.720 ; 
                RECT 43.320 149.400 65.400 149.720 ; 
                RECT 73.240 149.400 84.440 149.720 ; 
                RECT 243.240 149.400 247.960 149.720 ; 
                RECT 2.880 150.760 32.760 151.080 ; 
                RECT 43.320 150.760 65.400 151.080 ; 
                RECT 73.240 150.760 84.440 151.080 ; 
                RECT 243.240 150.760 247.960 151.080 ; 
                RECT 2.880 152.120 32.760 152.440 ; 
                RECT 43.320 152.120 65.400 152.440 ; 
                RECT 69.840 152.120 84.440 152.440 ; 
                RECT 243.240 152.120 247.960 152.440 ; 
                RECT 2.880 153.480 84.440 153.800 ; 
                RECT 243.240 153.480 247.960 153.800 ; 
                RECT 2.880 154.840 65.400 155.160 ; 
                RECT 73.240 154.840 84.440 155.160 ; 
                RECT 243.240 154.840 247.960 155.160 ; 
                RECT 2.880 156.200 65.400 156.520 ; 
                RECT 73.240 156.200 84.440 156.520 ; 
                RECT 243.240 156.200 247.960 156.520 ; 
                RECT 2.880 157.560 15.760 157.880 ; 
                RECT 28.360 157.560 41.600 157.880 ; 
                RECT 44.000 157.560 70.160 157.880 ; 
                RECT 73.240 157.560 84.440 157.880 ; 
                RECT 243.240 157.560 247.960 157.880 ; 
                RECT 2.880 158.920 15.080 159.240 ; 
                RECT 28.360 158.920 65.400 159.240 ; 
                RECT 73.240 158.920 84.440 159.240 ; 
                RECT 243.240 158.920 247.960 159.240 ; 
                RECT 2.880 160.280 14.400 160.600 ; 
                RECT 28.360 160.280 65.400 160.600 ; 
                RECT 70.520 160.280 84.440 160.600 ; 
                RECT 243.240 160.280 247.960 160.600 ; 
                RECT 2.880 161.640 13.720 161.960 ; 
                RECT 28.360 161.640 67.440 161.960 ; 
                RECT 73.240 161.640 84.440 161.960 ; 
                RECT 243.240 161.640 247.960 161.960 ; 
                RECT 2.880 163.000 65.400 163.320 ; 
                RECT 67.120 163.000 84.440 163.320 ; 
                RECT 243.240 163.000 247.960 163.320 ; 
                RECT 2.880 164.360 13.040 164.680 ; 
                RECT 28.360 164.360 65.400 164.680 ; 
                RECT 71.200 164.360 84.440 164.680 ; 
                RECT 243.240 164.360 247.960 164.680 ; 
                RECT 2.880 165.720 65.400 166.040 ; 
                RECT 73.240 165.720 84.440 166.040 ; 
                RECT 243.240 165.720 247.960 166.040 ; 
                RECT 2.880 167.080 12.360 167.400 ; 
                RECT 28.360 167.080 41.600 167.400 ; 
                RECT 47.400 167.080 65.400 167.400 ; 
                RECT 73.240 167.080 84.440 167.400 ; 
                RECT 243.240 167.080 247.960 167.400 ; 
                RECT 2.880 168.440 11.680 168.760 ; 
                RECT 28.360 168.440 41.600 168.760 ; 
                RECT 46.040 168.440 65.400 168.760 ; 
                RECT 71.880 168.440 84.440 168.760 ; 
                RECT 243.240 168.440 247.960 168.760 ; 
                RECT 2.880 169.800 11.000 170.120 ; 
                RECT 28.360 169.800 41.600 170.120 ; 
                RECT 45.360 169.800 69.480 170.120 ; 
                RECT 73.240 169.800 84.440 170.120 ; 
                RECT 243.240 169.800 247.960 170.120 ; 
                RECT 2.880 171.160 65.400 171.480 ; 
                RECT 73.240 171.160 84.440 171.480 ; 
                RECT 243.240 171.160 247.960 171.480 ; 
                RECT 2.880 172.520 10.320 172.840 ; 
                RECT 28.360 172.520 41.600 172.840 ; 
                RECT 44.680 172.520 65.400 172.840 ; 
                RECT 71.880 172.520 84.440 172.840 ; 
                RECT 243.240 172.520 247.960 172.840 ; 
                RECT 2.880 173.880 9.640 174.200 ; 
                RECT 28.360 173.880 41.600 174.200 ; 
                RECT 44.000 173.880 65.400 174.200 ; 
                RECT 67.120 173.880 84.440 174.200 ; 
                RECT 243.240 173.880 247.960 174.200 ; 
                RECT 2.880 175.240 65.400 175.560 ; 
                RECT 73.240 175.240 84.440 175.560 ; 
                RECT 243.240 175.240 247.960 175.560 ; 
                RECT 2.880 176.600 84.440 176.920 ; 
                RECT 243.240 176.600 247.960 176.920 ; 
                RECT 2.880 177.960 67.440 178.280 ; 
                RECT 73.240 177.960 84.440 178.280 ; 
                RECT 243.240 177.960 247.960 178.280 ; 
                RECT 2.880 179.320 68.120 179.640 ; 
                RECT 73.240 179.320 84.440 179.640 ; 
                RECT 243.240 179.320 247.960 179.640 ; 
                RECT 2.880 180.680 68.800 181.000 ; 
                RECT 73.240 180.680 84.440 181.000 ; 
                RECT 243.240 180.680 247.960 181.000 ; 
                RECT 2.880 182.040 68.800 182.360 ; 
                RECT 73.240 182.040 84.440 182.360 ; 
                RECT 243.240 182.040 247.960 182.360 ; 
                RECT 2.880 183.400 84.440 183.720 ; 
                RECT 243.240 183.400 247.960 183.720 ; 
                RECT 2.880 184.760 44.320 185.080 ; 
                RECT 53.520 184.760 84.440 185.080 ; 
                RECT 243.240 184.760 247.960 185.080 ; 
                RECT 2.880 186.120 42.960 186.440 ; 
                RECT 52.160 186.120 65.400 186.440 ; 
                RECT 73.240 186.120 84.440 186.440 ; 
                RECT 243.240 186.120 247.960 186.440 ; 
                RECT 2.880 187.480 65.400 187.800 ; 
                RECT 73.240 187.480 84.440 187.800 ; 
                RECT 243.240 187.480 247.960 187.800 ; 
                RECT 2.880 188.840 65.400 189.160 ; 
                RECT 73.240 188.840 84.440 189.160 ; 
                RECT 243.240 188.840 247.960 189.160 ; 
                RECT 2.880 190.200 65.400 190.520 ; 
                RECT 73.240 190.200 84.440 190.520 ; 
                RECT 243.240 190.200 247.960 190.520 ; 
                RECT 2.880 191.560 65.400 191.880 ; 
                RECT 68.480 191.560 84.440 191.880 ; 
                RECT 243.240 191.560 247.960 191.880 ; 
                RECT 2.880 192.920 84.440 193.240 ; 
                RECT 243.240 192.920 247.960 193.240 ; 
                RECT 2.880 194.280 67.440 194.600 ; 
                RECT 73.240 194.280 84.440 194.600 ; 
                RECT 243.240 194.280 247.960 194.600 ; 
                RECT 2.880 195.640 68.120 195.960 ; 
                RECT 73.240 195.640 84.440 195.960 ; 
                RECT 243.240 195.640 247.960 195.960 ; 
                RECT 2.880 197.000 68.800 197.320 ; 
                RECT 73.240 197.000 84.440 197.320 ; 
                RECT 243.240 197.000 247.960 197.320 ; 
                RECT 2.880 198.360 68.800 198.680 ; 
                RECT 73.240 198.360 84.440 198.680 ; 
                RECT 243.240 198.360 247.960 198.680 ; 
                RECT 2.880 199.720 84.440 200.040 ; 
                RECT 243.240 199.720 247.960 200.040 ; 
                RECT 2.880 201.080 69.480 201.400 ; 
                RECT 73.240 201.080 84.440 201.400 ; 
                RECT 243.240 201.080 247.960 201.400 ; 
                RECT 2.880 202.440 84.440 202.760 ; 
                RECT 243.240 202.440 247.960 202.760 ; 
                RECT 2.880 203.800 70.160 204.120 ; 
                RECT 73.240 203.800 84.440 204.120 ; 
                RECT 243.240 203.800 247.960 204.120 ; 
                RECT 2.880 205.160 70.160 205.480 ; 
                RECT 73.240 205.160 84.440 205.480 ; 
                RECT 243.240 205.160 247.960 205.480 ; 
                RECT 2.880 206.520 70.840 206.840 ; 
                RECT 73.240 206.520 84.440 206.840 ; 
                RECT 243.240 206.520 247.960 206.840 ; 
                RECT 2.880 207.880 84.440 208.200 ; 
                RECT 243.240 207.880 247.960 208.200 ; 
                RECT 2.880 209.240 84.440 209.560 ; 
                RECT 243.240 209.240 247.960 209.560 ; 
                RECT 2.880 210.600 125.920 210.920 ; 
                RECT 243.240 210.600 247.960 210.920 ; 
                RECT 2.880 211.960 125.920 212.280 ; 
                RECT 243.240 211.960 247.960 212.280 ; 
                RECT 2.880 213.320 247.960 213.640 ; 
                RECT 2.880 214.680 247.960 215.000 ; 
                RECT 2.880 216.040 247.960 216.360 ; 
                RECT 2.880 217.400 247.960 217.720 ; 
                RECT 2.880 218.760 247.960 219.080 ; 
                RECT 2.880 2.880 247.960 4.240 ; 
                RECT 2.880 220.080 247.960 221.440 ; 
                RECT 130.060 38.075 135.860 39.195 ; 
                RECT 233.160 38.075 238.960 39.195 ; 
                RECT 130.060 43.875 135.860 44.525 ; 
                RECT 233.160 43.875 238.960 44.525 ; 
                RECT 130.060 49.085 135.860 49.775 ; 
                RECT 233.160 49.085 238.960 49.775 ; 
                RECT 130.060 54.555 135.860 55.245 ; 
                RECT 233.160 54.555 238.960 55.245 ; 
                RECT 130.060 88.845 238.960 89.915 ; 
                RECT 130.060 82.510 238.960 83.310 ; 
                RECT 130.060 80.830 238.960 81.630 ; 
                RECT 130.060 68.770 238.960 70.570 ; 
                RECT 130.060 77.820 238.960 78.620 ; 
                RECT 130.060 107.565 238.960 107.855 ; 
                RECT 130.060 121.790 238.960 122.160 ; 
                RECT 130.060 85.720 238.960 86.520 ; 
                RECT 130.060 28.705 238.960 30.505 ; 
                RECT 85.170 144.355 87.090 209.135 ; 
                RECT 98.825 144.355 100.745 209.135 ; 
                RECT 102.665 144.355 104.585 209.135 ; 
                RECT 90.650 65.060 91.540 91.860 ; 
                RECT 97.410 65.060 98.300 91.860 ; 
                RECT 104.385 65.060 105.705 91.860 ; 
                RECT 92.885 119.500 93.995 137.720 ; 
                RECT 100.400 119.500 101.290 137.720 ; 
                RECT 107.160 119.500 108.050 137.720 ; 
                RECT 92.455 97.860 93.565 113.500 ; 
                RECT 99.970 97.860 100.860 113.500 ; 
                RECT 106.730 97.860 107.620 113.500 ; 
                RECT 107.180 55.480 108.070 59.060 ; 
                RECT 33.450 145.420 42.610 145.790 ; 
                RECT 33.450 148.755 42.610 149.645 ; 
                RECT 17.220 131.580 32.060 132.250 ; 
                RECT 17.220 132.930 32.060 133.940 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 250.840 224.320 ; 
        LAYER met2 ;
            RECT 0.000 0.000 250.840 224.320 ; 
    END 
END sram22_128x16m4w8 
END LIBRARY 

