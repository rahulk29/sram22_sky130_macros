VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_2048x8m8w1
    CLASS BLOCK  ;
    FOREIGN sram22_2048x8m8w1   ;
    SIZE 310.680 BY 760.160 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.142200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 212.950 0.000 213.090 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.142200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 223.850 0.000 223.990 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.142200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 234.750 0.000 234.890 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.142200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 245.650 0.000 245.790 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.142200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 256.550 0.000 256.690 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.142200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 267.450 0.000 267.590 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.142200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 278.350 0.000 278.490 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.142200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 289.250 0.000 289.390 0.140 ; 
        END 
    END dout[7] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.678800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.863800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 212.530 0.000 212.670 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.678800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.863800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 223.430 0.000 223.570 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.678800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.863800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 234.330 0.000 234.470 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.678800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.863800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 245.230 0.000 245.370 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.678800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.863800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 256.130 0.000 256.270 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.678800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.863800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 267.030 0.000 267.170 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.678800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.863800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 277.930 0.000 278.070 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.678800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.863800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 288.830 0.000 288.970 0.140 ; 
        END 
    END din[7] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.489200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 212.180 0.000 212.320 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.489200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 223.080 0.000 223.220 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.489200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 233.980 0.000 234.120 0.140 ; 
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.489200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 244.880 0.000 245.020 0.140 ; 
        END 
    END wmask[3] 
    PIN wmask[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.489200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 255.780 0.000 255.920 0.140 ; 
        END 
    END wmask[4] 
    PIN wmask[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.489200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 266.680 0.000 266.820 0.140 ; 
        END 
    END wmask[5] 
    PIN wmask[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.489200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 277.580 0.000 277.720 0.140 ; 
        END 
    END wmask[6] 
    PIN wmask[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.489200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 288.480 0.000 288.620 0.140 ; 
        END 
    END wmask[7] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 156.880 0.000 157.200 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 150.760 0.000 151.080 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 144.640 0.000 144.960 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 138.520 0.000 138.840 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 133.080 0.000 133.400 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 126.960 0.000 127.280 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 120.840 0.000 121.160 0.320 ; 
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 114.720 0.000 115.040 0.320 ; 
        END 
    END addr[7] 
    PIN addr[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 108.600 0.000 108.920 0.320 ; 
        END 
    END addr[8] 
    PIN addr[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 102.480 0.000 102.800 0.320 ; 
        END 
    END addr[9] 
    PIN addr[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 96.360 0.000 96.680 0.320 ; 
        END 
    END addr[10] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 169.120 0.000 169.440 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.848700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 163.000 0.000 163.320 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 10.881000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 172.520 0.000 172.840 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 14.787000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 173.200 0.000 173.520 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 212.280 6.240 ; 
                RECT 214.000 5.920 223.160 6.240 ; 
                RECT 224.880 5.920 234.040 6.240 ; 
                RECT 235.760 5.920 244.920 6.240 ; 
                RECT 246.640 5.920 255.800 6.240 ; 
                RECT 257.520 5.920 266.680 6.240 ; 
                RECT 268.400 5.920 277.560 6.240 ; 
                RECT 279.280 5.920 288.440 6.240 ; 
                RECT 290.160 5.920 310.520 6.240 ; 
                RECT 0.160 7.280 310.520 7.600 ; 
                RECT 0.160 8.640 310.520 8.960 ; 
                RECT 0.160 10.000 172.160 10.320 ; 
                RECT 205.840 10.000 310.520 10.320 ; 
                RECT 0.160 11.360 310.520 11.680 ; 
                RECT 0.160 12.720 310.520 13.040 ; 
                RECT 0.160 14.080 91.920 14.400 ; 
                RECT 173.880 14.080 310.520 14.400 ; 
                RECT 0.160 15.440 310.520 15.760 ; 
                RECT 0.160 16.800 310.520 17.120 ; 
                RECT 0.160 18.160 91.920 18.480 ; 
                RECT 173.200 18.160 310.520 18.480 ; 
                RECT 0.160 19.520 310.520 19.840 ; 
                RECT 0.160 20.880 310.520 21.200 ; 
                RECT 0.160 22.240 310.520 22.560 ; 
                RECT 0.160 23.600 199.360 23.920 ; 
                RECT 301.040 23.600 310.520 23.920 ; 
                RECT 0.160 24.960 199.360 25.280 ; 
                RECT 301.040 24.960 310.520 25.280 ; 
                RECT 0.160 26.320 199.360 26.640 ; 
                RECT 301.040 26.320 310.520 26.640 ; 
                RECT 0.160 27.680 199.360 28.000 ; 
                RECT 301.040 27.680 310.520 28.000 ; 
                RECT 0.160 29.040 199.360 29.360 ; 
                RECT 301.040 29.040 310.520 29.360 ; 
                RECT 0.160 30.400 199.360 30.720 ; 
                RECT 301.040 30.400 310.520 30.720 ; 
                RECT 0.160 31.760 199.360 32.080 ; 
                RECT 301.040 31.760 310.520 32.080 ; 
                RECT 0.160 33.120 199.360 33.440 ; 
                RECT 301.040 33.120 310.520 33.440 ; 
                RECT 0.160 34.480 199.360 34.800 ; 
                RECT 301.040 34.480 310.520 34.800 ; 
                RECT 0.160 35.840 199.360 36.160 ; 
                RECT 301.040 35.840 310.520 36.160 ; 
                RECT 0.160 37.200 104.840 37.520 ; 
                RECT 144.640 37.200 199.360 37.520 ; 
                RECT 301.040 37.200 310.520 37.520 ; 
                RECT 0.160 38.560 103.480 38.880 ; 
                RECT 150.760 38.560 199.360 38.880 ; 
                RECT 301.040 38.560 310.520 38.880 ; 
                RECT 0.160 39.920 102.120 40.240 ; 
                RECT 156.880 39.920 199.360 40.240 ; 
                RECT 301.040 39.920 310.520 40.240 ; 
                RECT 0.160 41.280 83.080 41.600 ; 
                RECT 173.880 41.280 198.680 41.600 ; 
                RECT 301.040 41.280 310.520 41.600 ; 
                RECT 0.160 42.640 81.720 42.960 ; 
                RECT 169.800 42.640 199.360 42.960 ; 
                RECT 301.040 42.640 310.520 42.960 ; 
                RECT 0.160 44.000 199.360 44.320 ; 
                RECT 301.040 44.000 310.520 44.320 ; 
                RECT 0.160 45.360 199.360 45.680 ; 
                RECT 301.040 45.360 310.520 45.680 ; 
                RECT 0.160 46.720 166.040 47.040 ; 
                RECT 171.840 46.720 199.360 47.040 ; 
                RECT 301.040 46.720 310.520 47.040 ; 
                RECT 0.160 48.080 166.040 48.400 ; 
                RECT 301.040 48.080 310.520 48.400 ; 
                RECT 0.160 49.440 166.040 49.760 ; 
                RECT 301.040 49.440 310.520 49.760 ; 
                RECT 0.160 50.800 100.760 51.120 ; 
                RECT 163.000 50.800 166.040 51.120 ; 
                RECT 171.840 50.800 199.360 51.120 ; 
                RECT 301.040 50.800 310.520 51.120 ; 
                RECT 0.160 52.160 199.360 52.480 ; 
                RECT 301.040 52.160 310.520 52.480 ; 
                RECT 0.160 53.520 199.360 53.840 ; 
                RECT 301.040 53.520 310.520 53.840 ; 
                RECT 0.160 54.880 199.360 55.200 ; 
                RECT 301.040 54.880 310.520 55.200 ; 
                RECT 0.160 56.240 199.360 56.560 ; 
                RECT 301.040 56.240 310.520 56.560 ; 
                RECT 0.160 57.600 102.120 57.920 ; 
                RECT 110.640 57.600 117.080 57.920 ; 
                RECT 171.160 57.600 199.360 57.920 ; 
                RECT 301.040 57.600 310.520 57.920 ; 
                RECT 0.160 58.960 103.480 59.280 ; 
                RECT 109.960 58.960 117.080 59.280 ; 
                RECT 180.680 58.960 199.360 59.280 ; 
                RECT 301.040 58.960 310.520 59.280 ; 
                RECT 0.160 60.320 104.840 60.640 ; 
                RECT 108.600 60.320 117.080 60.640 ; 
                RECT 180.680 60.320 199.360 60.640 ; 
                RECT 301.040 60.320 310.520 60.640 ; 
                RECT 0.160 61.680 117.080 62.000 ; 
                RECT 179.320 61.680 199.360 62.000 ; 
                RECT 301.040 61.680 310.520 62.000 ; 
                RECT 0.160 63.040 117.080 63.360 ; 
                RECT 180.680 63.040 199.360 63.360 ; 
                RECT 301.040 63.040 310.520 63.360 ; 
                RECT 0.160 64.400 117.080 64.720 ; 
                RECT 180.680 64.400 199.360 64.720 ; 
                RECT 301.040 64.400 310.520 64.720 ; 
                RECT 0.160 65.760 117.080 66.080 ; 
                RECT 179.320 65.760 199.360 66.080 ; 
                RECT 301.040 65.760 310.520 66.080 ; 
                RECT 0.160 67.120 117.080 67.440 ; 
                RECT 183.400 67.120 199.360 67.440 ; 
                RECT 301.040 67.120 310.520 67.440 ; 
                RECT 0.160 68.480 117.080 68.800 ; 
                RECT 182.040 68.480 199.360 68.800 ; 
                RECT 301.040 68.480 310.520 68.800 ; 
                RECT 0.160 69.840 117.080 70.160 ; 
                RECT 183.400 69.840 199.360 70.160 ; 
                RECT 301.040 69.840 310.520 70.160 ; 
                RECT 0.160 71.200 117.080 71.520 ; 
                RECT 183.400 71.200 199.360 71.520 ; 
                RECT 301.040 71.200 310.520 71.520 ; 
                RECT 0.160 72.560 117.080 72.880 ; 
                RECT 182.040 72.560 199.360 72.880 ; 
                RECT 301.040 72.560 310.520 72.880 ; 
                RECT 0.160 73.920 117.080 74.240 ; 
                RECT 183.400 73.920 199.360 74.240 ; 
                RECT 301.040 73.920 310.520 74.240 ; 
                RECT 0.160 75.280 117.080 75.600 ; 
                RECT 171.160 75.280 199.360 75.600 ; 
                RECT 301.040 75.280 310.520 75.600 ; 
                RECT 0.160 76.640 117.080 76.960 ; 
                RECT 186.120 76.640 199.360 76.960 ; 
                RECT 301.040 76.640 310.520 76.960 ; 
                RECT 0.160 78.000 117.080 78.320 ; 
                RECT 186.120 78.000 199.360 78.320 ; 
                RECT 301.040 78.000 310.520 78.320 ; 
                RECT 0.160 79.360 117.080 79.680 ; 
                RECT 171.160 79.360 199.360 79.680 ; 
                RECT 301.040 79.360 310.520 79.680 ; 
                RECT 0.160 80.720 117.080 81.040 ; 
                RECT 184.760 80.720 199.360 81.040 ; 
                RECT 301.040 80.720 310.520 81.040 ; 
                RECT 0.160 82.080 117.080 82.400 ; 
                RECT 186.120 82.080 199.360 82.400 ; 
                RECT 301.040 82.080 310.520 82.400 ; 
                RECT 0.160 83.440 117.080 83.760 ; 
                RECT 171.160 83.440 199.360 83.760 ; 
                RECT 301.040 83.440 310.520 83.760 ; 
                RECT 0.160 84.800 117.080 85.120 ; 
                RECT 188.840 84.800 199.360 85.120 ; 
                RECT 301.040 84.800 310.520 85.120 ; 
                RECT 0.160 86.160 117.080 86.480 ; 
                RECT 188.840 86.160 199.360 86.480 ; 
                RECT 301.040 86.160 310.520 86.480 ; 
                RECT 0.160 87.520 117.080 87.840 ; 
                RECT 187.480 87.520 199.360 87.840 ; 
                RECT 301.040 87.520 310.520 87.840 ; 
                RECT 0.160 88.880 117.080 89.200 ; 
                RECT 188.840 88.880 199.360 89.200 ; 
                RECT 301.040 88.880 310.520 89.200 ; 
                RECT 0.160 90.240 117.080 90.560 ; 
                RECT 188.840 90.240 199.360 90.560 ; 
                RECT 301.040 90.240 310.520 90.560 ; 
                RECT 0.160 91.600 117.080 91.920 ; 
                RECT 187.480 91.600 199.360 91.920 ; 
                RECT 301.040 91.600 310.520 91.920 ; 
                RECT 0.160 92.960 117.080 93.280 ; 
                RECT 191.560 92.960 199.360 93.280 ; 
                RECT 301.040 92.960 310.520 93.280 ; 
                RECT 0.160 94.320 117.080 94.640 ; 
                RECT 190.200 94.320 199.360 94.640 ; 
                RECT 301.040 94.320 310.520 94.640 ; 
                RECT 0.160 95.680 117.080 96.000 ; 
                RECT 191.560 95.680 199.360 96.000 ; 
                RECT 301.040 95.680 310.520 96.000 ; 
                RECT 0.160 97.040 117.080 97.360 ; 
                RECT 191.560 97.040 199.360 97.360 ; 
                RECT 301.040 97.040 310.520 97.360 ; 
                RECT 0.160 98.400 117.080 98.720 ; 
                RECT 190.200 98.400 199.360 98.720 ; 
                RECT 301.040 98.400 310.520 98.720 ; 
                RECT 0.160 99.760 117.080 100.080 ; 
                RECT 191.560 99.760 199.360 100.080 ; 
                RECT 301.040 99.760 310.520 100.080 ; 
                RECT 0.160 101.120 117.080 101.440 ; 
                RECT 171.160 101.120 199.360 101.440 ; 
                RECT 301.040 101.120 310.520 101.440 ; 
                RECT 0.160 102.480 117.080 102.800 ; 
                RECT 194.280 102.480 199.360 102.800 ; 
                RECT 301.040 102.480 310.520 102.800 ; 
                RECT 0.160 103.840 117.080 104.160 ; 
                RECT 194.280 103.840 199.360 104.160 ; 
                RECT 301.040 103.840 310.520 104.160 ; 
                RECT 0.160 105.200 117.080 105.520 ; 
                RECT 171.160 105.200 199.360 105.520 ; 
                RECT 301.040 105.200 310.520 105.520 ; 
                RECT 0.160 106.560 117.080 106.880 ; 
                RECT 192.920 106.560 199.360 106.880 ; 
                RECT 301.040 106.560 310.520 106.880 ; 
                RECT 0.160 107.920 117.080 108.240 ; 
                RECT 194.280 107.920 199.360 108.240 ; 
                RECT 301.040 107.920 310.520 108.240 ; 
                RECT 0.160 109.280 117.080 109.600 ; 
                RECT 171.160 109.280 199.360 109.600 ; 
                RECT 301.040 109.280 310.520 109.600 ; 
                RECT 0.160 110.640 117.080 110.960 ; 
                RECT 197.000 110.640 199.360 110.960 ; 
                RECT 301.040 110.640 310.520 110.960 ; 
                RECT 0.160 112.000 117.080 112.320 ; 
                RECT 197.000 112.000 199.360 112.320 ; 
                RECT 301.040 112.000 310.520 112.320 ; 
                RECT 0.160 113.360 117.080 113.680 ; 
                RECT 195.640 113.360 199.360 113.680 ; 
                RECT 301.040 113.360 310.520 113.680 ; 
                RECT 0.160 114.720 117.080 115.040 ; 
                RECT 197.000 114.720 199.360 115.040 ; 
                RECT 301.040 114.720 310.520 115.040 ; 
                RECT 0.160 116.080 117.080 116.400 ; 
                RECT 197.000 116.080 199.360 116.400 ; 
                RECT 301.040 116.080 310.520 116.400 ; 
                RECT 0.160 117.440 117.080 117.760 ; 
                RECT 195.640 117.440 199.360 117.760 ; 
                RECT 301.040 117.440 310.520 117.760 ; 
                RECT 0.160 118.800 117.080 119.120 ; 
                RECT 301.040 118.800 310.520 119.120 ; 
                RECT 0.160 120.160 117.080 120.480 ; 
                RECT 301.040 120.160 310.520 120.480 ; 
                RECT 0.160 121.520 117.080 121.840 ; 
                RECT 301.040 121.520 310.520 121.840 ; 
                RECT 0.160 122.880 117.080 123.200 ; 
                RECT 301.040 122.880 310.520 123.200 ; 
                RECT 0.160 124.240 117.080 124.560 ; 
                RECT 171.160 124.240 199.360 124.560 ; 
                RECT 301.040 124.240 310.520 124.560 ; 
                RECT 0.160 125.600 117.080 125.920 ; 
                RECT 301.040 125.600 310.520 125.920 ; 
                RECT 0.160 126.960 117.080 127.280 ; 
                RECT 171.160 126.960 199.360 127.280 ; 
                RECT 301.040 126.960 310.520 127.280 ; 
                RECT 0.160 128.320 199.360 128.640 ; 
                RECT 301.040 128.320 310.520 128.640 ; 
                RECT 0.160 129.680 174.880 130.000 ; 
                RECT 301.040 129.680 310.520 130.000 ; 
                RECT 0.160 131.040 196.640 131.360 ; 
                RECT 301.040 131.040 310.520 131.360 ; 
                RECT 0.160 132.400 193.920 132.720 ; 
                RECT 301.040 132.400 310.520 132.720 ; 
                RECT 0.160 133.760 191.200 134.080 ; 
                RECT 301.040 133.760 310.520 134.080 ; 
                RECT 0.160 135.120 188.480 135.440 ; 
                RECT 301.040 135.120 310.520 135.440 ; 
                RECT 0.160 136.480 78.320 136.800 ; 
                RECT 88.880 136.480 185.760 136.800 ; 
                RECT 301.040 136.480 310.520 136.800 ; 
                RECT 0.160 137.840 79.680 138.160 ; 
                RECT 82.080 137.840 183.040 138.160 ; 
                RECT 301.040 137.840 310.520 138.160 ; 
                RECT 0.160 139.200 81.040 139.520 ; 
                RECT 85.480 139.200 93.280 139.520 ; 
                RECT 95.680 139.200 180.320 139.520 ; 
                RECT 301.040 139.200 310.520 139.520 ; 
                RECT 0.160 140.560 81.040 140.880 ; 
                RECT 84.800 140.560 177.600 140.880 ; 
                RECT 301.040 140.560 310.520 140.880 ; 
                RECT 0.160 141.920 56.560 142.240 ; 
                RECT 75.280 141.920 87.160 142.240 ; 
                RECT 96.360 141.920 199.360 142.240 ; 
                RECT 301.040 141.920 310.520 142.240 ; 
                RECT 0.160 143.280 56.560 143.600 ; 
                RECT 75.280 143.280 83.080 143.600 ; 
                RECT 88.880 143.280 199.360 143.600 ; 
                RECT 301.040 143.280 310.520 143.600 ; 
                RECT 0.160 144.640 56.560 144.960 ; 
                RECT 75.280 144.640 80.360 144.960 ; 
                RECT 88.880 144.640 199.360 144.960 ; 
                RECT 301.040 144.640 310.520 144.960 ; 
                RECT 0.160 146.000 56.560 146.320 ; 
                RECT 75.280 146.000 199.360 146.320 ; 
                RECT 301.040 146.000 310.520 146.320 ; 
                RECT 0.160 147.360 56.560 147.680 ; 
                RECT 75.280 147.360 77.640 147.680 ; 
                RECT 88.880 147.360 199.360 147.680 ; 
                RECT 301.040 147.360 310.520 147.680 ; 
                RECT 0.160 148.720 56.560 149.040 ; 
                RECT 75.280 148.720 87.160 149.040 ; 
                RECT 95.000 148.720 199.360 149.040 ; 
                RECT 301.040 148.720 310.520 149.040 ; 
                RECT 0.160 150.080 56.560 150.400 ; 
                RECT 75.280 150.080 86.480 150.400 ; 
                RECT 88.880 150.080 199.360 150.400 ; 
                RECT 301.040 150.080 310.520 150.400 ; 
                RECT 0.160 151.440 56.560 151.760 ; 
                RECT 75.280 151.440 199.360 151.760 ; 
                RECT 301.040 151.440 310.520 151.760 ; 
                RECT 0.160 152.800 56.560 153.120 ; 
                RECT 75.280 152.800 87.160 153.120 ; 
                RECT 95.680 152.800 199.360 153.120 ; 
                RECT 301.040 152.800 310.520 153.120 ; 
                RECT 0.160 154.160 56.560 154.480 ; 
                RECT 75.280 154.160 84.440 154.480 ; 
                RECT 88.880 154.160 199.360 154.480 ; 
                RECT 301.040 154.160 310.520 154.480 ; 
                RECT 0.160 155.520 56.560 155.840 ; 
                RECT 75.280 155.520 86.480 155.840 ; 
                RECT 88.880 155.520 199.360 155.840 ; 
                RECT 301.040 155.520 310.520 155.840 ; 
                RECT 0.160 156.880 56.560 157.200 ; 
                RECT 75.280 156.880 199.360 157.200 ; 
                RECT 301.040 156.880 310.520 157.200 ; 
                RECT 0.160 158.240 56.560 158.560 ; 
                RECT 75.280 158.240 77.640 158.560 ; 
                RECT 100.440 158.240 199.360 158.560 ; 
                RECT 301.040 158.240 310.520 158.560 ; 
                RECT 0.160 159.600 56.560 159.920 ; 
                RECT 75.280 159.600 94.640 159.920 ; 
                RECT 101.800 159.600 199.360 159.920 ; 
                RECT 301.040 159.600 310.520 159.920 ; 
                RECT 0.160 160.960 56.560 161.280 ; 
                RECT 75.280 160.960 86.480 161.280 ; 
                RECT 88.880 160.960 98.720 161.280 ; 
                RECT 102.480 160.960 199.360 161.280 ; 
                RECT 301.040 160.960 310.520 161.280 ; 
                RECT 0.160 162.320 56.560 162.640 ; 
                RECT 75.280 162.320 78.320 162.640 ; 
                RECT 91.600 162.320 199.360 162.640 ; 
                RECT 301.040 162.320 310.520 162.640 ; 
                RECT 0.160 163.680 56.560 164.000 ; 
                RECT 75.280 163.680 87.160 164.000 ; 
                RECT 95.680 163.680 199.360 164.000 ; 
                RECT 301.040 163.680 310.520 164.000 ; 
                RECT 0.160 165.040 56.560 165.360 ; 
                RECT 75.280 165.040 84.440 165.360 ; 
                RECT 96.360 165.040 199.360 165.360 ; 
                RECT 301.040 165.040 310.520 165.360 ; 
                RECT 0.160 166.400 56.560 166.720 ; 
                RECT 75.280 166.400 199.360 166.720 ; 
                RECT 301.040 166.400 310.520 166.720 ; 
                RECT 0.160 167.760 56.560 168.080 ; 
                RECT 75.280 167.760 199.360 168.080 ; 
                RECT 301.040 167.760 310.520 168.080 ; 
                RECT 0.160 169.120 56.560 169.440 ; 
                RECT 75.280 169.120 80.360 169.440 ; 
                RECT 88.880 169.120 199.360 169.440 ; 
                RECT 301.040 169.120 310.520 169.440 ; 
                RECT 0.160 170.480 56.560 170.800 ; 
                RECT 75.280 170.480 80.360 170.800 ; 
                RECT 86.160 170.480 199.360 170.800 ; 
                RECT 301.040 170.480 310.520 170.800 ; 
                RECT 0.160 171.840 56.560 172.160 ; 
                RECT 75.280 171.840 199.360 172.160 ; 
                RECT 301.040 171.840 310.520 172.160 ; 
                RECT 0.160 173.200 56.560 173.520 ; 
                RECT 75.280 173.200 86.480 173.520 ; 
                RECT 88.880 173.200 199.360 173.520 ; 
                RECT 301.040 173.200 310.520 173.520 ; 
                RECT 0.160 174.560 56.560 174.880 ; 
                RECT 75.280 174.560 79.680 174.880 ; 
                RECT 95.000 174.560 199.360 174.880 ; 
                RECT 301.040 174.560 310.520 174.880 ; 
                RECT 0.160 175.920 56.560 176.240 ; 
                RECT 75.280 175.920 199.360 176.240 ; 
                RECT 301.040 175.920 310.520 176.240 ; 
                RECT 0.160 177.280 56.560 177.600 ; 
                RECT 75.280 177.280 86.480 177.600 ; 
                RECT 88.880 177.280 199.360 177.600 ; 
                RECT 301.040 177.280 310.520 177.600 ; 
                RECT 0.160 178.640 56.560 178.960 ; 
                RECT 75.280 178.640 81.720 178.960 ; 
                RECT 88.880 178.640 165.360 178.960 ; 
                RECT 171.160 178.640 199.360 178.960 ; 
                RECT 301.040 178.640 310.520 178.960 ; 
                RECT 0.160 180.000 56.560 180.320 ; 
                RECT 75.280 180.000 78.320 180.320 ; 
                RECT 85.480 180.000 87.160 180.320 ; 
                RECT 89.560 180.000 165.360 180.320 ; 
                RECT 171.160 180.000 199.360 180.320 ; 
                RECT 301.040 180.000 310.520 180.320 ; 
                RECT 0.160 181.360 56.560 181.680 ; 
                RECT 75.280 181.360 165.360 181.680 ; 
                RECT 171.160 181.360 199.360 181.680 ; 
                RECT 301.040 181.360 310.520 181.680 ; 
                RECT 0.160 182.720 56.560 183.040 ; 
                RECT 75.280 182.720 77.640 183.040 ; 
                RECT 95.680 182.720 165.360 183.040 ; 
                RECT 171.160 182.720 199.360 183.040 ; 
                RECT 301.040 182.720 310.520 183.040 ; 
                RECT 0.160 184.080 56.560 184.400 ; 
                RECT 88.200 184.080 199.360 184.400 ; 
                RECT 301.040 184.080 310.520 184.400 ; 
                RECT 0.160 185.440 56.560 185.760 ; 
                RECT 75.280 185.440 78.320 185.760 ; 
                RECT 91.600 185.440 199.360 185.760 ; 
                RECT 301.040 185.440 310.520 185.760 ; 
                RECT 0.160 186.800 56.560 187.120 ; 
                RECT 75.280 186.800 199.360 187.120 ; 
                RECT 301.040 186.800 310.520 187.120 ; 
                RECT 0.160 188.160 56.560 188.480 ; 
                RECT 75.280 188.160 199.360 188.480 ; 
                RECT 301.040 188.160 310.520 188.480 ; 
                RECT 0.160 189.520 56.560 189.840 ; 
                RECT 75.280 189.520 89.880 189.840 ; 
                RECT 96.360 189.520 130.680 189.840 ; 
                RECT 170.480 189.520 178.960 189.840 ; 
                RECT 301.040 189.520 310.520 189.840 ; 
                RECT 0.160 190.880 56.560 191.200 ; 
                RECT 75.280 190.880 93.280 191.200 ; 
                RECT 95.680 190.880 130.680 191.200 ; 
                RECT 170.480 190.880 178.960 191.200 ; 
                RECT 301.040 190.880 310.520 191.200 ; 
                RECT 0.160 192.240 56.560 192.560 ; 
                RECT 75.280 192.240 130.680 192.560 ; 
                RECT 170.480 192.240 181.680 192.560 ; 
                RECT 301.040 192.240 310.520 192.560 ; 
                RECT 0.160 193.600 56.560 193.920 ; 
                RECT 75.280 193.600 80.360 193.920 ; 
                RECT 83.440 193.600 130.680 193.920 ; 
                RECT 170.480 193.600 184.400 193.920 ; 
                RECT 301.040 193.600 310.520 193.920 ; 
                RECT 0.160 194.960 56.560 195.280 ; 
                RECT 75.280 194.960 77.640 195.280 ; 
                RECT 82.080 194.960 130.680 195.280 ; 
                RECT 170.480 194.960 187.120 195.280 ; 
                RECT 301.040 194.960 310.520 195.280 ; 
                RECT 0.160 196.320 56.560 196.640 ; 
                RECT 75.280 196.320 130.680 196.640 ; 
                RECT 170.480 196.320 192.560 196.640 ; 
                RECT 301.040 196.320 310.520 196.640 ; 
                RECT 0.160 197.680 56.560 198.000 ; 
                RECT 75.280 197.680 130.680 198.000 ; 
                RECT 170.480 197.680 195.280 198.000 ; 
                RECT 301.040 197.680 310.520 198.000 ; 
                RECT 0.160 199.040 56.560 199.360 ; 
                RECT 75.280 199.040 130.680 199.360 ; 
                RECT 170.480 199.040 198.000 199.360 ; 
                RECT 301.040 199.040 310.520 199.360 ; 
                RECT 0.160 200.400 56.560 200.720 ; 
                RECT 75.280 200.400 130.680 200.720 ; 
                RECT 301.040 200.400 310.520 200.720 ; 
                RECT 0.160 201.760 56.560 202.080 ; 
                RECT 75.280 201.760 83.080 202.080 ; 
                RECT 95.680 201.760 130.680 202.080 ; 
                RECT 170.480 201.760 199.360 202.080 ; 
                RECT 301.040 201.760 310.520 202.080 ; 
                RECT 0.160 203.120 56.560 203.440 ; 
                RECT 75.280 203.120 80.360 203.440 ; 
                RECT 84.800 203.120 130.680 203.440 ; 
                RECT 170.480 203.120 199.360 203.440 ; 
                RECT 301.040 203.120 310.520 203.440 ; 
                RECT 0.160 204.480 56.560 204.800 ; 
                RECT 75.280 204.480 130.680 204.800 ; 
                RECT 170.480 204.480 199.360 204.800 ; 
                RECT 301.040 204.480 310.520 204.800 ; 
                RECT 0.160 205.840 56.560 206.160 ; 
                RECT 75.280 205.840 130.680 206.160 ; 
                RECT 170.480 205.840 199.360 206.160 ; 
                RECT 301.040 205.840 310.520 206.160 ; 
                RECT 0.160 207.200 56.560 207.520 ; 
                RECT 75.280 207.200 130.680 207.520 ; 
                RECT 170.480 207.200 199.360 207.520 ; 
                RECT 301.040 207.200 310.520 207.520 ; 
                RECT 0.160 208.560 56.560 208.880 ; 
                RECT 75.280 208.560 83.080 208.880 ; 
                RECT 85.480 208.560 130.680 208.880 ; 
                RECT 170.480 208.560 199.360 208.880 ; 
                RECT 301.040 208.560 310.520 208.880 ; 
                RECT 0.160 209.920 56.560 210.240 ; 
                RECT 75.280 209.920 79.680 210.240 ; 
                RECT 82.760 209.920 93.280 210.240 ; 
                RECT 96.360 209.920 130.680 210.240 ; 
                RECT 170.480 209.920 199.360 210.240 ; 
                RECT 301.040 209.920 310.520 210.240 ; 
                RECT 0.160 211.280 56.560 211.600 ; 
                RECT 75.280 211.280 130.680 211.600 ; 
                RECT 170.480 211.280 199.360 211.600 ; 
                RECT 301.040 211.280 310.520 211.600 ; 
                RECT 0.160 212.640 56.560 212.960 ; 
                RECT 75.280 212.640 130.680 212.960 ; 
                RECT 170.480 212.640 199.360 212.960 ; 
                RECT 301.040 212.640 310.520 212.960 ; 
                RECT 0.160 214.000 56.560 214.320 ; 
                RECT 75.280 214.000 130.680 214.320 ; 
                RECT 170.480 214.000 199.360 214.320 ; 
                RECT 301.040 214.000 310.520 214.320 ; 
                RECT 0.160 215.360 56.560 215.680 ; 
                RECT 75.280 215.360 130.680 215.680 ; 
                RECT 170.480 215.360 199.360 215.680 ; 
                RECT 301.040 215.360 310.520 215.680 ; 
                RECT 0.160 216.720 130.680 217.040 ; 
                RECT 170.480 216.720 199.360 217.040 ; 
                RECT 301.040 216.720 310.520 217.040 ; 
                RECT 0.160 218.080 130.680 218.400 ; 
                RECT 170.480 218.080 199.360 218.400 ; 
                RECT 301.040 218.080 310.520 218.400 ; 
                RECT 0.160 219.440 81.720 219.760 ; 
                RECT 95.000 219.440 130.680 219.760 ; 
                RECT 170.480 219.440 199.360 219.760 ; 
                RECT 301.040 219.440 310.520 219.760 ; 
                RECT 0.160 220.800 35.480 221.120 ; 
                RECT 56.240 220.800 130.680 221.120 ; 
                RECT 170.480 220.800 199.360 221.120 ; 
                RECT 301.040 220.800 310.520 221.120 ; 
                RECT 0.160 222.160 35.480 222.480 ; 
                RECT 56.240 222.160 130.680 222.480 ; 
                RECT 170.480 222.160 199.360 222.480 ; 
                RECT 301.040 222.160 310.520 222.480 ; 
                RECT 0.160 223.520 35.480 223.840 ; 
                RECT 56.240 223.520 62.680 223.840 ; 
                RECT 69.840 223.520 130.680 223.840 ; 
                RECT 170.480 223.520 199.360 223.840 ; 
                RECT 301.040 223.520 310.520 223.840 ; 
                RECT 0.160 224.880 83.760 225.200 ; 
                RECT 89.560 224.880 130.680 225.200 ; 
                RECT 170.480 224.880 199.360 225.200 ; 
                RECT 301.040 224.880 310.520 225.200 ; 
                RECT 0.160 226.240 35.480 226.560 ; 
                RECT 56.240 226.240 57.240 226.560 ; 
                RECT 74.600 226.240 130.680 226.560 ; 
                RECT 170.480 226.240 199.360 226.560 ; 
                RECT 301.040 226.240 310.520 226.560 ; 
                RECT 0.160 227.600 35.480 227.920 ; 
                RECT 56.240 227.600 57.240 227.920 ; 
                RECT 74.600 227.600 130.680 227.920 ; 
                RECT 170.480 227.600 199.360 227.920 ; 
                RECT 301.040 227.600 310.520 227.920 ; 
                RECT 0.160 228.960 35.480 229.280 ; 
                RECT 56.240 228.960 130.680 229.280 ; 
                RECT 301.040 228.960 310.520 229.280 ; 
                RECT 0.160 230.320 21.200 230.640 ; 
                RECT 69.840 230.320 78.320 230.640 ; 
                RECT 88.200 230.320 130.680 230.640 ; 
                RECT 170.480 230.320 199.360 230.640 ; 
                RECT 301.040 230.320 310.520 230.640 ; 
                RECT 0.160 231.680 62.680 232.000 ; 
                RECT 82.760 231.680 310.520 232.000 ; 
                RECT 0.160 233.040 80.360 233.360 ; 
                RECT 84.120 233.040 310.520 233.360 ; 
                RECT 0.160 234.400 196.640 234.720 ; 
                RECT 303.760 234.400 310.520 234.720 ; 
                RECT 0.160 235.760 196.640 236.080 ; 
                RECT 303.760 235.760 310.520 236.080 ; 
                RECT 0.160 237.120 78.320 237.440 ; 
                RECT 84.800 237.120 155.840 237.440 ; 
                RECT 303.760 237.120 310.520 237.440 ; 
                RECT 0.160 238.480 76.280 238.800 ; 
                RECT 101.120 238.480 155.840 238.800 ; 
                RECT 303.760 238.480 310.520 238.800 ; 
                RECT 0.160 239.840 76.280 240.160 ; 
                RECT 99.760 239.840 112.320 240.160 ; 
                RECT 114.040 239.840 127.280 240.160 ; 
                RECT 145.320 239.840 155.840 240.160 ; 
                RECT 303.760 239.840 310.520 240.160 ; 
                RECT 0.160 241.200 112.320 241.520 ; 
                RECT 114.040 241.200 127.280 241.520 ; 
                RECT 145.320 241.200 155.840 241.520 ; 
                RECT 303.760 241.200 310.520 241.520 ; 
                RECT 0.160 242.560 76.280 242.880 ; 
                RECT 86.840 242.560 112.320 242.880 ; 
                RECT 117.440 242.560 127.280 242.880 ; 
                RECT 145.320 242.560 155.840 242.880 ; 
                RECT 303.760 242.560 310.520 242.880 ; 
                RECT 0.160 243.920 112.320 244.240 ; 
                RECT 117.440 243.920 127.280 244.240 ; 
                RECT 145.320 243.920 155.840 244.240 ; 
                RECT 303.760 243.920 310.520 244.240 ; 
                RECT 0.160 245.280 76.280 245.600 ; 
                RECT 86.840 245.280 112.320 245.600 ; 
                RECT 118.120 245.280 127.280 245.600 ; 
                RECT 145.320 245.280 155.840 245.600 ; 
                RECT 303.760 245.280 310.520 245.600 ; 
                RECT 0.160 246.640 76.280 246.960 ; 
                RECT 86.840 246.640 155.840 246.960 ; 
                RECT 303.760 246.640 310.520 246.960 ; 
                RECT 0.160 248.000 127.280 248.320 ; 
                RECT 145.320 248.000 155.840 248.320 ; 
                RECT 303.760 248.000 310.520 248.320 ; 
                RECT 0.160 249.360 127.280 249.680 ; 
                RECT 145.320 249.360 155.840 249.680 ; 
                RECT 303.760 249.360 310.520 249.680 ; 
                RECT 0.160 250.720 127.280 251.040 ; 
                RECT 145.320 250.720 155.840 251.040 ; 
                RECT 303.760 250.720 310.520 251.040 ; 
                RECT 0.160 252.080 20.520 252.400 ; 
                RECT 71.880 252.080 85.120 252.400 ; 
                RECT 88.200 252.080 127.280 252.400 ; 
                RECT 145.320 252.080 155.840 252.400 ; 
                RECT 303.760 252.080 310.520 252.400 ; 
                RECT 0.160 253.440 19.840 253.760 ; 
                RECT 71.880 253.440 89.880 253.760 ; 
                RECT 101.120 253.440 127.280 253.760 ; 
                RECT 138.520 253.440 155.840 253.760 ; 
                RECT 303.760 253.440 310.520 253.760 ; 
                RECT 0.160 254.800 19.160 255.120 ; 
                RECT 71.880 254.800 91.240 255.120 ; 
                RECT 100.440 254.800 139.520 255.120 ; 
                RECT 145.320 254.800 155.840 255.120 ; 
                RECT 303.760 254.800 310.520 255.120 ; 
                RECT 0.160 256.160 18.480 256.480 ; 
                RECT 71.880 256.160 112.320 256.480 ; 
                RECT 114.720 256.160 127.280 256.480 ; 
                RECT 145.320 256.160 155.840 256.480 ; 
                RECT 303.760 256.160 310.520 256.480 ; 
                RECT 0.160 257.520 112.320 257.840 ; 
                RECT 115.400 257.520 127.280 257.840 ; 
                RECT 145.320 257.520 155.840 257.840 ; 
                RECT 303.760 257.520 310.520 257.840 ; 
                RECT 0.160 258.880 17.800 259.200 ; 
                RECT 71.880 258.880 112.320 259.200 ; 
                RECT 115.400 258.880 127.280 259.200 ; 
                RECT 145.320 258.880 155.840 259.200 ; 
                RECT 303.760 258.880 310.520 259.200 ; 
                RECT 0.160 260.240 17.120 260.560 ; 
                RECT 71.880 260.240 112.320 260.560 ; 
                RECT 114.040 260.240 127.280 260.560 ; 
                RECT 145.320 260.240 155.840 260.560 ; 
                RECT 303.760 260.240 310.520 260.560 ; 
                RECT 0.160 261.600 112.320 261.920 ; 
                RECT 116.080 261.600 127.280 261.920 ; 
                RECT 138.520 261.600 155.840 261.920 ; 
                RECT 303.760 261.600 310.520 261.920 ; 
                RECT 0.160 262.960 16.440 263.280 ; 
                RECT 71.880 262.960 85.120 263.280 ; 
                RECT 92.280 262.960 127.280 263.280 ; 
                RECT 145.320 262.960 155.840 263.280 ; 
                RECT 303.760 262.960 310.520 263.280 ; 
                RECT 0.160 264.320 15.760 264.640 ; 
                RECT 71.880 264.320 85.120 264.640 ; 
                RECT 92.960 264.320 127.280 264.640 ; 
                RECT 145.320 264.320 155.840 264.640 ; 
                RECT 303.760 264.320 310.520 264.640 ; 
                RECT 0.160 265.680 127.280 266.000 ; 
                RECT 145.320 265.680 155.840 266.000 ; 
                RECT 303.760 265.680 310.520 266.000 ; 
                RECT 0.160 267.040 15.080 267.360 ; 
                RECT 71.880 267.040 85.120 267.360 ; 
                RECT 92.960 267.040 127.280 267.360 ; 
                RECT 145.320 267.040 155.840 267.360 ; 
                RECT 303.760 267.040 310.520 267.360 ; 
                RECT 0.160 268.400 14.400 268.720 ; 
                RECT 71.880 268.400 85.120 268.720 ; 
                RECT 92.280 268.400 127.280 268.720 ; 
                RECT 145.320 268.400 155.840 268.720 ; 
                RECT 303.760 268.400 310.520 268.720 ; 
                RECT 0.160 269.760 13.720 270.080 ; 
                RECT 71.880 269.760 155.840 270.080 ; 
                RECT 303.760 269.760 310.520 270.080 ; 
                RECT 0.160 271.120 13.040 271.440 ; 
                RECT 71.880 271.120 127.280 271.440 ; 
                RECT 145.320 271.120 155.840 271.440 ; 
                RECT 303.760 271.120 310.520 271.440 ; 
                RECT 0.160 272.480 127.280 272.800 ; 
                RECT 145.320 272.480 155.840 272.800 ; 
                RECT 303.760 272.480 310.520 272.800 ; 
                RECT 0.160 273.840 12.360 274.160 ; 
                RECT 71.880 273.840 127.280 274.160 ; 
                RECT 145.320 273.840 155.840 274.160 ; 
                RECT 303.760 273.840 310.520 274.160 ; 
                RECT 0.160 275.200 11.680 275.520 ; 
                RECT 71.880 275.200 127.280 275.520 ; 
                RECT 145.320 275.200 155.840 275.520 ; 
                RECT 303.760 275.200 310.520 275.520 ; 
                RECT 0.160 276.560 11.000 276.880 ; 
                RECT 71.880 276.560 127.280 276.880 ; 
                RECT 145.320 276.560 155.840 276.880 ; 
                RECT 303.760 276.560 310.520 276.880 ; 
                RECT 0.160 277.920 155.840 278.240 ; 
                RECT 303.760 277.920 310.520 278.240 ; 
                RECT 0.160 279.280 10.320 279.600 ; 
                RECT 71.880 279.280 85.120 279.600 ; 
                RECT 88.200 279.280 127.280 279.600 ; 
                RECT 145.320 279.280 155.840 279.600 ; 
                RECT 303.760 279.280 310.520 279.600 ; 
                RECT 0.160 280.640 127.280 280.960 ; 
                RECT 145.320 280.640 155.840 280.960 ; 
                RECT 303.760 280.640 310.520 280.960 ; 
                RECT 0.160 282.000 127.280 282.320 ; 
                RECT 145.320 282.000 155.840 282.320 ; 
                RECT 303.760 282.000 310.520 282.320 ; 
                RECT 0.160 283.360 127.280 283.680 ; 
                RECT 145.320 283.360 155.840 283.680 ; 
                RECT 303.760 283.360 310.520 283.680 ; 
                RECT 0.160 284.720 127.280 285.040 ; 
                RECT 145.320 284.720 155.840 285.040 ; 
                RECT 303.760 284.720 310.520 285.040 ; 
                RECT 0.160 286.080 155.840 286.400 ; 
                RECT 303.760 286.080 310.520 286.400 ; 
                RECT 0.160 287.440 127.280 287.760 ; 
                RECT 145.320 287.440 155.840 287.760 ; 
                RECT 303.760 287.440 310.520 287.760 ; 
                RECT 0.160 288.800 127.280 289.120 ; 
                RECT 145.320 288.800 155.840 289.120 ; 
                RECT 303.760 288.800 310.520 289.120 ; 
                RECT 0.160 290.160 127.280 290.480 ; 
                RECT 145.320 290.160 155.840 290.480 ; 
                RECT 303.760 290.160 310.520 290.480 ; 
                RECT 0.160 291.520 127.280 291.840 ; 
                RECT 145.320 291.520 155.840 291.840 ; 
                RECT 303.760 291.520 310.520 291.840 ; 
                RECT 0.160 292.880 127.280 293.200 ; 
                RECT 141.920 292.880 155.840 293.200 ; 
                RECT 303.760 292.880 310.520 293.200 ; 
                RECT 0.160 294.240 141.560 294.560 ; 
                RECT 145.320 294.240 155.840 294.560 ; 
                RECT 303.760 294.240 310.520 294.560 ; 
                RECT 0.160 295.600 127.280 295.920 ; 
                RECT 145.320 295.600 155.840 295.920 ; 
                RECT 303.760 295.600 310.520 295.920 ; 
                RECT 0.160 296.960 127.280 297.280 ; 
                RECT 145.320 296.960 155.840 297.280 ; 
                RECT 303.760 296.960 310.520 297.280 ; 
                RECT 0.160 298.320 127.280 298.640 ; 
                RECT 145.320 298.320 155.840 298.640 ; 
                RECT 303.760 298.320 310.520 298.640 ; 
                RECT 0.160 299.680 127.280 300.000 ; 
                RECT 145.320 299.680 155.840 300.000 ; 
                RECT 303.760 299.680 310.520 300.000 ; 
                RECT 0.160 301.040 127.280 301.360 ; 
                RECT 141.920 301.040 155.840 301.360 ; 
                RECT 303.760 301.040 310.520 301.360 ; 
                RECT 0.160 302.400 127.280 302.720 ; 
                RECT 145.320 302.400 155.840 302.720 ; 
                RECT 303.760 302.400 310.520 302.720 ; 
                RECT 0.160 303.760 127.280 304.080 ; 
                RECT 145.320 303.760 155.840 304.080 ; 
                RECT 303.760 303.760 310.520 304.080 ; 
                RECT 0.160 305.120 127.280 305.440 ; 
                RECT 145.320 305.120 155.840 305.440 ; 
                RECT 303.760 305.120 310.520 305.440 ; 
                RECT 0.160 306.480 127.280 306.800 ; 
                RECT 145.320 306.480 155.840 306.800 ; 
                RECT 303.760 306.480 310.520 306.800 ; 
                RECT 0.160 307.840 127.280 308.160 ; 
                RECT 145.320 307.840 155.840 308.160 ; 
                RECT 303.760 307.840 310.520 308.160 ; 
                RECT 0.160 309.200 155.840 309.520 ; 
                RECT 303.760 309.200 310.520 309.520 ; 
                RECT 0.160 310.560 127.280 310.880 ; 
                RECT 145.320 310.560 155.840 310.880 ; 
                RECT 303.760 310.560 310.520 310.880 ; 
                RECT 0.160 311.920 127.280 312.240 ; 
                RECT 145.320 311.920 155.840 312.240 ; 
                RECT 303.760 311.920 310.520 312.240 ; 
                RECT 0.160 313.280 127.280 313.600 ; 
                RECT 145.320 313.280 155.840 313.600 ; 
                RECT 303.760 313.280 310.520 313.600 ; 
                RECT 0.160 314.640 127.280 314.960 ; 
                RECT 145.320 314.640 155.840 314.960 ; 
                RECT 303.760 314.640 310.520 314.960 ; 
                RECT 0.160 316.000 127.280 316.320 ; 
                RECT 145.320 316.000 155.840 316.320 ; 
                RECT 303.760 316.000 310.520 316.320 ; 
                RECT 0.160 317.360 155.840 317.680 ; 
                RECT 303.760 317.360 310.520 317.680 ; 
                RECT 0.160 318.720 127.280 319.040 ; 
                RECT 145.320 318.720 155.840 319.040 ; 
                RECT 303.760 318.720 310.520 319.040 ; 
                RECT 0.160 320.080 127.280 320.400 ; 
                RECT 145.320 320.080 155.840 320.400 ; 
                RECT 303.760 320.080 310.520 320.400 ; 
                RECT 0.160 321.440 127.280 321.760 ; 
                RECT 145.320 321.440 155.840 321.760 ; 
                RECT 303.760 321.440 310.520 321.760 ; 
                RECT 0.160 322.800 127.280 323.120 ; 
                RECT 145.320 322.800 155.840 323.120 ; 
                RECT 303.760 322.800 310.520 323.120 ; 
                RECT 0.160 324.160 127.280 324.480 ; 
                RECT 145.320 324.160 155.840 324.480 ; 
                RECT 303.760 324.160 310.520 324.480 ; 
                RECT 0.160 325.520 155.840 325.840 ; 
                RECT 303.760 325.520 310.520 325.840 ; 
                RECT 0.160 326.880 127.280 327.200 ; 
                RECT 145.320 326.880 155.840 327.200 ; 
                RECT 303.760 326.880 310.520 327.200 ; 
                RECT 0.160 328.240 127.280 328.560 ; 
                RECT 145.320 328.240 155.840 328.560 ; 
                RECT 303.760 328.240 310.520 328.560 ; 
                RECT 0.160 329.600 127.280 329.920 ; 
                RECT 145.320 329.600 155.840 329.920 ; 
                RECT 303.760 329.600 310.520 329.920 ; 
                RECT 0.160 330.960 127.280 331.280 ; 
                RECT 145.320 330.960 155.840 331.280 ; 
                RECT 303.760 330.960 310.520 331.280 ; 
                RECT 0.160 332.320 127.280 332.640 ; 
                RECT 144.640 332.320 155.840 332.640 ; 
                RECT 303.760 332.320 310.520 332.640 ; 
                RECT 0.160 333.680 135.440 334.000 ; 
                RECT 145.320 333.680 155.840 334.000 ; 
                RECT 303.760 333.680 310.520 334.000 ; 
                RECT 0.160 335.040 129.320 335.360 ; 
                RECT 145.320 335.040 155.840 335.360 ; 
                RECT 303.760 335.040 310.520 335.360 ; 
                RECT 0.160 336.400 129.320 336.720 ; 
                RECT 145.320 336.400 155.840 336.720 ; 
                RECT 303.760 336.400 310.520 336.720 ; 
                RECT 0.160 337.760 129.320 338.080 ; 
                RECT 145.320 337.760 155.840 338.080 ; 
                RECT 303.760 337.760 310.520 338.080 ; 
                RECT 0.160 339.120 129.320 339.440 ; 
                RECT 145.320 339.120 155.840 339.440 ; 
                RECT 303.760 339.120 310.520 339.440 ; 
                RECT 0.160 340.480 91.920 340.800 ; 
                RECT 101.120 340.480 155.840 340.800 ; 
                RECT 303.760 340.480 310.520 340.800 ; 
                RECT 0.160 341.840 90.560 342.160 ; 
                RECT 100.440 341.840 112.320 342.160 ; 
                RECT 114.040 341.840 127.280 342.160 ; 
                RECT 145.320 341.840 155.840 342.160 ; 
                RECT 303.760 341.840 310.520 342.160 ; 
                RECT 0.160 343.200 112.320 343.520 ; 
                RECT 116.760 343.200 127.280 343.520 ; 
                RECT 145.320 343.200 155.840 343.520 ; 
                RECT 303.760 343.200 310.520 343.520 ; 
                RECT 0.160 344.560 112.320 344.880 ; 
                RECT 117.440 344.560 127.280 344.880 ; 
                RECT 145.320 344.560 155.840 344.880 ; 
                RECT 303.760 344.560 310.520 344.880 ; 
                RECT 0.160 345.920 112.320 346.240 ; 
                RECT 117.440 345.920 127.280 346.240 ; 
                RECT 145.320 345.920 155.840 346.240 ; 
                RECT 303.760 345.920 310.520 346.240 ; 
                RECT 0.160 347.280 112.320 347.600 ; 
                RECT 114.040 347.280 127.280 347.600 ; 
                RECT 145.320 347.280 155.840 347.600 ; 
                RECT 303.760 347.280 310.520 347.600 ; 
                RECT 0.160 348.640 155.840 348.960 ; 
                RECT 303.760 348.640 310.520 348.960 ; 
                RECT 0.160 350.000 127.280 350.320 ; 
                RECT 145.320 350.000 155.840 350.320 ; 
                RECT 303.760 350.000 310.520 350.320 ; 
                RECT 0.160 351.360 127.280 351.680 ; 
                RECT 145.320 351.360 155.840 351.680 ; 
                RECT 303.760 351.360 310.520 351.680 ; 
                RECT 0.160 352.720 127.280 353.040 ; 
                RECT 145.320 352.720 155.840 353.040 ; 
                RECT 303.760 352.720 310.520 353.040 ; 
                RECT 0.160 354.080 127.280 354.400 ; 
                RECT 145.320 354.080 155.840 354.400 ; 
                RECT 303.760 354.080 310.520 354.400 ; 
                RECT 0.160 355.440 127.280 355.760 ; 
                RECT 145.320 355.440 155.840 355.760 ; 
                RECT 303.760 355.440 310.520 355.760 ; 
                RECT 0.160 356.800 88.520 357.120 ; 
                RECT 101.120 356.800 155.840 357.120 ; 
                RECT 303.760 356.800 310.520 357.120 ; 
                RECT 0.160 358.160 87.160 358.480 ; 
                RECT 99.760 358.160 112.320 358.480 ; 
                RECT 114.040 358.160 127.280 358.480 ; 
                RECT 145.320 358.160 155.840 358.480 ; 
                RECT 303.760 358.160 310.520 358.480 ; 
                RECT 0.160 359.520 112.320 359.840 ; 
                RECT 114.720 359.520 127.280 359.840 ; 
                RECT 145.320 359.520 155.840 359.840 ; 
                RECT 303.760 359.520 310.520 359.840 ; 
                RECT 0.160 360.880 112.320 361.200 ; 
                RECT 115.400 360.880 127.280 361.200 ; 
                RECT 145.320 360.880 155.840 361.200 ; 
                RECT 303.760 360.880 310.520 361.200 ; 
                RECT 0.160 362.240 112.320 362.560 ; 
                RECT 115.400 362.240 127.280 362.560 ; 
                RECT 145.320 362.240 155.840 362.560 ; 
                RECT 303.760 362.240 310.520 362.560 ; 
                RECT 0.160 363.600 112.320 363.920 ; 
                RECT 116.080 363.600 127.280 363.920 ; 
                RECT 145.320 363.600 155.840 363.920 ; 
                RECT 303.760 363.600 310.520 363.920 ; 
                RECT 0.160 364.960 155.840 365.280 ; 
                RECT 303.760 364.960 310.520 365.280 ; 
                RECT 0.160 366.320 127.280 366.640 ; 
                RECT 145.320 366.320 155.840 366.640 ; 
                RECT 303.760 366.320 310.520 366.640 ; 
                RECT 0.160 367.680 127.280 368.000 ; 
                RECT 145.320 367.680 155.840 368.000 ; 
                RECT 303.760 367.680 310.520 368.000 ; 
                RECT 0.160 369.040 127.280 369.360 ; 
                RECT 145.320 369.040 155.840 369.360 ; 
                RECT 303.760 369.040 310.520 369.360 ; 
                RECT 0.160 370.400 127.280 370.720 ; 
                RECT 145.320 370.400 155.840 370.720 ; 
                RECT 303.760 370.400 310.520 370.720 ; 
                RECT 0.160 371.760 127.280 372.080 ; 
                RECT 132.400 371.760 155.840 372.080 ; 
                RECT 303.760 371.760 310.520 372.080 ; 
                RECT 0.160 373.120 155.840 373.440 ; 
                RECT 303.760 373.120 310.520 373.440 ; 
                RECT 0.160 374.480 127.280 374.800 ; 
                RECT 145.320 374.480 155.840 374.800 ; 
                RECT 303.760 374.480 310.520 374.800 ; 
                RECT 0.160 375.840 127.280 376.160 ; 
                RECT 145.320 375.840 155.840 376.160 ; 
                RECT 303.760 375.840 310.520 376.160 ; 
                RECT 0.160 377.200 127.280 377.520 ; 
                RECT 145.320 377.200 155.840 377.520 ; 
                RECT 303.760 377.200 310.520 377.520 ; 
                RECT 0.160 378.560 127.280 378.880 ; 
                RECT 145.320 378.560 155.840 378.880 ; 
                RECT 303.760 378.560 310.520 378.880 ; 
                RECT 0.160 379.920 127.280 380.240 ; 
                RECT 132.400 379.920 155.840 380.240 ; 
                RECT 303.760 379.920 310.520 380.240 ; 
                RECT 0.160 381.280 127.280 381.600 ; 
                RECT 145.320 381.280 155.840 381.600 ; 
                RECT 303.760 381.280 310.520 381.600 ; 
                RECT 0.160 382.640 127.280 382.960 ; 
                RECT 145.320 382.640 155.840 382.960 ; 
                RECT 303.760 382.640 310.520 382.960 ; 
                RECT 0.160 384.000 127.280 384.320 ; 
                RECT 145.320 384.000 155.840 384.320 ; 
                RECT 303.760 384.000 310.520 384.320 ; 
                RECT 0.160 385.360 127.280 385.680 ; 
                RECT 145.320 385.360 155.840 385.680 ; 
                RECT 303.760 385.360 310.520 385.680 ; 
                RECT 0.160 386.720 127.280 387.040 ; 
                RECT 145.320 386.720 155.840 387.040 ; 
                RECT 303.760 386.720 310.520 387.040 ; 
                RECT 0.160 388.080 127.280 388.400 ; 
                RECT 133.080 388.080 155.840 388.400 ; 
                RECT 303.760 388.080 310.520 388.400 ; 
                RECT 0.160 389.440 127.280 389.760 ; 
                RECT 145.320 389.440 155.840 389.760 ; 
                RECT 303.760 389.440 310.520 389.760 ; 
                RECT 0.160 390.800 127.280 391.120 ; 
                RECT 145.320 390.800 155.840 391.120 ; 
                RECT 303.760 390.800 310.520 391.120 ; 
                RECT 0.160 392.160 127.280 392.480 ; 
                RECT 145.320 392.160 155.840 392.480 ; 
                RECT 303.760 392.160 310.520 392.480 ; 
                RECT 0.160 393.520 127.280 393.840 ; 
                RECT 145.320 393.520 155.840 393.840 ; 
                RECT 303.760 393.520 310.520 393.840 ; 
                RECT 0.160 394.880 127.280 395.200 ; 
                RECT 145.320 394.880 155.840 395.200 ; 
                RECT 303.760 394.880 310.520 395.200 ; 
                RECT 0.160 396.240 155.840 396.560 ; 
                RECT 303.760 396.240 310.520 396.560 ; 
                RECT 0.160 397.600 127.280 397.920 ; 
                RECT 145.320 397.600 155.840 397.920 ; 
                RECT 303.760 397.600 310.520 397.920 ; 
                RECT 0.160 398.960 127.280 399.280 ; 
                RECT 145.320 398.960 155.840 399.280 ; 
                RECT 303.760 398.960 310.520 399.280 ; 
                RECT 0.160 400.320 127.280 400.640 ; 
                RECT 145.320 400.320 155.840 400.640 ; 
                RECT 303.760 400.320 310.520 400.640 ; 
                RECT 0.160 401.680 127.280 402.000 ; 
                RECT 145.320 401.680 155.840 402.000 ; 
                RECT 303.760 401.680 310.520 402.000 ; 
                RECT 0.160 403.040 127.280 403.360 ; 
                RECT 145.320 403.040 155.840 403.360 ; 
                RECT 303.760 403.040 310.520 403.360 ; 
                RECT 0.160 404.400 155.840 404.720 ; 
                RECT 303.760 404.400 310.520 404.720 ; 
                RECT 0.160 405.760 127.280 406.080 ; 
                RECT 145.320 405.760 155.840 406.080 ; 
                RECT 303.760 405.760 310.520 406.080 ; 
                RECT 0.160 407.120 127.280 407.440 ; 
                RECT 145.320 407.120 155.840 407.440 ; 
                RECT 303.760 407.120 310.520 407.440 ; 
                RECT 0.160 408.480 127.280 408.800 ; 
                RECT 145.320 408.480 155.840 408.800 ; 
                RECT 303.760 408.480 310.520 408.800 ; 
                RECT 0.160 409.840 127.280 410.160 ; 
                RECT 145.320 409.840 155.840 410.160 ; 
                RECT 303.760 409.840 310.520 410.160 ; 
                RECT 0.160 411.200 127.280 411.520 ; 
                RECT 145.320 411.200 155.840 411.520 ; 
                RECT 303.760 411.200 310.520 411.520 ; 
                RECT 0.160 412.560 155.840 412.880 ; 
                RECT 303.760 412.560 310.520 412.880 ; 
                RECT 0.160 413.920 127.280 414.240 ; 
                RECT 145.320 413.920 155.840 414.240 ; 
                RECT 303.760 413.920 310.520 414.240 ; 
                RECT 0.160 415.280 127.280 415.600 ; 
                RECT 145.320 415.280 155.840 415.600 ; 
                RECT 303.760 415.280 310.520 415.600 ; 
                RECT 0.160 416.640 127.280 416.960 ; 
                RECT 145.320 416.640 155.840 416.960 ; 
                RECT 303.760 416.640 310.520 416.960 ; 
                RECT 0.160 418.000 127.280 418.320 ; 
                RECT 145.320 418.000 155.840 418.320 ; 
                RECT 303.760 418.000 310.520 418.320 ; 
                RECT 0.160 419.360 127.280 419.680 ; 
                RECT 135.800 419.360 155.840 419.680 ; 
                RECT 303.760 419.360 310.520 419.680 ; 
                RECT 0.160 420.720 141.560 421.040 ; 
                RECT 145.320 420.720 155.840 421.040 ; 
                RECT 303.760 420.720 310.520 421.040 ; 
                RECT 0.160 422.080 127.280 422.400 ; 
                RECT 145.320 422.080 155.840 422.400 ; 
                RECT 303.760 422.080 310.520 422.400 ; 
                RECT 0.160 423.440 127.280 423.760 ; 
                RECT 145.320 423.440 155.840 423.760 ; 
                RECT 303.760 423.440 310.520 423.760 ; 
                RECT 0.160 424.800 127.280 425.120 ; 
                RECT 145.320 424.800 155.840 425.120 ; 
                RECT 303.760 424.800 310.520 425.120 ; 
                RECT 0.160 426.160 127.280 426.480 ; 
                RECT 145.320 426.160 155.840 426.480 ; 
                RECT 303.760 426.160 310.520 426.480 ; 
                RECT 0.160 427.520 127.280 427.840 ; 
                RECT 136.480 427.520 155.840 427.840 ; 
                RECT 303.760 427.520 310.520 427.840 ; 
                RECT 0.160 428.880 127.280 429.200 ; 
                RECT 145.320 428.880 155.840 429.200 ; 
                RECT 303.760 428.880 310.520 429.200 ; 
                RECT 0.160 430.240 127.280 430.560 ; 
                RECT 145.320 430.240 155.840 430.560 ; 
                RECT 303.760 430.240 310.520 430.560 ; 
                RECT 0.160 431.600 127.280 431.920 ; 
                RECT 145.320 431.600 155.840 431.920 ; 
                RECT 303.760 431.600 310.520 431.920 ; 
                RECT 0.160 432.960 127.280 433.280 ; 
                RECT 145.320 432.960 155.840 433.280 ; 
                RECT 303.760 432.960 310.520 433.280 ; 
                RECT 0.160 434.320 127.280 434.640 ; 
                RECT 145.320 434.320 155.840 434.640 ; 
                RECT 303.760 434.320 310.520 434.640 ; 
                RECT 0.160 435.680 155.840 436.000 ; 
                RECT 303.760 435.680 310.520 436.000 ; 
                RECT 0.160 437.040 130.680 437.360 ; 
                RECT 145.320 437.040 155.840 437.360 ; 
                RECT 303.760 437.040 310.520 437.360 ; 
                RECT 0.160 438.400 130.680 438.720 ; 
                RECT 145.320 438.400 155.840 438.720 ; 
                RECT 303.760 438.400 310.520 438.720 ; 
                RECT 0.160 439.760 138.840 440.080 ; 
                RECT 145.320 439.760 155.840 440.080 ; 
                RECT 303.760 439.760 310.520 440.080 ; 
                RECT 0.160 441.120 130.680 441.440 ; 
                RECT 145.320 441.120 155.840 441.440 ; 
                RECT 303.760 441.120 310.520 441.440 ; 
                RECT 0.160 442.480 130.680 442.800 ; 
                RECT 145.320 442.480 155.840 442.800 ; 
                RECT 303.760 442.480 310.520 442.800 ; 
                RECT 0.160 443.840 155.840 444.160 ; 
                RECT 303.760 443.840 310.520 444.160 ; 
                RECT 0.160 445.200 130.680 445.520 ; 
                RECT 145.320 445.200 155.840 445.520 ; 
                RECT 303.760 445.200 310.520 445.520 ; 
                RECT 0.160 446.560 130.680 446.880 ; 
                RECT 145.320 446.560 155.840 446.880 ; 
                RECT 303.760 446.560 310.520 446.880 ; 
                RECT 0.160 447.920 130.680 448.240 ; 
                RECT 145.320 447.920 155.840 448.240 ; 
                RECT 303.760 447.920 310.520 448.240 ; 
                RECT 0.160 449.280 140.880 449.600 ; 
                RECT 145.320 449.280 155.840 449.600 ; 
                RECT 303.760 449.280 310.520 449.600 ; 
                RECT 0.160 450.640 130.680 450.960 ; 
                RECT 145.320 450.640 155.840 450.960 ; 
                RECT 303.760 450.640 310.520 450.960 ; 
                RECT 0.160 452.000 155.840 452.320 ; 
                RECT 303.760 452.000 310.520 452.320 ; 
                RECT 0.160 453.360 130.680 453.680 ; 
                RECT 145.320 453.360 155.840 453.680 ; 
                RECT 303.760 453.360 310.520 453.680 ; 
                RECT 0.160 454.720 130.680 455.040 ; 
                RECT 145.320 454.720 155.840 455.040 ; 
                RECT 303.760 454.720 310.520 455.040 ; 
                RECT 0.160 456.080 130.680 456.400 ; 
                RECT 145.320 456.080 155.840 456.400 ; 
                RECT 303.760 456.080 310.520 456.400 ; 
                RECT 0.160 457.440 130.680 457.760 ; 
                RECT 145.320 457.440 155.840 457.760 ; 
                RECT 303.760 457.440 310.520 457.760 ; 
                RECT 0.160 458.800 155.840 459.120 ; 
                RECT 303.760 458.800 310.520 459.120 ; 
                RECT 0.160 460.160 135.440 460.480 ; 
                RECT 145.320 460.160 155.840 460.480 ; 
                RECT 303.760 460.160 310.520 460.480 ; 
                RECT 0.160 461.520 131.360 461.840 ; 
                RECT 145.320 461.520 155.840 461.840 ; 
                RECT 303.760 461.520 310.520 461.840 ; 
                RECT 0.160 462.880 131.360 463.200 ; 
                RECT 145.320 462.880 155.840 463.200 ; 
                RECT 303.760 462.880 310.520 463.200 ; 
                RECT 0.160 464.240 131.360 464.560 ; 
                RECT 145.320 464.240 155.840 464.560 ; 
                RECT 303.760 464.240 310.520 464.560 ; 
                RECT 0.160 465.600 131.360 465.920 ; 
                RECT 145.320 465.600 155.840 465.920 ; 
                RECT 303.760 465.600 310.520 465.920 ; 
                RECT 0.160 466.960 155.840 467.280 ; 
                RECT 303.760 466.960 310.520 467.280 ; 
                RECT 0.160 468.320 137.480 468.640 ; 
                RECT 145.320 468.320 155.840 468.640 ; 
                RECT 303.760 468.320 310.520 468.640 ; 
                RECT 0.160 469.680 131.360 470.000 ; 
                RECT 145.320 469.680 155.840 470.000 ; 
                RECT 303.760 469.680 310.520 470.000 ; 
                RECT 0.160 471.040 131.360 471.360 ; 
                RECT 145.320 471.040 155.840 471.360 ; 
                RECT 303.760 471.040 310.520 471.360 ; 
                RECT 0.160 472.400 131.360 472.720 ; 
                RECT 145.320 472.400 155.840 472.720 ; 
                RECT 303.760 472.400 310.520 472.720 ; 
                RECT 0.160 473.760 131.360 474.080 ; 
                RECT 145.320 473.760 155.840 474.080 ; 
                RECT 303.760 473.760 310.520 474.080 ; 
                RECT 0.160 475.120 155.840 475.440 ; 
                RECT 303.760 475.120 310.520 475.440 ; 
                RECT 0.160 476.480 131.360 476.800 ; 
                RECT 145.320 476.480 155.840 476.800 ; 
                RECT 303.760 476.480 310.520 476.800 ; 
                RECT 0.160 477.840 140.200 478.160 ; 
                RECT 145.320 477.840 155.840 478.160 ; 
                RECT 303.760 477.840 310.520 478.160 ; 
                RECT 0.160 479.200 140.200 479.520 ; 
                RECT 145.320 479.200 155.840 479.520 ; 
                RECT 303.760 479.200 310.520 479.520 ; 
                RECT 0.160 480.560 131.360 480.880 ; 
                RECT 145.320 480.560 155.840 480.880 ; 
                RECT 303.760 480.560 310.520 480.880 ; 
                RECT 0.160 481.920 131.360 482.240 ; 
                RECT 145.320 481.920 155.840 482.240 ; 
                RECT 303.760 481.920 310.520 482.240 ; 
                RECT 0.160 483.280 155.840 483.600 ; 
                RECT 303.760 483.280 310.520 483.600 ; 
                RECT 0.160 484.640 131.360 484.960 ; 
                RECT 145.320 484.640 155.840 484.960 ; 
                RECT 303.760 484.640 310.520 484.960 ; 
                RECT 0.160 486.000 131.360 486.320 ; 
                RECT 145.320 486.000 155.840 486.320 ; 
                RECT 303.760 486.000 310.520 486.320 ; 
                RECT 0.160 487.360 142.240 487.680 ; 
                RECT 145.320 487.360 155.840 487.680 ; 
                RECT 303.760 487.360 310.520 487.680 ; 
                RECT 0.160 488.720 142.920 489.040 ; 
                RECT 145.320 488.720 155.840 489.040 ; 
                RECT 303.760 488.720 310.520 489.040 ; 
                RECT 0.160 490.080 131.360 490.400 ; 
                RECT 145.320 490.080 155.840 490.400 ; 
                RECT 303.760 490.080 310.520 490.400 ; 
                RECT 0.160 491.440 155.840 491.760 ; 
                RECT 303.760 491.440 310.520 491.760 ; 
                RECT 0.160 492.800 132.040 493.120 ; 
                RECT 145.320 492.800 155.840 493.120 ; 
                RECT 303.760 492.800 310.520 493.120 ; 
                RECT 0.160 494.160 132.040 494.480 ; 
                RECT 145.320 494.160 155.840 494.480 ; 
                RECT 303.760 494.160 310.520 494.480 ; 
                RECT 0.160 495.520 132.040 495.840 ; 
                RECT 145.320 495.520 155.840 495.840 ; 
                RECT 303.760 495.520 310.520 495.840 ; 
                RECT 0.160 496.880 132.040 497.200 ; 
                RECT 145.320 496.880 155.840 497.200 ; 
                RECT 303.760 496.880 310.520 497.200 ; 
                RECT 0.160 498.240 155.840 498.560 ; 
                RECT 303.760 498.240 310.520 498.560 ; 
                RECT 0.160 499.600 137.480 499.920 ; 
                RECT 145.320 499.600 155.840 499.920 ; 
                RECT 303.760 499.600 310.520 499.920 ; 
                RECT 0.160 500.960 132.040 501.280 ; 
                RECT 145.320 500.960 155.840 501.280 ; 
                RECT 303.760 500.960 310.520 501.280 ; 
                RECT 0.160 502.320 132.040 502.640 ; 
                RECT 145.320 502.320 155.840 502.640 ; 
                RECT 303.760 502.320 310.520 502.640 ; 
                RECT 0.160 503.680 132.040 504.000 ; 
                RECT 145.320 503.680 155.840 504.000 ; 
                RECT 303.760 503.680 310.520 504.000 ; 
                RECT 0.160 505.040 132.040 505.360 ; 
                RECT 145.320 505.040 155.840 505.360 ; 
                RECT 303.760 505.040 310.520 505.360 ; 
                RECT 0.160 506.400 155.840 506.720 ; 
                RECT 303.760 506.400 310.520 506.720 ; 
                RECT 0.160 507.760 139.520 508.080 ; 
                RECT 145.320 507.760 155.840 508.080 ; 
                RECT 303.760 507.760 310.520 508.080 ; 
                RECT 0.160 509.120 132.040 509.440 ; 
                RECT 145.320 509.120 155.840 509.440 ; 
                RECT 303.760 509.120 310.520 509.440 ; 
                RECT 0.160 510.480 132.040 510.800 ; 
                RECT 145.320 510.480 155.840 510.800 ; 
                RECT 303.760 510.480 310.520 510.800 ; 
                RECT 0.160 511.840 132.040 512.160 ; 
                RECT 145.320 511.840 155.840 512.160 ; 
                RECT 303.760 511.840 310.520 512.160 ; 
                RECT 0.160 513.200 132.040 513.520 ; 
                RECT 145.320 513.200 155.840 513.520 ; 
                RECT 303.760 513.200 310.520 513.520 ; 
                RECT 0.160 514.560 155.840 514.880 ; 
                RECT 303.760 514.560 310.520 514.880 ; 
                RECT 0.160 515.920 132.040 516.240 ; 
                RECT 145.320 515.920 155.840 516.240 ; 
                RECT 303.760 515.920 310.520 516.240 ; 
                RECT 0.160 517.280 142.240 517.600 ; 
                RECT 145.320 517.280 155.840 517.600 ; 
                RECT 303.760 517.280 310.520 517.600 ; 
                RECT 0.160 518.640 132.040 518.960 ; 
                RECT 145.320 518.640 155.840 518.960 ; 
                RECT 303.760 518.640 310.520 518.960 ; 
                RECT 0.160 520.000 132.040 520.320 ; 
                RECT 145.320 520.000 155.840 520.320 ; 
                RECT 303.760 520.000 310.520 520.320 ; 
                RECT 0.160 521.360 132.040 521.680 ; 
                RECT 145.320 521.360 155.840 521.680 ; 
                RECT 303.760 521.360 310.520 521.680 ; 
                RECT 0.160 522.720 155.840 523.040 ; 
                RECT 303.760 522.720 310.520 523.040 ; 
                RECT 0.160 524.080 132.040 524.400 ; 
                RECT 145.320 524.080 155.840 524.400 ; 
                RECT 303.760 524.080 310.520 524.400 ; 
                RECT 0.160 525.440 132.040 525.760 ; 
                RECT 145.320 525.440 155.840 525.760 ; 
                RECT 303.760 525.440 310.520 525.760 ; 
                RECT 0.160 526.800 136.800 527.120 ; 
                RECT 145.320 526.800 155.840 527.120 ; 
                RECT 303.760 526.800 310.520 527.120 ; 
                RECT 0.160 528.160 132.040 528.480 ; 
                RECT 145.320 528.160 155.840 528.480 ; 
                RECT 303.760 528.160 310.520 528.480 ; 
                RECT 0.160 529.520 132.040 529.840 ; 
                RECT 145.320 529.520 155.840 529.840 ; 
                RECT 303.760 529.520 310.520 529.840 ; 
                RECT 0.160 530.880 155.840 531.200 ; 
                RECT 303.760 530.880 310.520 531.200 ; 
                RECT 0.160 532.240 132.040 532.560 ; 
                RECT 145.320 532.240 155.840 532.560 ; 
                RECT 303.760 532.240 310.520 532.560 ; 
                RECT 0.160 533.600 132.040 533.920 ; 
                RECT 145.320 533.600 155.840 533.920 ; 
                RECT 303.760 533.600 310.520 533.920 ; 
                RECT 0.160 534.960 132.040 535.280 ; 
                RECT 145.320 534.960 155.840 535.280 ; 
                RECT 303.760 534.960 310.520 535.280 ; 
                RECT 0.160 536.320 138.840 536.640 ; 
                RECT 145.320 536.320 155.840 536.640 ; 
                RECT 303.760 536.320 310.520 536.640 ; 
                RECT 0.160 537.680 155.840 538.000 ; 
                RECT 303.760 537.680 310.520 538.000 ; 
                RECT 0.160 539.040 139.520 539.360 ; 
                RECT 145.320 539.040 155.840 539.360 ; 
                RECT 303.760 539.040 310.520 539.360 ; 
                RECT 0.160 540.400 132.040 540.720 ; 
                RECT 145.320 540.400 155.840 540.720 ; 
                RECT 303.760 540.400 310.520 540.720 ; 
                RECT 0.160 541.760 132.040 542.080 ; 
                RECT 145.320 541.760 155.840 542.080 ; 
                RECT 303.760 541.760 310.520 542.080 ; 
                RECT 0.160 543.120 132.040 543.440 ; 
                RECT 145.320 543.120 155.840 543.440 ; 
                RECT 303.760 543.120 310.520 543.440 ; 
                RECT 0.160 544.480 132.040 544.800 ; 
                RECT 145.320 544.480 155.840 544.800 ; 
                RECT 303.760 544.480 310.520 544.800 ; 
                RECT 0.160 545.840 155.840 546.160 ; 
                RECT 303.760 545.840 310.520 546.160 ; 
                RECT 0.160 547.200 141.560 547.520 ; 
                RECT 145.320 547.200 155.840 547.520 ; 
                RECT 303.760 547.200 310.520 547.520 ; 
                RECT 0.160 548.560 132.040 548.880 ; 
                RECT 145.320 548.560 155.840 548.880 ; 
                RECT 303.760 548.560 310.520 548.880 ; 
                RECT 0.160 549.920 132.040 550.240 ; 
                RECT 145.320 549.920 155.840 550.240 ; 
                RECT 303.760 549.920 310.520 550.240 ; 
                RECT 0.160 551.280 132.040 551.600 ; 
                RECT 145.320 551.280 155.840 551.600 ; 
                RECT 303.760 551.280 310.520 551.600 ; 
                RECT 0.160 552.640 132.040 552.960 ; 
                RECT 145.320 552.640 155.840 552.960 ; 
                RECT 303.760 552.640 310.520 552.960 ; 
                RECT 0.160 554.000 155.840 554.320 ; 
                RECT 303.760 554.000 310.520 554.320 ; 
                RECT 0.160 555.360 132.720 555.680 ; 
                RECT 145.320 555.360 155.840 555.680 ; 
                RECT 303.760 555.360 310.520 555.680 ; 
                RECT 0.160 556.720 136.120 557.040 ; 
                RECT 145.320 556.720 155.840 557.040 ; 
                RECT 303.760 556.720 310.520 557.040 ; 
                RECT 0.160 558.080 132.720 558.400 ; 
                RECT 145.320 558.080 155.840 558.400 ; 
                RECT 303.760 558.080 310.520 558.400 ; 
                RECT 0.160 559.440 132.720 559.760 ; 
                RECT 145.320 559.440 155.840 559.760 ; 
                RECT 303.760 559.440 310.520 559.760 ; 
                RECT 0.160 560.800 132.720 561.120 ; 
                RECT 145.320 560.800 155.840 561.120 ; 
                RECT 303.760 560.800 310.520 561.120 ; 
                RECT 0.160 562.160 155.840 562.480 ; 
                RECT 303.760 562.160 310.520 562.480 ; 
                RECT 0.160 563.520 132.720 563.840 ; 
                RECT 145.320 563.520 155.840 563.840 ; 
                RECT 303.760 563.520 310.520 563.840 ; 
                RECT 0.160 564.880 132.720 565.200 ; 
                RECT 145.320 564.880 155.840 565.200 ; 
                RECT 303.760 564.880 310.520 565.200 ; 
                RECT 0.160 566.240 138.840 566.560 ; 
                RECT 145.320 566.240 155.840 566.560 ; 
                RECT 303.760 566.240 310.520 566.560 ; 
                RECT 0.160 567.600 132.720 567.920 ; 
                RECT 145.320 567.600 155.840 567.920 ; 
                RECT 303.760 567.600 310.520 567.920 ; 
                RECT 0.160 568.960 132.720 569.280 ; 
                RECT 145.320 568.960 155.840 569.280 ; 
                RECT 303.760 568.960 310.520 569.280 ; 
                RECT 0.160 570.320 155.840 570.640 ; 
                RECT 303.760 570.320 310.520 570.640 ; 
                RECT 0.160 571.680 132.720 572.000 ; 
                RECT 145.320 571.680 155.840 572.000 ; 
                RECT 303.760 571.680 310.520 572.000 ; 
                RECT 0.160 573.040 132.720 573.360 ; 
                RECT 145.320 573.040 155.840 573.360 ; 
                RECT 303.760 573.040 310.520 573.360 ; 
                RECT 0.160 574.400 132.720 574.720 ; 
                RECT 145.320 574.400 155.840 574.720 ; 
                RECT 303.760 574.400 310.520 574.720 ; 
                RECT 0.160 575.760 140.880 576.080 ; 
                RECT 145.320 575.760 155.840 576.080 ; 
                RECT 303.760 575.760 310.520 576.080 ; 
                RECT 0.160 577.120 132.720 577.440 ; 
                RECT 145.320 577.120 155.840 577.440 ; 
                RECT 303.760 577.120 310.520 577.440 ; 
                RECT 0.160 578.480 155.840 578.800 ; 
                RECT 303.760 578.480 310.520 578.800 ; 
                RECT 0.160 579.840 132.720 580.160 ; 
                RECT 145.320 579.840 155.840 580.160 ; 
                RECT 303.760 579.840 310.520 580.160 ; 
                RECT 0.160 581.200 132.720 581.520 ; 
                RECT 145.320 581.200 155.840 581.520 ; 
                RECT 303.760 581.200 310.520 581.520 ; 
                RECT 0.160 582.560 132.720 582.880 ; 
                RECT 145.320 582.560 155.840 582.880 ; 
                RECT 303.760 582.560 310.520 582.880 ; 
                RECT 0.160 583.920 132.720 584.240 ; 
                RECT 145.320 583.920 155.840 584.240 ; 
                RECT 303.760 583.920 310.520 584.240 ; 
                RECT 0.160 585.280 155.840 585.600 ; 
                RECT 303.760 585.280 310.520 585.600 ; 
                RECT 0.160 586.640 135.440 586.960 ; 
                RECT 145.320 586.640 155.840 586.960 ; 
                RECT 303.760 586.640 310.520 586.960 ; 
                RECT 0.160 588.000 133.400 588.320 ; 
                RECT 145.320 588.000 155.840 588.320 ; 
                RECT 303.760 588.000 310.520 588.320 ; 
                RECT 0.160 589.360 133.400 589.680 ; 
                RECT 145.320 589.360 155.840 589.680 ; 
                RECT 303.760 589.360 310.520 589.680 ; 
                RECT 0.160 590.720 133.400 591.040 ; 
                RECT 145.320 590.720 155.840 591.040 ; 
                RECT 303.760 590.720 310.520 591.040 ; 
                RECT 0.160 592.080 133.400 592.400 ; 
                RECT 145.320 592.080 155.840 592.400 ; 
                RECT 303.760 592.080 310.520 592.400 ; 
                RECT 0.160 593.440 155.840 593.760 ; 
                RECT 303.760 593.440 310.520 593.760 ; 
                RECT 0.160 594.800 137.480 595.120 ; 
                RECT 145.320 594.800 155.840 595.120 ; 
                RECT 303.760 594.800 310.520 595.120 ; 
                RECT 0.160 596.160 138.160 596.480 ; 
                RECT 145.320 596.160 155.840 596.480 ; 
                RECT 303.760 596.160 310.520 596.480 ; 
                RECT 0.160 597.520 133.400 597.840 ; 
                RECT 145.320 597.520 155.840 597.840 ; 
                RECT 303.760 597.520 310.520 597.840 ; 
                RECT 0.160 598.880 133.400 599.200 ; 
                RECT 145.320 598.880 155.840 599.200 ; 
                RECT 303.760 598.880 310.520 599.200 ; 
                RECT 0.160 600.240 133.400 600.560 ; 
                RECT 145.320 600.240 155.840 600.560 ; 
                RECT 303.760 600.240 310.520 600.560 ; 
                RECT 0.160 601.600 155.840 601.920 ; 
                RECT 303.760 601.600 310.520 601.920 ; 
                RECT 0.160 602.960 133.400 603.280 ; 
                RECT 145.320 602.960 155.840 603.280 ; 
                RECT 303.760 602.960 310.520 603.280 ; 
                RECT 0.160 604.320 133.400 604.640 ; 
                RECT 145.320 604.320 155.840 604.640 ; 
                RECT 303.760 604.320 310.520 604.640 ; 
                RECT 0.160 605.680 140.200 606.000 ; 
                RECT 145.320 605.680 155.840 606.000 ; 
                RECT 303.760 605.680 310.520 606.000 ; 
                RECT 0.160 607.040 133.400 607.360 ; 
                RECT 145.320 607.040 155.840 607.360 ; 
                RECT 303.760 607.040 310.520 607.360 ; 
                RECT 0.160 608.400 133.400 608.720 ; 
                RECT 145.320 608.400 155.840 608.720 ; 
                RECT 303.760 608.400 310.520 608.720 ; 
                RECT 0.160 609.760 155.840 610.080 ; 
                RECT 303.760 609.760 310.520 610.080 ; 
                RECT 0.160 611.120 133.400 611.440 ; 
                RECT 145.320 611.120 155.840 611.440 ; 
                RECT 303.760 611.120 310.520 611.440 ; 
                RECT 0.160 612.480 133.400 612.800 ; 
                RECT 145.320 612.480 155.840 612.800 ; 
                RECT 303.760 612.480 310.520 612.800 ; 
                RECT 0.160 613.840 133.400 614.160 ; 
                RECT 145.320 613.840 155.840 614.160 ; 
                RECT 303.760 613.840 310.520 614.160 ; 
                RECT 0.160 615.200 142.920 615.520 ; 
                RECT 145.320 615.200 155.840 615.520 ; 
                RECT 303.760 615.200 310.520 615.520 ; 
                RECT 0.160 616.560 133.400 616.880 ; 
                RECT 145.320 616.560 155.840 616.880 ; 
                RECT 303.760 616.560 310.520 616.880 ; 
                RECT 0.160 617.920 155.840 618.240 ; 
                RECT 303.760 617.920 310.520 618.240 ; 
                RECT 0.160 619.280 134.080 619.600 ; 
                RECT 145.320 619.280 155.840 619.600 ; 
                RECT 303.760 619.280 310.520 619.600 ; 
                RECT 0.160 620.640 134.080 620.960 ; 
                RECT 145.320 620.640 155.840 620.960 ; 
                RECT 303.760 620.640 310.520 620.960 ; 
                RECT 0.160 622.000 134.080 622.320 ; 
                RECT 145.320 622.000 155.840 622.320 ; 
                RECT 303.760 622.000 310.520 622.320 ; 
                RECT 0.160 623.360 134.080 623.680 ; 
                RECT 145.320 623.360 155.840 623.680 ; 
                RECT 303.760 623.360 310.520 623.680 ; 
                RECT 0.160 624.720 155.840 625.040 ; 
                RECT 303.760 624.720 310.520 625.040 ; 
                RECT 0.160 626.080 137.480 626.400 ; 
                RECT 145.320 626.080 155.840 626.400 ; 
                RECT 303.760 626.080 310.520 626.400 ; 
                RECT 0.160 627.440 134.080 627.760 ; 
                RECT 145.320 627.440 155.840 627.760 ; 
                RECT 303.760 627.440 310.520 627.760 ; 
                RECT 0.160 628.800 134.080 629.120 ; 
                RECT 145.320 628.800 155.840 629.120 ; 
                RECT 303.760 628.800 310.520 629.120 ; 
                RECT 0.160 630.160 134.080 630.480 ; 
                RECT 145.320 630.160 155.840 630.480 ; 
                RECT 303.760 630.160 310.520 630.480 ; 
                RECT 0.160 631.520 134.080 631.840 ; 
                RECT 145.320 631.520 155.840 631.840 ; 
                RECT 303.760 631.520 310.520 631.840 ; 
                RECT 0.160 632.880 155.840 633.200 ; 
                RECT 303.760 632.880 310.520 633.200 ; 
                RECT 0.160 634.240 139.520 634.560 ; 
                RECT 145.320 634.240 155.840 634.560 ; 
                RECT 303.760 634.240 310.520 634.560 ; 
                RECT 0.160 635.600 134.080 635.920 ; 
                RECT 145.320 635.600 155.840 635.920 ; 
                RECT 303.760 635.600 310.520 635.920 ; 
                RECT 0.160 636.960 134.080 637.280 ; 
                RECT 145.320 636.960 155.840 637.280 ; 
                RECT 303.760 636.960 310.520 637.280 ; 
                RECT 0.160 638.320 134.080 638.640 ; 
                RECT 145.320 638.320 155.840 638.640 ; 
                RECT 303.760 638.320 310.520 638.640 ; 
                RECT 0.160 639.680 134.080 640.000 ; 
                RECT 145.320 639.680 155.840 640.000 ; 
                RECT 303.760 639.680 310.520 640.000 ; 
                RECT 0.160 641.040 155.840 641.360 ; 
                RECT 303.760 641.040 310.520 641.360 ; 
                RECT 0.160 642.400 134.080 642.720 ; 
                RECT 145.320 642.400 155.840 642.720 ; 
                RECT 303.760 642.400 310.520 642.720 ; 
                RECT 0.160 643.760 142.240 644.080 ; 
                RECT 145.320 643.760 155.840 644.080 ; 
                RECT 303.760 643.760 310.520 644.080 ; 
                RECT 0.160 645.120 142.240 645.440 ; 
                RECT 145.320 645.120 155.840 645.440 ; 
                RECT 303.760 645.120 310.520 645.440 ; 
                RECT 0.160 646.480 134.080 646.800 ; 
                RECT 145.320 646.480 155.840 646.800 ; 
                RECT 303.760 646.480 310.520 646.800 ; 
                RECT 0.160 647.840 134.080 648.160 ; 
                RECT 145.320 647.840 155.840 648.160 ; 
                RECT 303.760 647.840 310.520 648.160 ; 
                RECT 0.160 649.200 155.840 649.520 ; 
                RECT 303.760 649.200 310.520 649.520 ; 
                RECT 0.160 650.560 134.080 650.880 ; 
                RECT 145.320 650.560 155.840 650.880 ; 
                RECT 303.760 650.560 310.520 650.880 ; 
                RECT 0.160 651.920 134.080 652.240 ; 
                RECT 145.320 651.920 155.840 652.240 ; 
                RECT 303.760 651.920 310.520 652.240 ; 
                RECT 0.160 653.280 134.080 653.600 ; 
                RECT 145.320 653.280 155.840 653.600 ; 
                RECT 303.760 653.280 310.520 653.600 ; 
                RECT 0.160 654.640 136.800 654.960 ; 
                RECT 145.320 654.640 155.840 654.960 ; 
                RECT 303.760 654.640 310.520 654.960 ; 
                RECT 0.160 656.000 134.080 656.320 ; 
                RECT 145.320 656.000 155.840 656.320 ; 
                RECT 303.760 656.000 310.520 656.320 ; 
                RECT 0.160 657.360 155.840 657.680 ; 
                RECT 303.760 657.360 310.520 657.680 ; 
                RECT 0.160 658.720 134.080 659.040 ; 
                RECT 145.320 658.720 155.840 659.040 ; 
                RECT 303.760 658.720 310.520 659.040 ; 
                RECT 0.160 660.080 134.080 660.400 ; 
                RECT 145.320 660.080 155.840 660.400 ; 
                RECT 303.760 660.080 310.520 660.400 ; 
                RECT 0.160 661.440 134.080 661.760 ; 
                RECT 145.320 661.440 155.840 661.760 ; 
                RECT 303.760 661.440 310.520 661.760 ; 
                RECT 0.160 662.800 134.080 663.120 ; 
                RECT 145.320 662.800 155.840 663.120 ; 
                RECT 303.760 662.800 310.520 663.120 ; 
                RECT 0.160 664.160 155.840 664.480 ; 
                RECT 303.760 664.160 310.520 664.480 ; 
                RECT 0.160 665.520 139.520 665.840 ; 
                RECT 145.320 665.520 155.840 665.840 ; 
                RECT 303.760 665.520 310.520 665.840 ; 
                RECT 0.160 666.880 134.080 667.200 ; 
                RECT 145.320 666.880 155.840 667.200 ; 
                RECT 303.760 666.880 310.520 667.200 ; 
                RECT 0.160 668.240 134.080 668.560 ; 
                RECT 145.320 668.240 155.840 668.560 ; 
                RECT 303.760 668.240 310.520 668.560 ; 
                RECT 0.160 669.600 134.080 669.920 ; 
                RECT 145.320 669.600 155.840 669.920 ; 
                RECT 303.760 669.600 310.520 669.920 ; 
                RECT 0.160 670.960 134.080 671.280 ; 
                RECT 145.320 670.960 155.840 671.280 ; 
                RECT 303.760 670.960 310.520 671.280 ; 
                RECT 0.160 672.320 155.840 672.640 ; 
                RECT 303.760 672.320 310.520 672.640 ; 
                RECT 0.160 673.680 141.560 674.000 ; 
                RECT 145.320 673.680 155.840 674.000 ; 
                RECT 303.760 673.680 310.520 674.000 ; 
                RECT 0.160 675.040 134.080 675.360 ; 
                RECT 145.320 675.040 155.840 675.360 ; 
                RECT 303.760 675.040 310.520 675.360 ; 
                RECT 0.160 676.400 134.080 676.720 ; 
                RECT 145.320 676.400 155.840 676.720 ; 
                RECT 303.760 676.400 310.520 676.720 ; 
                RECT 0.160 677.760 134.080 678.080 ; 
                RECT 145.320 677.760 155.840 678.080 ; 
                RECT 303.760 677.760 310.520 678.080 ; 
                RECT 0.160 679.120 134.080 679.440 ; 
                RECT 145.320 679.120 155.840 679.440 ; 
                RECT 303.760 679.120 310.520 679.440 ; 
                RECT 0.160 680.480 155.840 680.800 ; 
                RECT 303.760 680.480 310.520 680.800 ; 
                RECT 0.160 681.840 134.760 682.160 ; 
                RECT 145.320 681.840 155.840 682.160 ; 
                RECT 303.760 681.840 310.520 682.160 ; 
                RECT 0.160 683.200 136.120 683.520 ; 
                RECT 145.320 683.200 155.840 683.520 ; 
                RECT 303.760 683.200 310.520 683.520 ; 
                RECT 0.160 684.560 134.760 684.880 ; 
                RECT 145.320 684.560 155.840 684.880 ; 
                RECT 303.760 684.560 310.520 684.880 ; 
                RECT 0.160 685.920 134.760 686.240 ; 
                RECT 145.320 685.920 155.840 686.240 ; 
                RECT 303.760 685.920 310.520 686.240 ; 
                RECT 0.160 687.280 134.760 687.600 ; 
                RECT 145.320 687.280 155.840 687.600 ; 
                RECT 303.760 687.280 310.520 687.600 ; 
                RECT 0.160 688.640 155.840 688.960 ; 
                RECT 303.760 688.640 310.520 688.960 ; 
                RECT 0.160 690.000 134.760 690.320 ; 
                RECT 145.320 690.000 155.840 690.320 ; 
                RECT 303.760 690.000 310.520 690.320 ; 
                RECT 0.160 691.360 134.760 691.680 ; 
                RECT 145.320 691.360 155.840 691.680 ; 
                RECT 303.760 691.360 310.520 691.680 ; 
                RECT 0.160 692.720 138.840 693.040 ; 
                RECT 145.320 692.720 155.840 693.040 ; 
                RECT 303.760 692.720 310.520 693.040 ; 
                RECT 0.160 694.080 138.840 694.400 ; 
                RECT 145.320 694.080 155.840 694.400 ; 
                RECT 303.760 694.080 310.520 694.400 ; 
                RECT 0.160 695.440 134.760 695.760 ; 
                RECT 145.320 695.440 155.840 695.760 ; 
                RECT 303.760 695.440 310.520 695.760 ; 
                RECT 0.160 696.800 155.840 697.120 ; 
                RECT 303.760 696.800 310.520 697.120 ; 
                RECT 0.160 698.160 134.760 698.480 ; 
                RECT 145.320 698.160 155.840 698.480 ; 
                RECT 303.760 698.160 310.520 698.480 ; 
                RECT 0.160 699.520 134.760 699.840 ; 
                RECT 145.320 699.520 155.840 699.840 ; 
                RECT 303.760 699.520 310.520 699.840 ; 
                RECT 0.160 700.880 134.760 701.200 ; 
                RECT 145.320 700.880 155.840 701.200 ; 
                RECT 303.760 700.880 310.520 701.200 ; 
                RECT 0.160 702.240 140.880 702.560 ; 
                RECT 145.320 702.240 155.840 702.560 ; 
                RECT 303.760 702.240 310.520 702.560 ; 
                RECT 0.160 703.600 155.840 703.920 ; 
                RECT 303.760 703.600 310.520 703.920 ; 
                RECT 0.160 704.960 141.560 705.280 ; 
                RECT 145.320 704.960 155.840 705.280 ; 
                RECT 303.760 704.960 310.520 705.280 ; 
                RECT 0.160 706.320 134.760 706.640 ; 
                RECT 145.320 706.320 155.840 706.640 ; 
                RECT 303.760 706.320 310.520 706.640 ; 
                RECT 0.160 707.680 134.760 708.000 ; 
                RECT 145.320 707.680 155.840 708.000 ; 
                RECT 303.760 707.680 310.520 708.000 ; 
                RECT 0.160 709.040 134.760 709.360 ; 
                RECT 145.320 709.040 155.840 709.360 ; 
                RECT 303.760 709.040 310.520 709.360 ; 
                RECT 0.160 710.400 134.760 710.720 ; 
                RECT 145.320 710.400 155.840 710.720 ; 
                RECT 303.760 710.400 310.520 710.720 ; 
                RECT 0.160 711.760 155.840 712.080 ; 
                RECT 303.760 711.760 310.520 712.080 ; 
                RECT 0.160 713.120 135.440 713.440 ; 
                RECT 145.320 713.120 155.840 713.440 ; 
                RECT 303.760 713.120 310.520 713.440 ; 
                RECT 0.160 714.480 135.440 714.800 ; 
                RECT 145.320 714.480 155.840 714.800 ; 
                RECT 303.760 714.480 310.520 714.800 ; 
                RECT 0.160 715.840 135.440 716.160 ; 
                RECT 145.320 715.840 155.840 716.160 ; 
                RECT 303.760 715.840 310.520 716.160 ; 
                RECT 0.160 717.200 135.440 717.520 ; 
                RECT 145.320 717.200 155.840 717.520 ; 
                RECT 303.760 717.200 310.520 717.520 ; 
                RECT 0.160 718.560 135.440 718.880 ; 
                RECT 145.320 718.560 155.840 718.880 ; 
                RECT 303.760 718.560 310.520 718.880 ; 
                RECT 0.160 719.920 155.840 720.240 ; 
                RECT 303.760 719.920 310.520 720.240 ; 
                RECT 0.160 721.280 135.440 721.600 ; 
                RECT 145.320 721.280 155.840 721.600 ; 
                RECT 303.760 721.280 310.520 721.600 ; 
                RECT 0.160 722.640 138.160 722.960 ; 
                RECT 145.320 722.640 155.840 722.960 ; 
                RECT 303.760 722.640 310.520 722.960 ; 
                RECT 0.160 724.000 135.440 724.320 ; 
                RECT 145.320 724.000 155.840 724.320 ; 
                RECT 303.760 724.000 310.520 724.320 ; 
                RECT 0.160 725.360 135.440 725.680 ; 
                RECT 145.320 725.360 155.840 725.680 ; 
                RECT 303.760 725.360 310.520 725.680 ; 
                RECT 0.160 726.720 135.440 727.040 ; 
                RECT 145.320 726.720 155.840 727.040 ; 
                RECT 303.760 726.720 310.520 727.040 ; 
                RECT 0.160 728.080 155.840 728.400 ; 
                RECT 303.760 728.080 310.520 728.400 ; 
                RECT 0.160 729.440 135.440 729.760 ; 
                RECT 145.320 729.440 155.840 729.760 ; 
                RECT 303.760 729.440 310.520 729.760 ; 
                RECT 0.160 730.800 135.440 731.120 ; 
                RECT 145.320 730.800 155.840 731.120 ; 
                RECT 303.760 730.800 310.520 731.120 ; 
                RECT 0.160 732.160 140.200 732.480 ; 
                RECT 145.320 732.160 155.840 732.480 ; 
                RECT 303.760 732.160 310.520 732.480 ; 
                RECT 0.160 733.520 135.440 733.840 ; 
                RECT 145.320 733.520 155.840 733.840 ; 
                RECT 303.760 733.520 310.520 733.840 ; 
                RECT 0.160 734.880 135.440 735.200 ; 
                RECT 145.320 734.880 155.840 735.200 ; 
                RECT 303.760 734.880 310.520 735.200 ; 
                RECT 0.160 736.240 155.840 736.560 ; 
                RECT 303.760 736.240 310.520 736.560 ; 
                RECT 0.160 737.600 135.440 737.920 ; 
                RECT 145.320 737.600 155.840 737.920 ; 
                RECT 303.760 737.600 310.520 737.920 ; 
                RECT 0.160 738.960 135.440 739.280 ; 
                RECT 145.320 738.960 155.840 739.280 ; 
                RECT 303.760 738.960 310.520 739.280 ; 
                RECT 0.160 740.320 135.440 740.640 ; 
                RECT 145.320 740.320 155.840 740.640 ; 
                RECT 303.760 740.320 310.520 740.640 ; 
                RECT 0.160 741.680 142.920 742.000 ; 
                RECT 145.320 741.680 155.840 742.000 ; 
                RECT 303.760 741.680 310.520 742.000 ; 
                RECT 0.160 743.040 135.440 743.360 ; 
                RECT 145.320 743.040 155.840 743.360 ; 
                RECT 303.760 743.040 310.520 743.360 ; 
                RECT 0.160 744.400 155.840 744.720 ; 
                RECT 303.760 744.400 310.520 744.720 ; 
                RECT 0.160 745.760 196.640 746.080 ; 
                RECT 303.760 745.760 310.520 746.080 ; 
                RECT 0.160 747.120 196.640 747.440 ; 
                RECT 303.760 747.120 310.520 747.440 ; 
                RECT 0.160 748.480 196.640 748.800 ; 
                RECT 303.760 748.480 310.520 748.800 ; 
                RECT 0.160 749.840 310.520 750.160 ; 
                RECT 0.160 751.200 310.520 751.520 ; 
                RECT 0.160 752.560 310.520 752.880 ; 
                RECT 0.160 753.920 310.520 754.240 ; 
                RECT 0.160 0.160 310.520 1.520 ; 
                RECT 0.160 758.640 310.520 760.000 ; 
                RECT 200.780 45.420 206.580 46.790 ; 
                RECT 293.480 45.420 299.280 46.790 ; 
                RECT 200.780 50.465 206.580 51.855 ; 
                RECT 293.480 50.465 299.280 51.855 ; 
                RECT 200.780 55.615 206.580 57.055 ; 
                RECT 293.480 55.615 299.280 57.055 ; 
                RECT 200.780 60.845 206.580 62.285 ; 
                RECT 293.480 60.845 299.280 62.285 ; 
                RECT 200.780 106.210 299.280 109.810 ; 
                RECT 200.780 154.905 299.280 156.705 ; 
                RECT 200.780 116.015 299.280 116.305 ; 
                RECT 200.780 88.410 299.280 89.210 ; 
                RECT 200.780 216.045 299.280 219.645 ; 
                RECT 200.780 80.510 299.280 81.310 ; 
                RECT 200.780 83.520 299.280 84.320 ; 
                RECT 200.780 69.040 299.280 70.840 ; 
                RECT 200.780 29.665 299.280 31.465 ; 
                RECT 160.980 237.515 162.900 744.695 ; 
                RECT 164.820 237.515 166.740 744.695 ; 
                RECT 179.810 237.515 181.730 744.695 ; 
                RECT 183.650 237.515 185.570 744.695 ; 
                RECT 187.490 237.515 189.410 744.695 ; 
                RECT 191.330 237.515 193.250 744.695 ; 
                RECT 120.225 57.215 121.975 127.015 ; 
                RECT 126.685 57.215 128.605 127.015 ; 
                RECT 133.445 57.215 135.365 127.015 ; 
                RECT 141.940 57.215 143.860 127.015 ; 
                RECT 145.780 57.215 147.700 127.015 ; 
                RECT 157.330 57.215 159.250 127.015 ; 
                RECT 161.170 57.215 163.090 127.015 ; 
                RECT 165.010 57.215 166.930 127.015 ; 
                RECT 168.850 57.215 170.770 127.015 ; 
                RECT 134.310 189.120 136.230 230.880 ; 
                RECT 141.285 189.120 143.205 230.880 ; 
                RECT 147.915 189.120 149.665 230.880 ; 
                RECT 154.375 189.120 156.295 230.880 ; 
                RECT 164.160 189.120 166.080 230.880 ; 
                RECT 168.000 189.120 169.920 230.880 ; 
                RECT 168.875 177.960 170.795 183.120 ; 
                RECT 169.175 46.055 170.925 51.215 ; 
                RECT 77.080 239.785 86.240 240.535 ; 
                RECT 77.080 245.185 86.240 247.105 ; 
                RECT 57.740 225.795 73.780 227.445 ; 
                RECT 36.140 225.925 55.780 229.525 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 212.280 5.560 ; 
                RECT 214.000 5.240 223.160 5.560 ; 
                RECT 224.880 5.240 234.040 5.560 ; 
                RECT 235.760 5.240 244.920 5.560 ; 
                RECT 246.640 5.240 255.800 5.560 ; 
                RECT 257.520 5.240 266.680 5.560 ; 
                RECT 268.400 5.240 277.560 5.560 ; 
                RECT 279.280 5.240 288.440 5.560 ; 
                RECT 290.160 5.240 307.800 5.560 ; 
                RECT 2.880 6.600 307.800 6.920 ; 
                RECT 2.880 7.960 307.800 8.280 ; 
                RECT 2.880 9.320 172.840 9.640 ; 
                RECT 205.160 9.320 307.800 9.640 ; 
                RECT 2.880 10.680 307.800 11.000 ; 
                RECT 2.880 12.040 307.800 12.360 ; 
                RECT 2.880 13.400 91.920 13.720 ; 
                RECT 173.880 13.400 307.800 13.720 ; 
                RECT 2.880 14.760 307.800 15.080 ; 
                RECT 2.880 16.120 307.800 16.440 ; 
                RECT 2.880 17.480 91.920 17.800 ; 
                RECT 173.200 17.480 307.800 17.800 ; 
                RECT 2.880 18.840 307.800 19.160 ; 
                RECT 2.880 20.200 307.800 20.520 ; 
                RECT 2.880 21.560 307.800 21.880 ; 
                RECT 2.880 22.920 211.600 23.240 ; 
                RECT 289.480 22.920 307.800 23.240 ; 
                RECT 2.880 24.280 199.360 24.600 ; 
                RECT 301.040 24.280 307.800 24.600 ; 
                RECT 2.880 25.640 199.360 25.960 ; 
                RECT 301.040 25.640 307.800 25.960 ; 
                RECT 2.880 27.000 199.360 27.320 ; 
                RECT 301.040 27.000 307.800 27.320 ; 
                RECT 2.880 28.360 199.360 28.680 ; 
                RECT 301.040 28.360 307.800 28.680 ; 
                RECT 2.880 29.720 199.360 30.040 ; 
                RECT 301.040 29.720 307.800 30.040 ; 
                RECT 2.880 31.080 199.360 31.400 ; 
                RECT 301.040 31.080 307.800 31.400 ; 
                RECT 2.880 32.440 199.360 32.760 ; 
                RECT 301.040 32.440 307.800 32.760 ; 
                RECT 2.880 33.800 199.360 34.120 ; 
                RECT 301.040 33.800 307.800 34.120 ; 
                RECT 2.880 35.160 199.360 35.480 ; 
                RECT 301.040 35.160 307.800 35.480 ; 
                RECT 2.880 36.520 105.520 36.840 ; 
                RECT 146.000 36.520 199.360 36.840 ; 
                RECT 301.040 36.520 307.800 36.840 ; 
                RECT 2.880 37.880 104.160 38.200 ; 
                RECT 152.120 37.880 199.360 38.200 ; 
                RECT 301.040 37.880 307.800 38.200 ; 
                RECT 2.880 39.240 102.800 39.560 ; 
                RECT 158.240 39.240 199.360 39.560 ; 
                RECT 301.040 39.240 307.800 39.560 ; 
                RECT 2.880 40.600 80.360 40.920 ; 
                RECT 173.200 40.600 199.360 40.920 ; 
                RECT 301.040 40.600 307.800 40.920 ; 
                RECT 2.880 41.960 81.040 42.280 ; 
                RECT 163.680 41.960 198.680 42.280 ; 
                RECT 301.040 41.960 307.800 42.280 ; 
                RECT 2.880 43.320 199.360 43.640 ; 
                RECT 301.040 43.320 307.800 43.640 ; 
                RECT 2.880 44.680 199.360 45.000 ; 
                RECT 301.040 44.680 307.800 45.000 ; 
                RECT 2.880 46.040 166.040 46.360 ; 
                RECT 171.840 46.040 199.360 46.360 ; 
                RECT 301.040 46.040 307.800 46.360 ; 
                RECT 2.880 47.400 166.040 47.720 ; 
                RECT 301.040 47.400 307.800 47.720 ; 
                RECT 2.880 48.760 166.040 49.080 ; 
                RECT 301.040 48.760 307.800 49.080 ; 
                RECT 2.880 50.120 166.040 50.440 ; 
                RECT 171.840 50.120 199.360 50.440 ; 
                RECT 301.040 50.120 307.800 50.440 ; 
                RECT 2.880 51.480 166.040 51.800 ; 
                RECT 171.840 51.480 199.360 51.800 ; 
                RECT 301.040 51.480 307.800 51.800 ; 
                RECT 2.880 52.840 199.360 53.160 ; 
                RECT 301.040 52.840 307.800 53.160 ; 
                RECT 2.880 54.200 199.360 54.520 ; 
                RECT 301.040 54.200 307.800 54.520 ; 
                RECT 2.880 55.560 199.360 55.880 ; 
                RECT 301.040 55.560 307.800 55.880 ; 
                RECT 2.880 56.920 117.080 57.240 ; 
                RECT 171.160 56.920 199.360 57.240 ; 
                RECT 301.040 56.920 307.800 57.240 ; 
                RECT 2.880 58.280 102.800 58.600 ; 
                RECT 109.960 58.280 117.080 58.600 ; 
                RECT 171.160 58.280 199.360 58.600 ; 
                RECT 301.040 58.280 307.800 58.600 ; 
                RECT 2.880 59.640 104.160 59.960 ; 
                RECT 109.280 59.640 117.080 59.960 ; 
                RECT 180.680 59.640 199.360 59.960 ; 
                RECT 301.040 59.640 307.800 59.960 ; 
                RECT 2.880 61.000 105.520 61.320 ; 
                RECT 107.920 61.000 117.080 61.320 ; 
                RECT 180.680 61.000 199.360 61.320 ; 
                RECT 301.040 61.000 307.800 61.320 ; 
                RECT 2.880 62.360 117.080 62.680 ; 
                RECT 180.680 62.360 199.360 62.680 ; 
                RECT 301.040 62.360 307.800 62.680 ; 
                RECT 2.880 63.720 117.080 64.040 ; 
                RECT 179.320 63.720 199.360 64.040 ; 
                RECT 301.040 63.720 307.800 64.040 ; 
                RECT 2.880 65.080 117.080 65.400 ; 
                RECT 180.680 65.080 199.360 65.400 ; 
                RECT 301.040 65.080 307.800 65.400 ; 
                RECT 2.880 66.440 117.080 66.760 ; 
                RECT 171.160 66.440 199.360 66.760 ; 
                RECT 301.040 66.440 307.800 66.760 ; 
                RECT 2.880 67.800 117.080 68.120 ; 
                RECT 183.400 67.800 199.360 68.120 ; 
                RECT 301.040 67.800 307.800 68.120 ; 
                RECT 2.880 69.160 117.080 69.480 ; 
                RECT 183.400 69.160 199.360 69.480 ; 
                RECT 301.040 69.160 307.800 69.480 ; 
                RECT 2.880 70.520 117.080 70.840 ; 
                RECT 182.040 70.520 199.360 70.840 ; 
                RECT 301.040 70.520 307.800 70.840 ; 
                RECT 2.880 71.880 117.080 72.200 ; 
                RECT 183.400 71.880 199.360 72.200 ; 
                RECT 301.040 71.880 307.800 72.200 ; 
                RECT 2.880 73.240 117.080 73.560 ; 
                RECT 183.400 73.240 199.360 73.560 ; 
                RECT 301.040 73.240 307.800 73.560 ; 
                RECT 2.880 74.600 117.080 74.920 ; 
                RECT 171.160 74.600 199.360 74.920 ; 
                RECT 301.040 74.600 307.800 74.920 ; 
                RECT 2.880 75.960 117.080 76.280 ; 
                RECT 186.120 75.960 199.360 76.280 ; 
                RECT 301.040 75.960 307.800 76.280 ; 
                RECT 2.880 77.320 117.080 77.640 ; 
                RECT 184.760 77.320 199.360 77.640 ; 
                RECT 301.040 77.320 307.800 77.640 ; 
                RECT 2.880 78.680 117.080 79.000 ; 
                RECT 186.120 78.680 199.360 79.000 ; 
                RECT 301.040 78.680 307.800 79.000 ; 
                RECT 2.880 80.040 117.080 80.360 ; 
                RECT 186.120 80.040 199.360 80.360 ; 
                RECT 301.040 80.040 307.800 80.360 ; 
                RECT 2.880 81.400 117.080 81.720 ; 
                RECT 186.120 81.400 199.360 81.720 ; 
                RECT 301.040 81.400 307.800 81.720 ; 
                RECT 2.880 82.760 117.080 83.080 ; 
                RECT 184.760 82.760 199.360 83.080 ; 
                RECT 301.040 82.760 307.800 83.080 ; 
                RECT 2.880 84.120 117.080 84.440 ; 
                RECT 171.160 84.120 199.360 84.440 ; 
                RECT 301.040 84.120 307.800 84.440 ; 
                RECT 2.880 85.480 117.080 85.800 ; 
                RECT 187.480 85.480 199.360 85.800 ; 
                RECT 301.040 85.480 307.800 85.800 ; 
                RECT 2.880 86.840 117.080 87.160 ; 
                RECT 188.840 86.840 199.360 87.160 ; 
                RECT 301.040 86.840 307.800 87.160 ; 
                RECT 2.880 88.200 117.080 88.520 ; 
                RECT 188.840 88.200 199.360 88.520 ; 
                RECT 301.040 88.200 307.800 88.520 ; 
                RECT 2.880 89.560 117.080 89.880 ; 
                RECT 187.480 89.560 199.360 89.880 ; 
                RECT 301.040 89.560 307.800 89.880 ; 
                RECT 2.880 90.920 117.080 91.240 ; 
                RECT 188.840 90.920 199.360 91.240 ; 
                RECT 301.040 90.920 307.800 91.240 ; 
                RECT 2.880 92.280 117.080 92.600 ; 
                RECT 171.160 92.280 199.360 92.600 ; 
                RECT 301.040 92.280 307.800 92.600 ; 
                RECT 2.880 93.640 117.080 93.960 ; 
                RECT 191.560 93.640 199.360 93.960 ; 
                RECT 301.040 93.640 307.800 93.960 ; 
                RECT 2.880 95.000 117.080 95.320 ; 
                RECT 191.560 95.000 199.360 95.320 ; 
                RECT 301.040 95.000 307.800 95.320 ; 
                RECT 2.880 96.360 117.080 96.680 ; 
                RECT 190.200 96.360 199.360 96.680 ; 
                RECT 301.040 96.360 307.800 96.680 ; 
                RECT 2.880 97.720 117.080 98.040 ; 
                RECT 191.560 97.720 199.360 98.040 ; 
                RECT 301.040 97.720 307.800 98.040 ; 
                RECT 2.880 99.080 117.080 99.400 ; 
                RECT 191.560 99.080 199.360 99.400 ; 
                RECT 301.040 99.080 307.800 99.400 ; 
                RECT 2.880 100.440 117.080 100.760 ; 
                RECT 171.160 100.440 199.360 100.760 ; 
                RECT 301.040 100.440 307.800 100.760 ; 
                RECT 2.880 101.800 117.080 102.120 ; 
                RECT 194.280 101.800 199.360 102.120 ; 
                RECT 301.040 101.800 307.800 102.120 ; 
                RECT 2.880 103.160 117.080 103.480 ; 
                RECT 192.920 103.160 199.360 103.480 ; 
                RECT 301.040 103.160 307.800 103.480 ; 
                RECT 2.880 104.520 117.080 104.840 ; 
                RECT 194.280 104.520 199.360 104.840 ; 
                RECT 301.040 104.520 307.800 104.840 ; 
                RECT 2.880 105.880 117.080 106.200 ; 
                RECT 194.280 105.880 199.360 106.200 ; 
                RECT 301.040 105.880 307.800 106.200 ; 
                RECT 2.880 107.240 117.080 107.560 ; 
                RECT 194.280 107.240 199.360 107.560 ; 
                RECT 301.040 107.240 307.800 107.560 ; 
                RECT 2.880 108.600 117.080 108.920 ; 
                RECT 192.920 108.600 199.360 108.920 ; 
                RECT 301.040 108.600 307.800 108.920 ; 
                RECT 2.880 109.960 117.080 110.280 ; 
                RECT 171.160 109.960 199.360 110.280 ; 
                RECT 301.040 109.960 307.800 110.280 ; 
                RECT 2.880 111.320 117.080 111.640 ; 
                RECT 195.640 111.320 199.360 111.640 ; 
                RECT 301.040 111.320 307.800 111.640 ; 
                RECT 2.880 112.680 117.080 113.000 ; 
                RECT 197.000 112.680 199.360 113.000 ; 
                RECT 301.040 112.680 307.800 113.000 ; 
                RECT 2.880 114.040 117.080 114.360 ; 
                RECT 197.000 114.040 199.360 114.360 ; 
                RECT 301.040 114.040 307.800 114.360 ; 
                RECT 2.880 115.400 117.080 115.720 ; 
                RECT 195.640 115.400 199.360 115.720 ; 
                RECT 301.040 115.400 307.800 115.720 ; 
                RECT 2.880 116.760 117.080 117.080 ; 
                RECT 197.000 116.760 199.360 117.080 ; 
                RECT 301.040 116.760 307.800 117.080 ; 
                RECT 2.880 118.120 117.080 118.440 ; 
                RECT 171.160 118.120 199.360 118.440 ; 
                RECT 301.040 118.120 307.800 118.440 ; 
                RECT 2.880 119.480 117.080 119.800 ; 
                RECT 301.040 119.480 307.800 119.800 ; 
                RECT 2.880 120.840 117.080 121.160 ; 
                RECT 301.040 120.840 307.800 121.160 ; 
                RECT 2.880 122.200 117.080 122.520 ; 
                RECT 301.040 122.200 307.800 122.520 ; 
                RECT 2.880 123.560 117.080 123.880 ; 
                RECT 301.040 123.560 307.800 123.880 ; 
                RECT 2.880 124.920 117.080 125.240 ; 
                RECT 301.040 124.920 307.800 125.240 ; 
                RECT 2.880 126.280 117.080 126.600 ; 
                RECT 171.160 126.280 199.360 126.600 ; 
                RECT 301.040 126.280 307.800 126.600 ; 
                RECT 2.880 127.640 199.360 127.960 ; 
                RECT 301.040 127.640 307.800 127.960 ; 
                RECT 2.880 129.000 199.360 129.320 ; 
                RECT 301.040 129.000 307.800 129.320 ; 
                RECT 2.880 130.360 174.880 130.680 ; 
                RECT 301.040 130.360 307.800 130.680 ; 
                RECT 2.880 131.720 196.640 132.040 ; 
                RECT 301.040 131.720 307.800 132.040 ; 
                RECT 2.880 133.080 193.920 133.400 ; 
                RECT 301.040 133.080 307.800 133.400 ; 
                RECT 2.880 134.440 191.200 134.760 ; 
                RECT 301.040 134.440 307.800 134.760 ; 
                RECT 2.880 135.800 188.480 136.120 ; 
                RECT 301.040 135.800 307.800 136.120 ; 
                RECT 2.880 137.160 78.320 137.480 ; 
                RECT 88.880 137.160 183.040 137.480 ; 
                RECT 301.040 137.160 307.800 137.480 ; 
                RECT 2.880 138.520 79.680 138.840 ; 
                RECT 85.480 138.520 93.280 138.840 ; 
                RECT 95.680 138.520 180.320 138.840 ; 
                RECT 301.040 138.520 307.800 138.840 ; 
                RECT 2.880 139.880 81.040 140.200 ; 
                RECT 84.800 139.880 177.600 140.200 ; 
                RECT 301.040 139.880 307.800 140.200 ; 
                RECT 2.880 141.240 56.560 141.560 ; 
                RECT 75.280 141.240 177.600 141.560 ; 
                RECT 301.040 141.240 307.800 141.560 ; 
                RECT 2.880 142.600 56.560 142.920 ; 
                RECT 75.280 142.600 87.160 142.920 ; 
                RECT 96.360 142.600 199.360 142.920 ; 
                RECT 301.040 142.600 307.800 142.920 ; 
                RECT 2.880 143.960 56.560 144.280 ; 
                RECT 75.280 143.960 80.360 144.280 ; 
                RECT 88.880 143.960 199.360 144.280 ; 
                RECT 301.040 143.960 307.800 144.280 ; 
                RECT 2.880 145.320 56.560 145.640 ; 
                RECT 75.280 145.320 83.760 145.640 ; 
                RECT 88.880 145.320 199.360 145.640 ; 
                RECT 301.040 145.320 307.800 145.640 ; 
                RECT 2.880 146.680 56.560 147.000 ; 
                RECT 75.280 146.680 199.360 147.000 ; 
                RECT 301.040 146.680 307.800 147.000 ; 
                RECT 2.880 148.040 56.560 148.360 ; 
                RECT 75.280 148.040 77.640 148.360 ; 
                RECT 88.880 148.040 199.360 148.360 ; 
                RECT 301.040 148.040 307.800 148.360 ; 
                RECT 2.880 149.400 56.560 149.720 ; 
                RECT 75.280 149.400 86.480 149.720 ; 
                RECT 95.000 149.400 199.360 149.720 ; 
                RECT 301.040 149.400 307.800 149.720 ; 
                RECT 2.880 150.760 56.560 151.080 ; 
                RECT 75.280 150.760 199.360 151.080 ; 
                RECT 301.040 150.760 307.800 151.080 ; 
                RECT 2.880 152.120 56.560 152.440 ; 
                RECT 75.280 152.120 87.160 152.440 ; 
                RECT 92.960 152.120 199.360 152.440 ; 
                RECT 301.040 152.120 307.800 152.440 ; 
                RECT 2.880 153.480 56.560 153.800 ; 
                RECT 75.280 153.480 89.880 153.800 ; 
                RECT 95.680 153.480 199.360 153.800 ; 
                RECT 301.040 153.480 307.800 153.800 ; 
                RECT 2.880 154.840 56.560 155.160 ; 
                RECT 75.280 154.840 84.440 155.160 ; 
                RECT 88.880 154.840 199.360 155.160 ; 
                RECT 301.040 154.840 307.800 155.160 ; 
                RECT 2.880 156.200 56.560 156.520 ; 
                RECT 75.280 156.200 199.360 156.520 ; 
                RECT 301.040 156.200 307.800 156.520 ; 
                RECT 2.880 157.560 56.560 157.880 ; 
                RECT 75.280 157.560 77.640 157.880 ; 
                RECT 100.440 157.560 199.360 157.880 ; 
                RECT 301.040 157.560 307.800 157.880 ; 
                RECT 2.880 158.920 56.560 159.240 ; 
                RECT 75.280 158.920 87.160 159.240 ; 
                RECT 95.680 158.920 199.360 159.240 ; 
                RECT 301.040 158.920 307.800 159.240 ; 
                RECT 2.880 160.280 56.560 160.600 ; 
                RECT 75.280 160.280 86.480 160.600 ; 
                RECT 88.880 160.280 94.640 160.600 ; 
                RECT 102.480 160.280 199.360 160.600 ; 
                RECT 301.040 160.280 307.800 160.600 ; 
                RECT 2.880 161.640 56.560 161.960 ; 
                RECT 75.280 161.640 78.320 161.960 ; 
                RECT 91.600 161.640 199.360 161.960 ; 
                RECT 301.040 161.640 307.800 161.960 ; 
                RECT 2.880 163.000 56.560 163.320 ; 
                RECT 75.280 163.000 87.160 163.320 ; 
                RECT 95.680 163.000 199.360 163.320 ; 
                RECT 301.040 163.000 307.800 163.320 ; 
                RECT 2.880 164.360 56.560 164.680 ; 
                RECT 75.280 164.360 84.440 164.680 ; 
                RECT 88.880 164.360 199.360 164.680 ; 
                RECT 301.040 164.360 307.800 164.680 ; 
                RECT 2.880 165.720 56.560 166.040 ; 
                RECT 75.280 165.720 87.160 166.040 ; 
                RECT 96.360 165.720 199.360 166.040 ; 
                RECT 301.040 165.720 307.800 166.040 ; 
                RECT 2.880 167.080 56.560 167.400 ; 
                RECT 75.280 167.080 199.360 167.400 ; 
                RECT 301.040 167.080 307.800 167.400 ; 
                RECT 2.880 168.440 56.560 168.760 ; 
                RECT 75.280 168.440 80.360 168.760 ; 
                RECT 83.440 168.440 199.360 168.760 ; 
                RECT 301.040 168.440 307.800 168.760 ; 
                RECT 2.880 169.800 56.560 170.120 ; 
                RECT 75.280 169.800 80.360 170.120 ; 
                RECT 88.880 169.800 199.360 170.120 ; 
                RECT 301.040 169.800 307.800 170.120 ; 
                RECT 2.880 171.160 56.560 171.480 ; 
                RECT 75.280 171.160 199.360 171.480 ; 
                RECT 301.040 171.160 307.800 171.480 ; 
                RECT 2.880 172.520 56.560 172.840 ; 
                RECT 75.280 172.520 199.360 172.840 ; 
                RECT 301.040 172.520 307.800 172.840 ; 
                RECT 2.880 173.880 56.560 174.200 ; 
                RECT 75.280 173.880 86.480 174.200 ; 
                RECT 88.880 173.880 199.360 174.200 ; 
                RECT 301.040 173.880 307.800 174.200 ; 
                RECT 2.880 175.240 56.560 175.560 ; 
                RECT 75.280 175.240 79.680 175.560 ; 
                RECT 95.000 175.240 199.360 175.560 ; 
                RECT 301.040 175.240 307.800 175.560 ; 
                RECT 2.880 176.600 56.560 176.920 ; 
                RECT 75.280 176.600 86.480 176.920 ; 
                RECT 88.880 176.600 199.360 176.920 ; 
                RECT 301.040 176.600 307.800 176.920 ; 
                RECT 2.880 177.960 56.560 178.280 ; 
                RECT 75.280 177.960 101.440 178.280 ; 
                RECT 171.160 177.960 199.360 178.280 ; 
                RECT 301.040 177.960 307.800 178.280 ; 
                RECT 2.880 179.320 56.560 179.640 ; 
                RECT 75.280 179.320 81.720 179.640 ; 
                RECT 88.880 179.320 165.360 179.640 ; 
                RECT 171.160 179.320 199.360 179.640 ; 
                RECT 301.040 179.320 307.800 179.640 ; 
                RECT 2.880 180.680 56.560 181.000 ; 
                RECT 75.280 180.680 78.320 181.000 ; 
                RECT 89.560 180.680 165.360 181.000 ; 
                RECT 171.160 180.680 199.360 181.000 ; 
                RECT 301.040 180.680 307.800 181.000 ; 
                RECT 2.880 182.040 56.560 182.360 ; 
                RECT 75.280 182.040 83.760 182.360 ; 
                RECT 95.680 182.040 165.360 182.360 ; 
                RECT 171.160 182.040 199.360 182.360 ; 
                RECT 301.040 182.040 307.800 182.360 ; 
                RECT 2.880 183.400 56.560 183.720 ; 
                RECT 75.280 183.400 77.640 183.720 ; 
                RECT 85.480 183.400 165.360 183.720 ; 
                RECT 171.160 183.400 199.360 183.720 ; 
                RECT 301.040 183.400 307.800 183.720 ; 
                RECT 2.880 184.760 56.560 185.080 ; 
                RECT 91.600 184.760 199.360 185.080 ; 
                RECT 301.040 184.760 307.800 185.080 ; 
                RECT 2.880 186.120 56.560 186.440 ; 
                RECT 75.280 186.120 199.360 186.440 ; 
                RECT 301.040 186.120 307.800 186.440 ; 
                RECT 2.880 187.480 56.560 187.800 ; 
                RECT 75.280 187.480 199.360 187.800 ; 
                RECT 301.040 187.480 307.800 187.800 ; 
                RECT 2.880 188.840 56.560 189.160 ; 
                RECT 75.280 188.840 130.680 189.160 ; 
                RECT 170.480 188.840 199.360 189.160 ; 
                RECT 301.040 188.840 307.800 189.160 ; 
                RECT 2.880 190.200 56.560 190.520 ; 
                RECT 75.280 190.200 89.880 190.520 ; 
                RECT 96.360 190.200 130.680 190.520 ; 
                RECT 170.480 190.200 178.960 190.520 ; 
                RECT 301.040 190.200 307.800 190.520 ; 
                RECT 2.880 191.560 56.560 191.880 ; 
                RECT 75.280 191.560 130.680 191.880 ; 
                RECT 170.480 191.560 181.680 191.880 ; 
                RECT 301.040 191.560 307.800 191.880 ; 
                RECT 2.880 192.920 56.560 193.240 ; 
                RECT 75.280 192.920 130.680 193.240 ; 
                RECT 170.480 192.920 184.400 193.240 ; 
                RECT 301.040 192.920 307.800 193.240 ; 
                RECT 2.880 194.280 56.560 194.600 ; 
                RECT 75.280 194.280 77.640 194.600 ; 
                RECT 83.440 194.280 130.680 194.600 ; 
                RECT 170.480 194.280 187.120 194.600 ; 
                RECT 301.040 194.280 307.800 194.600 ; 
                RECT 2.880 195.640 56.560 195.960 ; 
                RECT 75.280 195.640 130.680 195.960 ; 
                RECT 170.480 195.640 189.840 195.960 ; 
                RECT 301.040 195.640 307.800 195.960 ; 
                RECT 2.880 197.000 56.560 197.320 ; 
                RECT 75.280 197.000 130.680 197.320 ; 
                RECT 170.480 197.000 192.560 197.320 ; 
                RECT 301.040 197.000 307.800 197.320 ; 
                RECT 2.880 198.360 56.560 198.680 ; 
                RECT 75.280 198.360 130.680 198.680 ; 
                RECT 170.480 198.360 195.280 198.680 ; 
                RECT 301.040 198.360 307.800 198.680 ; 
                RECT 2.880 199.720 56.560 200.040 ; 
                RECT 75.280 199.720 130.680 200.040 ; 
                RECT 301.040 199.720 307.800 200.040 ; 
                RECT 2.880 201.080 56.560 201.400 ; 
                RECT 75.280 201.080 83.080 201.400 ; 
                RECT 95.680 201.080 130.680 201.400 ; 
                RECT 301.040 201.080 307.800 201.400 ; 
                RECT 2.880 202.440 56.560 202.760 ; 
                RECT 75.280 202.440 130.680 202.760 ; 
                RECT 170.480 202.440 199.360 202.760 ; 
                RECT 301.040 202.440 307.800 202.760 ; 
                RECT 2.880 203.800 56.560 204.120 ; 
                RECT 75.280 203.800 80.360 204.120 ; 
                RECT 84.800 203.800 130.680 204.120 ; 
                RECT 170.480 203.800 199.360 204.120 ; 
                RECT 301.040 203.800 307.800 204.120 ; 
                RECT 2.880 205.160 56.560 205.480 ; 
                RECT 75.280 205.160 130.680 205.480 ; 
                RECT 170.480 205.160 199.360 205.480 ; 
                RECT 301.040 205.160 307.800 205.480 ; 
                RECT 2.880 206.520 56.560 206.840 ; 
                RECT 75.280 206.520 130.680 206.840 ; 
                RECT 170.480 206.520 199.360 206.840 ; 
                RECT 301.040 206.520 307.800 206.840 ; 
                RECT 2.880 207.880 56.560 208.200 ; 
                RECT 75.280 207.880 130.680 208.200 ; 
                RECT 170.480 207.880 199.360 208.200 ; 
                RECT 301.040 207.880 307.800 208.200 ; 
                RECT 2.880 209.240 56.560 209.560 ; 
                RECT 75.280 209.240 83.080 209.560 ; 
                RECT 85.480 209.240 130.680 209.560 ; 
                RECT 170.480 209.240 199.360 209.560 ; 
                RECT 301.040 209.240 307.800 209.560 ; 
                RECT 2.880 210.600 56.560 210.920 ; 
                RECT 75.280 210.600 79.680 210.920 ; 
                RECT 82.760 210.600 93.280 210.920 ; 
                RECT 96.360 210.600 130.680 210.920 ; 
                RECT 170.480 210.600 199.360 210.920 ; 
                RECT 301.040 210.600 307.800 210.920 ; 
                RECT 2.880 211.960 56.560 212.280 ; 
                RECT 75.280 211.960 130.680 212.280 ; 
                RECT 170.480 211.960 199.360 212.280 ; 
                RECT 301.040 211.960 307.800 212.280 ; 
                RECT 2.880 213.320 56.560 213.640 ; 
                RECT 75.280 213.320 130.680 213.640 ; 
                RECT 170.480 213.320 199.360 213.640 ; 
                RECT 301.040 213.320 307.800 213.640 ; 
                RECT 2.880 214.680 56.560 215.000 ; 
                RECT 75.280 214.680 130.680 215.000 ; 
                RECT 170.480 214.680 199.360 215.000 ; 
                RECT 301.040 214.680 307.800 215.000 ; 
                RECT 2.880 216.040 56.560 216.360 ; 
                RECT 75.280 216.040 130.680 216.360 ; 
                RECT 170.480 216.040 199.360 216.360 ; 
                RECT 301.040 216.040 307.800 216.360 ; 
                RECT 2.880 217.400 130.680 217.720 ; 
                RECT 170.480 217.400 199.360 217.720 ; 
                RECT 301.040 217.400 307.800 217.720 ; 
                RECT 2.880 218.760 86.480 219.080 ; 
                RECT 95.000 218.760 130.680 219.080 ; 
                RECT 170.480 218.760 199.360 219.080 ; 
                RECT 301.040 218.760 307.800 219.080 ; 
                RECT 2.880 220.120 35.480 220.440 ; 
                RECT 56.240 220.120 81.720 220.440 ; 
                RECT 85.480 220.120 130.680 220.440 ; 
                RECT 170.480 220.120 199.360 220.440 ; 
                RECT 301.040 220.120 307.800 220.440 ; 
                RECT 2.880 221.480 35.480 221.800 ; 
                RECT 56.240 221.480 130.680 221.800 ; 
                RECT 170.480 221.480 199.360 221.800 ; 
                RECT 301.040 221.480 307.800 221.800 ; 
                RECT 2.880 222.840 35.480 223.160 ; 
                RECT 56.240 222.840 130.680 223.160 ; 
                RECT 170.480 222.840 199.360 223.160 ; 
                RECT 301.040 222.840 307.800 223.160 ; 
                RECT 2.880 224.200 35.480 224.520 ; 
                RECT 56.240 224.200 62.680 224.520 ; 
                RECT 69.840 224.200 83.760 224.520 ; 
                RECT 89.560 224.200 130.680 224.520 ; 
                RECT 170.480 224.200 199.360 224.520 ; 
                RECT 301.040 224.200 307.800 224.520 ; 
                RECT 2.880 225.560 35.480 225.880 ; 
                RECT 56.240 225.560 57.240 225.880 ; 
                RECT 74.600 225.560 130.680 225.880 ; 
                RECT 170.480 225.560 199.360 225.880 ; 
                RECT 301.040 225.560 307.800 225.880 ; 
                RECT 2.880 226.920 35.480 227.240 ; 
                RECT 56.240 226.920 57.240 227.240 ; 
                RECT 74.600 226.920 130.680 227.240 ; 
                RECT 170.480 226.920 199.360 227.240 ; 
                RECT 301.040 226.920 307.800 227.240 ; 
                RECT 2.880 228.280 35.480 228.600 ; 
                RECT 56.240 228.280 130.680 228.600 ; 
                RECT 301.040 228.280 307.800 228.600 ; 
                RECT 2.880 229.640 35.480 229.960 ; 
                RECT 56.240 229.640 62.680 229.960 ; 
                RECT 69.840 229.640 78.320 229.960 ; 
                RECT 88.200 229.640 130.680 229.960 ; 
                RECT 301.040 229.640 307.800 229.960 ; 
                RECT 2.880 231.000 21.200 231.320 ; 
                RECT 69.160 231.000 130.680 231.320 ; 
                RECT 170.480 231.000 307.800 231.320 ; 
                RECT 2.880 232.360 68.800 232.680 ; 
                RECT 127.640 232.360 307.800 232.680 ; 
                RECT 2.880 233.720 196.640 234.040 ; 
                RECT 303.760 233.720 307.800 234.040 ; 
                RECT 2.880 235.080 196.640 235.400 ; 
                RECT 303.760 235.080 307.800 235.400 ; 
                RECT 2.880 236.440 196.640 236.760 ; 
                RECT 303.760 236.440 307.800 236.760 ; 
                RECT 2.880 237.800 78.320 238.120 ; 
                RECT 84.800 237.800 87.160 238.120 ; 
                RECT 101.120 237.800 155.840 238.120 ; 
                RECT 303.760 237.800 307.800 238.120 ; 
                RECT 2.880 239.160 76.280 239.480 ; 
                RECT 86.840 239.160 88.520 239.480 ; 
                RECT 100.440 239.160 112.320 239.480 ; 
                RECT 114.040 239.160 127.280 239.480 ; 
                RECT 145.320 239.160 155.840 239.480 ; 
                RECT 303.760 239.160 307.800 239.480 ; 
                RECT 2.880 240.520 76.280 240.840 ; 
                RECT 86.840 240.520 112.320 240.840 ; 
                RECT 116.760 240.520 127.280 240.840 ; 
                RECT 145.320 240.520 155.840 240.840 ; 
                RECT 303.760 240.520 307.800 240.840 ; 
                RECT 2.880 241.880 76.280 242.200 ; 
                RECT 86.840 241.880 112.320 242.200 ; 
                RECT 117.440 241.880 127.280 242.200 ; 
                RECT 145.320 241.880 155.840 242.200 ; 
                RECT 303.760 241.880 307.800 242.200 ; 
                RECT 2.880 243.240 76.280 243.560 ; 
                RECT 86.840 243.240 112.320 243.560 ; 
                RECT 117.440 243.240 127.280 243.560 ; 
                RECT 145.320 243.240 155.840 243.560 ; 
                RECT 303.760 243.240 307.800 243.560 ; 
                RECT 2.880 244.600 76.280 244.920 ; 
                RECT 86.840 244.600 112.320 244.920 ; 
                RECT 114.040 244.600 127.280 244.920 ; 
                RECT 145.320 244.600 155.840 244.920 ; 
                RECT 303.760 244.600 307.800 244.920 ; 
                RECT 2.880 245.960 76.280 246.280 ; 
                RECT 86.840 245.960 155.840 246.280 ; 
                RECT 303.760 245.960 307.800 246.280 ; 
                RECT 2.880 247.320 76.280 247.640 ; 
                RECT 86.840 247.320 127.280 247.640 ; 
                RECT 145.320 247.320 155.840 247.640 ; 
                RECT 303.760 247.320 307.800 247.640 ; 
                RECT 2.880 248.680 127.280 249.000 ; 
                RECT 145.320 248.680 155.840 249.000 ; 
                RECT 303.760 248.680 307.800 249.000 ; 
                RECT 2.880 250.040 127.280 250.360 ; 
                RECT 145.320 250.040 155.840 250.360 ; 
                RECT 303.760 250.040 307.800 250.360 ; 
                RECT 2.880 251.400 20.520 251.720 ; 
                RECT 71.880 251.400 127.280 251.720 ; 
                RECT 145.320 251.400 155.840 251.720 ; 
                RECT 303.760 251.400 307.800 251.720 ; 
                RECT 2.880 252.760 127.280 253.080 ; 
                RECT 145.320 252.760 155.840 253.080 ; 
                RECT 303.760 252.760 307.800 253.080 ; 
                RECT 2.880 254.120 19.840 254.440 ; 
                RECT 71.880 254.120 85.120 254.440 ; 
                RECT 101.120 254.120 155.840 254.440 ; 
                RECT 303.760 254.120 307.800 254.440 ; 
                RECT 2.880 255.480 19.160 255.800 ; 
                RECT 71.880 255.480 85.120 255.800 ; 
                RECT 99.760 255.480 112.320 255.800 ; 
                RECT 114.040 255.480 127.280 255.800 ; 
                RECT 145.320 255.480 155.840 255.800 ; 
                RECT 303.760 255.480 307.800 255.800 ; 
                RECT 2.880 256.840 18.480 257.160 ; 
                RECT 71.880 256.840 85.120 257.160 ; 
                RECT 90.240 256.840 112.320 257.160 ; 
                RECT 114.720 256.840 127.280 257.160 ; 
                RECT 145.320 256.840 155.840 257.160 ; 
                RECT 303.760 256.840 307.800 257.160 ; 
                RECT 2.880 258.200 112.320 258.520 ; 
                RECT 115.400 258.200 127.280 258.520 ; 
                RECT 145.320 258.200 155.840 258.520 ; 
                RECT 303.760 258.200 307.800 258.520 ; 
                RECT 2.880 259.560 17.800 259.880 ; 
                RECT 71.880 259.560 85.120 259.880 ; 
                RECT 90.920 259.560 112.320 259.880 ; 
                RECT 115.400 259.560 127.280 259.880 ; 
                RECT 145.320 259.560 155.840 259.880 ; 
                RECT 303.760 259.560 307.800 259.880 ; 
                RECT 2.880 260.920 17.120 261.240 ; 
                RECT 71.880 260.920 85.120 261.240 ; 
                RECT 91.600 260.920 112.320 261.240 ; 
                RECT 116.080 260.920 127.280 261.240 ; 
                RECT 145.320 260.920 155.840 261.240 ; 
                RECT 303.760 260.920 307.800 261.240 ; 
                RECT 2.880 262.280 16.440 262.600 ; 
                RECT 71.880 262.280 155.840 262.600 ; 
                RECT 303.760 262.280 307.800 262.600 ; 
                RECT 2.880 263.640 15.760 263.960 ; 
                RECT 71.880 263.640 127.280 263.960 ; 
                RECT 145.320 263.640 155.840 263.960 ; 
                RECT 303.760 263.640 307.800 263.960 ; 
                RECT 2.880 265.000 127.280 265.320 ; 
                RECT 145.320 265.000 155.840 265.320 ; 
                RECT 303.760 265.000 307.800 265.320 ; 
                RECT 2.880 266.360 15.080 266.680 ; 
                RECT 71.880 266.360 127.280 266.680 ; 
                RECT 145.320 266.360 155.840 266.680 ; 
                RECT 303.760 266.360 307.800 266.680 ; 
                RECT 2.880 267.720 14.400 268.040 ; 
                RECT 71.880 267.720 127.280 268.040 ; 
                RECT 145.320 267.720 155.840 268.040 ; 
                RECT 303.760 267.720 307.800 268.040 ; 
                RECT 2.880 269.080 127.280 269.400 ; 
                RECT 139.880 269.080 155.840 269.400 ; 
                RECT 303.760 269.080 307.800 269.400 ; 
                RECT 2.880 270.440 13.720 270.760 ; 
                RECT 71.880 270.440 85.120 270.760 ; 
                RECT 91.600 270.440 135.440 270.760 ; 
                RECT 145.320 270.440 155.840 270.760 ; 
                RECT 303.760 270.440 307.800 270.760 ; 
                RECT 2.880 271.800 13.040 272.120 ; 
                RECT 71.880 271.800 85.120 272.120 ; 
                RECT 90.920 271.800 127.280 272.120 ; 
                RECT 145.320 271.800 155.840 272.120 ; 
                RECT 303.760 271.800 307.800 272.120 ; 
                RECT 2.880 273.160 127.280 273.480 ; 
                RECT 145.320 273.160 155.840 273.480 ; 
                RECT 303.760 273.160 307.800 273.480 ; 
                RECT 2.880 274.520 12.360 274.840 ; 
                RECT 71.880 274.520 85.120 274.840 ; 
                RECT 90.240 274.520 127.280 274.840 ; 
                RECT 145.320 274.520 155.840 274.840 ; 
                RECT 303.760 274.520 307.800 274.840 ; 
                RECT 2.880 275.880 11.680 276.200 ; 
                RECT 71.880 275.880 85.120 276.200 ; 
                RECT 89.560 275.880 127.280 276.200 ; 
                RECT 145.320 275.880 155.840 276.200 ; 
                RECT 303.760 275.880 307.800 276.200 ; 
                RECT 2.880 277.240 11.000 277.560 ; 
                RECT 71.880 277.240 85.120 277.560 ; 
                RECT 88.880 277.240 127.280 277.560 ; 
                RECT 140.560 277.240 155.840 277.560 ; 
                RECT 303.760 277.240 307.800 277.560 ; 
                RECT 2.880 278.600 10.320 278.920 ; 
                RECT 71.880 278.600 127.280 278.920 ; 
                RECT 145.320 278.600 155.840 278.920 ; 
                RECT 303.760 278.600 307.800 278.920 ; 
                RECT 2.880 279.960 127.280 280.280 ; 
                RECT 145.320 279.960 155.840 280.280 ; 
                RECT 303.760 279.960 307.800 280.280 ; 
                RECT 2.880 281.320 127.280 281.640 ; 
                RECT 145.320 281.320 155.840 281.640 ; 
                RECT 303.760 281.320 307.800 281.640 ; 
                RECT 2.880 282.680 127.280 283.000 ; 
                RECT 145.320 282.680 155.840 283.000 ; 
                RECT 303.760 282.680 307.800 283.000 ; 
                RECT 2.880 284.040 127.280 284.360 ; 
                RECT 145.320 284.040 155.840 284.360 ; 
                RECT 303.760 284.040 307.800 284.360 ; 
                RECT 2.880 285.400 127.280 285.720 ; 
                RECT 140.560 285.400 155.840 285.720 ; 
                RECT 303.760 285.400 307.800 285.720 ; 
                RECT 2.880 286.760 127.280 287.080 ; 
                RECT 145.320 286.760 155.840 287.080 ; 
                RECT 303.760 286.760 307.800 287.080 ; 
                RECT 2.880 288.120 127.280 288.440 ; 
                RECT 145.320 288.120 155.840 288.440 ; 
                RECT 303.760 288.120 307.800 288.440 ; 
                RECT 2.880 289.480 127.280 289.800 ; 
                RECT 145.320 289.480 155.840 289.800 ; 
                RECT 303.760 289.480 307.800 289.800 ; 
                RECT 2.880 290.840 127.280 291.160 ; 
                RECT 145.320 290.840 155.840 291.160 ; 
                RECT 303.760 290.840 307.800 291.160 ; 
                RECT 2.880 292.200 127.280 292.520 ; 
                RECT 145.320 292.200 155.840 292.520 ; 
                RECT 303.760 292.200 307.800 292.520 ; 
                RECT 2.880 293.560 155.840 293.880 ; 
                RECT 303.760 293.560 307.800 293.880 ; 
                RECT 2.880 294.920 127.280 295.240 ; 
                RECT 145.320 294.920 155.840 295.240 ; 
                RECT 303.760 294.920 307.800 295.240 ; 
                RECT 2.880 296.280 127.280 296.600 ; 
                RECT 145.320 296.280 155.840 296.600 ; 
                RECT 303.760 296.280 307.800 296.600 ; 
                RECT 2.880 297.640 127.280 297.960 ; 
                RECT 145.320 297.640 155.840 297.960 ; 
                RECT 303.760 297.640 307.800 297.960 ; 
                RECT 2.880 299.000 127.280 299.320 ; 
                RECT 145.320 299.000 155.840 299.320 ; 
                RECT 303.760 299.000 307.800 299.320 ; 
                RECT 2.880 300.360 127.280 300.680 ; 
                RECT 145.320 300.360 155.840 300.680 ; 
                RECT 303.760 300.360 307.800 300.680 ; 
                RECT 2.880 301.720 155.840 302.040 ; 
                RECT 303.760 301.720 307.800 302.040 ; 
                RECT 2.880 303.080 127.280 303.400 ; 
                RECT 145.320 303.080 155.840 303.400 ; 
                RECT 303.760 303.080 307.800 303.400 ; 
                RECT 2.880 304.440 127.280 304.760 ; 
                RECT 145.320 304.440 155.840 304.760 ; 
                RECT 303.760 304.440 307.800 304.760 ; 
                RECT 2.880 305.800 127.280 306.120 ; 
                RECT 145.320 305.800 155.840 306.120 ; 
                RECT 303.760 305.800 307.800 306.120 ; 
                RECT 2.880 307.160 127.280 307.480 ; 
                RECT 145.320 307.160 155.840 307.480 ; 
                RECT 303.760 307.160 307.800 307.480 ; 
                RECT 2.880 308.520 127.280 308.840 ; 
                RECT 145.320 308.520 155.840 308.840 ; 
                RECT 303.760 308.520 307.800 308.840 ; 
                RECT 2.880 309.880 155.840 310.200 ; 
                RECT 303.760 309.880 307.800 310.200 ; 
                RECT 2.880 311.240 127.280 311.560 ; 
                RECT 145.320 311.240 155.840 311.560 ; 
                RECT 303.760 311.240 307.800 311.560 ; 
                RECT 2.880 312.600 127.280 312.920 ; 
                RECT 145.320 312.600 155.840 312.920 ; 
                RECT 303.760 312.600 307.800 312.920 ; 
                RECT 2.880 313.960 127.280 314.280 ; 
                RECT 145.320 313.960 155.840 314.280 ; 
                RECT 303.760 313.960 307.800 314.280 ; 
                RECT 2.880 315.320 127.280 315.640 ; 
                RECT 145.320 315.320 155.840 315.640 ; 
                RECT 303.760 315.320 307.800 315.640 ; 
                RECT 2.880 316.680 127.280 317.000 ; 
                RECT 143.960 316.680 155.840 317.000 ; 
                RECT 303.760 316.680 307.800 317.000 ; 
                RECT 2.880 318.040 139.520 318.360 ; 
                RECT 145.320 318.040 155.840 318.360 ; 
                RECT 303.760 318.040 307.800 318.360 ; 
                RECT 2.880 319.400 127.280 319.720 ; 
                RECT 145.320 319.400 155.840 319.720 ; 
                RECT 303.760 319.400 307.800 319.720 ; 
                RECT 2.880 320.760 127.280 321.080 ; 
                RECT 145.320 320.760 155.840 321.080 ; 
                RECT 303.760 320.760 307.800 321.080 ; 
                RECT 2.880 322.120 127.280 322.440 ; 
                RECT 145.320 322.120 155.840 322.440 ; 
                RECT 303.760 322.120 307.800 322.440 ; 
                RECT 2.880 323.480 127.280 323.800 ; 
                RECT 145.320 323.480 155.840 323.800 ; 
                RECT 303.760 323.480 307.800 323.800 ; 
                RECT 2.880 324.840 127.280 325.160 ; 
                RECT 143.960 324.840 155.840 325.160 ; 
                RECT 303.760 324.840 307.800 325.160 ; 
                RECT 2.880 326.200 127.280 326.520 ; 
                RECT 145.320 326.200 155.840 326.520 ; 
                RECT 303.760 326.200 307.800 326.520 ; 
                RECT 2.880 327.560 127.280 327.880 ; 
                RECT 145.320 327.560 155.840 327.880 ; 
                RECT 303.760 327.560 307.800 327.880 ; 
                RECT 2.880 328.920 127.280 329.240 ; 
                RECT 145.320 328.920 155.840 329.240 ; 
                RECT 303.760 328.920 307.800 329.240 ; 
                RECT 2.880 330.280 127.280 330.600 ; 
                RECT 145.320 330.280 155.840 330.600 ; 
                RECT 303.760 330.280 307.800 330.600 ; 
                RECT 2.880 331.640 127.280 331.960 ; 
                RECT 145.320 331.640 155.840 331.960 ; 
                RECT 303.760 331.640 307.800 331.960 ; 
                RECT 2.880 333.000 155.840 333.320 ; 
                RECT 303.760 333.000 307.800 333.320 ; 
                RECT 2.880 334.360 129.320 334.680 ; 
                RECT 145.320 334.360 155.840 334.680 ; 
                RECT 303.760 334.360 307.800 334.680 ; 
                RECT 2.880 335.720 129.320 336.040 ; 
                RECT 145.320 335.720 155.840 336.040 ; 
                RECT 303.760 335.720 307.800 336.040 ; 
                RECT 2.880 337.080 136.800 337.400 ; 
                RECT 145.320 337.080 155.840 337.400 ; 
                RECT 303.760 337.080 307.800 337.400 ; 
                RECT 2.880 338.440 129.320 338.760 ; 
                RECT 145.320 338.440 155.840 338.760 ; 
                RECT 303.760 338.440 307.800 338.760 ; 
                RECT 2.880 339.800 129.320 340.120 ; 
                RECT 145.320 339.800 155.840 340.120 ; 
                RECT 303.760 339.800 307.800 340.120 ; 
                RECT 2.880 341.160 91.240 341.480 ; 
                RECT 101.120 341.160 155.840 341.480 ; 
                RECT 303.760 341.160 307.800 341.480 ; 
                RECT 2.880 342.520 89.880 342.840 ; 
                RECT 99.760 342.520 112.320 342.840 ; 
                RECT 114.040 342.520 127.280 342.840 ; 
                RECT 145.320 342.520 155.840 342.840 ; 
                RECT 303.760 342.520 307.800 342.840 ; 
                RECT 2.880 343.880 112.320 344.200 ; 
                RECT 116.760 343.880 127.280 344.200 ; 
                RECT 145.320 343.880 155.840 344.200 ; 
                RECT 303.760 343.880 307.800 344.200 ; 
                RECT 2.880 345.240 112.320 345.560 ; 
                RECT 117.440 345.240 127.280 345.560 ; 
                RECT 145.320 345.240 155.840 345.560 ; 
                RECT 303.760 345.240 307.800 345.560 ; 
                RECT 2.880 346.600 112.320 346.920 ; 
                RECT 117.440 346.600 127.280 346.920 ; 
                RECT 145.320 346.600 155.840 346.920 ; 
                RECT 303.760 346.600 307.800 346.920 ; 
                RECT 2.880 347.960 112.320 348.280 ; 
                RECT 118.120 347.960 127.280 348.280 ; 
                RECT 145.320 347.960 155.840 348.280 ; 
                RECT 303.760 347.960 307.800 348.280 ; 
                RECT 2.880 349.320 155.840 349.640 ; 
                RECT 303.760 349.320 307.800 349.640 ; 
                RECT 2.880 350.680 127.280 351.000 ; 
                RECT 145.320 350.680 155.840 351.000 ; 
                RECT 303.760 350.680 307.800 351.000 ; 
                RECT 2.880 352.040 127.280 352.360 ; 
                RECT 145.320 352.040 155.840 352.360 ; 
                RECT 303.760 352.040 307.800 352.360 ; 
                RECT 2.880 353.400 127.280 353.720 ; 
                RECT 145.320 353.400 155.840 353.720 ; 
                RECT 303.760 353.400 307.800 353.720 ; 
                RECT 2.880 354.760 127.280 355.080 ; 
                RECT 145.320 354.760 155.840 355.080 ; 
                RECT 303.760 354.760 307.800 355.080 ; 
                RECT 2.880 356.120 89.200 356.440 ; 
                RECT 101.120 356.120 127.280 356.440 ; 
                RECT 130.360 356.120 155.840 356.440 ; 
                RECT 303.760 356.120 307.800 356.440 ; 
                RECT 2.880 357.480 87.840 357.800 ; 
                RECT 100.440 357.480 141.560 357.800 ; 
                RECT 145.320 357.480 155.840 357.800 ; 
                RECT 303.760 357.480 307.800 357.800 ; 
                RECT 2.880 358.840 112.320 359.160 ; 
                RECT 114.720 358.840 127.280 359.160 ; 
                RECT 145.320 358.840 155.840 359.160 ; 
                RECT 303.760 358.840 307.800 359.160 ; 
                RECT 2.880 360.200 112.320 360.520 ; 
                RECT 115.400 360.200 127.280 360.520 ; 
                RECT 145.320 360.200 155.840 360.520 ; 
                RECT 303.760 360.200 307.800 360.520 ; 
                RECT 2.880 361.560 112.320 361.880 ; 
                RECT 115.400 361.560 127.280 361.880 ; 
                RECT 145.320 361.560 155.840 361.880 ; 
                RECT 303.760 361.560 307.800 361.880 ; 
                RECT 2.880 362.920 112.320 363.240 ; 
                RECT 114.040 362.920 127.280 363.240 ; 
                RECT 145.320 362.920 155.840 363.240 ; 
                RECT 303.760 362.920 307.800 363.240 ; 
                RECT 2.880 364.280 112.320 364.600 ; 
                RECT 116.080 364.280 127.280 364.600 ; 
                RECT 131.040 364.280 155.840 364.600 ; 
                RECT 303.760 364.280 307.800 364.600 ; 
                RECT 2.880 365.640 127.280 365.960 ; 
                RECT 145.320 365.640 155.840 365.960 ; 
                RECT 303.760 365.640 307.800 365.960 ; 
                RECT 2.880 367.000 127.280 367.320 ; 
                RECT 145.320 367.000 155.840 367.320 ; 
                RECT 303.760 367.000 307.800 367.320 ; 
                RECT 2.880 368.360 127.280 368.680 ; 
                RECT 145.320 368.360 155.840 368.680 ; 
                RECT 303.760 368.360 307.800 368.680 ; 
                RECT 2.880 369.720 127.280 370.040 ; 
                RECT 145.320 369.720 155.840 370.040 ; 
                RECT 303.760 369.720 307.800 370.040 ; 
                RECT 2.880 371.080 127.280 371.400 ; 
                RECT 145.320 371.080 155.840 371.400 ; 
                RECT 303.760 371.080 307.800 371.400 ; 
                RECT 2.880 372.440 155.840 372.760 ; 
                RECT 303.760 372.440 307.800 372.760 ; 
                RECT 2.880 373.800 127.280 374.120 ; 
                RECT 145.320 373.800 155.840 374.120 ; 
                RECT 303.760 373.800 307.800 374.120 ; 
                RECT 2.880 375.160 127.280 375.480 ; 
                RECT 145.320 375.160 155.840 375.480 ; 
                RECT 303.760 375.160 307.800 375.480 ; 
                RECT 2.880 376.520 127.280 376.840 ; 
                RECT 145.320 376.520 155.840 376.840 ; 
                RECT 303.760 376.520 307.800 376.840 ; 
                RECT 2.880 377.880 127.280 378.200 ; 
                RECT 145.320 377.880 155.840 378.200 ; 
                RECT 303.760 377.880 307.800 378.200 ; 
                RECT 2.880 379.240 127.280 379.560 ; 
                RECT 145.320 379.240 155.840 379.560 ; 
                RECT 303.760 379.240 307.800 379.560 ; 
                RECT 2.880 380.600 155.840 380.920 ; 
                RECT 303.760 380.600 307.800 380.920 ; 
                RECT 2.880 381.960 127.280 382.280 ; 
                RECT 145.320 381.960 155.840 382.280 ; 
                RECT 303.760 381.960 307.800 382.280 ; 
                RECT 2.880 383.320 127.280 383.640 ; 
                RECT 145.320 383.320 155.840 383.640 ; 
                RECT 303.760 383.320 307.800 383.640 ; 
                RECT 2.880 384.680 127.280 385.000 ; 
                RECT 145.320 384.680 155.840 385.000 ; 
                RECT 303.760 384.680 307.800 385.000 ; 
                RECT 2.880 386.040 127.280 386.360 ; 
                RECT 145.320 386.040 155.840 386.360 ; 
                RECT 303.760 386.040 307.800 386.360 ; 
                RECT 2.880 387.400 127.280 387.720 ; 
                RECT 145.320 387.400 155.840 387.720 ; 
                RECT 303.760 387.400 307.800 387.720 ; 
                RECT 2.880 388.760 155.840 389.080 ; 
                RECT 303.760 388.760 307.800 389.080 ; 
                RECT 2.880 390.120 127.280 390.440 ; 
                RECT 145.320 390.120 155.840 390.440 ; 
                RECT 303.760 390.120 307.800 390.440 ; 
                RECT 2.880 391.480 127.280 391.800 ; 
                RECT 145.320 391.480 155.840 391.800 ; 
                RECT 303.760 391.480 307.800 391.800 ; 
                RECT 2.880 392.840 127.280 393.160 ; 
                RECT 145.320 392.840 155.840 393.160 ; 
                RECT 303.760 392.840 307.800 393.160 ; 
                RECT 2.880 394.200 127.280 394.520 ; 
                RECT 145.320 394.200 155.840 394.520 ; 
                RECT 303.760 394.200 307.800 394.520 ; 
                RECT 2.880 395.560 127.280 395.880 ; 
                RECT 133.760 395.560 155.840 395.880 ; 
                RECT 303.760 395.560 307.800 395.880 ; 
                RECT 2.880 396.920 135.440 397.240 ; 
                RECT 145.320 396.920 155.840 397.240 ; 
                RECT 303.760 396.920 307.800 397.240 ; 
                RECT 2.880 398.280 127.280 398.600 ; 
                RECT 145.320 398.280 155.840 398.600 ; 
                RECT 303.760 398.280 307.800 398.600 ; 
                RECT 2.880 399.640 127.280 399.960 ; 
                RECT 145.320 399.640 155.840 399.960 ; 
                RECT 303.760 399.640 307.800 399.960 ; 
                RECT 2.880 401.000 127.280 401.320 ; 
                RECT 145.320 401.000 155.840 401.320 ; 
                RECT 303.760 401.000 307.800 401.320 ; 
                RECT 2.880 402.360 127.280 402.680 ; 
                RECT 145.320 402.360 155.840 402.680 ; 
                RECT 303.760 402.360 307.800 402.680 ; 
                RECT 2.880 403.720 127.280 404.040 ; 
                RECT 134.440 403.720 155.840 404.040 ; 
                RECT 303.760 403.720 307.800 404.040 ; 
                RECT 2.880 405.080 127.280 405.400 ; 
                RECT 145.320 405.080 155.840 405.400 ; 
                RECT 303.760 405.080 307.800 405.400 ; 
                RECT 2.880 406.440 127.280 406.760 ; 
                RECT 145.320 406.440 155.840 406.760 ; 
                RECT 303.760 406.440 307.800 406.760 ; 
                RECT 2.880 407.800 127.280 408.120 ; 
                RECT 145.320 407.800 155.840 408.120 ; 
                RECT 303.760 407.800 307.800 408.120 ; 
                RECT 2.880 409.160 127.280 409.480 ; 
                RECT 145.320 409.160 155.840 409.480 ; 
                RECT 303.760 409.160 307.800 409.480 ; 
                RECT 2.880 410.520 127.280 410.840 ; 
                RECT 145.320 410.520 155.840 410.840 ; 
                RECT 303.760 410.520 307.800 410.840 ; 
                RECT 2.880 411.880 155.840 412.200 ; 
                RECT 303.760 411.880 307.800 412.200 ; 
                RECT 2.880 413.240 127.280 413.560 ; 
                RECT 145.320 413.240 155.840 413.560 ; 
                RECT 303.760 413.240 307.800 413.560 ; 
                RECT 2.880 414.600 127.280 414.920 ; 
                RECT 145.320 414.600 155.840 414.920 ; 
                RECT 303.760 414.600 307.800 414.920 ; 
                RECT 2.880 415.960 127.280 416.280 ; 
                RECT 145.320 415.960 155.840 416.280 ; 
                RECT 303.760 415.960 307.800 416.280 ; 
                RECT 2.880 417.320 127.280 417.640 ; 
                RECT 145.320 417.320 155.840 417.640 ; 
                RECT 303.760 417.320 307.800 417.640 ; 
                RECT 2.880 418.680 127.280 419.000 ; 
                RECT 145.320 418.680 155.840 419.000 ; 
                RECT 303.760 418.680 307.800 419.000 ; 
                RECT 2.880 420.040 155.840 420.360 ; 
                RECT 303.760 420.040 307.800 420.360 ; 
                RECT 2.880 421.400 127.280 421.720 ; 
                RECT 145.320 421.400 155.840 421.720 ; 
                RECT 303.760 421.400 307.800 421.720 ; 
                RECT 2.880 422.760 127.280 423.080 ; 
                RECT 145.320 422.760 155.840 423.080 ; 
                RECT 303.760 422.760 307.800 423.080 ; 
                RECT 2.880 424.120 127.280 424.440 ; 
                RECT 145.320 424.120 155.840 424.440 ; 
                RECT 303.760 424.120 307.800 424.440 ; 
                RECT 2.880 425.480 127.280 425.800 ; 
                RECT 145.320 425.480 155.840 425.800 ; 
                RECT 303.760 425.480 307.800 425.800 ; 
                RECT 2.880 426.840 127.280 427.160 ; 
                RECT 145.320 426.840 155.840 427.160 ; 
                RECT 303.760 426.840 307.800 427.160 ; 
                RECT 2.880 428.200 155.840 428.520 ; 
                RECT 303.760 428.200 307.800 428.520 ; 
                RECT 2.880 429.560 127.280 429.880 ; 
                RECT 145.320 429.560 155.840 429.880 ; 
                RECT 303.760 429.560 307.800 429.880 ; 
                RECT 2.880 430.920 127.280 431.240 ; 
                RECT 145.320 430.920 155.840 431.240 ; 
                RECT 303.760 430.920 307.800 431.240 ; 
                RECT 2.880 432.280 127.280 432.600 ; 
                RECT 145.320 432.280 155.840 432.600 ; 
                RECT 303.760 432.280 307.800 432.600 ; 
                RECT 2.880 433.640 127.280 433.960 ; 
                RECT 145.320 433.640 155.840 433.960 ; 
                RECT 303.760 433.640 307.800 433.960 ; 
                RECT 2.880 435.000 127.280 435.320 ; 
                RECT 137.160 435.000 155.840 435.320 ; 
                RECT 303.760 435.000 307.800 435.320 ; 
                RECT 2.880 436.360 137.480 436.680 ; 
                RECT 145.320 436.360 155.840 436.680 ; 
                RECT 303.760 436.360 307.800 436.680 ; 
                RECT 2.880 437.720 130.680 438.040 ; 
                RECT 145.320 437.720 155.840 438.040 ; 
                RECT 303.760 437.720 307.800 438.040 ; 
                RECT 2.880 439.080 130.680 439.400 ; 
                RECT 145.320 439.080 155.840 439.400 ; 
                RECT 303.760 439.080 307.800 439.400 ; 
                RECT 2.880 440.440 130.680 440.760 ; 
                RECT 145.320 440.440 155.840 440.760 ; 
                RECT 303.760 440.440 307.800 440.760 ; 
                RECT 2.880 441.800 130.680 442.120 ; 
                RECT 145.320 441.800 155.840 442.120 ; 
                RECT 303.760 441.800 307.800 442.120 ; 
                RECT 2.880 443.160 155.840 443.480 ; 
                RECT 303.760 443.160 307.800 443.480 ; 
                RECT 2.880 444.520 139.520 444.840 ; 
                RECT 145.320 444.520 155.840 444.840 ; 
                RECT 303.760 444.520 307.800 444.840 ; 
                RECT 2.880 445.880 130.680 446.200 ; 
                RECT 145.320 445.880 155.840 446.200 ; 
                RECT 303.760 445.880 307.800 446.200 ; 
                RECT 2.880 447.240 130.680 447.560 ; 
                RECT 145.320 447.240 155.840 447.560 ; 
                RECT 303.760 447.240 307.800 447.560 ; 
                RECT 2.880 448.600 130.680 448.920 ; 
                RECT 145.320 448.600 155.840 448.920 ; 
                RECT 303.760 448.600 307.800 448.920 ; 
                RECT 2.880 449.960 130.680 450.280 ; 
                RECT 145.320 449.960 155.840 450.280 ; 
                RECT 303.760 449.960 307.800 450.280 ; 
                RECT 2.880 451.320 155.840 451.640 ; 
                RECT 303.760 451.320 307.800 451.640 ; 
                RECT 2.880 452.680 130.680 453.000 ; 
                RECT 145.320 452.680 155.840 453.000 ; 
                RECT 303.760 452.680 307.800 453.000 ; 
                RECT 2.880 454.040 142.240 454.360 ; 
                RECT 145.320 454.040 155.840 454.360 ; 
                RECT 303.760 454.040 307.800 454.360 ; 
                RECT 2.880 455.400 130.680 455.720 ; 
                RECT 145.320 455.400 155.840 455.720 ; 
                RECT 303.760 455.400 307.800 455.720 ; 
                RECT 2.880 456.760 130.680 457.080 ; 
                RECT 145.320 456.760 155.840 457.080 ; 
                RECT 303.760 456.760 307.800 457.080 ; 
                RECT 2.880 458.120 130.680 458.440 ; 
                RECT 145.320 458.120 155.840 458.440 ; 
                RECT 303.760 458.120 307.800 458.440 ; 
                RECT 2.880 459.480 155.840 459.800 ; 
                RECT 303.760 459.480 307.800 459.800 ; 
                RECT 2.880 460.840 131.360 461.160 ; 
                RECT 145.320 460.840 155.840 461.160 ; 
                RECT 303.760 460.840 307.800 461.160 ; 
                RECT 2.880 462.200 131.360 462.520 ; 
                RECT 145.320 462.200 155.840 462.520 ; 
                RECT 303.760 462.200 307.800 462.520 ; 
                RECT 2.880 463.560 136.800 463.880 ; 
                RECT 145.320 463.560 155.840 463.880 ; 
                RECT 303.760 463.560 307.800 463.880 ; 
                RECT 2.880 464.920 131.360 465.240 ; 
                RECT 145.320 464.920 155.840 465.240 ; 
                RECT 303.760 464.920 307.800 465.240 ; 
                RECT 2.880 466.280 131.360 466.600 ; 
                RECT 145.320 466.280 155.840 466.600 ; 
                RECT 303.760 466.280 307.800 466.600 ; 
                RECT 2.880 467.640 155.840 467.960 ; 
                RECT 303.760 467.640 307.800 467.960 ; 
                RECT 2.880 469.000 131.360 469.320 ; 
                RECT 145.320 469.000 155.840 469.320 ; 
                RECT 303.760 469.000 307.800 469.320 ; 
                RECT 2.880 470.360 131.360 470.680 ; 
                RECT 145.320 470.360 155.840 470.680 ; 
                RECT 303.760 470.360 307.800 470.680 ; 
                RECT 2.880 471.720 131.360 472.040 ; 
                RECT 145.320 471.720 155.840 472.040 ; 
                RECT 303.760 471.720 307.800 472.040 ; 
                RECT 2.880 473.080 138.840 473.400 ; 
                RECT 145.320 473.080 155.840 473.400 ; 
                RECT 303.760 473.080 307.800 473.400 ; 
                RECT 2.880 474.440 131.360 474.760 ; 
                RECT 145.320 474.440 155.840 474.760 ; 
                RECT 303.760 474.440 307.800 474.760 ; 
                RECT 2.880 475.800 155.840 476.120 ; 
                RECT 303.760 475.800 307.800 476.120 ; 
                RECT 2.880 477.160 131.360 477.480 ; 
                RECT 145.320 477.160 155.840 477.480 ; 
                RECT 303.760 477.160 307.800 477.480 ; 
                RECT 2.880 478.520 131.360 478.840 ; 
                RECT 145.320 478.520 155.840 478.840 ; 
                RECT 303.760 478.520 307.800 478.840 ; 
                RECT 2.880 479.880 131.360 480.200 ; 
                RECT 145.320 479.880 155.840 480.200 ; 
                RECT 303.760 479.880 307.800 480.200 ; 
                RECT 2.880 481.240 131.360 481.560 ; 
                RECT 145.320 481.240 155.840 481.560 ; 
                RECT 303.760 481.240 307.800 481.560 ; 
                RECT 2.880 482.600 155.840 482.920 ; 
                RECT 303.760 482.600 307.800 482.920 ; 
                RECT 2.880 483.960 141.560 484.280 ; 
                RECT 145.320 483.960 155.840 484.280 ; 
                RECT 303.760 483.960 307.800 484.280 ; 
                RECT 2.880 485.320 131.360 485.640 ; 
                RECT 145.320 485.320 155.840 485.640 ; 
                RECT 303.760 485.320 307.800 485.640 ; 
                RECT 2.880 486.680 131.360 487.000 ; 
                RECT 145.320 486.680 155.840 487.000 ; 
                RECT 303.760 486.680 307.800 487.000 ; 
                RECT 2.880 488.040 131.360 488.360 ; 
                RECT 145.320 488.040 155.840 488.360 ; 
                RECT 303.760 488.040 307.800 488.360 ; 
                RECT 2.880 489.400 131.360 489.720 ; 
                RECT 145.320 489.400 155.840 489.720 ; 
                RECT 303.760 489.400 307.800 489.720 ; 
                RECT 2.880 490.760 155.840 491.080 ; 
                RECT 303.760 490.760 307.800 491.080 ; 
                RECT 2.880 492.120 132.040 492.440 ; 
                RECT 145.320 492.120 155.840 492.440 ; 
                RECT 303.760 492.120 307.800 492.440 ; 
                RECT 2.880 493.480 136.120 493.800 ; 
                RECT 145.320 493.480 155.840 493.800 ; 
                RECT 303.760 493.480 307.800 493.800 ; 
                RECT 2.880 494.840 132.040 495.160 ; 
                RECT 145.320 494.840 155.840 495.160 ; 
                RECT 303.760 494.840 307.800 495.160 ; 
                RECT 2.880 496.200 132.040 496.520 ; 
                RECT 145.320 496.200 155.840 496.520 ; 
                RECT 303.760 496.200 307.800 496.520 ; 
                RECT 2.880 497.560 132.040 497.880 ; 
                RECT 145.320 497.560 155.840 497.880 ; 
                RECT 303.760 497.560 307.800 497.880 ; 
                RECT 2.880 498.920 155.840 499.240 ; 
                RECT 303.760 498.920 307.800 499.240 ; 
                RECT 2.880 500.280 132.040 500.600 ; 
                RECT 145.320 500.280 155.840 500.600 ; 
                RECT 303.760 500.280 307.800 500.600 ; 
                RECT 2.880 501.640 132.040 501.960 ; 
                RECT 145.320 501.640 155.840 501.960 ; 
                RECT 303.760 501.640 307.800 501.960 ; 
                RECT 2.880 503.000 138.840 503.320 ; 
                RECT 145.320 503.000 155.840 503.320 ; 
                RECT 303.760 503.000 307.800 503.320 ; 
                RECT 2.880 504.360 132.040 504.680 ; 
                RECT 145.320 504.360 155.840 504.680 ; 
                RECT 303.760 504.360 307.800 504.680 ; 
                RECT 2.880 505.720 132.040 506.040 ; 
                RECT 145.320 505.720 155.840 506.040 ; 
                RECT 303.760 505.720 307.800 506.040 ; 
                RECT 2.880 507.080 155.840 507.400 ; 
                RECT 303.760 507.080 307.800 507.400 ; 
                RECT 2.880 508.440 132.040 508.760 ; 
                RECT 145.320 508.440 155.840 508.760 ; 
                RECT 303.760 508.440 307.800 508.760 ; 
                RECT 2.880 509.800 132.040 510.120 ; 
                RECT 145.320 509.800 155.840 510.120 ; 
                RECT 303.760 509.800 307.800 510.120 ; 
                RECT 2.880 511.160 132.040 511.480 ; 
                RECT 145.320 511.160 155.840 511.480 ; 
                RECT 303.760 511.160 307.800 511.480 ; 
                RECT 2.880 512.520 140.880 512.840 ; 
                RECT 145.320 512.520 155.840 512.840 ; 
                RECT 303.760 512.520 307.800 512.840 ; 
                RECT 2.880 513.880 132.040 514.200 ; 
                RECT 145.320 513.880 155.840 514.200 ; 
                RECT 303.760 513.880 307.800 514.200 ; 
                RECT 2.880 515.240 155.840 515.560 ; 
                RECT 303.760 515.240 307.800 515.560 ; 
                RECT 2.880 516.600 132.040 516.920 ; 
                RECT 145.320 516.600 155.840 516.920 ; 
                RECT 303.760 516.600 307.800 516.920 ; 
                RECT 2.880 517.960 132.040 518.280 ; 
                RECT 145.320 517.960 155.840 518.280 ; 
                RECT 303.760 517.960 307.800 518.280 ; 
                RECT 2.880 519.320 132.040 519.640 ; 
                RECT 145.320 519.320 155.840 519.640 ; 
                RECT 303.760 519.320 307.800 519.640 ; 
                RECT 2.880 520.680 132.040 521.000 ; 
                RECT 145.320 520.680 155.840 521.000 ; 
                RECT 303.760 520.680 307.800 521.000 ; 
                RECT 2.880 522.040 155.840 522.360 ; 
                RECT 303.760 522.040 307.800 522.360 ; 
                RECT 2.880 523.400 135.440 523.720 ; 
                RECT 145.320 523.400 155.840 523.720 ; 
                RECT 303.760 523.400 307.800 523.720 ; 
                RECT 2.880 524.760 132.040 525.080 ; 
                RECT 145.320 524.760 155.840 525.080 ; 
                RECT 303.760 524.760 307.800 525.080 ; 
                RECT 2.880 526.120 132.040 526.440 ; 
                RECT 145.320 526.120 155.840 526.440 ; 
                RECT 303.760 526.120 307.800 526.440 ; 
                RECT 2.880 527.480 132.040 527.800 ; 
                RECT 145.320 527.480 155.840 527.800 ; 
                RECT 303.760 527.480 307.800 527.800 ; 
                RECT 2.880 528.840 132.040 529.160 ; 
                RECT 145.320 528.840 155.840 529.160 ; 
                RECT 303.760 528.840 307.800 529.160 ; 
                RECT 2.880 530.200 155.840 530.520 ; 
                RECT 303.760 530.200 307.800 530.520 ; 
                RECT 2.880 531.560 137.480 531.880 ; 
                RECT 145.320 531.560 155.840 531.880 ; 
                RECT 303.760 531.560 307.800 531.880 ; 
                RECT 2.880 532.920 138.160 533.240 ; 
                RECT 145.320 532.920 155.840 533.240 ; 
                RECT 303.760 532.920 307.800 533.240 ; 
                RECT 2.880 534.280 132.040 534.600 ; 
                RECT 145.320 534.280 155.840 534.600 ; 
                RECT 303.760 534.280 307.800 534.600 ; 
                RECT 2.880 535.640 132.040 535.960 ; 
                RECT 145.320 535.640 155.840 535.960 ; 
                RECT 303.760 535.640 307.800 535.960 ; 
                RECT 2.880 537.000 132.040 537.320 ; 
                RECT 145.320 537.000 155.840 537.320 ; 
                RECT 303.760 537.000 307.800 537.320 ; 
                RECT 2.880 538.360 155.840 538.680 ; 
                RECT 303.760 538.360 307.800 538.680 ; 
                RECT 2.880 539.720 132.040 540.040 ; 
                RECT 145.320 539.720 155.840 540.040 ; 
                RECT 303.760 539.720 307.800 540.040 ; 
                RECT 2.880 541.080 140.200 541.400 ; 
                RECT 145.320 541.080 155.840 541.400 ; 
                RECT 303.760 541.080 307.800 541.400 ; 
                RECT 2.880 542.440 140.200 542.760 ; 
                RECT 145.320 542.440 155.840 542.760 ; 
                RECT 303.760 542.440 307.800 542.760 ; 
                RECT 2.880 543.800 132.040 544.120 ; 
                RECT 145.320 543.800 155.840 544.120 ; 
                RECT 303.760 543.800 307.800 544.120 ; 
                RECT 2.880 545.160 132.040 545.480 ; 
                RECT 145.320 545.160 155.840 545.480 ; 
                RECT 303.760 545.160 307.800 545.480 ; 
                RECT 2.880 546.520 155.840 546.840 ; 
                RECT 303.760 546.520 307.800 546.840 ; 
                RECT 2.880 547.880 132.040 548.200 ; 
                RECT 145.320 547.880 155.840 548.200 ; 
                RECT 303.760 547.880 307.800 548.200 ; 
                RECT 2.880 549.240 132.040 549.560 ; 
                RECT 145.320 549.240 155.840 549.560 ; 
                RECT 303.760 549.240 307.800 549.560 ; 
                RECT 2.880 550.600 132.040 550.920 ; 
                RECT 145.320 550.600 155.840 550.920 ; 
                RECT 303.760 550.600 307.800 550.920 ; 
                RECT 2.880 551.960 142.920 552.280 ; 
                RECT 145.320 551.960 155.840 552.280 ; 
                RECT 303.760 551.960 307.800 552.280 ; 
                RECT 2.880 553.320 132.040 553.640 ; 
                RECT 145.320 553.320 155.840 553.640 ; 
                RECT 303.760 553.320 307.800 553.640 ; 
                RECT 2.880 554.680 155.840 555.000 ; 
                RECT 303.760 554.680 307.800 555.000 ; 
                RECT 2.880 556.040 132.720 556.360 ; 
                RECT 145.320 556.040 155.840 556.360 ; 
                RECT 303.760 556.040 307.800 556.360 ; 
                RECT 2.880 557.400 132.720 557.720 ; 
                RECT 145.320 557.400 155.840 557.720 ; 
                RECT 303.760 557.400 307.800 557.720 ; 
                RECT 2.880 558.760 132.720 559.080 ; 
                RECT 145.320 558.760 155.840 559.080 ; 
                RECT 303.760 558.760 307.800 559.080 ; 
                RECT 2.880 560.120 132.720 560.440 ; 
                RECT 145.320 560.120 155.840 560.440 ; 
                RECT 303.760 560.120 307.800 560.440 ; 
                RECT 2.880 561.480 155.840 561.800 ; 
                RECT 303.760 561.480 307.800 561.800 ; 
                RECT 2.880 562.840 137.480 563.160 ; 
                RECT 145.320 562.840 155.840 563.160 ; 
                RECT 303.760 562.840 307.800 563.160 ; 
                RECT 2.880 564.200 132.720 564.520 ; 
                RECT 145.320 564.200 155.840 564.520 ; 
                RECT 303.760 564.200 307.800 564.520 ; 
                RECT 2.880 565.560 132.720 565.880 ; 
                RECT 145.320 565.560 155.840 565.880 ; 
                RECT 303.760 565.560 307.800 565.880 ; 
                RECT 2.880 566.920 132.720 567.240 ; 
                RECT 145.320 566.920 155.840 567.240 ; 
                RECT 303.760 566.920 307.800 567.240 ; 
                RECT 2.880 568.280 132.720 568.600 ; 
                RECT 145.320 568.280 155.840 568.600 ; 
                RECT 303.760 568.280 307.800 568.600 ; 
                RECT 2.880 569.640 155.840 569.960 ; 
                RECT 303.760 569.640 307.800 569.960 ; 
                RECT 2.880 571.000 139.520 571.320 ; 
                RECT 145.320 571.000 155.840 571.320 ; 
                RECT 303.760 571.000 307.800 571.320 ; 
                RECT 2.880 572.360 132.720 572.680 ; 
                RECT 145.320 572.360 155.840 572.680 ; 
                RECT 303.760 572.360 307.800 572.680 ; 
                RECT 2.880 573.720 132.720 574.040 ; 
                RECT 145.320 573.720 155.840 574.040 ; 
                RECT 303.760 573.720 307.800 574.040 ; 
                RECT 2.880 575.080 132.720 575.400 ; 
                RECT 145.320 575.080 155.840 575.400 ; 
                RECT 303.760 575.080 307.800 575.400 ; 
                RECT 2.880 576.440 132.720 576.760 ; 
                RECT 145.320 576.440 155.840 576.760 ; 
                RECT 303.760 576.440 307.800 576.760 ; 
                RECT 2.880 577.800 155.840 578.120 ; 
                RECT 303.760 577.800 307.800 578.120 ; 
                RECT 2.880 579.160 132.720 579.480 ; 
                RECT 145.320 579.160 155.840 579.480 ; 
                RECT 303.760 579.160 307.800 579.480 ; 
                RECT 2.880 580.520 142.240 580.840 ; 
                RECT 145.320 580.520 155.840 580.840 ; 
                RECT 303.760 580.520 307.800 580.840 ; 
                RECT 2.880 581.880 132.720 582.200 ; 
                RECT 145.320 581.880 155.840 582.200 ; 
                RECT 303.760 581.880 307.800 582.200 ; 
                RECT 2.880 583.240 132.720 583.560 ; 
                RECT 145.320 583.240 155.840 583.560 ; 
                RECT 303.760 583.240 307.800 583.560 ; 
                RECT 2.880 584.600 132.720 584.920 ; 
                RECT 145.320 584.600 155.840 584.920 ; 
                RECT 303.760 584.600 307.800 584.920 ; 
                RECT 2.880 585.960 155.840 586.280 ; 
                RECT 303.760 585.960 307.800 586.280 ; 
                RECT 2.880 587.320 133.400 587.640 ; 
                RECT 145.320 587.320 155.840 587.640 ; 
                RECT 303.760 587.320 307.800 587.640 ; 
                RECT 2.880 588.680 133.400 589.000 ; 
                RECT 145.320 588.680 155.840 589.000 ; 
                RECT 303.760 588.680 307.800 589.000 ; 
                RECT 2.880 590.040 136.800 590.360 ; 
                RECT 145.320 590.040 155.840 590.360 ; 
                RECT 303.760 590.040 307.800 590.360 ; 
                RECT 2.880 591.400 136.800 591.720 ; 
                RECT 145.320 591.400 155.840 591.720 ; 
                RECT 303.760 591.400 307.800 591.720 ; 
                RECT 2.880 592.760 133.400 593.080 ; 
                RECT 145.320 592.760 155.840 593.080 ; 
                RECT 303.760 592.760 307.800 593.080 ; 
                RECT 2.880 594.120 155.840 594.440 ; 
                RECT 303.760 594.120 307.800 594.440 ; 
                RECT 2.880 595.480 133.400 595.800 ; 
                RECT 145.320 595.480 155.840 595.800 ; 
                RECT 303.760 595.480 307.800 595.800 ; 
                RECT 2.880 596.840 133.400 597.160 ; 
                RECT 145.320 596.840 155.840 597.160 ; 
                RECT 303.760 596.840 307.800 597.160 ; 
                RECT 2.880 598.200 133.400 598.520 ; 
                RECT 145.320 598.200 155.840 598.520 ; 
                RECT 303.760 598.200 307.800 598.520 ; 
                RECT 2.880 599.560 133.400 599.880 ; 
                RECT 145.320 599.560 155.840 599.880 ; 
                RECT 303.760 599.560 307.800 599.880 ; 
                RECT 2.880 600.920 155.840 601.240 ; 
                RECT 303.760 600.920 307.800 601.240 ; 
                RECT 2.880 602.280 139.520 602.600 ; 
                RECT 145.320 602.280 155.840 602.600 ; 
                RECT 303.760 602.280 307.800 602.600 ; 
                RECT 2.880 603.640 133.400 603.960 ; 
                RECT 145.320 603.640 155.840 603.960 ; 
                RECT 303.760 603.640 307.800 603.960 ; 
                RECT 2.880 605.000 133.400 605.320 ; 
                RECT 145.320 605.000 155.840 605.320 ; 
                RECT 303.760 605.000 307.800 605.320 ; 
                RECT 2.880 606.360 133.400 606.680 ; 
                RECT 145.320 606.360 155.840 606.680 ; 
                RECT 303.760 606.360 307.800 606.680 ; 
                RECT 2.880 607.720 133.400 608.040 ; 
                RECT 145.320 607.720 155.840 608.040 ; 
                RECT 303.760 607.720 307.800 608.040 ; 
                RECT 2.880 609.080 155.840 609.400 ; 
                RECT 303.760 609.080 307.800 609.400 ; 
                RECT 2.880 610.440 141.560 610.760 ; 
                RECT 145.320 610.440 155.840 610.760 ; 
                RECT 303.760 610.440 307.800 610.760 ; 
                RECT 2.880 611.800 133.400 612.120 ; 
                RECT 145.320 611.800 155.840 612.120 ; 
                RECT 303.760 611.800 307.800 612.120 ; 
                RECT 2.880 613.160 133.400 613.480 ; 
                RECT 145.320 613.160 155.840 613.480 ; 
                RECT 303.760 613.160 307.800 613.480 ; 
                RECT 2.880 614.520 133.400 614.840 ; 
                RECT 145.320 614.520 155.840 614.840 ; 
                RECT 303.760 614.520 307.800 614.840 ; 
                RECT 2.880 615.880 133.400 616.200 ; 
                RECT 145.320 615.880 155.840 616.200 ; 
                RECT 303.760 615.880 307.800 616.200 ; 
                RECT 2.880 617.240 155.840 617.560 ; 
                RECT 303.760 617.240 307.800 617.560 ; 
                RECT 2.880 618.600 134.080 618.920 ; 
                RECT 145.320 618.600 155.840 618.920 ; 
                RECT 303.760 618.600 307.800 618.920 ; 
                RECT 2.880 619.960 136.120 620.280 ; 
                RECT 145.320 619.960 155.840 620.280 ; 
                RECT 303.760 619.960 307.800 620.280 ; 
                RECT 2.880 621.320 134.080 621.640 ; 
                RECT 145.320 621.320 155.840 621.640 ; 
                RECT 303.760 621.320 307.800 621.640 ; 
                RECT 2.880 622.680 134.080 623.000 ; 
                RECT 145.320 622.680 155.840 623.000 ; 
                RECT 303.760 622.680 307.800 623.000 ; 
                RECT 2.880 624.040 134.080 624.360 ; 
                RECT 145.320 624.040 155.840 624.360 ; 
                RECT 303.760 624.040 307.800 624.360 ; 
                RECT 2.880 625.400 155.840 625.720 ; 
                RECT 303.760 625.400 307.800 625.720 ; 
                RECT 2.880 626.760 134.080 627.080 ; 
                RECT 145.320 626.760 155.840 627.080 ; 
                RECT 303.760 626.760 307.800 627.080 ; 
                RECT 2.880 628.120 134.080 628.440 ; 
                RECT 145.320 628.120 155.840 628.440 ; 
                RECT 303.760 628.120 307.800 628.440 ; 
                RECT 2.880 629.480 138.840 629.800 ; 
                RECT 145.320 629.480 155.840 629.800 ; 
                RECT 303.760 629.480 307.800 629.800 ; 
                RECT 2.880 630.840 134.080 631.160 ; 
                RECT 145.320 630.840 155.840 631.160 ; 
                RECT 303.760 630.840 307.800 631.160 ; 
                RECT 2.880 632.200 134.080 632.520 ; 
                RECT 145.320 632.200 155.840 632.520 ; 
                RECT 303.760 632.200 307.800 632.520 ; 
                RECT 2.880 633.560 155.840 633.880 ; 
                RECT 303.760 633.560 307.800 633.880 ; 
                RECT 2.880 634.920 134.080 635.240 ; 
                RECT 145.320 634.920 155.840 635.240 ; 
                RECT 303.760 634.920 307.800 635.240 ; 
                RECT 2.880 636.280 134.080 636.600 ; 
                RECT 145.320 636.280 155.840 636.600 ; 
                RECT 303.760 636.280 307.800 636.600 ; 
                RECT 2.880 637.640 134.080 637.960 ; 
                RECT 145.320 637.640 155.840 637.960 ; 
                RECT 303.760 637.640 307.800 637.960 ; 
                RECT 2.880 639.000 140.880 639.320 ; 
                RECT 145.320 639.000 155.840 639.320 ; 
                RECT 303.760 639.000 307.800 639.320 ; 
                RECT 2.880 640.360 155.840 640.680 ; 
                RECT 303.760 640.360 307.800 640.680 ; 
                RECT 2.880 641.720 155.840 642.040 ; 
                RECT 303.760 641.720 307.800 642.040 ; 
                RECT 2.880 643.080 134.080 643.400 ; 
                RECT 145.320 643.080 155.840 643.400 ; 
                RECT 303.760 643.080 307.800 643.400 ; 
                RECT 2.880 644.440 134.080 644.760 ; 
                RECT 145.320 644.440 155.840 644.760 ; 
                RECT 303.760 644.440 307.800 644.760 ; 
                RECT 2.880 645.800 134.080 646.120 ; 
                RECT 145.320 645.800 155.840 646.120 ; 
                RECT 303.760 645.800 307.800 646.120 ; 
                RECT 2.880 647.160 134.080 647.480 ; 
                RECT 145.320 647.160 155.840 647.480 ; 
                RECT 303.760 647.160 307.800 647.480 ; 
                RECT 2.880 648.520 155.840 648.840 ; 
                RECT 303.760 648.520 307.800 648.840 ; 
                RECT 2.880 649.880 135.440 650.200 ; 
                RECT 145.320 649.880 155.840 650.200 ; 
                RECT 303.760 649.880 307.800 650.200 ; 
                RECT 2.880 651.240 134.080 651.560 ; 
                RECT 145.320 651.240 155.840 651.560 ; 
                RECT 303.760 651.240 307.800 651.560 ; 
                RECT 2.880 652.600 134.080 652.920 ; 
                RECT 145.320 652.600 155.840 652.920 ; 
                RECT 303.760 652.600 307.800 652.920 ; 
                RECT 2.880 653.960 134.080 654.280 ; 
                RECT 145.320 653.960 155.840 654.280 ; 
                RECT 303.760 653.960 307.800 654.280 ; 
                RECT 2.880 655.320 134.080 655.640 ; 
                RECT 145.320 655.320 155.840 655.640 ; 
                RECT 303.760 655.320 307.800 655.640 ; 
                RECT 2.880 656.680 155.840 657.000 ; 
                RECT 303.760 656.680 307.800 657.000 ; 
                RECT 2.880 658.040 134.080 658.360 ; 
                RECT 145.320 658.040 155.840 658.360 ; 
                RECT 303.760 658.040 307.800 658.360 ; 
                RECT 2.880 659.400 138.160 659.720 ; 
                RECT 145.320 659.400 155.840 659.720 ; 
                RECT 303.760 659.400 307.800 659.720 ; 
                RECT 2.880 660.760 134.080 661.080 ; 
                RECT 145.320 660.760 155.840 661.080 ; 
                RECT 303.760 660.760 307.800 661.080 ; 
                RECT 2.880 662.120 134.080 662.440 ; 
                RECT 145.320 662.120 155.840 662.440 ; 
                RECT 303.760 662.120 307.800 662.440 ; 
                RECT 2.880 663.480 134.080 663.800 ; 
                RECT 145.320 663.480 155.840 663.800 ; 
                RECT 303.760 663.480 307.800 663.800 ; 
                RECT 2.880 664.840 155.840 665.160 ; 
                RECT 303.760 664.840 307.800 665.160 ; 
                RECT 2.880 666.200 134.080 666.520 ; 
                RECT 145.320 666.200 155.840 666.520 ; 
                RECT 303.760 666.200 307.800 666.520 ; 
                RECT 2.880 667.560 134.080 667.880 ; 
                RECT 145.320 667.560 155.840 667.880 ; 
                RECT 303.760 667.560 307.800 667.880 ; 
                RECT 2.880 668.920 140.200 669.240 ; 
                RECT 145.320 668.920 155.840 669.240 ; 
                RECT 303.760 668.920 307.800 669.240 ; 
                RECT 2.880 670.280 134.080 670.600 ; 
                RECT 145.320 670.280 155.840 670.600 ; 
                RECT 303.760 670.280 307.800 670.600 ; 
                RECT 2.880 671.640 134.080 671.960 ; 
                RECT 145.320 671.640 155.840 671.960 ; 
                RECT 303.760 671.640 307.800 671.960 ; 
                RECT 2.880 673.000 155.840 673.320 ; 
                RECT 303.760 673.000 307.800 673.320 ; 
                RECT 2.880 674.360 134.080 674.680 ; 
                RECT 145.320 674.360 155.840 674.680 ; 
                RECT 303.760 674.360 307.800 674.680 ; 
                RECT 2.880 675.720 134.080 676.040 ; 
                RECT 145.320 675.720 155.840 676.040 ; 
                RECT 303.760 675.720 307.800 676.040 ; 
                RECT 2.880 677.080 134.080 677.400 ; 
                RECT 145.320 677.080 155.840 677.400 ; 
                RECT 303.760 677.080 307.800 677.400 ; 
                RECT 2.880 678.440 142.920 678.760 ; 
                RECT 145.320 678.440 155.840 678.760 ; 
                RECT 303.760 678.440 307.800 678.760 ; 
                RECT 2.880 679.800 134.080 680.120 ; 
                RECT 145.320 679.800 155.840 680.120 ; 
                RECT 303.760 679.800 307.800 680.120 ; 
                RECT 2.880 681.160 155.840 681.480 ; 
                RECT 303.760 681.160 307.800 681.480 ; 
                RECT 2.880 682.520 134.760 682.840 ; 
                RECT 145.320 682.520 155.840 682.840 ; 
                RECT 303.760 682.520 307.800 682.840 ; 
                RECT 2.880 683.880 134.760 684.200 ; 
                RECT 145.320 683.880 155.840 684.200 ; 
                RECT 303.760 683.880 307.800 684.200 ; 
                RECT 2.880 685.240 134.760 685.560 ; 
                RECT 145.320 685.240 155.840 685.560 ; 
                RECT 303.760 685.240 307.800 685.560 ; 
                RECT 2.880 686.600 134.760 686.920 ; 
                RECT 145.320 686.600 155.840 686.920 ; 
                RECT 303.760 686.600 307.800 686.920 ; 
                RECT 2.880 687.960 155.840 688.280 ; 
                RECT 303.760 687.960 307.800 688.280 ; 
                RECT 2.880 689.320 137.480 689.640 ; 
                RECT 145.320 689.320 155.840 689.640 ; 
                RECT 303.760 689.320 307.800 689.640 ; 
                RECT 2.880 690.680 134.760 691.000 ; 
                RECT 145.320 690.680 155.840 691.000 ; 
                RECT 303.760 690.680 307.800 691.000 ; 
                RECT 2.880 692.040 134.760 692.360 ; 
                RECT 145.320 692.040 155.840 692.360 ; 
                RECT 303.760 692.040 307.800 692.360 ; 
                RECT 2.880 693.400 134.760 693.720 ; 
                RECT 145.320 693.400 155.840 693.720 ; 
                RECT 303.760 693.400 307.800 693.720 ; 
                RECT 2.880 694.760 134.760 695.080 ; 
                RECT 145.320 694.760 155.840 695.080 ; 
                RECT 303.760 694.760 307.800 695.080 ; 
                RECT 2.880 696.120 155.840 696.440 ; 
                RECT 303.760 696.120 307.800 696.440 ; 
                RECT 2.880 697.480 139.520 697.800 ; 
                RECT 145.320 697.480 155.840 697.800 ; 
                RECT 303.760 697.480 307.800 697.800 ; 
                RECT 2.880 698.840 140.200 699.160 ; 
                RECT 145.320 698.840 155.840 699.160 ; 
                RECT 303.760 698.840 307.800 699.160 ; 
                RECT 2.880 700.200 134.760 700.520 ; 
                RECT 145.320 700.200 155.840 700.520 ; 
                RECT 303.760 700.200 307.800 700.520 ; 
                RECT 2.880 701.560 134.760 701.880 ; 
                RECT 145.320 701.560 155.840 701.880 ; 
                RECT 303.760 701.560 307.800 701.880 ; 
                RECT 2.880 702.920 134.760 703.240 ; 
                RECT 145.320 702.920 155.840 703.240 ; 
                RECT 303.760 702.920 307.800 703.240 ; 
                RECT 2.880 704.280 155.840 704.600 ; 
                RECT 303.760 704.280 307.800 704.600 ; 
                RECT 2.880 705.640 134.760 705.960 ; 
                RECT 145.320 705.640 155.840 705.960 ; 
                RECT 303.760 705.640 307.800 705.960 ; 
                RECT 2.880 707.000 134.760 707.320 ; 
                RECT 145.320 707.000 155.840 707.320 ; 
                RECT 303.760 707.000 307.800 707.320 ; 
                RECT 2.880 708.360 142.240 708.680 ; 
                RECT 145.320 708.360 155.840 708.680 ; 
                RECT 303.760 708.360 307.800 708.680 ; 
                RECT 2.880 709.720 134.760 710.040 ; 
                RECT 145.320 709.720 155.840 710.040 ; 
                RECT 303.760 709.720 307.800 710.040 ; 
                RECT 2.880 711.080 134.760 711.400 ; 
                RECT 145.320 711.080 155.840 711.400 ; 
                RECT 303.760 711.080 307.800 711.400 ; 
                RECT 2.880 712.440 155.840 712.760 ; 
                RECT 303.760 712.440 307.800 712.760 ; 
                RECT 2.880 713.800 135.440 714.120 ; 
                RECT 145.320 713.800 155.840 714.120 ; 
                RECT 303.760 713.800 307.800 714.120 ; 
                RECT 2.880 715.160 135.440 715.480 ; 
                RECT 145.320 715.160 155.840 715.480 ; 
                RECT 303.760 715.160 307.800 715.480 ; 
                RECT 2.880 716.520 135.440 716.840 ; 
                RECT 145.320 716.520 155.840 716.840 ; 
                RECT 303.760 716.520 307.800 716.840 ; 
                RECT 2.880 717.880 136.800 718.200 ; 
                RECT 145.320 717.880 155.840 718.200 ; 
                RECT 303.760 717.880 307.800 718.200 ; 
                RECT 2.880 719.240 135.440 719.560 ; 
                RECT 145.320 719.240 155.840 719.560 ; 
                RECT 303.760 719.240 307.800 719.560 ; 
                RECT 2.880 720.600 155.840 720.920 ; 
                RECT 303.760 720.600 307.800 720.920 ; 
                RECT 2.880 721.960 135.440 722.280 ; 
                RECT 145.320 721.960 155.840 722.280 ; 
                RECT 303.760 721.960 307.800 722.280 ; 
                RECT 2.880 723.320 135.440 723.640 ; 
                RECT 145.320 723.320 155.840 723.640 ; 
                RECT 303.760 723.320 307.800 723.640 ; 
                RECT 2.880 724.680 135.440 725.000 ; 
                RECT 145.320 724.680 155.840 725.000 ; 
                RECT 303.760 724.680 307.800 725.000 ; 
                RECT 2.880 726.040 135.440 726.360 ; 
                RECT 145.320 726.040 155.840 726.360 ; 
                RECT 303.760 726.040 307.800 726.360 ; 
                RECT 2.880 727.400 155.840 727.720 ; 
                RECT 303.760 727.400 307.800 727.720 ; 
                RECT 2.880 728.760 139.520 729.080 ; 
                RECT 145.320 728.760 155.840 729.080 ; 
                RECT 303.760 728.760 307.800 729.080 ; 
                RECT 2.880 730.120 135.440 730.440 ; 
                RECT 145.320 730.120 155.840 730.440 ; 
                RECT 303.760 730.120 307.800 730.440 ; 
                RECT 2.880 731.480 135.440 731.800 ; 
                RECT 145.320 731.480 155.840 731.800 ; 
                RECT 303.760 731.480 307.800 731.800 ; 
                RECT 2.880 732.840 135.440 733.160 ; 
                RECT 145.320 732.840 155.840 733.160 ; 
                RECT 303.760 732.840 307.800 733.160 ; 
                RECT 2.880 734.200 135.440 734.520 ; 
                RECT 145.320 734.200 155.840 734.520 ; 
                RECT 303.760 734.200 307.800 734.520 ; 
                RECT 2.880 735.560 155.840 735.880 ; 
                RECT 303.760 735.560 307.800 735.880 ; 
                RECT 2.880 736.920 141.560 737.240 ; 
                RECT 145.320 736.920 155.840 737.240 ; 
                RECT 303.760 736.920 307.800 737.240 ; 
                RECT 2.880 738.280 135.440 738.600 ; 
                RECT 145.320 738.280 155.840 738.600 ; 
                RECT 303.760 738.280 307.800 738.600 ; 
                RECT 2.880 739.640 135.440 739.960 ; 
                RECT 145.320 739.640 155.840 739.960 ; 
                RECT 303.760 739.640 307.800 739.960 ; 
                RECT 2.880 741.000 135.440 741.320 ; 
                RECT 145.320 741.000 155.840 741.320 ; 
                RECT 303.760 741.000 307.800 741.320 ; 
                RECT 2.880 742.360 135.440 742.680 ; 
                RECT 145.320 742.360 155.840 742.680 ; 
                RECT 303.760 742.360 307.800 742.680 ; 
                RECT 2.880 743.720 155.840 744.040 ; 
                RECT 303.760 743.720 307.800 744.040 ; 
                RECT 2.880 745.080 196.640 745.400 ; 
                RECT 303.760 745.080 307.800 745.400 ; 
                RECT 2.880 746.440 196.640 746.760 ; 
                RECT 303.760 746.440 307.800 746.760 ; 
                RECT 2.880 747.800 196.640 748.120 ; 
                RECT 303.760 747.800 307.800 748.120 ; 
                RECT 2.880 749.160 307.800 749.480 ; 
                RECT 2.880 750.520 307.800 750.840 ; 
                RECT 2.880 751.880 307.800 752.200 ; 
                RECT 2.880 753.240 307.800 753.560 ; 
                RECT 2.880 754.600 307.800 754.920 ; 
                RECT 2.880 2.880 307.800 4.240 ; 
                RECT 2.880 755.920 307.800 757.280 ; 
                RECT 200.780 42.775 206.580 43.895 ; 
                RECT 293.480 42.775 299.280 43.895 ; 
                RECT 200.780 48.565 206.580 49.185 ; 
                RECT 293.480 48.565 299.280 49.185 ; 
                RECT 200.780 53.645 206.580 54.295 ; 
                RECT 293.480 53.645 299.280 54.295 ; 
                RECT 200.780 58.875 206.580 59.525 ; 
                RECT 293.480 58.875 299.280 59.525 ; 
                RECT 200.780 95.840 299.280 99.440 ; 
                RECT 200.780 72.780 299.280 74.580 ; 
                RECT 200.780 89.730 299.280 90.530 ; 
                RECT 200.780 179.010 299.280 180.810 ; 
                RECT 200.780 84.840 299.280 85.640 ; 
                RECT 200.780 128.575 299.280 128.865 ; 
                RECT 200.780 86.520 299.280 87.320 ; 
                RECT 200.780 81.830 299.280 82.630 ; 
                RECT 200.780 33.405 299.280 35.205 ; 
                RECT 156.620 237.515 158.370 744.695 ; 
                RECT 169.975 237.515 171.895 744.695 ; 
                RECT 173.815 237.515 175.735 744.695 ; 
                RECT 117.730 57.215 118.620 127.015 ; 
                RECT 124.060 57.215 124.950 127.015 ; 
                RECT 130.820 57.215 131.710 127.015 ; 
                RECT 138.010 57.215 139.760 127.015 ; 
                RECT 151.780 57.215 153.700 127.015 ; 
                RECT 131.145 189.120 132.255 230.880 ; 
                RECT 138.660 189.120 139.550 230.880 ; 
                RECT 145.420 189.120 146.310 230.880 ; 
                RECT 151.750 189.120 152.640 230.880 ; 
                RECT 159.070 189.120 160.990 230.880 ; 
                RECT 166.250 177.960 167.140 183.120 ; 
                RECT 166.680 46.055 167.570 51.215 ; 
                RECT 77.080 238.580 86.240 238.950 ; 
                RECT 77.080 242.020 86.240 243.130 ; 
                RECT 36.140 220.240 55.780 220.910 ; 
                RECT 36.140 221.470 55.780 224.520 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 310.680 760.160 ; 
        LAYER met2 ;
            RECT 0.000 0.000 310.680 760.160 ; 
    END 
END sram22_2048x8m8w1 
END LIBRARY 

