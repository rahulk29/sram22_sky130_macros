VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sramgen_sram_32x32m2w8_replica_v1
  CLASS BLOCK ;
  ORIGIN 52.415 146.21 ;
  FOREIGN sramgen_sram_32x32m2w8_replica_v1 -52.415 -146.21 ;
  SIZE 234.875 BY 157.925 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -46.6 -145.81 -46.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -145.81 -44.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.4 -145.81 -43 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -145.81 -41.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.2 -98.9 -39.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -109.5 -38.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -145.81 -38.2 -138.54 ;
    END
    PORT
      LAYER met3 ;
        RECT -37 -145.81 -36.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -105.26 -35 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -145.81 -35 -113.1 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.8 -110.56 -33.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.2 -145.81 -31.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -104.2 -30.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -145.81 -30.2 -113.1 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -104.2 -28.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -145.81 -28.6 -112.04 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -109.5 -27 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -145.81 -27 -138.54 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.8 -145.81 -25.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -103.14 -23.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -145.81 -23.8 -113.1 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.6 -110.56 -22.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -109.5 -20.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -145.81 -20.6 -138.54 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.4 -145.81 -19 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -102.08 -17.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -145.81 -17.4 -113.1 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.2 -110.56 -15.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.6 -145.81 -14.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -101.02 -12.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -145.81 -12.6 -113.1 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -102.08 -11 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -145.81 -11 -112.04 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -109.5 -9.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -145.81 -9.4 -138.54 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.2 -145.81 -7.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -96.78 -6.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -145.81 -6.2 -112.04 ;
    END
    PORT
      LAYER met3 ;
        RECT -5 -145.81 -4.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.4 -145.81 -3 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 2.86 -1.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 -145.81 -1.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 2.86 0.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 -145.81 0.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 2.86 1.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 -145.81 1.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 2.86 3.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 -74.52 3.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 -145.81 3.4 -78.12 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 2.86 5 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 -145.81 5 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 2.86 6.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 -44.84 6.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 -111.62 6.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 2.86 8.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 -44.84 8.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 -116.92 8.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 2.86 9.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 -132.82 9.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 2.86 11.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 -44.84 11.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 2.86 13 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 -44.84 13 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 -145.81 13 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 2.86 14.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 -145.81 14.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 2.86 16.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 -44.84 16.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 -111.62 16.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 2.86 17.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 -44.84 17.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 2.86 19.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 -145.81 19.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 2.86 21 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 -44.84 21 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 -111.62 21 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 2.86 22.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 -44.84 22.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 -145.81 22.6 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 2.86 24.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 -145.81 24.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 2.86 25.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 -44.84 25.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 -111.62 25.8 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 2.86 27.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 -44.84 27.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 2.86 29 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 -116.92 29 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 -145.81 29 -138.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 2.86 30.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 -44.84 30.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 -111.62 30.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 2.86 32.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 -52.26 32.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 -145.81 32.2 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 2.86 33.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -145.81 33.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 2.86 35.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 -145.81 35.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 2.86 37 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 -52.26 37 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 2.86 38.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 -44.84 38.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 -116.92 38.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 2.86 40.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 -145.81 40.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 2.86 41.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 -52.26 41.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 -145.81 41.8 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 2.86 43.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 -44.84 43.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 -145.81 43.4 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 2.86 45 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 -145.81 45 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 2.86 46.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 -44.84 46.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 -111.62 46.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 2.86 48.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 -44.84 48.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 -116.92 48.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 2.86 49.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 -132.82 49.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 2.86 51.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 -44.84 51.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 2.86 53 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 -44.84 53 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 -145.81 53 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 2.86 54.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 -145.81 54.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 2.86 56.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 -44.84 56.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 -111.62 56.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 2.86 57.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 -44.84 57.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 2.86 59.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 -145.81 59.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 2.86 61 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 -44.84 61 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 -111.62 61 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 2.86 62.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 -44.84 62.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 -145.81 62.6 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 2.86 64.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 -145.81 64.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 2.86 65.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 -44.84 65.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 -111.62 65.8 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 2.86 67.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 -44.84 67.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 2.86 69 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 -116.92 69 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 -145.81 69 -138.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 2.86 70.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 -44.84 70.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 -111.62 70.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 2.86 72.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 -52.26 72.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 -145.81 72.2 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 2.86 73.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -145.81 73.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 2.86 75.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 -145.81 75.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 2.86 77 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 -52.26 77 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 2.86 78.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 -44.84 78.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 -116.92 78.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 2.86 80.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 -145.81 80.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 2.86 81.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 -52.26 81.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 -145.81 81.8 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 2.86 83.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 -44.84 83.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 -145.81 83.4 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 2.86 85 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 -145.81 85 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 2.86 86.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 -44.84 86.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 -111.62 86.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 2.86 88.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 -44.84 88.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 -116.92 88.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 2.86 89.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 -132.82 89.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 2.86 91.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 -44.84 91.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 2.86 93 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 -44.84 93 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 -145.81 93 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 2.86 94.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 -145.81 94.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 2.86 96.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 -44.84 96.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 -111.62 96.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 2.86 97.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 -44.84 97.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 2.86 99.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 -145.81 99.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 2.86 101 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 -44.84 101 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 -111.62 101 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 2.86 102.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 -44.84 102.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 -145.81 102.6 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 2.86 104.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 -145.81 104.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 2.86 105.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 -44.84 105.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 -111.62 105.8 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 2.86 107.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 -44.84 107.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 2.86 109 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 -116.92 109 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 -145.81 109 -138.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 2.86 110.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 -44.84 110.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 -111.62 110.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 2.86 112.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 -52.26 112.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 -145.81 112.2 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 2.86 113.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -145.81 113.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 2.86 115.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 -145.81 115.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 2.86 117 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 -52.26 117 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 2.86 118.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 -44.84 118.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 -116.92 118.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 2.86 120.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 -145.81 120.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 2.86 121.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 -52.26 121.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 -145.81 121.8 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 2.86 123.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 -44.84 123.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 -145.81 123.4 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 2.86 125 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 -145.81 125 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 2.86 126.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 -44.84 126.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 -111.62 126.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 2.86 128.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 -44.84 128.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 -116.92 128.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 2.86 129.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 -132.82 129.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 2.86 131.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 -44.84 131.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 2.86 133 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 -44.84 133 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 -145.81 133 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 2.86 134.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 -145.81 134.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 2.86 136.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 -44.84 136.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 -111.62 136.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 2.86 137.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 -44.84 137.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 2.86 139.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 -145.81 139.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 2.86 141 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 -44.84 141 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 -111.62 141 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 2.86 142.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 -44.84 142.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 -145.81 142.6 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 2.86 144.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 -145.81 144.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 2.86 145.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 -44.84 145.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 -111.62 145.8 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 2.86 147.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 -44.84 147.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 2.86 149 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 -116.92 149 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 -145.81 149 -138.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 2.86 150.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 -44.84 150.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 -111.62 150.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 2.86 152.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 -52.26 152.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 -145.81 152.2 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 2.86 153.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -145.81 153.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 2.86 155.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 -145.81 155.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 2.86 157 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 -52.26 157 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 2.86 158.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 -44.84 158.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 -116.92 158.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 2.86 160.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 -145.81 160.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 2.86 161.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 -52.26 161.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 -145.81 161.8 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 2.86 163.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 -44.84 163.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 -145.81 163.4 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 2.86 165 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 -145.81 165 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 2.86 166.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 -145.81 166.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 2.86 168.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 -145.81 168.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 2.86 169.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 -145.81 169.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 171 -145.81 171.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 -145.81 173 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 -145.81 174.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.8 -145.81 176.2 11.315 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -47.4 -144.27 -47 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.8 -144.27 -45.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -144.27 -43.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.6 -144.27 -42.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -98.9 -40.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.4 -109.5 -39 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.8 -144.27 -37.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -105.26 -35.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -144.27 -35.8 -113.1 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.6 -105.26 -34.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -109.5 -32.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -144.27 -32.6 -138.54 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.4 -144.27 -31 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -104.2 -29.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -144.27 -29.4 -113.1 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.2 -110.56 -27.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -109.5 -26.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -144.27 -26.2 -138.54 ;
    END
    PORT
      LAYER met3 ;
        RECT -25 -144.27 -24.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -103.14 -23 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -144.27 -23 -112.04 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.8 -109.5 -21.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.2 -144.27 -19.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -102.08 -18.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -144.27 -18.2 -113.1 ;
    END
    PORT
      LAYER met3 ;
        RECT -17 -35.3 -16.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -17 -103.14 -16.6 -80.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -109.5 -15 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -144.27 -15 -138.54 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.8 -144.27 -13.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -101.02 -11.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -144.27 -11.8 -113.1 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -110.56 -10.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -109.5 -8.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -144.27 -8.6 -138.54 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.4 -144.27 -7 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -96.78 -5.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -144.27 -5.4 -112.04 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.2 -144.27 -3.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.6 -144.27 -2.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 2.86 -0.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 -144.27 -0.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 2.86 1 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 -144.27 1 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 2.86 2.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 -144.27 2.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 2.86 4.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 -74.52 4.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 -144.27 4.2 -78.12 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 2.86 5.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 -44.84 5.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 -111.62 5.8 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 2.86 7.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 -44.84 7.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 2.86 9 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 -116.92 9 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 2.86 10.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 -44.84 10.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 -111.62 10.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 2.86 12.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 -52.26 12.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 -144.27 12.2 -135.36 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 2.86 13.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -144.27 13.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 2.86 15.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 -144.27 15.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 2.86 17 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 -52.26 17 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 2.86 18.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 -44.84 18.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 -116.92 18.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 2.86 20.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 -144.27 20.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 2.86 21.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 -52.26 21.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 -144.27 21.8 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 2.86 23.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 -44.84 23.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 -144.27 23.4 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 2.86 25 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 -144.27 25 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 2.86 26.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 -44.84 26.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 -111.62 26.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 2.86 28.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 -44.84 28.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 -116.92 28.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 2.86 29.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 -144.27 29.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 2.86 31.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 -44.84 31.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 -111.62 31.4 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 2.86 33 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 -44.84 33 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 -144.27 33 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 2.86 34.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 -144.27 34.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 2.86 36.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 -44.84 36.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 -111.62 36.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 2.86 37.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 -44.84 37.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 2.86 39.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 -144.27 39.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 2.86 41 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 -44.84 41 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 -111.62 41 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 2.86 42.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 -44.84 42.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 -144.27 42.6 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 2.86 44.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 -144.27 44.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 2.86 45.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 -44.84 45.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 -111.62 45.8 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 2.86 47.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 -44.84 47.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 2.86 49 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 -116.92 49 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 2.86 50.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 -44.84 50.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 -111.62 50.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 2.86 52.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 -52.26 52.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 -144.27 52.2 -135.36 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 2.86 53.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -144.27 53.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 2.86 55.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 -144.27 55.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 2.86 57 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 -52.26 57 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 2.86 58.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 -44.84 58.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 -116.92 58.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 2.86 60.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 -144.27 60.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 2.86 61.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 -52.26 61.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 -144.27 61.8 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 2.86 63.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 -44.84 63.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 -144.27 63.4 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 2.86 65 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 -144.27 65 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 2.86 66.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 -44.84 66.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 -111.62 66.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 2.86 68.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 -44.84 68.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 -116.92 68.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 2.86 69.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 -144.27 69.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 2.86 71.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 -44.84 71.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 -111.62 71.4 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 2.86 73 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 -44.84 73 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 -144.27 73 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 2.86 74.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 -144.27 74.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 2.86 76.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 -44.84 76.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 -111.62 76.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 2.86 77.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 -44.84 77.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 2.86 79.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 -144.27 79.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 2.86 81 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 -44.84 81 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 -111.62 81 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 2.86 82.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 -44.84 82.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 -144.27 82.6 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 2.86 84.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 -144.27 84.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 2.86 85.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 -44.84 85.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 -111.62 85.8 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 2.86 87.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 -44.84 87.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 2.86 89 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 -116.92 89 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 2.86 90.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 -44.84 90.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 -111.62 90.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 2.86 92.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 -52.26 92.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 -144.27 92.2 -135.36 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 2.86 93.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -144.27 93.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 2.86 95.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 -144.27 95.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 2.86 97 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 -52.26 97 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 2.86 98.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 -44.84 98.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 -116.92 98.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 2.86 100.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 -144.27 100.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 2.86 101.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 -52.26 101.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 -144.27 101.8 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 2.86 103.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 -44.84 103.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 -144.27 103.4 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 2.86 105 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 -144.27 105 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 2.86 106.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 -44.84 106.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 -111.62 106.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 2.86 108.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 -44.84 108.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 -116.92 108.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 2.86 109.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 -144.27 109.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 2.86 111.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 -44.84 111.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 -111.62 111.4 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 2.86 113 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 -44.84 113 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 -144.27 113 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 2.86 114.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 -144.27 114.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 2.86 116.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 -44.84 116.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 -111.62 116.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 2.86 117.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 -44.84 117.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 2.86 119.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 -144.27 119.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 2.86 121 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 -44.84 121 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 -111.62 121 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 2.86 122.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 -44.84 122.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 -144.27 122.6 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 2.86 124.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 -144.27 124.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 2.86 125.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 -44.84 125.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 -111.62 125.8 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 2.86 127.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 -44.84 127.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 2.86 129 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 -116.92 129 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 2.86 130.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 -44.84 130.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 -111.62 130.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 2.86 132.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 -52.26 132.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 -144.27 132.2 -135.36 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 2.86 133.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -144.27 133.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 2.86 135.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 -144.27 135.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 2.86 137 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 -52.26 137 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 2.86 138.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 -44.84 138.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 -116.92 138.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 2.86 140.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 -144.27 140.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 2.86 141.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 -52.26 141.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 -144.27 141.8 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 2.86 143.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 -44.84 143.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 -144.27 143.4 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 2.86 145 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 -144.27 145 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 2.86 146.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 -44.84 146.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 -111.62 146.6 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 2.86 148.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 -44.84 148.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 -116.92 148.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 2.86 149.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 -144.27 149.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 2.86 151.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 -44.84 151.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 -111.62 151.4 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 2.86 153 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 -44.84 153 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 -144.27 153 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 2.86 154.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 -144.27 154.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 2.86 156.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 -44.84 156.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 -111.62 156.2 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 2.86 157.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 -44.84 157.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 2.86 159.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 -144.27 159.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 2.86 161 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 -44.84 161 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 -111.62 161 -102.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 2.86 162.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 -44.84 162.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 -144.27 162.6 -125.82 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 2.86 164.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 -144.27 164.2 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 2.86 165.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 -144.27 165.8 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 2.86 167.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 -144.27 167.4 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 2.86 169 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 -144.27 169 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 2.86 170.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 -144.27 170.6 -34.66 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.8 -144.27 172.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 -144.27 173.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 -144.27 175.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.6 -144.27 177 9.775 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -16.46 -146.21 -16.16 -145.91 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -22.3 -146.21 -22 -145.91 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -28.14 -146.21 -27.84 -145.91 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -33.98 -146.21 -33.68 -145.91 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -39.82 -146.21 -39.52 -145.91 ;
    END
  END addr[4]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -40.84 -146.21 -40.42 -145.79 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 7.015 -146.21 7.315 -145.91 ;
    END
  END din[0]
  PIN din[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 57.015 -146.21 57.315 -145.91 ;
    END
  END din[10]
  PIN din[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 57.63 -146.21 57.93 -145.91 ;
    END
  END din[11]
  PIN din[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.015 -146.21 67.315 -145.91 ;
    END
  END din[12]
  PIN din[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 67.63 -146.21 67.93 -145.91 ;
    END
  END din[13]
  PIN din[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 77.015 -146.21 77.315 -145.91 ;
    END
  END din[14]
  PIN din[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 77.63 -146.21 77.93 -145.91 ;
    END
  END din[15]
  PIN din[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 87.015 -146.21 87.315 -145.91 ;
    END
  END din[16]
  PIN din[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 87.63 -146.21 87.93 -145.91 ;
    END
  END din[17]
  PIN din[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 97.015 -146.21 97.315 -145.91 ;
    END
  END din[18]
  PIN din[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 97.63 -146.21 97.93 -145.91 ;
    END
  END din[19]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 7.63 -146.21 7.93 -145.91 ;
    END
  END din[1]
  PIN din[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.015 -146.21 107.315 -145.91 ;
    END
  END din[20]
  PIN din[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 107.63 -146.21 107.93 -145.91 ;
    END
  END din[21]
  PIN din[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.015 -146.21 117.315 -145.91 ;
    END
  END din[22]
  PIN din[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 117.63 -146.21 117.93 -145.91 ;
    END
  END din[23]
  PIN din[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 127.015 -146.21 127.315 -145.91 ;
    END
  END din[24]
  PIN din[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 127.63 -146.21 127.93 -145.91 ;
    END
  END din[25]
  PIN din[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 137.015 -146.21 137.315 -145.91 ;
    END
  END din[26]
  PIN din[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 137.63 -146.21 137.93 -145.91 ;
    END
  END din[27]
  PIN din[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 147.015 -146.21 147.315 -145.91 ;
    END
  END din[28]
  PIN din[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 147.63 -146.21 147.93 -145.91 ;
    END
  END din[29]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.015 -146.21 17.315 -145.91 ;
    END
  END din[2]
  PIN din[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 157.015 -146.21 157.315 -145.91 ;
    END
  END din[30]
  PIN din[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 157.63 -146.21 157.93 -145.91 ;
    END
  END din[31]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.63 -146.21 17.93 -145.91 ;
    END
  END din[3]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 27.015 -146.21 27.315 -145.91 ;
    END
  END din[4]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 27.63 -146.21 27.93 -145.91 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 37.015 -146.21 37.315 -145.91 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 37.63 -146.21 37.93 -145.91 ;
    END
  END din[7]
  PIN din[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 47.015 -146.21 47.315 -145.91 ;
    END
  END din[8]
  PIN din[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 47.63 -146.21 47.93 -145.91 ;
    END
  END din[9]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.785 -146.21 6.085 -145.91 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 55.785 -146.21 56.085 -145.91 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.785 -146.21 61.085 -145.91 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 65.785 -146.21 66.085 -145.91 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 70.785 -146.21 71.085 -145.91 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.785 -146.21 76.085 -145.91 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.785 -146.21 81.085 -145.91 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 85.785 -146.21 86.085 -145.91 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 90.785 -146.21 91.085 -145.91 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 95.785 -146.21 96.085 -145.91 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 100.785 -146.21 101.085 -145.91 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 10.785 -146.21 11.085 -145.91 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 105.785 -146.21 106.085 -145.91 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 110.785 -146.21 111.085 -145.91 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 115.785 -146.21 116.085 -145.91 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 120.785 -146.21 121.085 -145.91 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 125.785 -146.21 126.085 -145.91 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 130.785 -146.21 131.085 -145.91 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 135.785 -146.21 136.085 -145.91 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 140.785 -146.21 141.085 -145.91 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 145.785 -146.21 146.085 -145.91 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 150.785 -146.21 151.085 -145.91 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 15.785 -146.21 16.085 -145.91 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 155.785 -146.21 156.085 -145.91 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 160.785 -146.21 161.085 -145.91 ;
    END
  END dout[31]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 20.785 -146.21 21.085 -145.91 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.785 -146.21 26.085 -145.91 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 30.785 -146.21 31.085 -145.91 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 35.785 -146.21 36.085 -145.91 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 40.785 -146.21 41.085 -145.91 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 45.785 -146.21 46.085 -145.91 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 50.785 -146.21 51.085 -145.91 ;
    END
  END dout[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -10.62 -146.21 -10.32 -145.91 ;
    END
  END we
  PIN wmask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 9.125 -146.21 9.425 -145.91 ;
    END
  END wmask[0]
  PIN wmask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 49.125 -146.21 49.425 -145.91 ;
    END
  END wmask[1]
  PIN wmask[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 89.125 -146.21 89.425 -145.91 ;
    END
  END wmask[2]
  PIN wmask[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 129.125 -146.21 129.425 -145.91 ;
    END
  END wmask[3]
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -52.415 -146.21 182.46 11.715 ;
    LAYER met2 SPACING 0.14 ;
      RECT -52.415 -146.21 182.46 11.715 ;
    LAYER met3 SPACING 0.3 ;
      RECT 162.615 -85.91 162.945 -85.58 ;
      RECT 162.63 -101.34 162.93 -85.58 ;
      RECT 162.615 -101.34 162.945 -101.01 ;
      RECT 162.63 -82.125 162.93 -45.52 ;
      RECT 162.615 -47.495 162.945 -47.165 ;
      RECT 162.615 -81.715 162.945 -81.385 ;
      RECT 162.015 -125.23 162.315 -53.42 ;
      RECT 162 -53.795 162.33 -53.465 ;
      RECT 162 -69.495 162.33 -69.165 ;
      RECT 162 -125.23 162.33 -124.9 ;
      RECT 160.77 -112.315 161.1 -111.985 ;
      RECT 160.785 -145.42 161.085 -111.985 ;
      RECT 160.77 -86.37 161.1 -86.04 ;
      RECT 160.785 -101.34 161.085 -86.04 ;
      RECT 160.77 -101.34 161.1 -101.01 ;
      RECT 160.785 -82.145 161.085 -45.52 ;
      RECT 160.77 -45.895 161.1 -45.565 ;
      RECT 160.77 -82.145 161.1 -81.815 ;
      RECT 158.245 -117.705 158.575 -117.375 ;
      RECT 158.26 -138.15 158.56 -117.375 ;
      RECT 158.245 -124.945 158.575 -124.615 ;
      RECT 158.245 -138.105 158.575 -137.775 ;
      RECT 157.615 -124.145 157.945 -123.815 ;
      RECT 157.63 -145.42 157.93 -123.815 ;
      RECT 157.615 -85.91 157.945 -85.58 ;
      RECT 157.63 -101.34 157.93 -85.58 ;
      RECT 157.615 -101.34 157.945 -101.01 ;
      RECT 157.63 -82.125 157.93 -45.52 ;
      RECT 157.615 -47.495 157.945 -47.165 ;
      RECT 157.615 -81.715 157.945 -81.385 ;
      RECT 157 -118.505 157.33 -118.175 ;
      RECT 157.015 -145.42 157.315 -118.175 ;
      RECT 157.015 -117.22 157.315 -53.42 ;
      RECT 157 -53.795 157.33 -53.465 ;
      RECT 157 -69.495 157.33 -69.165 ;
      RECT 157 -117.22 157.33 -116.89 ;
      RECT 155.77 -112.315 156.1 -111.985 ;
      RECT 155.785 -145.42 156.085 -111.985 ;
      RECT 155.77 -86.37 156.1 -86.04 ;
      RECT 155.785 -101.34 156.085 -86.04 ;
      RECT 155.77 -101.34 156.1 -101.01 ;
      RECT 155.785 -82.145 156.085 -45.52 ;
      RECT 155.77 -45.895 156.1 -45.565 ;
      RECT 155.77 -82.145 156.1 -81.815 ;
      RECT 152.615 -85.91 152.945 -85.58 ;
      RECT 152.63 -101.34 152.93 -85.58 ;
      RECT 152.615 -101.34 152.945 -101.01 ;
      RECT 152.63 -82.125 152.93 -45.52 ;
      RECT 152.615 -47.495 152.945 -47.165 ;
      RECT 152.615 -81.715 152.945 -81.385 ;
      RECT 152.015 -125.23 152.315 -53.42 ;
      RECT 152 -53.795 152.33 -53.465 ;
      RECT 152 -69.495 152.33 -69.165 ;
      RECT 152 -125.23 152.33 -124.9 ;
      RECT 150.77 -112.315 151.1 -111.985 ;
      RECT 150.785 -145.42 151.085 -111.985 ;
      RECT 150.77 -86.37 151.1 -86.04 ;
      RECT 150.785 -101.34 151.085 -86.04 ;
      RECT 150.77 -101.34 151.1 -101.01 ;
      RECT 150.785 -82.145 151.085 -45.52 ;
      RECT 150.77 -45.895 151.1 -45.565 ;
      RECT 150.77 -82.145 151.1 -81.815 ;
      RECT 148.245 -117.705 148.575 -117.375 ;
      RECT 148.26 -138.15 148.56 -117.375 ;
      RECT 148.245 -124.945 148.575 -124.615 ;
      RECT 148.245 -138.105 148.575 -137.775 ;
      RECT 147.615 -124.145 147.945 -123.815 ;
      RECT 147.63 -145.42 147.93 -123.815 ;
      RECT 147.615 -85.91 147.945 -85.58 ;
      RECT 147.63 -101.34 147.93 -85.58 ;
      RECT 147.615 -101.34 147.945 -101.01 ;
      RECT 147.63 -82.125 147.93 -45.52 ;
      RECT 147.615 -47.495 147.945 -47.165 ;
      RECT 147.615 -81.715 147.945 -81.385 ;
      RECT 147 -118.505 147.33 -118.175 ;
      RECT 147.015 -145.42 147.315 -118.175 ;
      RECT 147.015 -117.22 147.315 -53.42 ;
      RECT 147 -53.795 147.33 -53.465 ;
      RECT 147 -69.495 147.33 -69.165 ;
      RECT 147 -117.22 147.33 -116.89 ;
      RECT 145.77 -112.315 146.1 -111.985 ;
      RECT 145.785 -145.42 146.085 -111.985 ;
      RECT 145.77 -86.37 146.1 -86.04 ;
      RECT 145.785 -101.34 146.085 -86.04 ;
      RECT 145.77 -101.34 146.1 -101.01 ;
      RECT 145.785 -82.145 146.085 -45.52 ;
      RECT 145.77 -45.895 146.1 -45.565 ;
      RECT 145.77 -82.145 146.1 -81.815 ;
      RECT 142.615 -85.91 142.945 -85.58 ;
      RECT 142.63 -101.34 142.93 -85.58 ;
      RECT 142.615 -101.34 142.945 -101.01 ;
      RECT 142.63 -82.125 142.93 -45.52 ;
      RECT 142.615 -47.495 142.945 -47.165 ;
      RECT 142.615 -81.715 142.945 -81.385 ;
      RECT 142.015 -125.23 142.315 -53.42 ;
      RECT 142 -53.795 142.33 -53.465 ;
      RECT 142 -69.495 142.33 -69.165 ;
      RECT 142 -125.23 142.33 -124.9 ;
      RECT 140.77 -112.315 141.1 -111.985 ;
      RECT 140.785 -145.42 141.085 -111.985 ;
      RECT 140.77 -86.37 141.1 -86.04 ;
      RECT 140.785 -101.34 141.085 -86.04 ;
      RECT 140.77 -101.34 141.1 -101.01 ;
      RECT 140.785 -82.145 141.085 -45.52 ;
      RECT 140.77 -45.895 141.1 -45.565 ;
      RECT 140.77 -82.145 141.1 -81.815 ;
      RECT 138.245 -117.705 138.575 -117.375 ;
      RECT 138.26 -138.15 138.56 -117.375 ;
      RECT 138.245 -124.945 138.575 -124.615 ;
      RECT 138.245 -138.105 138.575 -137.775 ;
      RECT 137.615 -124.145 137.945 -123.815 ;
      RECT 137.63 -145.42 137.93 -123.815 ;
      RECT 137.615 -85.91 137.945 -85.58 ;
      RECT 137.63 -101.34 137.93 -85.58 ;
      RECT 137.615 -101.34 137.945 -101.01 ;
      RECT 137.63 -82.125 137.93 -45.52 ;
      RECT 137.615 -47.495 137.945 -47.165 ;
      RECT 137.615 -81.715 137.945 -81.385 ;
      RECT 137 -118.505 137.33 -118.175 ;
      RECT 137.015 -145.42 137.315 -118.175 ;
      RECT 137.015 -117.22 137.315 -53.42 ;
      RECT 137 -53.795 137.33 -53.465 ;
      RECT 137 -69.495 137.33 -69.165 ;
      RECT 137 -117.22 137.33 -116.89 ;
      RECT 135.77 -112.315 136.1 -111.985 ;
      RECT 135.785 -145.42 136.085 -111.985 ;
      RECT 135.77 -86.37 136.1 -86.04 ;
      RECT 135.785 -101.34 136.085 -86.04 ;
      RECT 135.77 -101.34 136.1 -101.01 ;
      RECT 135.785 -82.145 136.085 -45.52 ;
      RECT 135.77 -45.895 136.1 -45.565 ;
      RECT 135.77 -82.145 136.1 -81.815 ;
      RECT 132.615 -85.91 132.945 -85.58 ;
      RECT 132.63 -101.34 132.93 -85.58 ;
      RECT 132.615 -101.34 132.945 -101.01 ;
      RECT 132.63 -82.125 132.93 -45.52 ;
      RECT 132.615 -47.495 132.945 -47.165 ;
      RECT 132.615 -81.715 132.945 -81.385 ;
      RECT 132.015 -125.23 132.315 -53.42 ;
      RECT 132 -53.795 132.33 -53.465 ;
      RECT 132 -69.495 132.33 -69.165 ;
      RECT 132 -125.23 132.33 -124.9 ;
      RECT 131.4 -134.07 131.7 -58.145 ;
      RECT 131.385 -58.52 131.715 -58.19 ;
      RECT 131.385 -134.07 131.715 -133.74 ;
      RECT 130.77 -112.315 131.1 -111.985 ;
      RECT 130.785 -145.42 131.085 -111.985 ;
      RECT 130.77 -86.37 131.1 -86.04 ;
      RECT 130.785 -101.34 131.085 -86.04 ;
      RECT 130.77 -101.34 131.1 -101.01 ;
      RECT 130.785 -82.145 131.085 -45.52 ;
      RECT 130.77 -45.895 131.1 -45.565 ;
      RECT 130.77 -82.145 131.1 -81.815 ;
      RECT 129.11 -134.445 129.44 -134.115 ;
      RECT 129.125 -145.42 129.425 -134.115 ;
      RECT 128.245 -117.705 128.575 -117.375 ;
      RECT 128.26 -138.15 128.56 -117.375 ;
      RECT 128.245 -124.945 128.575 -124.615 ;
      RECT 128.245 -133.645 128.575 -133.315 ;
      RECT 128.245 -138.105 128.575 -137.775 ;
      RECT 127.615 -124.145 127.945 -123.815 ;
      RECT 127.63 -145.42 127.93 -123.815 ;
      RECT 127.615 -85.91 127.945 -85.58 ;
      RECT 127.63 -101.34 127.93 -85.58 ;
      RECT 127.615 -101.34 127.945 -101.01 ;
      RECT 127.63 -82.125 127.93 -45.52 ;
      RECT 127.615 -47.495 127.945 -47.165 ;
      RECT 127.615 -81.715 127.945 -81.385 ;
      RECT 127 -118.505 127.33 -118.175 ;
      RECT 127.015 -145.42 127.315 -118.175 ;
      RECT 127.015 -117.22 127.315 -53.42 ;
      RECT 127 -53.795 127.33 -53.465 ;
      RECT 127 -69.495 127.33 -69.165 ;
      RECT 127 -117.22 127.33 -116.89 ;
      RECT 125.77 -112.315 126.1 -111.985 ;
      RECT 125.785 -145.42 126.085 -111.985 ;
      RECT 125.77 -86.37 126.1 -86.04 ;
      RECT 125.785 -101.34 126.085 -86.04 ;
      RECT 125.77 -101.34 126.1 -101.01 ;
      RECT 125.785 -82.145 126.085 -45.52 ;
      RECT 125.77 -45.895 126.1 -45.565 ;
      RECT 125.77 -82.145 126.1 -81.815 ;
      RECT 122.615 -85.91 122.945 -85.58 ;
      RECT 122.63 -101.34 122.93 -85.58 ;
      RECT 122.615 -101.34 122.945 -101.01 ;
      RECT 122.63 -82.125 122.93 -45.52 ;
      RECT 122.615 -47.495 122.945 -47.165 ;
      RECT 122.615 -81.715 122.945 -81.385 ;
      RECT 122.015 -125.23 122.315 -53.42 ;
      RECT 122 -53.795 122.33 -53.465 ;
      RECT 122 -69.495 122.33 -69.165 ;
      RECT 122 -125.23 122.33 -124.9 ;
      RECT 120.77 -112.315 121.1 -111.985 ;
      RECT 120.785 -145.42 121.085 -111.985 ;
      RECT 120.77 -86.37 121.1 -86.04 ;
      RECT 120.785 -101.34 121.085 -86.04 ;
      RECT 120.77 -101.34 121.1 -101.01 ;
      RECT 120.785 -82.145 121.085 -45.52 ;
      RECT 120.77 -45.895 121.1 -45.565 ;
      RECT 120.77 -82.145 121.1 -81.815 ;
      RECT 118.245 -117.705 118.575 -117.375 ;
      RECT 118.26 -138.15 118.56 -117.375 ;
      RECT 118.245 -124.945 118.575 -124.615 ;
      RECT 118.245 -138.105 118.575 -137.775 ;
      RECT 117.615 -124.145 117.945 -123.815 ;
      RECT 117.63 -145.42 117.93 -123.815 ;
      RECT 117.615 -85.91 117.945 -85.58 ;
      RECT 117.63 -101.34 117.93 -85.58 ;
      RECT 117.615 -101.34 117.945 -101.01 ;
      RECT 117.63 -82.125 117.93 -45.52 ;
      RECT 117.615 -47.495 117.945 -47.165 ;
      RECT 117.615 -81.715 117.945 -81.385 ;
      RECT 117 -118.505 117.33 -118.175 ;
      RECT 117.015 -145.42 117.315 -118.175 ;
      RECT 117.015 -117.22 117.315 -53.42 ;
      RECT 117 -53.795 117.33 -53.465 ;
      RECT 117 -69.495 117.33 -69.165 ;
      RECT 117 -117.22 117.33 -116.89 ;
      RECT 115.77 -112.315 116.1 -111.985 ;
      RECT 115.785 -145.42 116.085 -111.985 ;
      RECT 115.77 -86.37 116.1 -86.04 ;
      RECT 115.785 -101.34 116.085 -86.04 ;
      RECT 115.77 -101.34 116.1 -101.01 ;
      RECT 115.785 -82.145 116.085 -45.52 ;
      RECT 115.77 -45.895 116.1 -45.565 ;
      RECT 115.77 -82.145 116.1 -81.815 ;
      RECT 112.615 -85.91 112.945 -85.58 ;
      RECT 112.63 -101.34 112.93 -85.58 ;
      RECT 112.615 -101.34 112.945 -101.01 ;
      RECT 112.63 -82.125 112.93 -45.52 ;
      RECT 112.615 -47.495 112.945 -47.165 ;
      RECT 112.615 -81.715 112.945 -81.385 ;
      RECT 112.015 -125.23 112.315 -53.42 ;
      RECT 112 -53.795 112.33 -53.465 ;
      RECT 112 -69.495 112.33 -69.165 ;
      RECT 112 -125.23 112.33 -124.9 ;
      RECT 110.77 -112.315 111.1 -111.985 ;
      RECT 110.785 -145.42 111.085 -111.985 ;
      RECT 110.77 -86.37 111.1 -86.04 ;
      RECT 110.785 -101.34 111.085 -86.04 ;
      RECT 110.77 -101.34 111.1 -101.01 ;
      RECT 110.785 -82.145 111.085 -45.52 ;
      RECT 110.77 -45.895 111.1 -45.565 ;
      RECT 110.77 -82.145 111.1 -81.815 ;
      RECT 108.245 -117.705 108.575 -117.375 ;
      RECT 108.26 -138.15 108.56 -117.375 ;
      RECT 108.245 -124.945 108.575 -124.615 ;
      RECT 108.245 -138.105 108.575 -137.775 ;
      RECT 107.615 -124.145 107.945 -123.815 ;
      RECT 107.63 -145.42 107.93 -123.815 ;
      RECT 107.615 -85.91 107.945 -85.58 ;
      RECT 107.63 -101.34 107.93 -85.58 ;
      RECT 107.615 -101.34 107.945 -101.01 ;
      RECT 107.63 -82.125 107.93 -45.52 ;
      RECT 107.615 -47.495 107.945 -47.165 ;
      RECT 107.615 -81.715 107.945 -81.385 ;
      RECT 107 -118.505 107.33 -118.175 ;
      RECT 107.015 -145.42 107.315 -118.175 ;
      RECT 107.015 -117.22 107.315 -53.42 ;
      RECT 107 -53.795 107.33 -53.465 ;
      RECT 107 -69.495 107.33 -69.165 ;
      RECT 107 -117.22 107.33 -116.89 ;
      RECT 105.77 -112.315 106.1 -111.985 ;
      RECT 105.785 -145.42 106.085 -111.985 ;
      RECT 105.77 -86.37 106.1 -86.04 ;
      RECT 105.785 -101.34 106.085 -86.04 ;
      RECT 105.77 -101.34 106.1 -101.01 ;
      RECT 105.785 -82.145 106.085 -45.52 ;
      RECT 105.77 -45.895 106.1 -45.565 ;
      RECT 105.77 -82.145 106.1 -81.815 ;
      RECT 102.615 -85.91 102.945 -85.58 ;
      RECT 102.63 -101.34 102.93 -85.58 ;
      RECT 102.615 -101.34 102.945 -101.01 ;
      RECT 102.63 -82.125 102.93 -45.52 ;
      RECT 102.615 -47.495 102.945 -47.165 ;
      RECT 102.615 -81.715 102.945 -81.385 ;
      RECT 102.015 -125.23 102.315 -53.42 ;
      RECT 102 -53.795 102.33 -53.465 ;
      RECT 102 -69.495 102.33 -69.165 ;
      RECT 102 -125.23 102.33 -124.9 ;
      RECT 100.77 -112.315 101.1 -111.985 ;
      RECT 100.785 -145.42 101.085 -111.985 ;
      RECT 100.77 -86.37 101.1 -86.04 ;
      RECT 100.785 -101.34 101.085 -86.04 ;
      RECT 100.77 -101.34 101.1 -101.01 ;
      RECT 100.785 -82.145 101.085 -45.52 ;
      RECT 100.77 -45.895 101.1 -45.565 ;
      RECT 100.77 -82.145 101.1 -81.815 ;
      RECT 98.245 -117.705 98.575 -117.375 ;
      RECT 98.26 -138.15 98.56 -117.375 ;
      RECT 98.245 -124.945 98.575 -124.615 ;
      RECT 98.245 -138.105 98.575 -137.775 ;
      RECT 97.615 -124.145 97.945 -123.815 ;
      RECT 97.63 -145.42 97.93 -123.815 ;
      RECT 97.615 -85.91 97.945 -85.58 ;
      RECT 97.63 -101.34 97.93 -85.58 ;
      RECT 97.615 -101.34 97.945 -101.01 ;
      RECT 97.63 -82.125 97.93 -45.52 ;
      RECT 97.615 -47.495 97.945 -47.165 ;
      RECT 97.615 -81.715 97.945 -81.385 ;
      RECT 97 -118.505 97.33 -118.175 ;
      RECT 97.015 -145.42 97.315 -118.175 ;
      RECT 97.015 -117.22 97.315 -53.42 ;
      RECT 97 -53.795 97.33 -53.465 ;
      RECT 97 -69.495 97.33 -69.165 ;
      RECT 97 -117.22 97.33 -116.89 ;
      RECT 95.77 -112.315 96.1 -111.985 ;
      RECT 95.785 -145.42 96.085 -111.985 ;
      RECT 95.77 -86.37 96.1 -86.04 ;
      RECT 95.785 -101.34 96.085 -86.04 ;
      RECT 95.77 -101.34 96.1 -101.01 ;
      RECT 95.785 -82.145 96.085 -45.52 ;
      RECT 95.77 -45.895 96.1 -45.565 ;
      RECT 95.77 -82.145 96.1 -81.815 ;
      RECT 92.615 -85.91 92.945 -85.58 ;
      RECT 92.63 -101.34 92.93 -85.58 ;
      RECT 92.615 -101.34 92.945 -101.01 ;
      RECT 92.63 -82.125 92.93 -45.52 ;
      RECT 92.615 -47.495 92.945 -47.165 ;
      RECT 92.615 -81.715 92.945 -81.385 ;
      RECT 92.015 -125.23 92.315 -53.42 ;
      RECT 92 -53.795 92.33 -53.465 ;
      RECT 92 -69.495 92.33 -69.165 ;
      RECT 92 -125.23 92.33 -124.9 ;
      RECT 91.4 -134.07 91.7 -58.145 ;
      RECT 91.385 -58.52 91.715 -58.19 ;
      RECT 91.385 -134.07 91.715 -133.74 ;
      RECT 90.77 -112.315 91.1 -111.985 ;
      RECT 90.785 -145.42 91.085 -111.985 ;
      RECT 90.77 -86.37 91.1 -86.04 ;
      RECT 90.785 -101.34 91.085 -86.04 ;
      RECT 90.77 -101.34 91.1 -101.01 ;
      RECT 90.785 -82.145 91.085 -45.52 ;
      RECT 90.77 -45.895 91.1 -45.565 ;
      RECT 90.77 -82.145 91.1 -81.815 ;
      RECT 89.11 -134.445 89.44 -134.115 ;
      RECT 89.125 -145.42 89.425 -134.115 ;
      RECT 88.245 -117.705 88.575 -117.375 ;
      RECT 88.26 -138.15 88.56 -117.375 ;
      RECT 88.245 -124.945 88.575 -124.615 ;
      RECT 88.245 -133.645 88.575 -133.315 ;
      RECT 88.245 -138.105 88.575 -137.775 ;
      RECT 87.615 -124.145 87.945 -123.815 ;
      RECT 87.63 -145.42 87.93 -123.815 ;
      RECT 87.615 -85.91 87.945 -85.58 ;
      RECT 87.63 -101.34 87.93 -85.58 ;
      RECT 87.615 -101.34 87.945 -101.01 ;
      RECT 87.63 -82.125 87.93 -45.52 ;
      RECT 87.615 -47.495 87.945 -47.165 ;
      RECT 87.615 -81.715 87.945 -81.385 ;
      RECT 87 -118.505 87.33 -118.175 ;
      RECT 87.015 -145.42 87.315 -118.175 ;
      RECT 87.015 -117.22 87.315 -53.42 ;
      RECT 87 -53.795 87.33 -53.465 ;
      RECT 87 -69.495 87.33 -69.165 ;
      RECT 87 -117.22 87.33 -116.89 ;
      RECT 85.77 -112.315 86.1 -111.985 ;
      RECT 85.785 -145.42 86.085 -111.985 ;
      RECT 85.77 -86.37 86.1 -86.04 ;
      RECT 85.785 -101.34 86.085 -86.04 ;
      RECT 85.77 -101.34 86.1 -101.01 ;
      RECT 85.785 -82.145 86.085 -45.52 ;
      RECT 85.77 -45.895 86.1 -45.565 ;
      RECT 85.77 -82.145 86.1 -81.815 ;
      RECT 82.615 -85.91 82.945 -85.58 ;
      RECT 82.63 -101.34 82.93 -85.58 ;
      RECT 82.615 -101.34 82.945 -101.01 ;
      RECT 82.63 -82.125 82.93 -45.52 ;
      RECT 82.615 -47.495 82.945 -47.165 ;
      RECT 82.615 -81.715 82.945 -81.385 ;
      RECT 82.015 -125.23 82.315 -53.42 ;
      RECT 82 -53.795 82.33 -53.465 ;
      RECT 82 -69.495 82.33 -69.165 ;
      RECT 82 -125.23 82.33 -124.9 ;
      RECT 80.77 -112.315 81.1 -111.985 ;
      RECT 80.785 -145.42 81.085 -111.985 ;
      RECT 80.77 -86.37 81.1 -86.04 ;
      RECT 80.785 -101.34 81.085 -86.04 ;
      RECT 80.77 -101.34 81.1 -101.01 ;
      RECT 80.785 -82.145 81.085 -45.52 ;
      RECT 80.77 -45.895 81.1 -45.565 ;
      RECT 80.77 -82.145 81.1 -81.815 ;
      RECT 78.245 -117.705 78.575 -117.375 ;
      RECT 78.26 -138.15 78.56 -117.375 ;
      RECT 78.245 -124.945 78.575 -124.615 ;
      RECT 78.245 -138.105 78.575 -137.775 ;
      RECT 77.615 -124.145 77.945 -123.815 ;
      RECT 77.63 -145.42 77.93 -123.815 ;
      RECT 77.615 -85.91 77.945 -85.58 ;
      RECT 77.63 -101.34 77.93 -85.58 ;
      RECT 77.615 -101.34 77.945 -101.01 ;
      RECT 77.63 -82.125 77.93 -45.52 ;
      RECT 77.615 -47.495 77.945 -47.165 ;
      RECT 77.615 -81.715 77.945 -81.385 ;
      RECT 77 -118.505 77.33 -118.175 ;
      RECT 77.015 -145.42 77.315 -118.175 ;
      RECT 77.015 -117.22 77.315 -53.42 ;
      RECT 77 -53.795 77.33 -53.465 ;
      RECT 77 -69.495 77.33 -69.165 ;
      RECT 77 -117.22 77.33 -116.89 ;
      RECT 75.77 -112.315 76.1 -111.985 ;
      RECT 75.785 -145.42 76.085 -111.985 ;
      RECT 75.77 -86.37 76.1 -86.04 ;
      RECT 75.785 -101.34 76.085 -86.04 ;
      RECT 75.77 -101.34 76.1 -101.01 ;
      RECT 75.785 -82.145 76.085 -45.52 ;
      RECT 75.77 -45.895 76.1 -45.565 ;
      RECT 75.77 -82.145 76.1 -81.815 ;
      RECT 72.615 -85.91 72.945 -85.58 ;
      RECT 72.63 -101.34 72.93 -85.58 ;
      RECT 72.615 -101.34 72.945 -101.01 ;
      RECT 72.63 -82.125 72.93 -45.52 ;
      RECT 72.615 -47.495 72.945 -47.165 ;
      RECT 72.615 -81.715 72.945 -81.385 ;
      RECT 72.015 -125.23 72.315 -53.42 ;
      RECT 72 -53.795 72.33 -53.465 ;
      RECT 72 -69.495 72.33 -69.165 ;
      RECT 72 -125.23 72.33 -124.9 ;
      RECT 70.77 -112.315 71.1 -111.985 ;
      RECT 70.785 -145.42 71.085 -111.985 ;
      RECT 70.77 -86.37 71.1 -86.04 ;
      RECT 70.785 -101.34 71.085 -86.04 ;
      RECT 70.77 -101.34 71.1 -101.01 ;
      RECT 70.785 -82.145 71.085 -45.52 ;
      RECT 70.77 -45.895 71.1 -45.565 ;
      RECT 70.77 -82.145 71.1 -81.815 ;
      RECT 68.245 -117.705 68.575 -117.375 ;
      RECT 68.26 -138.15 68.56 -117.375 ;
      RECT 68.245 -124.945 68.575 -124.615 ;
      RECT 68.245 -138.105 68.575 -137.775 ;
      RECT 67.615 -124.145 67.945 -123.815 ;
      RECT 67.63 -145.42 67.93 -123.815 ;
      RECT 67.615 -85.91 67.945 -85.58 ;
      RECT 67.63 -101.34 67.93 -85.58 ;
      RECT 67.615 -101.34 67.945 -101.01 ;
      RECT 67.63 -82.125 67.93 -45.52 ;
      RECT 67.615 -47.495 67.945 -47.165 ;
      RECT 67.615 -81.715 67.945 -81.385 ;
      RECT 67 -118.505 67.33 -118.175 ;
      RECT 67.015 -145.42 67.315 -118.175 ;
      RECT 67.015 -117.22 67.315 -53.42 ;
      RECT 67 -53.795 67.33 -53.465 ;
      RECT 67 -69.495 67.33 -69.165 ;
      RECT 67 -117.22 67.33 -116.89 ;
      RECT 65.77 -112.315 66.1 -111.985 ;
      RECT 65.785 -145.42 66.085 -111.985 ;
      RECT 65.77 -86.37 66.1 -86.04 ;
      RECT 65.785 -101.34 66.085 -86.04 ;
      RECT 65.77 -101.34 66.1 -101.01 ;
      RECT 65.785 -82.145 66.085 -45.52 ;
      RECT 65.77 -45.895 66.1 -45.565 ;
      RECT 65.77 -82.145 66.1 -81.815 ;
      RECT 62.615 -85.91 62.945 -85.58 ;
      RECT 62.63 -101.34 62.93 -85.58 ;
      RECT 62.615 -101.34 62.945 -101.01 ;
      RECT 62.63 -82.125 62.93 -45.52 ;
      RECT 62.615 -47.495 62.945 -47.165 ;
      RECT 62.615 -81.715 62.945 -81.385 ;
      RECT 62.015 -125.23 62.315 -53.42 ;
      RECT 62 -53.795 62.33 -53.465 ;
      RECT 62 -69.495 62.33 -69.165 ;
      RECT 62 -125.23 62.33 -124.9 ;
      RECT 60.77 -112.315 61.1 -111.985 ;
      RECT 60.785 -145.42 61.085 -111.985 ;
      RECT 60.77 -86.37 61.1 -86.04 ;
      RECT 60.785 -101.34 61.085 -86.04 ;
      RECT 60.77 -101.34 61.1 -101.01 ;
      RECT 60.785 -82.145 61.085 -45.52 ;
      RECT 60.77 -45.895 61.1 -45.565 ;
      RECT 60.77 -82.145 61.1 -81.815 ;
      RECT 58.245 -117.705 58.575 -117.375 ;
      RECT 58.26 -138.15 58.56 -117.375 ;
      RECT 58.245 -124.945 58.575 -124.615 ;
      RECT 58.245 -138.105 58.575 -137.775 ;
      RECT 57.615 -124.145 57.945 -123.815 ;
      RECT 57.63 -145.42 57.93 -123.815 ;
      RECT 57.615 -85.91 57.945 -85.58 ;
      RECT 57.63 -101.34 57.93 -85.58 ;
      RECT 57.615 -101.34 57.945 -101.01 ;
      RECT 57.63 -82.125 57.93 -45.52 ;
      RECT 57.615 -47.495 57.945 -47.165 ;
      RECT 57.615 -81.715 57.945 -81.385 ;
      RECT 57 -118.505 57.33 -118.175 ;
      RECT 57.015 -145.42 57.315 -118.175 ;
      RECT 57.015 -117.22 57.315 -53.42 ;
      RECT 57 -53.795 57.33 -53.465 ;
      RECT 57 -69.495 57.33 -69.165 ;
      RECT 57 -117.22 57.33 -116.89 ;
      RECT 55.77 -112.315 56.1 -111.985 ;
      RECT 55.785 -145.42 56.085 -111.985 ;
      RECT 55.77 -86.37 56.1 -86.04 ;
      RECT 55.785 -101.34 56.085 -86.04 ;
      RECT 55.77 -101.34 56.1 -101.01 ;
      RECT 55.785 -82.145 56.085 -45.52 ;
      RECT 55.77 -45.895 56.1 -45.565 ;
      RECT 55.77 -82.145 56.1 -81.815 ;
      RECT 52.615 -85.91 52.945 -85.58 ;
      RECT 52.63 -101.34 52.93 -85.58 ;
      RECT 52.615 -101.34 52.945 -101.01 ;
      RECT 52.63 -82.125 52.93 -45.52 ;
      RECT 52.615 -47.495 52.945 -47.165 ;
      RECT 52.615 -81.715 52.945 -81.385 ;
      RECT 52.015 -125.23 52.315 -53.42 ;
      RECT 52 -53.795 52.33 -53.465 ;
      RECT 52 -69.495 52.33 -69.165 ;
      RECT 52 -125.23 52.33 -124.9 ;
      RECT 51.4 -134.07 51.7 -58.145 ;
      RECT 51.385 -58.52 51.715 -58.19 ;
      RECT 51.385 -134.07 51.715 -133.74 ;
      RECT 50.77 -112.315 51.1 -111.985 ;
      RECT 50.785 -145.42 51.085 -111.985 ;
      RECT 50.77 -86.37 51.1 -86.04 ;
      RECT 50.785 -101.34 51.085 -86.04 ;
      RECT 50.77 -101.34 51.1 -101.01 ;
      RECT 50.785 -82.145 51.085 -45.52 ;
      RECT 50.77 -45.895 51.1 -45.565 ;
      RECT 50.77 -82.145 51.1 -81.815 ;
      RECT 49.11 -134.445 49.44 -134.115 ;
      RECT 49.125 -145.42 49.425 -134.115 ;
      RECT 48.245 -117.705 48.575 -117.375 ;
      RECT 48.26 -138.15 48.56 -117.375 ;
      RECT 48.245 -124.945 48.575 -124.615 ;
      RECT 48.245 -133.645 48.575 -133.315 ;
      RECT 48.245 -138.105 48.575 -137.775 ;
      RECT 47.615 -124.145 47.945 -123.815 ;
      RECT 47.63 -145.42 47.93 -123.815 ;
      RECT 47.615 -85.91 47.945 -85.58 ;
      RECT 47.63 -101.34 47.93 -85.58 ;
      RECT 47.615 -101.34 47.945 -101.01 ;
      RECT 47.63 -82.125 47.93 -45.52 ;
      RECT 47.615 -47.495 47.945 -47.165 ;
      RECT 47.615 -81.715 47.945 -81.385 ;
      RECT 47 -118.505 47.33 -118.175 ;
      RECT 47.015 -145.42 47.315 -118.175 ;
      RECT 47.015 -117.22 47.315 -53.42 ;
      RECT 47 -53.795 47.33 -53.465 ;
      RECT 47 -69.495 47.33 -69.165 ;
      RECT 47 -117.22 47.33 -116.89 ;
      RECT 45.77 -112.315 46.1 -111.985 ;
      RECT 45.785 -145.42 46.085 -111.985 ;
      RECT 45.77 -86.37 46.1 -86.04 ;
      RECT 45.785 -101.34 46.085 -86.04 ;
      RECT 45.77 -101.34 46.1 -101.01 ;
      RECT 45.785 -82.145 46.085 -45.52 ;
      RECT 45.77 -45.895 46.1 -45.565 ;
      RECT 45.77 -82.145 46.1 -81.815 ;
      RECT 42.615 -85.91 42.945 -85.58 ;
      RECT 42.63 -101.34 42.93 -85.58 ;
      RECT 42.615 -101.34 42.945 -101.01 ;
      RECT 42.63 -82.125 42.93 -45.52 ;
      RECT 42.615 -47.495 42.945 -47.165 ;
      RECT 42.615 -81.715 42.945 -81.385 ;
      RECT 42.015 -125.23 42.315 -53.42 ;
      RECT 42 -53.795 42.33 -53.465 ;
      RECT 42 -69.495 42.33 -69.165 ;
      RECT 42 -125.23 42.33 -124.9 ;
      RECT 40.77 -112.315 41.1 -111.985 ;
      RECT 40.785 -145.42 41.085 -111.985 ;
      RECT 40.77 -86.37 41.1 -86.04 ;
      RECT 40.785 -101.34 41.085 -86.04 ;
      RECT 40.77 -101.34 41.1 -101.01 ;
      RECT 40.785 -82.145 41.085 -45.52 ;
      RECT 40.77 -45.895 41.1 -45.565 ;
      RECT 40.77 -82.145 41.1 -81.815 ;
      RECT 38.245 -117.705 38.575 -117.375 ;
      RECT 38.26 -138.15 38.56 -117.375 ;
      RECT 38.245 -124.945 38.575 -124.615 ;
      RECT 38.245 -138.105 38.575 -137.775 ;
      RECT 37.615 -124.145 37.945 -123.815 ;
      RECT 37.63 -145.42 37.93 -123.815 ;
      RECT 37.615 -85.91 37.945 -85.58 ;
      RECT 37.63 -101.34 37.93 -85.58 ;
      RECT 37.615 -101.34 37.945 -101.01 ;
      RECT 37.63 -82.125 37.93 -45.52 ;
      RECT 37.615 -47.495 37.945 -47.165 ;
      RECT 37.615 -81.715 37.945 -81.385 ;
      RECT 37 -118.505 37.33 -118.175 ;
      RECT 37.015 -145.42 37.315 -118.175 ;
      RECT 37.015 -117.22 37.315 -53.42 ;
      RECT 37 -53.795 37.33 -53.465 ;
      RECT 37 -69.495 37.33 -69.165 ;
      RECT 37 -117.22 37.33 -116.89 ;
      RECT 35.77 -112.315 36.1 -111.985 ;
      RECT 35.785 -145.42 36.085 -111.985 ;
      RECT 35.77 -86.37 36.1 -86.04 ;
      RECT 35.785 -101.34 36.085 -86.04 ;
      RECT 35.77 -101.34 36.1 -101.01 ;
      RECT 35.785 -82.145 36.085 -45.52 ;
      RECT 35.77 -45.895 36.1 -45.565 ;
      RECT 35.77 -82.145 36.1 -81.815 ;
      RECT 32.615 -85.91 32.945 -85.58 ;
      RECT 32.63 -101.34 32.93 -85.58 ;
      RECT 32.615 -101.34 32.945 -101.01 ;
      RECT 32.63 -82.125 32.93 -45.52 ;
      RECT 32.615 -47.495 32.945 -47.165 ;
      RECT 32.615 -81.715 32.945 -81.385 ;
      RECT 32.015 -125.23 32.315 -53.42 ;
      RECT 32 -53.795 32.33 -53.465 ;
      RECT 32 -69.495 32.33 -69.165 ;
      RECT 32 -125.23 32.33 -124.9 ;
      RECT 30.77 -112.315 31.1 -111.985 ;
      RECT 30.785 -145.42 31.085 -111.985 ;
      RECT 30.77 -86.37 31.1 -86.04 ;
      RECT 30.785 -101.34 31.085 -86.04 ;
      RECT 30.77 -101.34 31.1 -101.01 ;
      RECT 30.785 -82.145 31.085 -45.52 ;
      RECT 30.77 -45.895 31.1 -45.565 ;
      RECT 30.77 -82.145 31.1 -81.815 ;
      RECT 28.245 -117.705 28.575 -117.375 ;
      RECT 28.26 -138.15 28.56 -117.375 ;
      RECT 28.245 -124.945 28.575 -124.615 ;
      RECT 28.245 -138.105 28.575 -137.775 ;
      RECT 27.615 -124.145 27.945 -123.815 ;
      RECT 27.63 -145.42 27.93 -123.815 ;
      RECT 27.615 -85.91 27.945 -85.58 ;
      RECT 27.63 -101.34 27.93 -85.58 ;
      RECT 27.615 -101.34 27.945 -101.01 ;
      RECT 27.63 -82.125 27.93 -45.52 ;
      RECT 27.615 -47.495 27.945 -47.165 ;
      RECT 27.615 -81.715 27.945 -81.385 ;
      RECT 27 -118.505 27.33 -118.175 ;
      RECT 27.015 -145.42 27.315 -118.175 ;
      RECT 27.015 -117.22 27.315 -53.42 ;
      RECT 27 -53.795 27.33 -53.465 ;
      RECT 27 -69.495 27.33 -69.165 ;
      RECT 27 -117.22 27.33 -116.89 ;
      RECT 25.77 -112.315 26.1 -111.985 ;
      RECT 25.785 -145.42 26.085 -111.985 ;
      RECT 25.77 -86.37 26.1 -86.04 ;
      RECT 25.785 -101.34 26.085 -86.04 ;
      RECT 25.77 -101.34 26.1 -101.01 ;
      RECT 25.785 -82.145 26.085 -45.52 ;
      RECT 25.77 -45.895 26.1 -45.565 ;
      RECT 25.77 -82.145 26.1 -81.815 ;
      RECT 22.615 -85.91 22.945 -85.58 ;
      RECT 22.63 -101.34 22.93 -85.58 ;
      RECT 22.615 -101.34 22.945 -101.01 ;
      RECT 22.63 -82.125 22.93 -45.52 ;
      RECT 22.615 -47.495 22.945 -47.165 ;
      RECT 22.615 -81.715 22.945 -81.385 ;
      RECT 22.015 -125.23 22.315 -53.42 ;
      RECT 22 -53.795 22.33 -53.465 ;
      RECT 22 -69.495 22.33 -69.165 ;
      RECT 22 -125.23 22.33 -124.9 ;
      RECT 20.77 -112.315 21.1 -111.985 ;
      RECT 20.785 -145.42 21.085 -111.985 ;
      RECT 20.77 -86.37 21.1 -86.04 ;
      RECT 20.785 -101.34 21.085 -86.04 ;
      RECT 20.77 -101.34 21.1 -101.01 ;
      RECT 20.785 -82.145 21.085 -45.52 ;
      RECT 20.77 -45.895 21.1 -45.565 ;
      RECT 20.77 -82.145 21.1 -81.815 ;
      RECT 18.245 -117.705 18.575 -117.375 ;
      RECT 18.26 -138.15 18.56 -117.375 ;
      RECT 18.245 -124.945 18.575 -124.615 ;
      RECT 18.245 -138.105 18.575 -137.775 ;
      RECT 17.615 -124.145 17.945 -123.815 ;
      RECT 17.63 -145.42 17.93 -123.815 ;
      RECT 17.615 -85.91 17.945 -85.58 ;
      RECT 17.63 -101.34 17.93 -85.58 ;
      RECT 17.615 -101.34 17.945 -101.01 ;
      RECT 17.63 -82.125 17.93 -45.52 ;
      RECT 17.615 -47.495 17.945 -47.165 ;
      RECT 17.615 -81.715 17.945 -81.385 ;
      RECT 17 -118.505 17.33 -118.175 ;
      RECT 17.015 -145.42 17.315 -118.175 ;
      RECT 17.015 -117.22 17.315 -53.42 ;
      RECT 17 -53.795 17.33 -53.465 ;
      RECT 17 -69.495 17.33 -69.165 ;
      RECT 17 -117.22 17.33 -116.89 ;
      RECT 15.77 -112.315 16.1 -111.985 ;
      RECT 15.785 -145.42 16.085 -111.985 ;
      RECT 15.77 -86.37 16.1 -86.04 ;
      RECT 15.785 -101.34 16.085 -86.04 ;
      RECT 15.77 -101.34 16.1 -101.01 ;
      RECT 15.785 -82.145 16.085 -45.52 ;
      RECT 15.77 -45.895 16.1 -45.565 ;
      RECT 15.77 -82.145 16.1 -81.815 ;
      RECT 12.615 -85.91 12.945 -85.58 ;
      RECT 12.63 -101.34 12.93 -85.58 ;
      RECT 12.615 -101.34 12.945 -101.01 ;
      RECT 12.63 -82.125 12.93 -45.52 ;
      RECT 12.615 -47.495 12.945 -47.165 ;
      RECT 12.615 -81.715 12.945 -81.385 ;
      RECT 12.015 -125.23 12.315 -53.42 ;
      RECT 12 -53.795 12.33 -53.465 ;
      RECT 12 -69.495 12.33 -69.165 ;
      RECT 12 -125.23 12.33 -124.9 ;
      RECT 11.4 -134.07 11.7 -58.145 ;
      RECT 11.385 -58.52 11.715 -58.19 ;
      RECT 11.385 -134.07 11.715 -133.74 ;
      RECT 10.77 -112.315 11.1 -111.985 ;
      RECT 10.785 -145.42 11.085 -111.985 ;
      RECT 10.77 -86.37 11.1 -86.04 ;
      RECT 10.785 -101.34 11.085 -86.04 ;
      RECT 10.77 -101.34 11.1 -101.01 ;
      RECT 10.785 -82.145 11.085 -45.52 ;
      RECT 10.77 -45.895 11.1 -45.565 ;
      RECT 10.77 -82.145 11.1 -81.815 ;
      RECT 9.11 -134.445 9.44 -134.115 ;
      RECT 9.125 -145.42 9.425 -134.115 ;
      RECT 8.245 -117.705 8.575 -117.375 ;
      RECT 8.26 -138.15 8.56 -117.375 ;
      RECT 8.245 -124.945 8.575 -124.615 ;
      RECT 8.245 -133.645 8.575 -133.315 ;
      RECT 8.245 -138.105 8.575 -137.775 ;
      RECT 7.615 -124.145 7.945 -123.815 ;
      RECT 7.63 -145.42 7.93 -123.815 ;
      RECT 7.615 -85.91 7.945 -85.58 ;
      RECT 7.63 -101.34 7.93 -85.58 ;
      RECT 7.615 -101.34 7.945 -101.01 ;
      RECT 7.63 -82.125 7.93 -45.52 ;
      RECT 7.615 -47.495 7.945 -47.165 ;
      RECT 7.615 -81.715 7.945 -81.385 ;
      RECT 7 -118.505 7.33 -118.175 ;
      RECT 7.015 -145.42 7.315 -118.175 ;
      RECT 7.015 -117.22 7.315 -53.42 ;
      RECT 7 -53.795 7.33 -53.465 ;
      RECT 7 -69.495 7.33 -69.165 ;
      RECT 7 -117.22 7.33 -116.89 ;
      RECT 5.77 -112.315 6.1 -111.985 ;
      RECT 5.785 -145.42 6.085 -111.985 ;
      RECT 5.77 -86.37 6.1 -86.04 ;
      RECT 5.785 -101.34 6.085 -86.04 ;
      RECT 5.77 -101.34 6.1 -101.01 ;
      RECT 5.785 -82.145 6.085 -45.52 ;
      RECT 5.77 -45.895 6.1 -45.565 ;
      RECT 5.77 -82.145 6.1 -81.815 ;
      RECT 3.505 -76.13 3.835 -75.8 ;
      RECT 3.52 -77.605 3.82 -75.8 ;
      RECT 3.505 -77.605 3.835 -77.275 ;
      RECT -5.91 -98.04 -5.58 -97.71 ;
      RECT -5.895 -111.475 -5.595 -97.71 ;
      RECT -5.91 -111.475 -5.58 -111.145 ;
      RECT -9.505 -111.03 -9.175 -110.7 ;
      RECT -9.49 -138.15 -9.19 -110.7 ;
      RECT -9.505 -138.105 -9.175 -137.775 ;
      RECT -10.635 -111.83 -10.305 -111.5 ;
      RECT -10.62 -145.42 -10.32 -111.5 ;
      RECT -11.75 -102.805 -11.42 -102.475 ;
      RECT -11.735 -111.475 -11.435 -102.475 ;
      RECT -11.75 -111.475 -11.42 -111.145 ;
      RECT -12.385 -102.305 -12.055 -101.975 ;
      RECT -12.37 -112.23 -12.07 -101.975 ;
      RECT -12.385 -112.23 -12.055 -111.9 ;
      RECT -15.345 -111.03 -15.015 -110.7 ;
      RECT -15.33 -138.15 -15.03 -110.7 ;
      RECT -15.345 -138.105 -15.015 -137.775 ;
      RECT -16.475 -111.83 -16.145 -111.5 ;
      RECT -16.46 -145.42 -16.16 -111.5 ;
      RECT -17 -36.06 -16.67 -35.73 ;
      RECT -16.985 -79.395 -16.685 -35.73 ;
      RECT -17 -79.395 -16.67 -79.065 ;
      RECT -17.59 -103.805 -17.26 -103.475 ;
      RECT -17.575 -111.475 -17.275 -103.475 ;
      RECT -17.59 -111.475 -17.26 -111.145 ;
      RECT -18.225 -103.305 -17.895 -102.975 ;
      RECT -18.21 -112.23 -17.91 -102.975 ;
      RECT -18.225 -112.23 -17.895 -111.9 ;
      RECT -21.185 -111.03 -20.855 -110.7 ;
      RECT -21.17 -138.15 -20.87 -110.7 ;
      RECT -21.185 -138.105 -20.855 -137.775 ;
      RECT -22.315 -111.83 -21.985 -111.5 ;
      RECT -22.3 -145.42 -22 -111.5 ;
      RECT -23.43 -104.805 -23.1 -104.475 ;
      RECT -23.415 -111.475 -23.115 -104.475 ;
      RECT -23.43 -111.475 -23.1 -111.145 ;
      RECT -24.065 -104.305 -23.735 -103.975 ;
      RECT -24.05 -112.23 -23.75 -103.975 ;
      RECT -24.065 -112.23 -23.735 -111.9 ;
      RECT -27.025 -111.03 -26.695 -110.7 ;
      RECT -27.01 -138.15 -26.71 -110.7 ;
      RECT -27.025 -138.105 -26.695 -137.775 ;
      RECT -28.155 -111.83 -27.825 -111.5 ;
      RECT -28.14 -145.42 -27.84 -111.5 ;
      RECT -29.27 -105.805 -28.94 -105.475 ;
      RECT -29.255 -111.475 -28.955 -105.475 ;
      RECT -29.27 -111.475 -28.94 -111.145 ;
      RECT -29.905 -105.305 -29.575 -104.975 ;
      RECT -29.89 -112.23 -29.59 -104.975 ;
      RECT -29.905 -112.23 -29.575 -111.9 ;
      RECT -32.865 -111.03 -32.535 -110.7 ;
      RECT -32.85 -138.15 -32.55 -110.7 ;
      RECT -32.865 -138.105 -32.535 -137.775 ;
      RECT -33.995 -111.83 -33.665 -111.5 ;
      RECT -33.98 -145.42 -33.68 -111.5 ;
      RECT -35.11 -106.805 -34.78 -106.475 ;
      RECT -35.095 -111.475 -34.795 -106.475 ;
      RECT -35.11 -111.475 -34.78 -111.145 ;
      RECT -35.745 -106.305 -35.415 -105.975 ;
      RECT -35.73 -112.23 -35.43 -105.975 ;
      RECT -35.745 -112.23 -35.415 -111.9 ;
      RECT -38.705 -111.03 -38.375 -110.7 ;
      RECT -38.69 -138.15 -38.39 -110.7 ;
      RECT -38.705 -138.105 -38.375 -137.775 ;
      RECT -39.835 -111.83 -39.505 -111.5 ;
      RECT -39.82 -145.42 -39.52 -111.5 ;
      RECT -40.7 -138.15 -40.3 -99.35 ;
      RECT -40.84 -145.3 -40.42 -137.73 ;
  END
END sramgen_sram_32x32m2w8_replica_v1

END LIBRARY
