VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_2048x64m8w8
    CLASS BLOCK  ;
    FOREIGN sram22_2048x64m8w8   ;
    SIZE 1126.000 BY 796.200 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 417.630 0.000 417.770 0.140 ;
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 428.530 0.000 428.670 0.140 ;
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 439.430 0.000 439.570 0.140 ;
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 450.330 0.000 450.470 0.140 ;
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 461.230 0.000 461.370 0.140 ;
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 472.130 0.000 472.270 0.140 ;
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 483.030 0.000 483.170 0.140 ;
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 493.930 0.000 494.070 0.140 ;
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 504.830 0.000 504.970 0.140 ;
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 515.730 0.000 515.870 0.140 ;
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 526.630 0.000 526.770 0.140 ;
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 537.530 0.000 537.670 0.140 ;
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 548.430 0.000 548.570 0.140 ;
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 559.330 0.000 559.470 0.140 ;
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 570.230 0.000 570.370 0.140 ;
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 581.130 0.000 581.270 0.140 ;
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 592.030 0.000 592.170 0.140 ;
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 602.930 0.000 603.070 0.140 ;
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 613.830 0.000 613.970 0.140 ;
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 624.730 0.000 624.870 0.140 ;
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 635.630 0.000 635.770 0.140 ;
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 646.530 0.000 646.670 0.140 ;
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 657.430 0.000 657.570 0.140 ;
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 668.330 0.000 668.470 0.140 ;
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 679.230 0.000 679.370 0.140 ;
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 690.130 0.000 690.270 0.140 ;
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 701.030 0.000 701.170 0.140 ;
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 711.930 0.000 712.070 0.140 ;
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 722.830 0.000 722.970 0.140 ;
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 733.730 0.000 733.870 0.140 ;
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 744.630 0.000 744.770 0.140 ;
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 755.530 0.000 755.670 0.140 ;
        END 
    END dout[31] 
    PIN dout[32] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 766.430 0.000 766.570 0.140 ;
        END 
    END dout[32] 
    PIN dout[33] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 777.330 0.000 777.470 0.140 ;
        END 
    END dout[33] 
    PIN dout[34] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 788.230 0.000 788.370 0.140 ;
        END 
    END dout[34] 
    PIN dout[35] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 799.130 0.000 799.270 0.140 ;
        END 
    END dout[35] 
    PIN dout[36] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 810.030 0.000 810.170 0.140 ;
        END 
    END dout[36] 
    PIN dout[37] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 820.930 0.000 821.070 0.140 ;
        END 
    END dout[37] 
    PIN dout[38] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 831.830 0.000 831.970 0.140 ;
        END 
    END dout[38] 
    PIN dout[39] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 842.730 0.000 842.870 0.140 ;
        END 
    END dout[39] 
    PIN dout[40] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 853.630 0.000 853.770 0.140 ;
        END 
    END dout[40] 
    PIN dout[41] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 864.530 0.000 864.670 0.140 ;
        END 
    END dout[41] 
    PIN dout[42] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 875.430 0.000 875.570 0.140 ;
        END 
    END dout[42] 
    PIN dout[43] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 886.330 0.000 886.470 0.140 ;
        END 
    END dout[43] 
    PIN dout[44] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 897.230 0.000 897.370 0.140 ;
        END 
    END dout[44] 
    PIN dout[45] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 908.130 0.000 908.270 0.140 ;
        END 
    END dout[45] 
    PIN dout[46] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 919.030 0.000 919.170 0.140 ;
        END 
    END dout[46] 
    PIN dout[47] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 929.930 0.000 930.070 0.140 ;
        END 
    END dout[47] 
    PIN dout[48] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 940.830 0.000 940.970 0.140 ;
        END 
    END dout[48] 
    PIN dout[49] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 951.730 0.000 951.870 0.140 ;
        END 
    END dout[49] 
    PIN dout[50] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 962.630 0.000 962.770 0.140 ;
        END 
    END dout[50] 
    PIN dout[51] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 973.530 0.000 973.670 0.140 ;
        END 
    END dout[51] 
    PIN dout[52] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 984.430 0.000 984.570 0.140 ;
        END 
    END dout[52] 
    PIN dout[53] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 995.330 0.000 995.470 0.140 ;
        END 
    END dout[53] 
    PIN dout[54] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1006.230 0.000 1006.370 0.140 ;
        END 
    END dout[54] 
    PIN dout[55] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1017.130 0.000 1017.270 0.140 ;
        END 
    END dout[55] 
    PIN dout[56] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1028.030 0.000 1028.170 0.140 ;
        END 
    END dout[56] 
    PIN dout[57] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1038.930 0.000 1039.070 0.140 ;
        END 
    END dout[57] 
    PIN dout[58] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1049.830 0.000 1049.970 0.140 ;
        END 
    END dout[58] 
    PIN dout[59] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1060.730 0.000 1060.870 0.140 ;
        END 
    END dout[59] 
    PIN dout[60] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1071.630 0.000 1071.770 0.140 ;
        END 
    END dout[60] 
    PIN dout[61] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1082.530 0.000 1082.670 0.140 ;
        END 
    END dout[61] 
    PIN dout[62] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1093.430 0.000 1093.570 0.140 ;
        END 
    END dout[62] 
    PIN dout[63] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 10.096200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1104.330 0.000 1104.470 0.140 ;
        END 
    END dout[63] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 417.210 0.000 417.350 0.140 ;
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 428.110 0.000 428.250 0.140 ;
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 439.010 0.000 439.150 0.140 ;
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 449.910 0.000 450.050 0.140 ;
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 460.810 0.000 460.950 0.140 ;
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 471.710 0.000 471.850 0.140 ;
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 482.610 0.000 482.750 0.140 ;
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 493.510 0.000 493.650 0.140 ;
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 504.410 0.000 504.550 0.140 ;
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 515.310 0.000 515.450 0.140 ;
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 526.210 0.000 526.350 0.140 ;
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 537.110 0.000 537.250 0.140 ;
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 548.010 0.000 548.150 0.140 ;
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 558.910 0.000 559.050 0.140 ;
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 569.810 0.000 569.950 0.140 ;
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 580.710 0.000 580.850 0.140 ;
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 591.610 0.000 591.750 0.140 ;
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 602.510 0.000 602.650 0.140 ;
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 613.410 0.000 613.550 0.140 ;
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 624.310 0.000 624.450 0.140 ;
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 635.210 0.000 635.350 0.140 ;
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 646.110 0.000 646.250 0.140 ;
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 657.010 0.000 657.150 0.140 ;
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 667.910 0.000 668.050 0.140 ;
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 678.810 0.000 678.950 0.140 ;
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 689.710 0.000 689.850 0.140 ;
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 700.610 0.000 700.750 0.140 ;
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 711.510 0.000 711.650 0.140 ;
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 722.410 0.000 722.550 0.140 ;
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 733.310 0.000 733.450 0.140 ;
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 744.210 0.000 744.350 0.140 ;
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 755.110 0.000 755.250 0.140 ;
        END 
    END din[31] 
    PIN din[32] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 766.010 0.000 766.150 0.140 ;
        END 
    END din[32] 
    PIN din[33] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 776.910 0.000 777.050 0.140 ;
        END 
    END din[33] 
    PIN din[34] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 787.810 0.000 787.950 0.140 ;
        END 
    END din[34] 
    PIN din[35] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 798.710 0.000 798.850 0.140 ;
        END 
    END din[35] 
    PIN din[36] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 809.610 0.000 809.750 0.140 ;
        END 
    END din[36] 
    PIN din[37] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 820.510 0.000 820.650 0.140 ;
        END 
    END din[37] 
    PIN din[38] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 831.410 0.000 831.550 0.140 ;
        END 
    END din[38] 
    PIN din[39] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 842.310 0.000 842.450 0.140 ;
        END 
    END din[39] 
    PIN din[40] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 853.210 0.000 853.350 0.140 ;
        END 
    END din[40] 
    PIN din[41] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 864.110 0.000 864.250 0.140 ;
        END 
    END din[41] 
    PIN din[42] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 875.010 0.000 875.150 0.140 ;
        END 
    END din[42] 
    PIN din[43] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 885.910 0.000 886.050 0.140 ;
        END 
    END din[43] 
    PIN din[44] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 896.810 0.000 896.950 0.140 ;
        END 
    END din[44] 
    PIN din[45] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 907.710 0.000 907.850 0.140 ;
        END 
    END din[45] 
    PIN din[46] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 918.610 0.000 918.750 0.140 ;
        END 
    END din[46] 
    PIN din[47] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 929.510 0.000 929.650 0.140 ;
        END 
    END din[47] 
    PIN din[48] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 940.410 0.000 940.550 0.140 ;
        END 
    END din[48] 
    PIN din[49] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 951.310 0.000 951.450 0.140 ;
        END 
    END din[49] 
    PIN din[50] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 962.210 0.000 962.350 0.140 ;
        END 
    END din[50] 
    PIN din[51] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 973.110 0.000 973.250 0.140 ;
        END 
    END din[51] 
    PIN din[52] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 984.010 0.000 984.150 0.140 ;
        END 
    END din[52] 
    PIN din[53] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 994.910 0.000 995.050 0.140 ;
        END 
    END din[53] 
    PIN din[54] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1005.810 0.000 1005.950 0.140 ;
        END 
    END din[54] 
    PIN din[55] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1016.710 0.000 1016.850 0.140 ;
        END 
    END din[55] 
    PIN din[56] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1027.610 0.000 1027.750 0.140 ;
        END 
    END din[56] 
    PIN din[57] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1038.510 0.000 1038.650 0.140 ;
        END 
    END din[57] 
    PIN din[58] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1049.410 0.000 1049.550 0.140 ;
        END 
    END din[58] 
    PIN din[59] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1060.310 0.000 1060.450 0.140 ;
        END 
    END din[59] 
    PIN din[60] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1071.210 0.000 1071.350 0.140 ;
        END 
    END din[60] 
    PIN din[61] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1082.110 0.000 1082.250 0.140 ;
        END 
    END din[61] 
    PIN din[62] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1093.010 0.000 1093.150 0.140 ;
        END 
    END din[62] 
    PIN din[63] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.196200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.817800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1103.910 0.000 1104.050 0.140 ;
        END 
    END din[63] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.006600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 416.860 0.000 417.000 0.140 ;
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.006600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 504.060 0.000 504.200 0.140 ;
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.006600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 591.260 0.000 591.400 0.140 ;
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.006600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 678.460 0.000 678.600 0.140 ;
        END 
    END wmask[3] 
    PIN wmask[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.006600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 765.660 0.000 765.800 0.140 ;
        END 
    END wmask[4] 
    PIN wmask[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.006600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 852.860 0.000 853.000 0.140 ;
        END 
    END wmask[5] 
    PIN wmask[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.006600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 940.060 0.000 940.200 0.140 ;
        END 
    END wmask[6] 
    PIN wmask[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.006600 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1027.260 0.000 1027.400 0.140 ;
        END 
    END wmask[7] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 335.040 0.000 335.360 0.320 ;
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 328.920 0.000 329.240 0.320 ;
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 322.800 0.000 323.120 0.320 ;
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 316.680 0.000 317.000 0.320 ;
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 310.560 0.000 310.880 0.320 ;
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 304.440 0.000 304.760 0.320 ;
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 298.320 0.000 298.640 0.320 ;
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 292.200 0.000 292.520 0.320 ;
        END 
    END addr[7] 
    PIN addr[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 286.760 0.000 287.080 0.320 ;
        END 
    END addr[8] 
    PIN addr[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 280.640 0.000 280.960 0.320 ;
        END 
    END addr[9] 
    PIN addr[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 274.520 0.000 274.840 0.320 ;
        END 
    END addr[10] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 347.280 0.000 347.600 0.320 ;
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.835900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 341.160 0.000 341.480 0.320 ;
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 42.129000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 350.680 0.000 351.000 0.320 ;
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 46.035000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 351.360 0.000 351.680 0.320 ;
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 416.960 6.240 ;
                RECT 418.680 5.920 427.840 6.240 ;
                RECT 429.560 5.920 438.720 6.240 ;
                RECT 440.440 5.920 449.600 6.240 ;
                RECT 451.320 5.920 460.480 6.240 ;
                RECT 462.200 5.920 471.360 6.240 ;
                RECT 473.080 5.920 482.240 6.240 ;
                RECT 483.960 5.920 493.120 6.240 ;
                RECT 494.840 5.920 504.000 6.240 ;
                RECT 505.720 5.920 514.880 6.240 ;
                RECT 516.600 5.920 525.760 6.240 ;
                RECT 527.480 5.920 536.640 6.240 ;
                RECT 538.360 5.920 547.520 6.240 ;
                RECT 549.240 5.920 558.400 6.240 ;
                RECT 560.120 5.920 569.280 6.240 ;
                RECT 571.000 5.920 580.160 6.240 ;
                RECT 581.880 5.920 591.040 6.240 ;
                RECT 592.760 5.920 601.920 6.240 ;
                RECT 603.640 5.920 612.800 6.240 ;
                RECT 614.520 5.920 624.360 6.240 ;
                RECT 625.400 5.920 635.240 6.240 ;
                RECT 636.280 5.920 646.120 6.240 ;
                RECT 647.160 5.920 657.000 6.240 ;
                RECT 658.040 5.920 667.880 6.240 ;
                RECT 668.920 5.920 678.760 6.240 ;
                RECT 679.800 5.920 689.640 6.240 ;
                RECT 690.680 5.920 700.520 6.240 ;
                RECT 701.560 5.920 711.400 6.240 ;
                RECT 712.440 5.920 722.280 6.240 ;
                RECT 724.000 5.920 733.160 6.240 ;
                RECT 734.880 5.920 744.040 6.240 ;
                RECT 745.760 5.920 754.920 6.240 ;
                RECT 756.640 5.920 765.800 6.240 ;
                RECT 767.520 5.920 776.680 6.240 ;
                RECT 778.400 5.920 787.560 6.240 ;
                RECT 789.280 5.920 798.440 6.240 ;
                RECT 800.160 5.920 809.320 6.240 ;
                RECT 811.040 5.920 820.200 6.240 ;
                RECT 821.920 5.920 831.080 6.240 ;
                RECT 832.800 5.920 841.960 6.240 ;
                RECT 843.680 5.920 852.840 6.240 ;
                RECT 854.560 5.920 863.720 6.240 ;
                RECT 865.440 5.920 874.600 6.240 ;
                RECT 876.320 5.920 885.480 6.240 ;
                RECT 887.200 5.920 896.360 6.240 ;
                RECT 898.080 5.920 907.240 6.240 ;
                RECT 908.960 5.920 918.120 6.240 ;
                RECT 919.840 5.920 929.000 6.240 ;
                RECT 930.720 5.920 939.880 6.240 ;
                RECT 941.600 5.920 950.760 6.240 ;
                RECT 952.480 5.920 961.640 6.240 ;
                RECT 963.360 5.920 972.520 6.240 ;
                RECT 974.240 5.920 983.400 6.240 ;
                RECT 985.120 5.920 994.960 6.240 ;
                RECT 996.000 5.920 1005.840 6.240 ;
                RECT 1006.880 5.920 1016.720 6.240 ;
                RECT 1017.760 5.920 1027.600 6.240 ;
                RECT 1028.640 5.920 1038.480 6.240 ;
                RECT 1039.520 5.920 1049.360 6.240 ;
                RECT 1050.400 5.920 1060.240 6.240 ;
                RECT 1061.280 5.920 1071.120 6.240 ;
                RECT 1072.160 5.920 1082.000 6.240 ;
                RECT 1083.040 5.920 1092.880 6.240 ;
                RECT 1094.600 5.920 1103.760 6.240 ;
                RECT 1105.480 5.920 1125.840 6.240 ;
                RECT 0.160 7.280 1125.840 7.600 ;
                RECT 0.160 8.640 1125.840 8.960 ;
                RECT 0.160 10.000 350.320 10.320 ;
                RECT 410.520 10.000 1125.840 10.320 ;
                RECT 0.160 11.360 1125.840 11.680 ;
                RECT 0.160 12.720 404.040 13.040 ;
                RECT 1116.360 12.720 1125.840 13.040 ;
                RECT 0.160 14.080 270.080 14.400 ;
                RECT 352.040 14.080 404.040 14.400 ;
                RECT 1116.360 14.080 1125.840 14.400 ;
                RECT 0.160 15.440 404.040 15.760 ;
                RECT 1116.360 15.440 1125.840 15.760 ;
                RECT 0.160 16.800 404.040 17.120 ;
                RECT 1116.360 16.800 1125.840 17.120 ;
                RECT 0.160 18.160 270.080 18.480 ;
                RECT 351.360 18.160 404.040 18.480 ;
                RECT 1116.360 18.160 1125.840 18.480 ;
                RECT 0.160 19.520 404.040 19.840 ;
                RECT 1116.360 19.520 1125.840 19.840 ;
                RECT 0.160 20.880 404.040 21.200 ;
                RECT 1116.360 20.880 1125.840 21.200 ;
                RECT 0.160 22.240 404.040 22.560 ;
                RECT 1116.360 22.240 1125.840 22.560 ;
                RECT 0.160 23.600 404.040 23.920 ;
                RECT 1116.360 23.600 1125.840 23.920 ;
                RECT 0.160 24.960 404.040 25.280 ;
                RECT 1116.360 24.960 1125.840 25.280 ;
                RECT 0.160 26.320 404.040 26.640 ;
                RECT 1116.360 26.320 1125.840 26.640 ;
                RECT 0.160 27.680 404.040 28.000 ;
                RECT 1116.360 27.680 1125.840 28.000 ;
                RECT 0.160 29.040 404.040 29.360 ;
                RECT 1116.360 29.040 1125.840 29.360 ;
                RECT 0.160 30.400 403.360 30.720 ;
                RECT 1116.360 30.400 1125.840 30.720 ;
                RECT 0.160 31.760 404.040 32.080 ;
                RECT 1116.360 31.760 1125.840 32.080 ;
                RECT 0.160 33.120 404.040 33.440 ;
                RECT 1116.360 33.120 1125.840 33.440 ;
                RECT 0.160 34.480 404.040 34.800 ;
                RECT 1116.360 34.480 1125.840 34.800 ;
                RECT 0.160 35.840 404.040 36.160 ;
                RECT 1116.360 35.840 1125.840 36.160 ;
                RECT 0.160 37.200 113.000 37.520 ;
                RECT 322.800 37.200 404.040 37.520 ;
                RECT 1116.360 37.200 1125.840 37.520 ;
                RECT 0.160 38.560 111.640 38.880 ;
                RECT 328.920 38.560 404.040 38.880 ;
                RECT 1116.360 38.560 1125.840 38.880 ;
                RECT 0.160 39.920 110.280 40.240 ;
                RECT 335.040 39.920 404.040 40.240 ;
                RECT 1116.360 39.920 1125.840 40.240 ;
                RECT 0.160 41.280 90.560 41.600 ;
                RECT 352.040 41.280 404.040 41.600 ;
                RECT 1116.360 41.280 1125.840 41.600 ;
                RECT 0.160 42.640 89.880 42.960 ;
                RECT 347.960 42.640 404.040 42.960 ;
                RECT 1116.360 42.640 1125.840 42.960 ;
                RECT 0.160 44.000 404.040 44.320 ;
                RECT 1116.360 44.000 1125.840 44.320 ;
                RECT 0.160 45.360 344.200 45.680 ;
                RECT 350.000 45.360 404.040 45.680 ;
                RECT 1116.360 45.360 1125.840 45.680 ;
                RECT 0.160 46.720 344.200 47.040 ;
                RECT 350.000 46.720 404.040 47.040 ;
                RECT 1116.360 46.720 1125.840 47.040 ;
                RECT 0.160 48.080 344.200 48.400 ;
                RECT 1116.360 48.080 1125.840 48.400 ;
                RECT 0.160 49.440 344.200 49.760 ;
                RECT 1116.360 49.440 1125.840 49.760 ;
                RECT 0.160 50.800 108.920 51.120 ;
                RECT 341.160 50.800 344.200 51.120 ;
                RECT 350.000 50.800 404.040 51.120 ;
                RECT 1116.360 50.800 1125.840 51.120 ;
                RECT 0.160 52.160 404.040 52.480 ;
                RECT 1116.360 52.160 1125.840 52.480 ;
                RECT 0.160 53.520 404.040 53.840 ;
                RECT 1116.360 53.520 1125.840 53.840 ;
                RECT 0.160 54.880 404.040 55.200 ;
                RECT 1116.360 54.880 1125.840 55.200 ;
                RECT 0.160 56.240 404.040 56.560 ;
                RECT 1116.360 56.240 1125.840 56.560 ;
                RECT 0.160 57.600 110.280 57.920 ;
                RECT 118.800 57.600 125.240 57.920 ;
                RECT 348.640 57.600 404.040 57.920 ;
                RECT 1116.360 57.600 1125.840 57.920 ;
                RECT 0.160 58.960 111.640 59.280 ;
                RECT 117.440 58.960 125.240 59.280 ;
                RECT 365.640 58.960 404.040 59.280 ;
                RECT 1116.360 58.960 1125.840 59.280 ;
                RECT 0.160 60.320 113.000 60.640 ;
                RECT 116.760 60.320 125.240 60.640 ;
                RECT 365.640 60.320 404.040 60.640 ;
                RECT 1116.360 60.320 1125.840 60.640 ;
                RECT 0.160 61.680 125.240 62.000 ;
                RECT 362.920 61.680 404.040 62.000 ;
                RECT 1116.360 61.680 1125.840 62.000 ;
                RECT 0.160 63.040 125.240 63.360 ;
                RECT 365.640 63.040 404.040 63.360 ;
                RECT 1116.360 63.040 1125.840 63.360 ;
                RECT 0.160 64.400 125.240 64.720 ;
                RECT 365.640 64.400 404.040 64.720 ;
                RECT 1116.360 64.400 1125.840 64.720 ;
                RECT 0.160 65.760 125.240 66.080 ;
                RECT 362.920 65.760 404.040 66.080 ;
                RECT 1116.360 65.760 1125.840 66.080 ;
                RECT 0.160 67.120 125.240 67.440 ;
                RECT 371.080 67.120 404.040 67.440 ;
                RECT 1116.360 67.120 1125.840 67.440 ;
                RECT 0.160 68.480 125.240 68.800 ;
                RECT 368.360 68.480 404.040 68.800 ;
                RECT 1116.360 68.480 1125.840 68.800 ;
                RECT 0.160 69.840 125.240 70.160 ;
                RECT 371.080 69.840 404.040 70.160 ;
                RECT 1116.360 69.840 1125.840 70.160 ;
                RECT 0.160 71.200 125.240 71.520 ;
                RECT 371.080 71.200 404.040 71.520 ;
                RECT 1116.360 71.200 1125.840 71.520 ;
                RECT 0.160 72.560 125.240 72.880 ;
                RECT 368.360 72.560 404.040 72.880 ;
                RECT 1116.360 72.560 1125.840 72.880 ;
                RECT 0.160 73.920 125.240 74.240 ;
                RECT 371.080 73.920 404.040 74.240 ;
                RECT 1116.360 73.920 1125.840 74.240 ;
                RECT 0.160 75.280 125.240 75.600 ;
                RECT 348.640 75.280 404.040 75.600 ;
                RECT 1116.360 75.280 1125.840 75.600 ;
                RECT 0.160 76.640 125.240 76.960 ;
                RECT 376.520 76.640 404.040 76.960 ;
                RECT 1116.360 76.640 1125.840 76.960 ;
                RECT 0.160 78.000 125.240 78.320 ;
                RECT 376.520 78.000 404.040 78.320 ;
                RECT 1116.360 78.000 1125.840 78.320 ;
                RECT 0.160 79.360 125.240 79.680 ;
                RECT 348.640 79.360 404.040 79.680 ;
                RECT 1116.360 79.360 1125.840 79.680 ;
                RECT 0.160 80.720 125.240 81.040 ;
                RECT 373.800 80.720 404.040 81.040 ;
                RECT 1116.360 80.720 1125.840 81.040 ;
                RECT 0.160 82.080 125.240 82.400 ;
                RECT 376.520 82.080 404.040 82.400 ;
                RECT 1116.360 82.080 1125.840 82.400 ;
                RECT 0.160 83.440 125.240 83.760 ;
                RECT 348.640 83.440 404.040 83.760 ;
                RECT 1116.360 83.440 1125.840 83.760 ;
                RECT 0.160 84.800 125.240 85.120 ;
                RECT 381.960 84.800 404.040 85.120 ;
                RECT 1116.360 84.800 1125.840 85.120 ;
                RECT 0.160 86.160 125.240 86.480 ;
                RECT 381.960 86.160 404.040 86.480 ;
                RECT 1116.360 86.160 1125.840 86.480 ;
                RECT 0.160 87.520 125.240 87.840 ;
                RECT 379.240 87.520 404.040 87.840 ;
                RECT 1116.360 87.520 1125.840 87.840 ;
                RECT 0.160 88.880 125.240 89.200 ;
                RECT 381.960 88.880 404.040 89.200 ;
                RECT 1116.360 88.880 1125.840 89.200 ;
                RECT 0.160 90.240 125.240 90.560 ;
                RECT 381.960 90.240 404.040 90.560 ;
                RECT 1116.360 90.240 1125.840 90.560 ;
                RECT 0.160 91.600 125.240 91.920 ;
                RECT 379.240 91.600 404.040 91.920 ;
                RECT 1116.360 91.600 1125.840 91.920 ;
                RECT 0.160 92.960 125.240 93.280 ;
                RECT 387.400 92.960 404.040 93.280 ;
                RECT 1116.360 92.960 1125.840 93.280 ;
                RECT 0.160 94.320 125.240 94.640 ;
                RECT 384.680 94.320 404.040 94.640 ;
                RECT 1116.360 94.320 1125.840 94.640 ;
                RECT 0.160 95.680 125.240 96.000 ;
                RECT 387.400 95.680 404.040 96.000 ;
                RECT 1116.360 95.680 1125.840 96.000 ;
                RECT 0.160 97.040 125.240 97.360 ;
                RECT 387.400 97.040 404.040 97.360 ;
                RECT 1116.360 97.040 1125.840 97.360 ;
                RECT 0.160 98.400 125.240 98.720 ;
                RECT 348.640 98.400 404.040 98.720 ;
                RECT 1116.360 98.400 1125.840 98.720 ;
                RECT 0.160 99.760 125.240 100.080 ;
                RECT 384.680 99.760 404.040 100.080 ;
                RECT 1116.360 99.760 1125.840 100.080 ;
                RECT 0.160 101.120 125.240 101.440 ;
                RECT 348.640 101.120 404.040 101.440 ;
                RECT 1116.360 101.120 1125.840 101.440 ;
                RECT 0.160 102.480 125.240 102.800 ;
                RECT 392.840 102.480 404.040 102.800 ;
                RECT 1116.360 102.480 1125.840 102.800 ;
                RECT 0.160 103.840 125.240 104.160 ;
                RECT 392.840 103.840 404.040 104.160 ;
                RECT 1116.360 103.840 1125.840 104.160 ;
                RECT 0.160 105.200 125.240 105.520 ;
                RECT 392.840 105.200 404.040 105.520 ;
                RECT 1116.360 105.200 1125.840 105.520 ;
                RECT 0.160 106.560 125.240 106.880 ;
                RECT 390.120 106.560 404.040 106.880 ;
                RECT 1116.360 106.560 1125.840 106.880 ;
                RECT 0.160 107.920 125.240 108.240 ;
                RECT 392.840 107.920 404.040 108.240 ;
                RECT 1116.360 107.920 1125.840 108.240 ;
                RECT 0.160 109.280 125.240 109.600 ;
                RECT 348.640 109.280 404.040 109.600 ;
                RECT 1116.360 109.280 1125.840 109.600 ;
                RECT 0.160 110.640 125.240 110.960 ;
                RECT 398.280 110.640 404.040 110.960 ;
                RECT 1116.360 110.640 1125.840 110.960 ;
                RECT 0.160 112.000 125.240 112.320 ;
                RECT 398.280 112.000 404.040 112.320 ;
                RECT 1116.360 112.000 1125.840 112.320 ;
                RECT 0.160 113.360 125.240 113.680 ;
                RECT 395.560 113.360 404.040 113.680 ;
                RECT 1116.360 113.360 1125.840 113.680 ;
                RECT 0.160 114.720 125.240 115.040 ;
                RECT 398.280 114.720 404.040 115.040 ;
                RECT 1116.360 114.720 1125.840 115.040 ;
                RECT 0.160 116.080 125.240 116.400 ;
                RECT 398.280 116.080 404.040 116.400 ;
                RECT 1116.360 116.080 1125.840 116.400 ;
                RECT 0.160 117.440 125.240 117.760 ;
                RECT 395.560 117.440 404.040 117.760 ;
                RECT 1116.360 117.440 1125.840 117.760 ;
                RECT 0.160 118.800 125.240 119.120 ;
                RECT 1116.360 118.800 1125.840 119.120 ;
                RECT 0.160 120.160 125.240 120.480 ;
                RECT 1116.360 120.160 1125.840 120.480 ;
                RECT 0.160 121.520 125.240 121.840 ;
                RECT 1116.360 121.520 1125.840 121.840 ;
                RECT 0.160 122.880 125.240 123.200 ;
                RECT 1116.360 122.880 1125.840 123.200 ;
                RECT 0.160 124.240 125.240 124.560 ;
                RECT 348.640 124.240 404.040 124.560 ;
                RECT 1116.360 124.240 1125.840 124.560 ;
                RECT 0.160 125.600 125.240 125.920 ;
                RECT 1116.360 125.600 1125.840 125.920 ;
                RECT 0.160 126.960 125.240 127.280 ;
                RECT 348.640 126.960 404.040 127.280 ;
                RECT 1116.360 126.960 1125.840 127.280 ;
                RECT 0.160 128.320 404.040 128.640 ;
                RECT 1116.360 128.320 1125.840 128.640 ;
                RECT 0.160 129.680 357.120 130.000 ;
                RECT 1116.360 129.680 1125.840 130.000 ;
                RECT 0.160 131.040 397.920 131.360 ;
                RECT 1116.360 131.040 1125.840 131.360 ;
                RECT 0.160 132.400 397.920 132.720 ;
                RECT 1116.360 132.400 1125.840 132.720 ;
                RECT 0.160 133.760 392.480 134.080 ;
                RECT 1116.360 133.760 1125.840 134.080 ;
                RECT 0.160 135.120 392.480 135.440 ;
                RECT 1116.360 135.120 1125.840 135.440 ;
                RECT 0.160 136.480 392.480 136.800 ;
                RECT 1116.360 136.480 1125.840 136.800 ;
                RECT 0.160 137.840 387.040 138.160 ;
                RECT 1116.360 137.840 1125.840 138.160 ;
                RECT 0.160 139.200 387.040 139.520 ;
                RECT 1116.360 139.200 1125.840 139.520 ;
                RECT 0.160 140.560 381.600 140.880 ;
                RECT 1116.360 140.560 1125.840 140.880 ;
                RECT 0.160 141.920 381.600 142.240 ;
                RECT 1116.360 141.920 1125.840 142.240 ;
                RECT 0.160 143.280 376.160 143.600 ;
                RECT 1116.360 143.280 1125.840 143.600 ;
                RECT 0.160 144.640 376.160 144.960 ;
                RECT 1116.360 144.640 1125.840 144.960 ;
                RECT 0.160 146.000 370.720 146.320 ;
                RECT 1116.360 146.000 1125.840 146.320 ;
                RECT 0.160 147.360 370.720 147.680 ;
                RECT 1116.360 147.360 1125.840 147.680 ;
                RECT 0.160 148.720 86.480 149.040 ;
                RECT 97.040 148.720 365.280 149.040 ;
                RECT 1116.360 148.720 1125.840 149.040 ;
                RECT 0.160 150.080 87.840 150.400 ;
                RECT 93.640 150.080 100.760 150.400 ;
                RECT 103.840 150.080 365.280 150.400 ;
                RECT 1116.360 150.080 1125.840 150.400 ;
                RECT 0.160 151.440 89.200 151.760 ;
                RECT 92.280 151.440 359.840 151.760 ;
                RECT 1116.360 151.440 1125.840 151.760 ;
                RECT 0.160 152.800 95.320 153.120 ;
                RECT 102.480 152.800 359.840 153.120 ;
                RECT 1116.360 152.800 1125.840 153.120 ;
                RECT 0.160 154.160 90.560 154.480 ;
                RECT 103.840 154.160 359.840 154.480 ;
                RECT 1116.360 154.160 1125.840 154.480 ;
                RECT 0.160 155.520 87.840 155.840 ;
                RECT 97.040 155.520 404.040 155.840 ;
                RECT 1116.360 155.520 1125.840 155.840 ;
                RECT 0.160 156.880 404.040 157.200 ;
                RECT 1116.360 156.880 1125.840 157.200 ;
                RECT 0.160 158.240 87.840 158.560 ;
                RECT 90.240 158.240 404.040 158.560 ;
                RECT 1116.360 158.240 1125.840 158.560 ;
                RECT 0.160 159.600 87.840 159.920 ;
                RECT 103.160 159.600 404.040 159.920 ;
                RECT 1116.360 159.600 1125.840 159.920 ;
                RECT 0.160 160.960 94.640 161.280 ;
                RECT 97.040 160.960 404.040 161.280 ;
                RECT 1116.360 160.960 1125.840 161.280 ;
                RECT 0.160 162.320 404.040 162.640 ;
                RECT 1116.360 162.320 1125.840 162.640 ;
                RECT 0.160 163.680 95.320 164.000 ;
                RECT 103.840 163.680 404.040 164.000 ;
                RECT 1116.360 163.680 1125.840 164.000 ;
                RECT 0.160 165.040 92.600 165.360 ;
                RECT 97.040 165.040 404.040 165.360 ;
                RECT 1116.360 165.040 1125.840 165.360 ;
                RECT 0.160 166.400 94.640 166.720 ;
                RECT 97.040 166.400 404.040 166.720 ;
                RECT 1116.360 166.400 1125.840 166.720 ;
                RECT 0.160 167.760 404.040 168.080 ;
                RECT 1116.360 167.760 1125.840 168.080 ;
                RECT 0.160 169.120 85.800 169.440 ;
                RECT 108.600 169.120 404.040 169.440 ;
                RECT 1116.360 169.120 1125.840 169.440 ;
                RECT 0.160 170.480 102.800 170.800 ;
                RECT 109.960 170.480 404.040 170.800 ;
                RECT 1116.360 170.480 1125.840 170.800 ;
                RECT 0.160 171.840 94.640 172.160 ;
                RECT 97.040 171.840 106.880 172.160 ;
                RECT 110.640 171.840 404.040 172.160 ;
                RECT 1116.360 171.840 1125.840 172.160 ;
                RECT 0.160 173.200 86.480 173.520 ;
                RECT 99.760 173.200 404.040 173.520 ;
                RECT 1116.360 173.200 1125.840 173.520 ;
                RECT 0.160 174.560 95.320 174.880 ;
                RECT 103.840 174.560 404.040 174.880 ;
                RECT 1116.360 174.560 1125.840 174.880 ;
                RECT 0.160 175.920 92.600 176.240 ;
                RECT 97.040 175.920 404.040 176.240 ;
                RECT 1116.360 175.920 1125.840 176.240 ;
                RECT 0.160 177.280 64.720 177.600 ;
                RECT 82.760 177.280 95.320 177.600 ;
                RECT 103.840 177.280 404.040 177.600 ;
                RECT 1116.360 177.280 1125.840 177.600 ;
                RECT 0.160 178.640 64.720 178.960 ;
                RECT 82.760 178.640 404.040 178.960 ;
                RECT 1116.360 178.640 1125.840 178.960 ;
                RECT 0.160 180.000 64.720 180.320 ;
                RECT 82.760 180.000 88.520 180.320 ;
                RECT 90.920 180.000 404.040 180.320 ;
                RECT 1116.360 180.000 1125.840 180.320 ;
                RECT 0.160 181.360 64.720 181.680 ;
                RECT 82.760 181.360 92.600 181.680 ;
                RECT 97.040 181.360 404.040 181.680 ;
                RECT 1116.360 181.360 1125.840 181.680 ;
                RECT 0.160 182.720 64.720 183.040 ;
                RECT 82.760 182.720 404.040 183.040 ;
                RECT 1116.360 182.720 1125.840 183.040 ;
                RECT 0.160 184.080 64.720 184.400 ;
                RECT 82.760 184.080 94.640 184.400 ;
                RECT 97.040 184.080 404.040 184.400 ;
                RECT 1116.360 184.080 1125.840 184.400 ;
                RECT 0.160 185.440 64.720 185.760 ;
                RECT 82.760 185.440 95.320 185.760 ;
                RECT 97.720 185.440 404.040 185.760 ;
                RECT 1116.360 185.440 1125.840 185.760 ;
                RECT 0.160 186.800 64.720 187.120 ;
                RECT 82.760 186.800 404.040 187.120 ;
                RECT 1116.360 186.800 1125.840 187.120 ;
                RECT 0.160 188.160 64.720 188.480 ;
                RECT 82.760 188.160 94.640 188.480 ;
                RECT 97.040 188.160 404.040 188.480 ;
                RECT 1116.360 188.160 1125.840 188.480 ;
                RECT 0.160 189.520 64.720 189.840 ;
                RECT 82.760 189.520 85.120 189.840 ;
                RECT 97.040 189.520 404.040 189.840 ;
                RECT 1116.360 189.520 1125.840 189.840 ;
                RECT 0.160 190.880 64.720 191.200 ;
                RECT 82.760 190.880 95.320 191.200 ;
                RECT 97.720 190.880 404.040 191.200 ;
                RECT 1116.360 190.880 1125.840 191.200 ;
                RECT 0.160 192.240 64.720 192.560 ;
                RECT 82.760 192.240 404.040 192.560 ;
                RECT 1116.360 192.240 1125.840 192.560 ;
                RECT 0.160 193.600 64.720 193.920 ;
                RECT 82.760 193.600 404.040 193.920 ;
                RECT 1116.360 193.600 1125.840 193.920 ;
                RECT 0.160 194.960 64.720 195.280 ;
                RECT 96.360 194.960 404.040 195.280 ;
                RECT 1116.360 194.960 1125.840 195.280 ;
                RECT 0.160 196.320 64.720 196.640 ;
                RECT 82.760 196.320 92.600 196.640 ;
                RECT 99.760 196.320 404.040 196.640 ;
                RECT 1116.360 196.320 1125.840 196.640 ;
                RECT 0.160 197.680 64.720 198.000 ;
                RECT 82.760 197.680 274.160 198.000 ;
                RECT 347.960 197.680 404.040 198.000 ;
                RECT 1116.360 197.680 1125.840 198.000 ;
                RECT 0.160 199.040 64.720 199.360 ;
                RECT 82.760 199.040 87.840 199.360 ;
                RECT 92.280 199.040 274.160 199.360 ;
                RECT 347.960 199.040 404.040 199.360 ;
                RECT 1116.360 199.040 1125.840 199.360 ;
                RECT 0.160 200.400 64.720 200.720 ;
                RECT 82.760 200.400 87.840 200.720 ;
                RECT 104.520 200.400 274.160 200.720 ;
                RECT 347.960 200.400 404.040 200.720 ;
                RECT 1116.360 200.400 1125.840 200.720 ;
                RECT 0.160 201.760 64.720 202.080 ;
                RECT 82.760 201.760 274.160 202.080 ;
                RECT 347.960 201.760 404.040 202.080 ;
                RECT 1116.360 201.760 1125.840 202.080 ;
                RECT 0.160 203.120 64.720 203.440 ;
                RECT 82.760 203.120 91.920 203.440 ;
                RECT 103.840 203.120 274.160 203.440 ;
                RECT 347.960 203.120 362.560 203.440 ;
                RECT 1116.360 203.120 1125.840 203.440 ;
                RECT 0.160 204.480 64.720 204.800 ;
                RECT 82.760 204.480 89.200 204.800 ;
                RECT 103.840 204.480 362.560 204.800 ;
                RECT 1116.360 204.480 1125.840 204.800 ;
                RECT 0.160 205.840 64.720 206.160 ;
                RECT 82.760 205.840 85.800 206.160 ;
                RECT 89.560 205.840 368.000 206.160 ;
                RECT 1116.360 205.840 1125.840 206.160 ;
                RECT 0.160 207.200 64.720 207.520 ;
                RECT 82.760 207.200 368.000 207.520 ;
                RECT 1116.360 207.200 1125.840 207.520 ;
                RECT 0.160 208.560 64.720 208.880 ;
                RECT 82.760 208.560 219.080 208.880 ;
                RECT 349.320 208.560 368.000 208.880 ;
                RECT 1116.360 208.560 1125.840 208.880 ;
                RECT 0.160 209.920 64.720 210.240 ;
                RECT 82.760 209.920 86.480 210.240 ;
                RECT 93.640 209.920 219.080 210.240 ;
                RECT 349.320 209.920 373.440 210.240 ;
                RECT 1116.360 209.920 1125.840 210.240 ;
                RECT 0.160 211.280 64.720 211.600 ;
                RECT 82.760 211.280 219.080 211.600 ;
                RECT 349.320 211.280 373.440 211.600 ;
                RECT 1116.360 211.280 1125.840 211.600 ;
                RECT 0.160 212.640 64.720 212.960 ;
                RECT 82.760 212.640 91.920 212.960 ;
                RECT 96.360 212.640 219.080 212.960 ;
                RECT 349.320 212.640 378.880 212.960 ;
                RECT 1116.360 212.640 1125.840 212.960 ;
                RECT 0.160 214.000 64.720 214.320 ;
                RECT 83.440 214.000 219.080 214.320 ;
                RECT 349.320 214.000 378.880 214.320 ;
                RECT 1116.360 214.000 1125.840 214.320 ;
                RECT 0.160 215.360 64.720 215.680 ;
                RECT 82.760 215.360 87.840 215.680 ;
                RECT 103.840 215.360 219.080 215.680 ;
                RECT 349.320 215.360 384.320 215.680 ;
                RECT 1116.360 215.360 1125.840 215.680 ;
                RECT 0.160 216.720 64.720 217.040 ;
                RECT 82.760 216.720 219.080 217.040 ;
                RECT 349.320 216.720 384.320 217.040 ;
                RECT 1116.360 216.720 1125.840 217.040 ;
                RECT 0.160 218.080 64.720 218.400 ;
                RECT 82.760 218.080 219.080 218.400 ;
                RECT 349.320 218.080 389.760 218.400 ;
                RECT 1116.360 218.080 1125.840 218.400 ;
                RECT 0.160 219.440 64.720 219.760 ;
                RECT 82.760 219.440 219.080 219.760 ;
                RECT 349.320 219.440 389.760 219.760 ;
                RECT 1116.360 219.440 1125.840 219.760 ;
                RECT 0.160 220.800 64.720 221.120 ;
                RECT 82.760 220.800 219.080 221.120 ;
                RECT 349.320 220.800 395.200 221.120 ;
                RECT 1116.360 220.800 1125.840 221.120 ;
                RECT 0.160 222.160 64.720 222.480 ;
                RECT 82.760 222.160 89.200 222.480 ;
                RECT 90.920 222.160 219.080 222.480 ;
                RECT 349.320 222.160 395.200 222.480 ;
                RECT 1116.360 222.160 1125.840 222.480 ;
                RECT 0.160 223.520 64.720 223.840 ;
                RECT 82.760 223.520 219.080 223.840 ;
                RECT 349.320 223.520 400.640 223.840 ;
                RECT 1116.360 223.520 1125.840 223.840 ;
                RECT 0.160 224.880 64.720 225.200 ;
                RECT 82.760 224.880 101.440 225.200 ;
                RECT 103.840 224.880 219.080 225.200 ;
                RECT 349.320 224.880 400.640 225.200 ;
                RECT 1116.360 224.880 1125.840 225.200 ;
                RECT 0.160 226.240 64.720 226.560 ;
                RECT 82.760 226.240 219.080 226.560 ;
                RECT 349.320 226.240 400.640 226.560 ;
                RECT 1116.360 226.240 1125.840 226.560 ;
                RECT 0.160 227.600 64.720 227.920 ;
                RECT 82.760 227.600 219.080 227.920 ;
                RECT 1116.360 227.600 1125.840 227.920 ;
                RECT 0.160 228.960 64.720 229.280 ;
                RECT 82.760 228.960 219.080 229.280 ;
                RECT 1116.360 228.960 1125.840 229.280 ;
                RECT 0.160 230.320 64.720 230.640 ;
                RECT 82.760 230.320 219.080 230.640 ;
                RECT 1116.360 230.320 1125.840 230.640 ;
                RECT 0.160 231.680 64.720 232.000 ;
                RECT 82.760 231.680 219.080 232.000 ;
                RECT 1116.360 231.680 1125.840 232.000 ;
                RECT 0.160 233.040 64.720 233.360 ;
                RECT 82.760 233.040 94.640 233.360 ;
                RECT 103.160 233.040 219.080 233.360 ;
                RECT 1116.360 233.040 1125.840 233.360 ;
                RECT 0.160 234.400 64.720 234.720 ;
                RECT 82.760 234.400 219.080 234.720 ;
                RECT 349.320 234.400 404.040 234.720 ;
                RECT 1116.360 234.400 1125.840 234.720 ;
                RECT 0.160 235.760 64.720 236.080 ;
                RECT 82.760 235.760 219.080 236.080 ;
                RECT 349.320 235.760 404.040 236.080 ;
                RECT 1116.360 235.760 1125.840 236.080 ;
                RECT 0.160 237.120 64.720 237.440 ;
                RECT 82.760 237.120 219.080 237.440 ;
                RECT 349.320 237.120 404.040 237.440 ;
                RECT 1116.360 237.120 1125.840 237.440 ;
                RECT 0.160 238.480 64.720 238.800 ;
                RECT 82.760 238.480 219.080 238.800 ;
                RECT 349.320 238.480 404.040 238.800 ;
                RECT 1116.360 238.480 1125.840 238.800 ;
                RECT 0.160 239.840 64.720 240.160 ;
                RECT 82.760 239.840 219.080 240.160 ;
                RECT 349.320 239.840 404.040 240.160 ;
                RECT 1116.360 239.840 1125.840 240.160 ;
                RECT 0.160 241.200 64.720 241.520 ;
                RECT 82.760 241.200 219.080 241.520 ;
                RECT 349.320 241.200 404.040 241.520 ;
                RECT 1116.360 241.200 1125.840 241.520 ;
                RECT 0.160 242.560 64.720 242.880 ;
                RECT 82.760 242.560 219.080 242.880 ;
                RECT 349.320 242.560 404.040 242.880 ;
                RECT 1116.360 242.560 1125.840 242.880 ;
                RECT 0.160 243.920 64.720 244.240 ;
                RECT 82.760 243.920 219.080 244.240 ;
                RECT 349.320 243.920 404.040 244.240 ;
                RECT 1116.360 243.920 1125.840 244.240 ;
                RECT 0.160 245.280 64.720 245.600 ;
                RECT 82.760 245.280 90.560 245.600 ;
                RECT 93.640 245.280 219.080 245.600 ;
                RECT 349.320 245.280 404.040 245.600 ;
                RECT 1116.360 245.280 1125.840 245.600 ;
                RECT 0.160 246.640 64.720 246.960 ;
                RECT 82.760 246.640 219.080 246.960 ;
                RECT 349.320 246.640 404.040 246.960 ;
                RECT 1116.360 246.640 1125.840 246.960 ;
                RECT 0.160 248.000 64.720 248.320 ;
                RECT 82.760 248.000 219.080 248.320 ;
                RECT 349.320 248.000 404.040 248.320 ;
                RECT 1116.360 248.000 1125.840 248.320 ;
                RECT 0.160 249.360 64.720 249.680 ;
                RECT 82.760 249.360 219.080 249.680 ;
                RECT 349.320 249.360 404.040 249.680 ;
                RECT 1116.360 249.360 1125.840 249.680 ;
                RECT 0.160 250.720 64.720 251.040 ;
                RECT 82.760 250.720 219.080 251.040 ;
                RECT 349.320 250.720 404.040 251.040 ;
                RECT 1116.360 250.720 1125.840 251.040 ;
                RECT 0.160 252.080 64.720 252.400 ;
                RECT 82.760 252.080 219.080 252.400 ;
                RECT 349.320 252.080 404.040 252.400 ;
                RECT 1116.360 252.080 1125.840 252.400 ;
                RECT 0.160 253.440 219.080 253.760 ;
                RECT 349.320 253.440 404.040 253.760 ;
                RECT 1116.360 253.440 1125.840 253.760 ;
                RECT 0.160 254.800 219.080 255.120 ;
                RECT 349.320 254.800 404.040 255.120 ;
                RECT 1116.360 254.800 1125.840 255.120 ;
                RECT 0.160 256.160 43.640 256.480 ;
                RECT 64.400 256.160 87.840 256.480 ;
                RECT 93.640 256.160 219.080 256.480 ;
                RECT 349.320 256.160 404.040 256.480 ;
                RECT 1116.360 256.160 1125.840 256.480 ;
                RECT 0.160 257.520 43.640 257.840 ;
                RECT 64.400 257.520 219.080 257.840 ;
                RECT 349.320 257.520 404.040 257.840 ;
                RECT 1116.360 257.520 1125.840 257.840 ;
                RECT 0.160 258.880 43.640 259.200 ;
                RECT 64.400 258.880 219.080 259.200 ;
                RECT 349.320 258.880 404.040 259.200 ;
                RECT 1116.360 258.880 1125.840 259.200 ;
                RECT 0.160 260.240 43.640 260.560 ;
                RECT 64.400 260.240 70.840 260.560 ;
                RECT 78.000 260.240 91.920 260.560 ;
                RECT 97.720 260.240 219.080 260.560 ;
                RECT 1116.360 260.240 1125.840 260.560 ;
                RECT 0.160 261.600 43.640 261.920 ;
                RECT 64.400 261.600 65.400 261.920 ;
                RECT 82.760 261.600 219.080 261.920 ;
                RECT 1116.360 261.600 1125.840 261.920 ;
                RECT 0.160 262.960 43.640 263.280 ;
                RECT 64.400 262.960 65.400 263.280 ;
                RECT 82.760 262.960 219.080 263.280 ;
                RECT 1116.360 262.960 1125.840 263.280 ;
                RECT 0.160 264.320 43.640 264.640 ;
                RECT 64.400 264.320 219.080 264.640 ;
                RECT 1116.360 264.320 1125.840 264.640 ;
                RECT 0.160 265.680 43.640 266.000 ;
                RECT 64.400 265.680 70.840 266.000 ;
                RECT 78.000 265.680 85.120 266.000 ;
                RECT 96.360 265.680 219.080 266.000 ;
                RECT 1116.360 265.680 1125.840 266.000 ;
                RECT 0.160 267.040 21.880 267.360 ;
                RECT 77.320 267.040 219.080 267.360 ;
                RECT 349.320 267.040 1125.840 267.360 ;
                RECT 0.160 268.400 76.960 268.720 ;
                RECT 216.720 268.400 1125.840 268.720 ;
                RECT 0.160 269.760 401.320 270.080 ;
                RECT 1118.400 269.760 1125.840 270.080 ;
                RECT 0.160 271.120 401.320 271.440 ;
                RECT 1118.400 271.120 1125.840 271.440 ;
                RECT 0.160 272.480 401.320 272.800 ;
                RECT 1118.400 272.480 1125.840 272.800 ;
                RECT 0.160 273.840 125.920 274.160 ;
                RECT 132.400 273.840 134.080 274.160 ;
                RECT 148.720 273.840 202.760 274.160 ;
                RECT 1118.400 273.840 1125.840 274.160 ;
                RECT 0.160 275.200 123.880 275.520 ;
                RECT 147.360 275.200 159.920 275.520 ;
                RECT 161.640 275.200 174.880 275.520 ;
                RECT 192.240 275.200 202.760 275.520 ;
                RECT 1118.400 275.200 1125.840 275.520 ;
                RECT 0.160 276.560 123.880 276.880 ;
                RECT 134.440 276.560 159.920 276.880 ;
                RECT 163.680 276.560 174.880 276.880 ;
                RECT 192.240 276.560 202.760 276.880 ;
                RECT 1118.400 276.560 1125.840 276.880 ;
                RECT 0.160 277.920 123.880 278.240 ;
                RECT 134.440 277.920 159.920 278.240 ;
                RECT 164.360 277.920 174.880 278.240 ;
                RECT 192.240 277.920 202.760 278.240 ;
                RECT 1118.400 277.920 1125.840 278.240 ;
                RECT 0.160 279.280 123.880 279.600 ;
                RECT 134.440 279.280 159.920 279.600 ;
                RECT 165.040 279.280 174.880 279.600 ;
                RECT 192.240 279.280 202.760 279.600 ;
                RECT 1118.400 279.280 1125.840 279.600 ;
                RECT 0.160 280.640 123.880 280.960 ;
                RECT 134.440 280.640 159.920 280.960 ;
                RECT 161.640 280.640 174.880 280.960 ;
                RECT 192.240 280.640 202.760 280.960 ;
                RECT 1118.400 280.640 1125.840 280.960 ;
                RECT 0.160 282.000 123.880 282.320 ;
                RECT 134.440 282.000 202.760 282.320 ;
                RECT 1118.400 282.000 1125.840 282.320 ;
                RECT 0.160 283.360 123.880 283.680 ;
                RECT 134.440 283.360 174.880 283.680 ;
                RECT 192.240 283.360 202.760 283.680 ;
                RECT 1118.400 283.360 1125.840 283.680 ;
                RECT 0.160 284.720 174.880 285.040 ;
                RECT 192.240 284.720 202.760 285.040 ;
                RECT 1118.400 284.720 1125.840 285.040 ;
                RECT 0.160 286.080 174.880 286.400 ;
                RECT 192.240 286.080 202.760 286.400 ;
                RECT 1118.400 286.080 1125.840 286.400 ;
                RECT 0.160 287.440 21.200 287.760 ;
                RECT 119.480 287.440 174.880 287.760 ;
                RECT 192.240 287.440 202.760 287.760 ;
                RECT 1118.400 287.440 1125.840 287.760 ;
                RECT 0.160 288.800 174.880 289.120 ;
                RECT 192.240 288.800 202.760 289.120 ;
                RECT 1118.400 288.800 1125.840 289.120 ;
                RECT 0.160 290.160 20.520 290.480 ;
                RECT 119.480 290.160 132.720 290.480 ;
                RECT 148.040 290.160 202.760 290.480 ;
                RECT 1118.400 290.160 1125.840 290.480 ;
                RECT 0.160 291.520 19.840 291.840 ;
                RECT 119.480 291.520 132.720 291.840 ;
                RECT 147.360 291.520 159.920 291.840 ;
                RECT 161.640 291.520 174.880 291.840 ;
                RECT 192.240 291.520 202.760 291.840 ;
                RECT 1118.400 291.520 1125.840 291.840 ;
                RECT 0.160 292.880 19.160 293.200 ;
                RECT 119.480 292.880 132.720 293.200 ;
                RECT 137.160 292.880 159.920 293.200 ;
                RECT 162.320 292.880 174.880 293.200 ;
                RECT 192.240 292.880 202.760 293.200 ;
                RECT 1118.400 292.880 1125.840 293.200 ;
                RECT 0.160 294.240 159.920 294.560 ;
                RECT 162.320 294.240 174.880 294.560 ;
                RECT 192.240 294.240 202.760 294.560 ;
                RECT 1118.400 294.240 1125.840 294.560 ;
                RECT 0.160 295.600 18.480 295.920 ;
                RECT 119.480 295.600 132.720 295.920 ;
                RECT 137.840 295.600 159.920 295.920 ;
                RECT 163.000 295.600 174.880 295.920 ;
                RECT 192.240 295.600 202.760 295.920 ;
                RECT 1118.400 295.600 1125.840 295.920 ;
                RECT 0.160 296.960 17.800 297.280 ;
                RECT 119.480 296.960 132.720 297.280 ;
                RECT 138.520 296.960 159.920 297.280 ;
                RECT 163.680 296.960 174.880 297.280 ;
                RECT 192.240 296.960 202.760 297.280 ;
                RECT 1118.400 296.960 1125.840 297.280 ;
                RECT 0.160 298.320 17.120 298.640 ;
                RECT 119.480 298.320 202.760 298.640 ;
                RECT 1118.400 298.320 1125.840 298.640 ;
                RECT 0.160 299.680 16.440 300.000 ;
                RECT 119.480 299.680 174.880 300.000 ;
                RECT 192.240 299.680 202.760 300.000 ;
                RECT 1118.400 299.680 1125.840 300.000 ;
                RECT 0.160 301.040 174.880 301.360 ;
                RECT 192.240 301.040 202.760 301.360 ;
                RECT 1118.400 301.040 1125.840 301.360 ;
                RECT 0.160 302.400 15.760 302.720 ;
                RECT 119.480 302.400 174.880 302.720 ;
                RECT 192.240 302.400 202.760 302.720 ;
                RECT 1118.400 302.400 1125.840 302.720 ;
                RECT 0.160 303.760 15.080 304.080 ;
                RECT 119.480 303.760 174.880 304.080 ;
                RECT 192.240 303.760 202.760 304.080 ;
                RECT 1118.400 303.760 1125.840 304.080 ;
                RECT 0.160 305.120 174.880 305.440 ;
                RECT 186.800 305.120 202.760 305.440 ;
                RECT 1118.400 305.120 1125.840 305.440 ;
                RECT 0.160 306.480 14.400 306.800 ;
                RECT 119.480 306.480 132.720 306.800 ;
                RECT 138.520 306.480 183.040 306.800 ;
                RECT 192.240 306.480 202.760 306.800 ;
                RECT 1118.400 306.480 1125.840 306.800 ;
                RECT 0.160 307.840 13.720 308.160 ;
                RECT 119.480 307.840 132.720 308.160 ;
                RECT 137.840 307.840 174.880 308.160 ;
                RECT 192.240 307.840 202.760 308.160 ;
                RECT 1118.400 307.840 1125.840 308.160 ;
                RECT 0.160 309.200 174.880 309.520 ;
                RECT 192.240 309.200 202.760 309.520 ;
                RECT 1118.400 309.200 1125.840 309.520 ;
                RECT 0.160 310.560 13.040 310.880 ;
                RECT 119.480 310.560 132.720 310.880 ;
                RECT 137.160 310.560 174.880 310.880 ;
                RECT 192.240 310.560 202.760 310.880 ;
                RECT 1118.400 310.560 1125.840 310.880 ;
                RECT 0.160 311.920 12.360 312.240 ;
                RECT 119.480 311.920 132.720 312.240 ;
                RECT 136.480 311.920 174.880 312.240 ;
                RECT 192.240 311.920 202.760 312.240 ;
                RECT 1118.400 311.920 1125.840 312.240 ;
                RECT 0.160 313.280 11.680 313.600 ;
                RECT 119.480 313.280 132.720 313.600 ;
                RECT 135.800 313.280 174.880 313.600 ;
                RECT 187.480 313.280 202.760 313.600 ;
                RECT 1118.400 313.280 1125.840 313.600 ;
                RECT 0.160 314.640 11.000 314.960 ;
                RECT 119.480 314.640 174.880 314.960 ;
                RECT 192.240 314.640 202.760 314.960 ;
                RECT 1118.400 314.640 1125.840 314.960 ;
                RECT 0.160 316.000 174.880 316.320 ;
                RECT 192.240 316.000 202.760 316.320 ;
                RECT 1118.400 316.000 1125.840 316.320 ;
                RECT 0.160 317.360 174.880 317.680 ;
                RECT 192.240 317.360 202.760 317.680 ;
                RECT 1118.400 317.360 1125.840 317.680 ;
                RECT 0.160 318.720 174.880 319.040 ;
                RECT 192.240 318.720 202.760 319.040 ;
                RECT 1118.400 318.720 1125.840 319.040 ;
                RECT 0.160 320.080 174.880 320.400 ;
                RECT 192.240 320.080 202.760 320.400 ;
                RECT 1118.400 320.080 1125.840 320.400 ;
                RECT 0.160 321.440 174.880 321.760 ;
                RECT 188.160 321.440 202.760 321.760 ;
                RECT 1118.400 321.440 1125.840 321.760 ;
                RECT 0.160 322.800 174.880 323.120 ;
                RECT 192.240 322.800 202.760 323.120 ;
                RECT 1118.400 322.800 1125.840 323.120 ;
                RECT 0.160 324.160 174.880 324.480 ;
                RECT 192.240 324.160 202.760 324.480 ;
                RECT 1118.400 324.160 1125.840 324.480 ;
                RECT 0.160 325.520 174.880 325.840 ;
                RECT 192.240 325.520 202.760 325.840 ;
                RECT 1118.400 325.520 1125.840 325.840 ;
                RECT 0.160 326.880 174.880 327.200 ;
                RECT 192.240 326.880 202.760 327.200 ;
                RECT 1118.400 326.880 1125.840 327.200 ;
                RECT 0.160 328.240 174.880 328.560 ;
                RECT 192.240 328.240 202.760 328.560 ;
                RECT 1118.400 328.240 1125.840 328.560 ;
                RECT 0.160 329.600 202.760 329.920 ;
                RECT 1118.400 329.600 1125.840 329.920 ;
                RECT 0.160 330.960 174.880 331.280 ;
                RECT 192.240 330.960 202.760 331.280 ;
                RECT 1118.400 330.960 1125.840 331.280 ;
                RECT 0.160 332.320 174.880 332.640 ;
                RECT 192.240 332.320 202.760 332.640 ;
                RECT 1118.400 332.320 1125.840 332.640 ;
                RECT 0.160 333.680 174.880 334.000 ;
                RECT 192.240 333.680 202.760 334.000 ;
                RECT 1118.400 333.680 1125.840 334.000 ;
                RECT 0.160 335.040 174.880 335.360 ;
                RECT 192.240 335.040 202.760 335.360 ;
                RECT 1118.400 335.040 1125.840 335.360 ;
                RECT 0.160 336.400 174.880 336.720 ;
                RECT 192.240 336.400 202.760 336.720 ;
                RECT 1118.400 336.400 1125.840 336.720 ;
                RECT 0.160 337.760 202.760 338.080 ;
                RECT 1118.400 337.760 1125.840 338.080 ;
                RECT 0.160 339.120 174.880 339.440 ;
                RECT 192.240 339.120 202.760 339.440 ;
                RECT 1118.400 339.120 1125.840 339.440 ;
                RECT 0.160 340.480 174.880 340.800 ;
                RECT 192.240 340.480 202.760 340.800 ;
                RECT 1118.400 340.480 1125.840 340.800 ;
                RECT 0.160 341.840 174.880 342.160 ;
                RECT 192.240 341.840 202.760 342.160 ;
                RECT 1118.400 341.840 1125.840 342.160 ;
                RECT 0.160 343.200 174.880 343.520 ;
                RECT 192.240 343.200 202.760 343.520 ;
                RECT 1118.400 343.200 1125.840 343.520 ;
                RECT 0.160 344.560 174.880 344.880 ;
                RECT 192.240 344.560 202.760 344.880 ;
                RECT 1118.400 344.560 1125.840 344.880 ;
                RECT 0.160 345.920 202.760 346.240 ;
                RECT 1118.400 345.920 1125.840 346.240 ;
                RECT 0.160 347.280 174.880 347.600 ;
                RECT 192.240 347.280 202.760 347.600 ;
                RECT 1118.400 347.280 1125.840 347.600 ;
                RECT 0.160 348.640 174.880 348.960 ;
                RECT 192.240 348.640 202.760 348.960 ;
                RECT 1118.400 348.640 1125.840 348.960 ;
                RECT 0.160 350.000 174.880 350.320 ;
                RECT 192.240 350.000 202.760 350.320 ;
                RECT 1118.400 350.000 1125.840 350.320 ;
                RECT 0.160 351.360 174.880 351.680 ;
                RECT 192.240 351.360 202.760 351.680 ;
                RECT 1118.400 351.360 1125.840 351.680 ;
                RECT 0.160 352.720 174.880 353.040 ;
                RECT 190.880 352.720 202.760 353.040 ;
                RECT 1118.400 352.720 1125.840 353.040 ;
                RECT 0.160 354.080 187.120 354.400 ;
                RECT 192.240 354.080 202.760 354.400 ;
                RECT 1118.400 354.080 1125.840 354.400 ;
                RECT 0.160 355.440 174.880 355.760 ;
                RECT 192.240 355.440 202.760 355.760 ;
                RECT 1118.400 355.440 1125.840 355.760 ;
                RECT 0.160 356.800 174.880 357.120 ;
                RECT 192.240 356.800 202.760 357.120 ;
                RECT 1118.400 356.800 1125.840 357.120 ;
                RECT 0.160 358.160 174.880 358.480 ;
                RECT 192.240 358.160 202.760 358.480 ;
                RECT 1118.400 358.160 1125.840 358.480 ;
                RECT 0.160 359.520 174.880 359.840 ;
                RECT 192.240 359.520 202.760 359.840 ;
                RECT 1118.400 359.520 1125.840 359.840 ;
                RECT 0.160 360.880 174.880 361.200 ;
                RECT 191.560 360.880 202.760 361.200 ;
                RECT 1118.400 360.880 1125.840 361.200 ;
                RECT 0.160 362.240 174.880 362.560 ;
                RECT 192.240 362.240 202.760 362.560 ;
                RECT 1118.400 362.240 1125.840 362.560 ;
                RECT 0.160 363.600 174.880 363.920 ;
                RECT 192.240 363.600 202.760 363.920 ;
                RECT 1118.400 363.600 1125.840 363.920 ;
                RECT 0.160 364.960 174.880 365.280 ;
                RECT 192.240 364.960 202.760 365.280 ;
                RECT 1118.400 364.960 1125.840 365.280 ;
                RECT 0.160 366.320 174.880 366.640 ;
                RECT 192.240 366.320 202.760 366.640 ;
                RECT 1118.400 366.320 1125.840 366.640 ;
                RECT 0.160 367.680 174.880 368.000 ;
                RECT 192.240 367.680 202.760 368.000 ;
                RECT 1118.400 367.680 1125.840 368.000 ;
                RECT 0.160 369.040 202.760 369.360 ;
                RECT 1118.400 369.040 1125.840 369.360 ;
                RECT 0.160 370.400 176.920 370.720 ;
                RECT 192.240 370.400 202.760 370.720 ;
                RECT 1118.400 370.400 1125.840 370.720 ;
                RECT 0.160 371.760 176.920 372.080 ;
                RECT 192.240 371.760 202.760 372.080 ;
                RECT 1118.400 371.760 1125.840 372.080 ;
                RECT 0.160 373.120 183.720 373.440 ;
                RECT 192.240 373.120 202.760 373.440 ;
                RECT 1118.400 373.120 1125.840 373.440 ;
                RECT 0.160 374.480 176.920 374.800 ;
                RECT 192.240 374.480 202.760 374.800 ;
                RECT 1118.400 374.480 1125.840 374.800 ;
                RECT 0.160 375.840 176.920 376.160 ;
                RECT 192.240 375.840 202.760 376.160 ;
                RECT 1118.400 375.840 1125.840 376.160 ;
                RECT 0.160 377.200 138.160 377.520 ;
                RECT 148.040 377.200 202.760 377.520 ;
                RECT 1118.400 377.200 1125.840 377.520 ;
                RECT 0.160 378.560 136.800 378.880 ;
                RECT 147.360 378.560 159.920 378.880 ;
                RECT 161.640 378.560 174.880 378.880 ;
                RECT 192.240 378.560 202.760 378.880 ;
                RECT 1118.400 378.560 1125.840 378.880 ;
                RECT 0.160 379.920 159.920 380.240 ;
                RECT 163.680 379.920 174.880 380.240 ;
                RECT 192.240 379.920 202.760 380.240 ;
                RECT 1118.400 379.920 1125.840 380.240 ;
                RECT 0.160 381.280 159.920 381.600 ;
                RECT 164.360 381.280 174.880 381.600 ;
                RECT 192.240 381.280 202.760 381.600 ;
                RECT 1118.400 381.280 1125.840 381.600 ;
                RECT 0.160 382.640 159.920 382.960 ;
                RECT 165.040 382.640 174.880 382.960 ;
                RECT 192.240 382.640 202.760 382.960 ;
                RECT 1118.400 382.640 1125.840 382.960 ;
                RECT 0.160 384.000 159.920 384.320 ;
                RECT 165.720 384.000 174.880 384.320 ;
                RECT 192.240 384.000 202.760 384.320 ;
                RECT 1118.400 384.000 1125.840 384.320 ;
                RECT 0.160 385.360 202.760 385.680 ;
                RECT 1118.400 385.360 1125.840 385.680 ;
                RECT 0.160 386.720 174.880 387.040 ;
                RECT 192.240 386.720 202.760 387.040 ;
                RECT 1118.400 386.720 1125.840 387.040 ;
                RECT 0.160 388.080 174.880 388.400 ;
                RECT 192.240 388.080 202.760 388.400 ;
                RECT 1118.400 388.080 1125.840 388.400 ;
                RECT 0.160 389.440 174.880 389.760 ;
                RECT 192.240 389.440 202.760 389.760 ;
                RECT 1118.400 389.440 1125.840 389.760 ;
                RECT 0.160 390.800 174.880 391.120 ;
                RECT 192.240 390.800 202.760 391.120 ;
                RECT 1118.400 390.800 1125.840 391.120 ;
                RECT 0.160 392.160 136.120 392.480 ;
                RECT 148.720 392.160 174.880 392.480 ;
                RECT 177.960 392.160 202.760 392.480 ;
                RECT 1118.400 392.160 1125.840 392.480 ;
                RECT 0.160 393.520 134.760 393.840 ;
                RECT 147.360 393.520 188.480 393.840 ;
                RECT 192.240 393.520 202.760 393.840 ;
                RECT 1118.400 393.520 1125.840 393.840 ;
                RECT 0.160 394.880 159.920 395.200 ;
                RECT 162.320 394.880 174.880 395.200 ;
                RECT 192.240 394.880 202.760 395.200 ;
                RECT 1118.400 394.880 1125.840 395.200 ;
                RECT 0.160 396.240 159.920 396.560 ;
                RECT 162.320 396.240 174.880 396.560 ;
                RECT 192.240 396.240 202.760 396.560 ;
                RECT 1118.400 396.240 1125.840 396.560 ;
                RECT 0.160 397.600 159.920 397.920 ;
                RECT 163.000 397.600 174.880 397.920 ;
                RECT 192.240 397.600 202.760 397.920 ;
                RECT 1118.400 397.600 1125.840 397.920 ;
                RECT 0.160 398.960 159.920 399.280 ;
                RECT 161.640 398.960 174.880 399.280 ;
                RECT 192.240 398.960 202.760 399.280 ;
                RECT 1118.400 398.960 1125.840 399.280 ;
                RECT 0.160 400.320 159.920 400.640 ;
                RECT 163.680 400.320 174.880 400.640 ;
                RECT 178.640 400.320 202.760 400.640 ;
                RECT 1118.400 400.320 1125.840 400.640 ;
                RECT 0.160 401.680 174.880 402.000 ;
                RECT 192.240 401.680 202.760 402.000 ;
                RECT 1118.400 401.680 1125.840 402.000 ;
                RECT 0.160 403.040 174.880 403.360 ;
                RECT 192.240 403.040 202.760 403.360 ;
                RECT 1118.400 403.040 1125.840 403.360 ;
                RECT 0.160 404.400 174.880 404.720 ;
                RECT 192.240 404.400 202.760 404.720 ;
                RECT 1118.400 404.400 1125.840 404.720 ;
                RECT 0.160 405.760 174.880 406.080 ;
                RECT 192.240 405.760 202.760 406.080 ;
                RECT 1118.400 405.760 1125.840 406.080 ;
                RECT 0.160 407.120 174.880 407.440 ;
                RECT 192.240 407.120 202.760 407.440 ;
                RECT 1118.400 407.120 1125.840 407.440 ;
                RECT 0.160 408.480 202.760 408.800 ;
                RECT 1118.400 408.480 1125.840 408.800 ;
                RECT 0.160 409.840 174.880 410.160 ;
                RECT 192.240 409.840 202.760 410.160 ;
                RECT 1118.400 409.840 1125.840 410.160 ;
                RECT 0.160 411.200 174.880 411.520 ;
                RECT 192.240 411.200 202.760 411.520 ;
                RECT 1118.400 411.200 1125.840 411.520 ;
                RECT 0.160 412.560 174.880 412.880 ;
                RECT 192.240 412.560 202.760 412.880 ;
                RECT 1118.400 412.560 1125.840 412.880 ;
                RECT 0.160 413.920 174.880 414.240 ;
                RECT 192.240 413.920 202.760 414.240 ;
                RECT 1118.400 413.920 1125.840 414.240 ;
                RECT 0.160 415.280 174.880 415.600 ;
                RECT 192.240 415.280 202.760 415.600 ;
                RECT 1118.400 415.280 1125.840 415.600 ;
                RECT 0.160 416.640 202.760 416.960 ;
                RECT 1118.400 416.640 1125.840 416.960 ;
                RECT 0.160 418.000 174.880 418.320 ;
                RECT 192.240 418.000 202.760 418.320 ;
                RECT 1118.400 418.000 1125.840 418.320 ;
                RECT 0.160 419.360 174.880 419.680 ;
                RECT 192.240 419.360 202.760 419.680 ;
                RECT 1118.400 419.360 1125.840 419.680 ;
                RECT 0.160 420.720 174.880 421.040 ;
                RECT 192.240 420.720 202.760 421.040 ;
                RECT 1118.400 420.720 1125.840 421.040 ;
                RECT 0.160 422.080 174.880 422.400 ;
                RECT 192.240 422.080 202.760 422.400 ;
                RECT 1118.400 422.080 1125.840 422.400 ;
                RECT 0.160 423.440 174.880 423.760 ;
                RECT 192.240 423.440 202.760 423.760 ;
                RECT 1118.400 423.440 1125.840 423.760 ;
                RECT 0.160 424.800 202.760 425.120 ;
                RECT 1118.400 424.800 1125.840 425.120 ;
                RECT 0.160 426.160 174.880 426.480 ;
                RECT 192.240 426.160 202.760 426.480 ;
                RECT 1118.400 426.160 1125.840 426.480 ;
                RECT 0.160 427.520 174.880 427.840 ;
                RECT 192.240 427.520 202.760 427.840 ;
                RECT 1118.400 427.520 1125.840 427.840 ;
                RECT 0.160 428.880 174.880 429.200 ;
                RECT 192.240 428.880 202.760 429.200 ;
                RECT 1118.400 428.880 1125.840 429.200 ;
                RECT 0.160 430.240 174.880 430.560 ;
                RECT 192.240 430.240 202.760 430.560 ;
                RECT 1118.400 430.240 1125.840 430.560 ;
                RECT 0.160 431.600 174.880 431.920 ;
                RECT 181.360 431.600 202.760 431.920 ;
                RECT 1118.400 431.600 1125.840 431.920 ;
                RECT 0.160 432.960 183.040 433.280 ;
                RECT 192.240 432.960 202.760 433.280 ;
                RECT 1118.400 432.960 1125.840 433.280 ;
                RECT 0.160 434.320 174.880 434.640 ;
                RECT 192.240 434.320 202.760 434.640 ;
                RECT 1118.400 434.320 1125.840 434.640 ;
                RECT 0.160 435.680 174.880 436.000 ;
                RECT 192.240 435.680 202.760 436.000 ;
                RECT 1118.400 435.680 1125.840 436.000 ;
                RECT 0.160 437.040 174.880 437.360 ;
                RECT 192.240 437.040 202.760 437.360 ;
                RECT 1118.400 437.040 1125.840 437.360 ;
                RECT 0.160 438.400 174.880 438.720 ;
                RECT 192.240 438.400 202.760 438.720 ;
                RECT 1118.400 438.400 1125.840 438.720 ;
                RECT 0.160 439.760 174.880 440.080 ;
                RECT 182.040 439.760 202.760 440.080 ;
                RECT 1118.400 439.760 1125.840 440.080 ;
                RECT 0.160 441.120 174.880 441.440 ;
                RECT 192.240 441.120 202.760 441.440 ;
                RECT 1118.400 441.120 1125.840 441.440 ;
                RECT 0.160 442.480 174.880 442.800 ;
                RECT 192.240 442.480 202.760 442.800 ;
                RECT 1118.400 442.480 1125.840 442.800 ;
                RECT 0.160 443.840 174.880 444.160 ;
                RECT 192.240 443.840 202.760 444.160 ;
                RECT 1118.400 443.840 1125.840 444.160 ;
                RECT 0.160 445.200 174.880 445.520 ;
                RECT 192.240 445.200 202.760 445.520 ;
                RECT 1118.400 445.200 1125.840 445.520 ;
                RECT 0.160 446.560 174.880 446.880 ;
                RECT 192.240 446.560 202.760 446.880 ;
                RECT 1118.400 446.560 1125.840 446.880 ;
                RECT 0.160 447.920 202.760 448.240 ;
                RECT 1118.400 447.920 1125.840 448.240 ;
                RECT 0.160 449.280 174.880 449.600 ;
                RECT 192.240 449.280 202.760 449.600 ;
                RECT 1118.400 449.280 1125.840 449.600 ;
                RECT 0.160 450.640 174.880 450.960 ;
                RECT 192.240 450.640 202.760 450.960 ;
                RECT 1118.400 450.640 1125.840 450.960 ;
                RECT 0.160 452.000 174.880 452.320 ;
                RECT 192.240 452.000 202.760 452.320 ;
                RECT 1118.400 452.000 1125.840 452.320 ;
                RECT 0.160 453.360 174.880 453.680 ;
                RECT 192.240 453.360 202.760 453.680 ;
                RECT 1118.400 453.360 1125.840 453.680 ;
                RECT 0.160 454.720 174.880 455.040 ;
                RECT 192.240 454.720 202.760 455.040 ;
                RECT 1118.400 454.720 1125.840 455.040 ;
                RECT 0.160 456.080 202.760 456.400 ;
                RECT 1118.400 456.080 1125.840 456.400 ;
                RECT 0.160 457.440 174.880 457.760 ;
                RECT 192.240 457.440 202.760 457.760 ;
                RECT 1118.400 457.440 1125.840 457.760 ;
                RECT 0.160 458.800 174.880 459.120 ;
                RECT 192.240 458.800 202.760 459.120 ;
                RECT 1118.400 458.800 1125.840 459.120 ;
                RECT 0.160 460.160 174.880 460.480 ;
                RECT 192.240 460.160 202.760 460.480 ;
                RECT 1118.400 460.160 1125.840 460.480 ;
                RECT 0.160 461.520 174.880 461.840 ;
                RECT 192.240 461.520 202.760 461.840 ;
                RECT 1118.400 461.520 1125.840 461.840 ;
                RECT 0.160 462.880 174.880 463.200 ;
                RECT 192.240 462.880 202.760 463.200 ;
                RECT 1118.400 462.880 1125.840 463.200 ;
                RECT 0.160 464.240 202.760 464.560 ;
                RECT 1118.400 464.240 1125.840 464.560 ;
                RECT 0.160 465.600 174.880 465.920 ;
                RECT 192.240 465.600 202.760 465.920 ;
                RECT 1118.400 465.600 1125.840 465.920 ;
                RECT 0.160 466.960 174.880 467.280 ;
                RECT 192.240 466.960 202.760 467.280 ;
                RECT 1118.400 466.960 1125.840 467.280 ;
                RECT 0.160 468.320 174.880 468.640 ;
                RECT 192.240 468.320 202.760 468.640 ;
                RECT 1118.400 468.320 1125.840 468.640 ;
                RECT 0.160 469.680 174.880 470.000 ;
                RECT 192.240 469.680 202.760 470.000 ;
                RECT 1118.400 469.680 1125.840 470.000 ;
                RECT 0.160 471.040 174.880 471.360 ;
                RECT 184.080 471.040 202.760 471.360 ;
                RECT 1118.400 471.040 1125.840 471.360 ;
                RECT 0.160 472.400 185.080 472.720 ;
                RECT 192.240 472.400 202.760 472.720 ;
                RECT 1118.400 472.400 1125.840 472.720 ;
                RECT 0.160 473.760 178.280 474.080 ;
                RECT 192.240 473.760 202.760 474.080 ;
                RECT 1118.400 473.760 1125.840 474.080 ;
                RECT 0.160 475.120 178.280 475.440 ;
                RECT 192.240 475.120 202.760 475.440 ;
                RECT 1118.400 475.120 1125.840 475.440 ;
                RECT 0.160 476.480 178.280 476.800 ;
                RECT 192.240 476.480 202.760 476.800 ;
                RECT 1118.400 476.480 1125.840 476.800 ;
                RECT 0.160 477.840 178.280 478.160 ;
                RECT 192.240 477.840 202.760 478.160 ;
                RECT 1118.400 477.840 1125.840 478.160 ;
                RECT 0.160 479.200 202.760 479.520 ;
                RECT 1118.400 479.200 1125.840 479.520 ;
                RECT 0.160 480.560 187.120 480.880 ;
                RECT 192.240 480.560 202.760 480.880 ;
                RECT 1118.400 480.560 1125.840 480.880 ;
                RECT 0.160 481.920 178.280 482.240 ;
                RECT 192.240 481.920 202.760 482.240 ;
                RECT 1118.400 481.920 1125.840 482.240 ;
                RECT 0.160 483.280 178.280 483.600 ;
                RECT 192.240 483.280 202.760 483.600 ;
                RECT 1118.400 483.280 1125.840 483.600 ;
                RECT 0.160 484.640 178.280 484.960 ;
                RECT 192.240 484.640 202.760 484.960 ;
                RECT 1118.400 484.640 1125.840 484.960 ;
                RECT 0.160 486.000 178.280 486.320 ;
                RECT 192.240 486.000 202.760 486.320 ;
                RECT 1118.400 486.000 1125.840 486.320 ;
                RECT 0.160 487.360 202.760 487.680 ;
                RECT 1118.400 487.360 1125.840 487.680 ;
                RECT 0.160 488.720 178.280 489.040 ;
                RECT 192.240 488.720 202.760 489.040 ;
                RECT 1118.400 488.720 1125.840 489.040 ;
                RECT 0.160 490.080 189.160 490.400 ;
                RECT 192.240 490.080 202.760 490.400 ;
                RECT 1118.400 490.080 1125.840 490.400 ;
                RECT 0.160 491.440 178.280 491.760 ;
                RECT 192.240 491.440 202.760 491.760 ;
                RECT 1118.400 491.440 1125.840 491.760 ;
                RECT 0.160 492.800 178.280 493.120 ;
                RECT 192.240 492.800 202.760 493.120 ;
                RECT 1118.400 492.800 1125.840 493.120 ;
                RECT 0.160 494.160 178.280 494.480 ;
                RECT 192.240 494.160 202.760 494.480 ;
                RECT 1118.400 494.160 1125.840 494.480 ;
                RECT 0.160 495.520 202.760 495.840 ;
                RECT 1118.400 495.520 1125.840 495.840 ;
                RECT 0.160 496.880 178.960 497.200 ;
                RECT 192.240 496.880 202.760 497.200 ;
                RECT 1118.400 496.880 1125.840 497.200 ;
                RECT 0.160 498.240 178.960 498.560 ;
                RECT 192.240 498.240 202.760 498.560 ;
                RECT 1118.400 498.240 1125.840 498.560 ;
                RECT 0.160 499.600 183.720 499.920 ;
                RECT 192.240 499.600 202.760 499.920 ;
                RECT 1118.400 499.600 1125.840 499.920 ;
                RECT 0.160 500.960 178.960 501.280 ;
                RECT 192.240 500.960 202.760 501.280 ;
                RECT 1118.400 500.960 1125.840 501.280 ;
                RECT 0.160 502.320 178.960 502.640 ;
                RECT 192.240 502.320 202.760 502.640 ;
                RECT 1118.400 502.320 1125.840 502.640 ;
                RECT 0.160 503.680 202.760 504.000 ;
                RECT 1118.400 503.680 1125.840 504.000 ;
                RECT 0.160 505.040 178.960 505.360 ;
                RECT 192.240 505.040 202.760 505.360 ;
                RECT 1118.400 505.040 1125.840 505.360 ;
                RECT 0.160 506.400 178.960 506.720 ;
                RECT 192.240 506.400 202.760 506.720 ;
                RECT 1118.400 506.400 1125.840 506.720 ;
                RECT 0.160 507.760 178.960 508.080 ;
                RECT 192.240 507.760 202.760 508.080 ;
                RECT 1118.400 507.760 1125.840 508.080 ;
                RECT 0.160 509.120 186.440 509.440 ;
                RECT 192.240 509.120 202.760 509.440 ;
                RECT 1118.400 509.120 1125.840 509.440 ;
                RECT 0.160 510.480 178.960 510.800 ;
                RECT 192.240 510.480 202.760 510.800 ;
                RECT 1118.400 510.480 1125.840 510.800 ;
                RECT 0.160 511.840 202.760 512.160 ;
                RECT 1118.400 511.840 1125.840 512.160 ;
                RECT 0.160 513.200 178.960 513.520 ;
                RECT 192.240 513.200 202.760 513.520 ;
                RECT 1118.400 513.200 1125.840 513.520 ;
                RECT 0.160 514.560 178.960 514.880 ;
                RECT 192.240 514.560 202.760 514.880 ;
                RECT 1118.400 514.560 1125.840 514.880 ;
                RECT 0.160 515.920 178.960 516.240 ;
                RECT 192.240 515.920 202.760 516.240 ;
                RECT 1118.400 515.920 1125.840 516.240 ;
                RECT 0.160 517.280 178.960 517.600 ;
                RECT 192.240 517.280 202.760 517.600 ;
                RECT 1118.400 517.280 1125.840 517.600 ;
                RECT 0.160 518.640 202.760 518.960 ;
                RECT 1118.400 518.640 1125.840 518.960 ;
                RECT 0.160 520.000 188.480 520.320 ;
                RECT 192.240 520.000 202.760 520.320 ;
                RECT 1118.400 520.000 1125.840 520.320 ;
                RECT 0.160 521.360 178.960 521.680 ;
                RECT 192.240 521.360 202.760 521.680 ;
                RECT 1118.400 521.360 1125.840 521.680 ;
                RECT 0.160 522.720 178.960 523.040 ;
                RECT 192.240 522.720 202.760 523.040 ;
                RECT 1118.400 522.720 1125.840 523.040 ;
                RECT 0.160 524.080 178.960 524.400 ;
                RECT 192.240 524.080 202.760 524.400 ;
                RECT 1118.400 524.080 1125.840 524.400 ;
                RECT 0.160 525.440 178.960 525.760 ;
                RECT 192.240 525.440 202.760 525.760 ;
                RECT 1118.400 525.440 1125.840 525.760 ;
                RECT 0.160 526.800 202.760 527.120 ;
                RECT 1118.400 526.800 1125.840 527.120 ;
                RECT 0.160 528.160 178.960 528.480 ;
                RECT 192.240 528.160 202.760 528.480 ;
                RECT 1118.400 528.160 1125.840 528.480 ;
                RECT 0.160 529.520 183.720 529.840 ;
                RECT 192.240 529.520 202.760 529.840 ;
                RECT 1118.400 529.520 1125.840 529.840 ;
                RECT 0.160 530.880 178.960 531.200 ;
                RECT 192.240 530.880 202.760 531.200 ;
                RECT 1118.400 530.880 1125.840 531.200 ;
                RECT 0.160 532.240 178.960 532.560 ;
                RECT 192.240 532.240 202.760 532.560 ;
                RECT 1118.400 532.240 1125.840 532.560 ;
                RECT 0.160 533.600 178.960 533.920 ;
                RECT 192.240 533.600 202.760 533.920 ;
                RECT 1118.400 533.600 1125.840 533.920 ;
                RECT 0.160 534.960 202.760 535.280 ;
                RECT 1118.400 534.960 1125.840 535.280 ;
                RECT 0.160 536.320 178.960 536.640 ;
                RECT 192.240 536.320 202.760 536.640 ;
                RECT 1118.400 536.320 1125.840 536.640 ;
                RECT 0.160 537.680 178.960 538.000 ;
                RECT 192.240 537.680 202.760 538.000 ;
                RECT 1118.400 537.680 1125.840 538.000 ;
                RECT 0.160 539.040 185.760 539.360 ;
                RECT 192.240 539.040 202.760 539.360 ;
                RECT 1118.400 539.040 1125.840 539.360 ;
                RECT 0.160 540.400 178.960 540.720 ;
                RECT 192.240 540.400 202.760 540.720 ;
                RECT 1118.400 540.400 1125.840 540.720 ;
                RECT 0.160 541.760 178.960 542.080 ;
                RECT 192.240 541.760 202.760 542.080 ;
                RECT 1118.400 541.760 1125.840 542.080 ;
                RECT 0.160 543.120 202.760 543.440 ;
                RECT 1118.400 543.120 1125.840 543.440 ;
                RECT 0.160 544.480 178.960 544.800 ;
                RECT 192.240 544.480 202.760 544.800 ;
                RECT 1118.400 544.480 1125.840 544.800 ;
                RECT 0.160 545.840 178.960 546.160 ;
                RECT 192.240 545.840 202.760 546.160 ;
                RECT 1118.400 545.840 1125.840 546.160 ;
                RECT 0.160 547.200 178.960 547.520 ;
                RECT 192.240 547.200 202.760 547.520 ;
                RECT 1118.400 547.200 1125.840 547.520 ;
                RECT 0.160 548.560 188.480 548.880 ;
                RECT 192.240 548.560 202.760 548.880 ;
                RECT 1118.400 548.560 1125.840 548.880 ;
                RECT 0.160 549.920 178.960 550.240 ;
                RECT 192.240 549.920 202.760 550.240 ;
                RECT 1118.400 549.920 1125.840 550.240 ;
                RECT 0.160 551.280 202.760 551.600 ;
                RECT 1118.400 551.280 1125.840 551.600 ;
                RECT 0.160 552.640 178.960 552.960 ;
                RECT 192.240 552.640 202.760 552.960 ;
                RECT 1118.400 552.640 1125.840 552.960 ;
                RECT 0.160 554.000 178.960 554.320 ;
                RECT 192.240 554.000 202.760 554.320 ;
                RECT 1118.400 554.000 1125.840 554.320 ;
                RECT 0.160 555.360 178.960 555.680 ;
                RECT 192.240 555.360 202.760 555.680 ;
                RECT 1118.400 555.360 1125.840 555.680 ;
                RECT 0.160 556.720 178.960 557.040 ;
                RECT 192.240 556.720 202.760 557.040 ;
                RECT 1118.400 556.720 1125.840 557.040 ;
                RECT 0.160 558.080 202.760 558.400 ;
                RECT 1118.400 558.080 1125.840 558.400 ;
                RECT 0.160 559.440 183.040 559.760 ;
                RECT 192.240 559.440 202.760 559.760 ;
                RECT 1118.400 559.440 1125.840 559.760 ;
                RECT 0.160 560.800 179.640 561.120 ;
                RECT 192.240 560.800 202.760 561.120 ;
                RECT 1118.400 560.800 1125.840 561.120 ;
                RECT 0.160 562.160 179.640 562.480 ;
                RECT 192.240 562.160 202.760 562.480 ;
                RECT 1118.400 562.160 1125.840 562.480 ;
                RECT 0.160 563.520 179.640 563.840 ;
                RECT 192.240 563.520 202.760 563.840 ;
                RECT 1118.400 563.520 1125.840 563.840 ;
                RECT 0.160 564.880 179.640 565.200 ;
                RECT 192.240 564.880 202.760 565.200 ;
                RECT 1118.400 564.880 1125.840 565.200 ;
                RECT 0.160 566.240 202.760 566.560 ;
                RECT 1118.400 566.240 1125.840 566.560 ;
                RECT 0.160 567.600 185.080 567.920 ;
                RECT 192.240 567.600 202.760 567.920 ;
                RECT 1118.400 567.600 1125.840 567.920 ;
                RECT 0.160 568.960 185.080 569.280 ;
                RECT 192.240 568.960 202.760 569.280 ;
                RECT 1118.400 568.960 1125.840 569.280 ;
                RECT 0.160 570.320 179.640 570.640 ;
                RECT 192.240 570.320 202.760 570.640 ;
                RECT 1118.400 570.320 1125.840 570.640 ;
                RECT 0.160 571.680 179.640 572.000 ;
                RECT 192.240 571.680 202.760 572.000 ;
                RECT 1118.400 571.680 1125.840 572.000 ;
                RECT 0.160 573.040 179.640 573.360 ;
                RECT 192.240 573.040 202.760 573.360 ;
                RECT 1118.400 573.040 1125.840 573.360 ;
                RECT 0.160 574.400 202.760 574.720 ;
                RECT 1118.400 574.400 1125.840 574.720 ;
                RECT 0.160 575.760 179.640 576.080 ;
                RECT 192.240 575.760 202.760 576.080 ;
                RECT 1118.400 575.760 1125.840 576.080 ;
                RECT 0.160 577.120 187.120 577.440 ;
                RECT 192.240 577.120 202.760 577.440 ;
                RECT 1118.400 577.120 1125.840 577.440 ;
                RECT 0.160 578.480 187.800 578.800 ;
                RECT 192.240 578.480 202.760 578.800 ;
                RECT 1118.400 578.480 1125.840 578.800 ;
                RECT 0.160 579.840 179.640 580.160 ;
                RECT 192.240 579.840 202.760 580.160 ;
                RECT 1118.400 579.840 1125.840 580.160 ;
                RECT 0.160 581.200 179.640 581.520 ;
                RECT 192.240 581.200 202.760 581.520 ;
                RECT 1118.400 581.200 1125.840 581.520 ;
                RECT 0.160 582.560 202.760 582.880 ;
                RECT 1118.400 582.560 1125.840 582.880 ;
                RECT 0.160 583.920 179.640 584.240 ;
                RECT 192.240 583.920 202.760 584.240 ;
                RECT 1118.400 583.920 1125.840 584.240 ;
                RECT 0.160 585.280 179.640 585.600 ;
                RECT 192.240 585.280 202.760 585.600 ;
                RECT 1118.400 585.280 1125.840 585.600 ;
                RECT 0.160 586.640 179.640 586.960 ;
                RECT 192.240 586.640 202.760 586.960 ;
                RECT 1118.400 586.640 1125.840 586.960 ;
                RECT 0.160 588.000 190.520 588.320 ;
                RECT 192.240 588.000 202.760 588.320 ;
                RECT 1118.400 588.000 1125.840 588.320 ;
                RECT 0.160 589.360 179.640 589.680 ;
                RECT 192.240 589.360 202.760 589.680 ;
                RECT 1118.400 589.360 1125.840 589.680 ;
                RECT 0.160 590.720 202.760 591.040 ;
                RECT 1118.400 590.720 1125.840 591.040 ;
                RECT 0.160 592.080 180.320 592.400 ;
                RECT 192.240 592.080 202.760 592.400 ;
                RECT 1118.400 592.080 1125.840 592.400 ;
                RECT 0.160 593.440 180.320 593.760 ;
                RECT 192.240 593.440 202.760 593.760 ;
                RECT 1118.400 593.440 1125.840 593.760 ;
                RECT 0.160 594.800 180.320 595.120 ;
                RECT 192.240 594.800 202.760 595.120 ;
                RECT 1118.400 594.800 1125.840 595.120 ;
                RECT 0.160 596.160 180.320 596.480 ;
                RECT 192.240 596.160 202.760 596.480 ;
                RECT 1118.400 596.160 1125.840 596.480 ;
                RECT 0.160 597.520 202.760 597.840 ;
                RECT 1118.400 597.520 1125.840 597.840 ;
                RECT 0.160 598.880 185.080 599.200 ;
                RECT 192.240 598.880 202.760 599.200 ;
                RECT 1118.400 598.880 1125.840 599.200 ;
                RECT 0.160 600.240 180.320 600.560 ;
                RECT 192.240 600.240 202.760 600.560 ;
                RECT 1118.400 600.240 1125.840 600.560 ;
                RECT 0.160 601.600 180.320 601.920 ;
                RECT 192.240 601.600 202.760 601.920 ;
                RECT 1118.400 601.600 1125.840 601.920 ;
                RECT 0.160 602.960 180.320 603.280 ;
                RECT 192.240 602.960 202.760 603.280 ;
                RECT 1118.400 602.960 1125.840 603.280 ;
                RECT 0.160 604.320 180.320 604.640 ;
                RECT 192.240 604.320 202.760 604.640 ;
                RECT 1118.400 604.320 1125.840 604.640 ;
                RECT 0.160 605.680 202.760 606.000 ;
                RECT 1118.400 605.680 1125.840 606.000 ;
                RECT 0.160 607.040 187.120 607.360 ;
                RECT 192.240 607.040 202.760 607.360 ;
                RECT 1118.400 607.040 1125.840 607.360 ;
                RECT 0.160 608.400 180.320 608.720 ;
                RECT 192.240 608.400 202.760 608.720 ;
                RECT 1118.400 608.400 1125.840 608.720 ;
                RECT 0.160 609.760 180.320 610.080 ;
                RECT 192.240 609.760 202.760 610.080 ;
                RECT 1118.400 609.760 1125.840 610.080 ;
                RECT 0.160 611.120 180.320 611.440 ;
                RECT 192.240 611.120 202.760 611.440 ;
                RECT 1118.400 611.120 1125.840 611.440 ;
                RECT 0.160 612.480 180.320 612.800 ;
                RECT 192.240 612.480 202.760 612.800 ;
                RECT 1118.400 612.480 1125.840 612.800 ;
                RECT 0.160 613.840 202.760 614.160 ;
                RECT 1118.400 613.840 1125.840 614.160 ;
                RECT 0.160 615.200 180.320 615.520 ;
                RECT 192.240 615.200 202.760 615.520 ;
                RECT 1118.400 615.200 1125.840 615.520 ;
                RECT 0.160 616.560 189.160 616.880 ;
                RECT 192.240 616.560 202.760 616.880 ;
                RECT 1118.400 616.560 1125.840 616.880 ;
                RECT 0.160 617.920 180.320 618.240 ;
                RECT 192.240 617.920 202.760 618.240 ;
                RECT 1118.400 617.920 1125.840 618.240 ;
                RECT 0.160 619.280 180.320 619.600 ;
                RECT 192.240 619.280 202.760 619.600 ;
                RECT 1118.400 619.280 1125.840 619.600 ;
                RECT 0.160 620.640 180.320 620.960 ;
                RECT 192.240 620.640 202.760 620.960 ;
                RECT 1118.400 620.640 1125.840 620.960 ;
                RECT 0.160 622.000 202.760 622.320 ;
                RECT 1118.400 622.000 1125.840 622.320 ;
                RECT 0.160 623.360 180.320 623.680 ;
                RECT 192.240 623.360 202.760 623.680 ;
                RECT 1118.400 623.360 1125.840 623.680 ;
                RECT 0.160 624.720 180.320 625.040 ;
                RECT 192.240 624.720 202.760 625.040 ;
                RECT 1118.400 624.720 1125.840 625.040 ;
                RECT 0.160 626.080 183.720 626.400 ;
                RECT 192.240 626.080 202.760 626.400 ;
                RECT 1118.400 626.080 1125.840 626.400 ;
                RECT 0.160 627.440 184.400 627.760 ;
                RECT 192.240 627.440 202.760 627.760 ;
                RECT 1118.400 627.440 1125.840 627.760 ;
                RECT 0.160 628.800 180.320 629.120 ;
                RECT 192.240 628.800 202.760 629.120 ;
                RECT 1118.400 628.800 1125.840 629.120 ;
                RECT 0.160 630.160 202.760 630.480 ;
                RECT 1118.400 630.160 1125.840 630.480 ;
                RECT 0.160 631.520 180.320 631.840 ;
                RECT 192.240 631.520 202.760 631.840 ;
                RECT 1118.400 631.520 1125.840 631.840 ;
                RECT 0.160 632.880 180.320 633.200 ;
                RECT 192.240 632.880 202.760 633.200 ;
                RECT 1118.400 632.880 1125.840 633.200 ;
                RECT 0.160 634.240 180.320 634.560 ;
                RECT 192.240 634.240 202.760 634.560 ;
                RECT 1118.400 634.240 1125.840 634.560 ;
                RECT 0.160 635.600 180.320 635.920 ;
                RECT 192.240 635.600 202.760 635.920 ;
                RECT 1118.400 635.600 1125.840 635.920 ;
                RECT 0.160 636.960 202.760 637.280 ;
                RECT 1118.400 636.960 1125.840 637.280 ;
                RECT 0.160 638.320 187.120 638.640 ;
                RECT 192.240 638.320 202.760 638.640 ;
                RECT 1118.400 638.320 1125.840 638.640 ;
                RECT 0.160 639.680 180.320 640.000 ;
                RECT 192.240 639.680 202.760 640.000 ;
                RECT 1118.400 639.680 1125.840 640.000 ;
                RECT 0.160 641.040 180.320 641.360 ;
                RECT 192.240 641.040 202.760 641.360 ;
                RECT 1118.400 641.040 1125.840 641.360 ;
                RECT 0.160 642.400 180.320 642.720 ;
                RECT 192.240 642.400 202.760 642.720 ;
                RECT 1118.400 642.400 1125.840 642.720 ;
                RECT 0.160 643.760 180.320 644.080 ;
                RECT 192.240 643.760 202.760 644.080 ;
                RECT 1118.400 643.760 1125.840 644.080 ;
                RECT 0.160 645.120 202.760 645.440 ;
                RECT 1118.400 645.120 1125.840 645.440 ;
                RECT 0.160 646.480 188.480 646.800 ;
                RECT 192.240 646.480 202.760 646.800 ;
                RECT 1118.400 646.480 1125.840 646.800 ;
                RECT 0.160 647.840 180.320 648.160 ;
                RECT 192.240 647.840 202.760 648.160 ;
                RECT 1118.400 647.840 1125.840 648.160 ;
                RECT 0.160 649.200 180.320 649.520 ;
                RECT 192.240 649.200 202.760 649.520 ;
                RECT 1118.400 649.200 1125.840 649.520 ;
                RECT 0.160 650.560 180.320 650.880 ;
                RECT 192.240 650.560 202.760 650.880 ;
                RECT 1118.400 650.560 1125.840 650.880 ;
                RECT 0.160 651.920 180.320 652.240 ;
                RECT 192.240 651.920 202.760 652.240 ;
                RECT 1118.400 651.920 1125.840 652.240 ;
                RECT 0.160 653.280 202.760 653.600 ;
                RECT 1118.400 653.280 1125.840 653.600 ;
                RECT 0.160 654.640 181.000 654.960 ;
                RECT 192.240 654.640 202.760 654.960 ;
                RECT 1118.400 654.640 1125.840 654.960 ;
                RECT 0.160 656.000 183.720 656.320 ;
                RECT 192.240 656.000 202.760 656.320 ;
                RECT 1118.400 656.000 1125.840 656.320 ;
                RECT 0.160 657.360 181.000 657.680 ;
                RECT 192.240 657.360 202.760 657.680 ;
                RECT 1118.400 657.360 1125.840 657.680 ;
                RECT 0.160 658.720 181.000 659.040 ;
                RECT 192.240 658.720 202.760 659.040 ;
                RECT 1118.400 658.720 1125.840 659.040 ;
                RECT 0.160 660.080 181.000 660.400 ;
                RECT 192.240 660.080 202.760 660.400 ;
                RECT 1118.400 660.080 1125.840 660.400 ;
                RECT 0.160 661.440 202.760 661.760 ;
                RECT 1118.400 661.440 1125.840 661.760 ;
                RECT 0.160 662.800 181.000 663.120 ;
                RECT 192.240 662.800 202.760 663.120 ;
                RECT 1118.400 662.800 1125.840 663.120 ;
                RECT 0.160 664.160 181.000 664.480 ;
                RECT 192.240 664.160 202.760 664.480 ;
                RECT 1118.400 664.160 1125.840 664.480 ;
                RECT 0.160 665.520 185.760 665.840 ;
                RECT 192.240 665.520 202.760 665.840 ;
                RECT 1118.400 665.520 1125.840 665.840 ;
                RECT 0.160 666.880 181.000 667.200 ;
                RECT 192.240 666.880 202.760 667.200 ;
                RECT 1118.400 666.880 1125.840 667.200 ;
                RECT 0.160 668.240 181.000 668.560 ;
                RECT 192.240 668.240 202.760 668.560 ;
                RECT 1118.400 668.240 1125.840 668.560 ;
                RECT 0.160 669.600 202.760 669.920 ;
                RECT 1118.400 669.600 1125.840 669.920 ;
                RECT 0.160 670.960 181.000 671.280 ;
                RECT 192.240 670.960 202.760 671.280 ;
                RECT 1118.400 670.960 1125.840 671.280 ;
                RECT 0.160 672.320 181.000 672.640 ;
                RECT 192.240 672.320 202.760 672.640 ;
                RECT 1118.400 672.320 1125.840 672.640 ;
                RECT 0.160 673.680 181.000 674.000 ;
                RECT 192.240 673.680 202.760 674.000 ;
                RECT 1118.400 673.680 1125.840 674.000 ;
                RECT 0.160 675.040 188.480 675.360 ;
                RECT 192.240 675.040 202.760 675.360 ;
                RECT 1118.400 675.040 1125.840 675.360 ;
                RECT 0.160 676.400 202.760 676.720 ;
                RECT 1118.400 676.400 1125.840 676.720 ;
                RECT 0.160 677.760 202.760 678.080 ;
                RECT 1118.400 677.760 1125.840 678.080 ;
                RECT 0.160 679.120 181.000 679.440 ;
                RECT 192.240 679.120 202.760 679.440 ;
                RECT 1118.400 679.120 1125.840 679.440 ;
                RECT 0.160 680.480 181.000 680.800 ;
                RECT 192.240 680.480 202.760 680.800 ;
                RECT 1118.400 680.480 1125.840 680.800 ;
                RECT 0.160 681.840 181.000 682.160 ;
                RECT 192.240 681.840 202.760 682.160 ;
                RECT 1118.400 681.840 1125.840 682.160 ;
                RECT 0.160 683.200 181.000 683.520 ;
                RECT 192.240 683.200 202.760 683.520 ;
                RECT 1118.400 683.200 1125.840 683.520 ;
                RECT 0.160 684.560 202.760 684.880 ;
                RECT 1118.400 684.560 1125.840 684.880 ;
                RECT 0.160 685.920 183.040 686.240 ;
                RECT 192.240 685.920 202.760 686.240 ;
                RECT 1118.400 685.920 1125.840 686.240 ;
                RECT 0.160 687.280 181.680 687.600 ;
                RECT 192.240 687.280 202.760 687.600 ;
                RECT 1118.400 687.280 1125.840 687.600 ;
                RECT 0.160 688.640 181.680 688.960 ;
                RECT 192.240 688.640 202.760 688.960 ;
                RECT 1118.400 688.640 1125.840 688.960 ;
                RECT 0.160 690.000 181.680 690.320 ;
                RECT 192.240 690.000 202.760 690.320 ;
                RECT 1118.400 690.000 1125.840 690.320 ;
                RECT 0.160 691.360 181.680 691.680 ;
                RECT 192.240 691.360 202.760 691.680 ;
                RECT 1118.400 691.360 1125.840 691.680 ;
                RECT 0.160 692.720 202.760 693.040 ;
                RECT 1118.400 692.720 1125.840 693.040 ;
                RECT 0.160 694.080 181.680 694.400 ;
                RECT 192.240 694.080 202.760 694.400 ;
                RECT 1118.400 694.080 1125.840 694.400 ;
                RECT 0.160 695.440 185.080 695.760 ;
                RECT 192.240 695.440 202.760 695.760 ;
                RECT 1118.400 695.440 1125.840 695.760 ;
                RECT 0.160 696.800 181.680 697.120 ;
                RECT 192.240 696.800 202.760 697.120 ;
                RECT 1118.400 696.800 1125.840 697.120 ;
                RECT 0.160 698.160 181.680 698.480 ;
                RECT 192.240 698.160 202.760 698.480 ;
                RECT 1118.400 698.160 1125.840 698.480 ;
                RECT 0.160 699.520 181.680 699.840 ;
                RECT 192.240 699.520 202.760 699.840 ;
                RECT 1118.400 699.520 1125.840 699.840 ;
                RECT 0.160 700.880 202.760 701.200 ;
                RECT 1118.400 700.880 1125.840 701.200 ;
                RECT 0.160 702.240 181.680 702.560 ;
                RECT 192.240 702.240 202.760 702.560 ;
                RECT 1118.400 702.240 1125.840 702.560 ;
                RECT 0.160 703.600 181.680 703.920 ;
                RECT 192.240 703.600 202.760 703.920 ;
                RECT 1118.400 703.600 1125.840 703.920 ;
                RECT 0.160 704.960 187.800 705.280 ;
                RECT 192.240 704.960 202.760 705.280 ;
                RECT 1118.400 704.960 1125.840 705.280 ;
                RECT 0.160 706.320 181.680 706.640 ;
                RECT 192.240 706.320 202.760 706.640 ;
                RECT 1118.400 706.320 1125.840 706.640 ;
                RECT 0.160 707.680 181.680 708.000 ;
                RECT 192.240 707.680 202.760 708.000 ;
                RECT 1118.400 707.680 1125.840 708.000 ;
                RECT 0.160 709.040 202.760 709.360 ;
                RECT 1118.400 709.040 1125.840 709.360 ;
                RECT 0.160 710.400 181.680 710.720 ;
                RECT 192.240 710.400 202.760 710.720 ;
                RECT 1118.400 710.400 1125.840 710.720 ;
                RECT 0.160 711.760 181.680 712.080 ;
                RECT 192.240 711.760 202.760 712.080 ;
                RECT 1118.400 711.760 1125.840 712.080 ;
                RECT 0.160 713.120 181.680 713.440 ;
                RECT 192.240 713.120 202.760 713.440 ;
                RECT 1118.400 713.120 1125.840 713.440 ;
                RECT 0.160 714.480 190.520 714.800 ;
                RECT 192.240 714.480 202.760 714.800 ;
                RECT 1118.400 714.480 1125.840 714.800 ;
                RECT 0.160 715.840 181.680 716.160 ;
                RECT 192.240 715.840 202.760 716.160 ;
                RECT 1118.400 715.840 1125.840 716.160 ;
                RECT 0.160 717.200 202.760 717.520 ;
                RECT 1118.400 717.200 1125.840 717.520 ;
                RECT 0.160 718.560 182.360 718.880 ;
                RECT 192.240 718.560 202.760 718.880 ;
                RECT 1118.400 718.560 1125.840 718.880 ;
                RECT 0.160 719.920 182.360 720.240 ;
                RECT 192.240 719.920 202.760 720.240 ;
                RECT 1118.400 719.920 1125.840 720.240 ;
                RECT 0.160 721.280 182.360 721.600 ;
                RECT 192.240 721.280 202.760 721.600 ;
                RECT 1118.400 721.280 1125.840 721.600 ;
                RECT 0.160 722.640 182.360 722.960 ;
                RECT 192.240 722.640 202.760 722.960 ;
                RECT 1118.400 722.640 1125.840 722.960 ;
                RECT 0.160 724.000 202.760 724.320 ;
                RECT 1118.400 724.000 1125.840 724.320 ;
                RECT 0.160 725.360 185.080 725.680 ;
                RECT 192.240 725.360 202.760 725.680 ;
                RECT 1118.400 725.360 1125.840 725.680 ;
                RECT 0.160 726.720 182.360 727.040 ;
                RECT 192.240 726.720 202.760 727.040 ;
                RECT 1118.400 726.720 1125.840 727.040 ;
                RECT 0.160 728.080 182.360 728.400 ;
                RECT 192.240 728.080 202.760 728.400 ;
                RECT 1118.400 728.080 1125.840 728.400 ;
                RECT 0.160 729.440 182.360 729.760 ;
                RECT 192.240 729.440 202.760 729.760 ;
                RECT 1118.400 729.440 1125.840 729.760 ;
                RECT 0.160 730.800 182.360 731.120 ;
                RECT 192.240 730.800 202.760 731.120 ;
                RECT 1118.400 730.800 1125.840 731.120 ;
                RECT 0.160 732.160 202.760 732.480 ;
                RECT 1118.400 732.160 1125.840 732.480 ;
                RECT 0.160 733.520 187.120 733.840 ;
                RECT 192.240 733.520 202.760 733.840 ;
                RECT 1118.400 733.520 1125.840 733.840 ;
                RECT 0.160 734.880 187.120 735.200 ;
                RECT 192.240 734.880 202.760 735.200 ;
                RECT 1118.400 734.880 1125.840 735.200 ;
                RECT 0.160 736.240 182.360 736.560 ;
                RECT 192.240 736.240 202.760 736.560 ;
                RECT 1118.400 736.240 1125.840 736.560 ;
                RECT 0.160 737.600 182.360 737.920 ;
                RECT 192.240 737.600 202.760 737.920 ;
                RECT 1118.400 737.600 1125.840 737.920 ;
                RECT 0.160 738.960 182.360 739.280 ;
                RECT 192.240 738.960 202.760 739.280 ;
                RECT 1118.400 738.960 1125.840 739.280 ;
                RECT 0.160 740.320 202.760 740.640 ;
                RECT 1118.400 740.320 1125.840 740.640 ;
                RECT 0.160 741.680 182.360 742.000 ;
                RECT 192.240 741.680 202.760 742.000 ;
                RECT 1118.400 741.680 1125.840 742.000 ;
                RECT 0.160 743.040 182.360 743.360 ;
                RECT 192.240 743.040 202.760 743.360 ;
                RECT 1118.400 743.040 1125.840 743.360 ;
                RECT 0.160 744.400 189.840 744.720 ;
                RECT 192.240 744.400 202.760 744.720 ;
                RECT 1118.400 744.400 1125.840 744.720 ;
                RECT 0.160 745.760 182.360 746.080 ;
                RECT 192.240 745.760 202.760 746.080 ;
                RECT 1118.400 745.760 1125.840 746.080 ;
                RECT 0.160 747.120 182.360 747.440 ;
                RECT 192.240 747.120 202.760 747.440 ;
                RECT 1118.400 747.120 1125.840 747.440 ;
                RECT 0.160 748.480 202.760 748.800 ;
                RECT 1118.400 748.480 1125.840 748.800 ;
                RECT 0.160 749.840 182.360 750.160 ;
                RECT 192.240 749.840 202.760 750.160 ;
                RECT 1118.400 749.840 1125.840 750.160 ;
                RECT 0.160 751.200 182.360 751.520 ;
                RECT 192.240 751.200 202.760 751.520 ;
                RECT 1118.400 751.200 1125.840 751.520 ;
                RECT 0.160 752.560 182.360 752.880 ;
                RECT 192.240 752.560 202.760 752.880 ;
                RECT 1118.400 752.560 1125.840 752.880 ;
                RECT 0.160 753.920 184.400 754.240 ;
                RECT 192.240 753.920 202.760 754.240 ;
                RECT 1118.400 753.920 1125.840 754.240 ;
                RECT 0.160 755.280 182.360 755.600 ;
                RECT 192.240 755.280 202.760 755.600 ;
                RECT 1118.400 755.280 1125.840 755.600 ;
                RECT 0.160 756.640 202.760 756.960 ;
                RECT 1118.400 756.640 1125.840 756.960 ;
                RECT 0.160 758.000 182.360 758.320 ;
                RECT 192.240 758.000 202.760 758.320 ;
                RECT 1118.400 758.000 1125.840 758.320 ;
                RECT 0.160 759.360 182.360 759.680 ;
                RECT 192.240 759.360 202.760 759.680 ;
                RECT 1118.400 759.360 1125.840 759.680 ;
                RECT 0.160 760.720 182.360 761.040 ;
                RECT 192.240 760.720 202.760 761.040 ;
                RECT 1118.400 760.720 1125.840 761.040 ;
                RECT 0.160 762.080 182.360 762.400 ;
                RECT 192.240 762.080 202.760 762.400 ;
                RECT 1118.400 762.080 1125.840 762.400 ;
                RECT 0.160 763.440 202.760 763.760 ;
                RECT 1118.400 763.440 1125.840 763.760 ;
                RECT 0.160 764.800 187.120 765.120 ;
                RECT 192.240 764.800 202.760 765.120 ;
                RECT 1118.400 764.800 1125.840 765.120 ;
                RECT 0.160 766.160 182.360 766.480 ;
                RECT 192.240 766.160 202.760 766.480 ;
                RECT 1118.400 766.160 1125.840 766.480 ;
                RECT 0.160 767.520 182.360 767.840 ;
                RECT 192.240 767.520 202.760 767.840 ;
                RECT 1118.400 767.520 1125.840 767.840 ;
                RECT 0.160 768.880 182.360 769.200 ;
                RECT 192.240 768.880 202.760 769.200 ;
                RECT 1118.400 768.880 1125.840 769.200 ;
                RECT 0.160 770.240 182.360 770.560 ;
                RECT 192.240 770.240 202.760 770.560 ;
                RECT 1118.400 770.240 1125.840 770.560 ;
                RECT 0.160 771.600 202.760 771.920 ;
                RECT 1118.400 771.600 1125.840 771.920 ;
                RECT 0.160 772.960 188.480 773.280 ;
                RECT 192.240 772.960 202.760 773.280 ;
                RECT 1118.400 772.960 1125.840 773.280 ;
                RECT 0.160 774.320 182.360 774.640 ;
                RECT 192.240 774.320 202.760 774.640 ;
                RECT 1118.400 774.320 1125.840 774.640 ;
                RECT 0.160 775.680 182.360 776.000 ;
                RECT 192.240 775.680 202.760 776.000 ;
                RECT 1118.400 775.680 1125.840 776.000 ;
                RECT 0.160 777.040 182.360 777.360 ;
                RECT 192.240 777.040 202.760 777.360 ;
                RECT 1118.400 777.040 1125.840 777.360 ;
                RECT 0.160 778.400 182.360 778.720 ;
                RECT 192.240 778.400 202.760 778.720 ;
                RECT 1118.400 778.400 1125.840 778.720 ;
                RECT 0.160 779.760 202.760 780.080 ;
                RECT 1118.400 779.760 1125.840 780.080 ;
                RECT 0.160 781.120 401.320 781.440 ;
                RECT 1118.400 781.120 1125.840 781.440 ;
                RECT 0.160 782.480 401.320 782.800 ;
                RECT 1118.400 782.480 1125.840 782.800 ;
                RECT 0.160 783.840 401.320 784.160 ;
                RECT 1118.400 783.840 1125.840 784.160 ;
                RECT 0.160 785.200 1125.840 785.520 ;
                RECT 0.160 786.560 1125.840 786.880 ;
                RECT 0.160 787.920 1125.840 788.240 ;
                RECT 0.160 789.280 1125.840 789.600 ;
                RECT 0.160 790.640 1125.840 790.960 ;
                RECT 0.160 0.160 1125.840 1.520 ;
                RECT 0.160 794.680 1125.840 796.040 ;
                RECT 405.460 34.830 411.260 36.200 ;
                RECT 1108.560 34.830 1114.360 36.200 ;
                RECT 405.460 40.085 411.260 41.635 ;
                RECT 1108.560 40.085 1114.360 41.635 ;
                RECT 405.460 45.940 411.260 47.740 ;
                RECT 1108.560 45.940 1114.360 47.740 ;
                RECT 405.460 51.470 411.260 52.720 ;
                RECT 1108.560 51.470 1114.360 52.720 ;
                RECT 405.460 56.230 411.260 57.520 ;
                RECT 1108.560 56.230 1114.360 57.520 ;
                RECT 405.460 61.050 411.260 62.340 ;
                RECT 1108.560 61.050 1114.360 62.340 ;
                RECT 405.460 168.125 1114.360 169.925 ;
                RECT 405.460 69.000 1114.360 70.800 ;
                RECT 405.460 106.170 1114.360 109.770 ;
                RECT 405.460 88.370 1114.360 89.170 ;
                RECT 405.460 83.480 1114.360 84.280 ;
                RECT 405.460 115.975 1114.360 116.265 ;
                RECT 405.460 247.965 1114.360 251.565 ;
                RECT 405.460 80.470 1114.360 81.270 ;
                RECT 405.460 19.075 1114.360 20.875 ;
                RECT 207.660 273.555 209.580 780.735 ;
                RECT 211.500 273.555 213.420 780.735 ;
                RECT 223.910 273.555 225.830 780.735 ;
                RECT 227.750 273.555 229.670 780.735 ;
                RECT 231.590 273.555 233.510 780.735 ;
                RECT 235.430 273.555 237.350 780.735 ;
                RECT 256.115 273.555 258.035 780.735 ;
                RECT 259.955 273.555 261.875 780.735 ;
                RECT 263.795 273.555 265.715 780.735 ;
                RECT 267.635 273.555 269.555 780.735 ;
                RECT 271.475 273.555 273.395 780.735 ;
                RECT 275.315 273.555 277.235 780.735 ;
                RECT 279.155 273.555 281.075 780.735 ;
                RECT 282.995 273.555 284.915 780.735 ;
                RECT 286.835 273.555 288.755 780.735 ;
                RECT 324.315 273.555 326.235 780.735 ;
                RECT 328.155 273.555 330.075 780.735 ;
                RECT 331.995 273.555 333.915 780.735 ;
                RECT 335.835 273.555 337.755 780.735 ;
                RECT 339.675 273.555 341.595 780.735 ;
                RECT 343.515 273.555 345.435 780.735 ;
                RECT 347.355 273.555 349.275 780.735 ;
                RECT 351.195 273.555 353.115 780.735 ;
                RECT 355.035 273.555 356.955 780.735 ;
                RECT 358.875 273.555 360.795 780.735 ;
                RECT 362.715 273.555 364.635 780.735 ;
                RECT 366.555 273.555 368.475 780.735 ;
                RECT 370.395 273.555 372.315 780.735 ;
                RECT 374.235 273.555 376.155 780.735 ;
                RECT 378.075 273.555 379.995 780.735 ;
                RECT 381.915 273.555 383.835 780.735 ;
                RECT 385.755 273.555 387.675 780.735 ;
                RECT 389.595 273.555 391.515 780.735 ;
                RECT 393.435 273.555 395.355 780.735 ;
                RECT 397.275 273.555 399.195 780.735 ;
                RECT 128.265 57.175 130.015 126.975 ;
                RECT 134.725 57.175 136.645 126.975 ;
                RECT 141.485 57.175 143.405 126.975 ;
                RECT 150.195 57.175 152.115 126.975 ;
                RECT 154.035 57.175 155.955 126.975 ;
                RECT 166.875 57.175 168.795 126.975 ;
                RECT 170.715 57.175 172.635 126.975 ;
                RECT 174.555 57.175 176.475 126.975 ;
                RECT 178.395 57.175 180.315 126.975 ;
                RECT 199.295 57.175 201.215 126.975 ;
                RECT 203.135 57.175 205.055 126.975 ;
                RECT 206.975 57.175 208.895 126.975 ;
                RECT 210.815 57.175 212.735 126.975 ;
                RECT 214.655 57.175 216.575 126.975 ;
                RECT 218.495 57.175 220.415 126.975 ;
                RECT 222.335 57.175 224.255 126.975 ;
                RECT 226.175 57.175 228.095 126.975 ;
                RECT 230.015 57.175 231.935 126.975 ;
                RECT 269.445 57.175 271.365 126.975 ;
                RECT 273.285 57.175 275.205 126.975 ;
                RECT 277.125 57.175 279.045 126.975 ;
                RECT 280.965 57.175 282.885 126.975 ;
                RECT 284.805 57.175 286.725 126.975 ;
                RECT 288.645 57.175 290.565 126.975 ;
                RECT 292.485 57.175 294.405 126.975 ;
                RECT 296.325 57.175 298.245 126.975 ;
                RECT 300.165 57.175 302.085 126.975 ;
                RECT 304.005 57.175 305.925 126.975 ;
                RECT 307.845 57.175 309.765 126.975 ;
                RECT 311.685 57.175 313.605 126.975 ;
                RECT 315.525 57.175 317.445 126.975 ;
                RECT 319.365 57.175 321.285 126.975 ;
                RECT 323.205 57.175 325.125 126.975 ;
                RECT 327.045 57.175 328.965 126.975 ;
                RECT 330.885 57.175 332.805 126.975 ;
                RECT 334.725 57.175 336.645 126.975 ;
                RECT 338.565 57.175 340.485 126.975 ;
                RECT 342.405 57.175 344.325 126.975 ;
                RECT 346.245 57.175 348.165 126.975 ;
                RECT 223.405 208.940 225.325 266.920 ;
                RECT 230.595 208.940 232.515 266.920 ;
                RECT 237.225 208.940 238.975 266.920 ;
                RECT 243.555 208.940 245.305 266.920 ;
                RECT 252.810 208.940 254.730 266.920 ;
                RECT 267.785 208.940 269.705 266.920 ;
                RECT 271.625 208.940 273.545 266.920 ;
                RECT 275.465 208.940 277.385 266.920 ;
                RECT 279.305 208.940 281.225 266.920 ;
                RECT 304.550 208.940 306.470 266.920 ;
                RECT 308.390 208.940 310.310 266.920 ;
                RECT 312.230 208.940 314.150 266.920 ;
                RECT 316.070 208.940 317.990 266.920 ;
                RECT 319.910 208.940 321.830 266.920 ;
                RECT 323.750 208.940 325.670 266.920 ;
                RECT 327.590 208.940 329.510 266.920 ;
                RECT 331.430 208.940 333.350 266.920 ;
                RECT 335.270 208.940 337.190 266.920 ;
                RECT 339.110 208.940 341.030 266.920 ;
                RECT 342.950 208.940 344.870 266.920 ;
                RECT 346.790 208.940 348.710 266.920 ;
                RECT 277.405 197.780 279.155 202.940 ;
                RECT 287.965 197.780 289.885 202.940 ;
                RECT 291.805 197.780 293.725 202.940 ;
                RECT 314.825 197.780 316.745 202.940 ;
                RECT 318.665 197.780 320.585 202.940 ;
                RECT 322.505 197.780 324.425 202.940 ;
                RECT 326.345 197.780 328.265 202.940 ;
                RECT 330.185 197.780 332.105 202.940 ;
                RECT 334.025 197.780 335.945 202.940 ;
                RECT 337.865 197.780 339.785 202.940 ;
                RECT 341.705 197.780 343.625 202.940 ;
                RECT 345.545 197.780 347.465 202.940 ;
                RECT 347.255 46.015 349.005 51.175 ;
                RECT 124.420 275.825 133.580 276.575 ;
                RECT 124.420 281.225 133.580 283.145 ;
                RECT 65.780 261.835 81.820 263.485 ;
                RECT 44.180 261.965 63.820 265.565 ;
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 416.960 5.560 ;
                RECT 418.680 5.240 427.840 5.560 ;
                RECT 429.560 5.240 438.720 5.560 ;
                RECT 440.440 5.240 449.600 5.560 ;
                RECT 451.320 5.240 460.480 5.560 ;
                RECT 462.200 5.240 471.360 5.560 ;
                RECT 473.080 5.240 482.240 5.560 ;
                RECT 483.960 5.240 493.120 5.560 ;
                RECT 494.840 5.240 504.000 5.560 ;
                RECT 505.720 5.240 514.880 5.560 ;
                RECT 516.600 5.240 525.760 5.560 ;
                RECT 527.480 5.240 536.640 5.560 ;
                RECT 538.360 5.240 547.520 5.560 ;
                RECT 549.240 5.240 558.400 5.560 ;
                RECT 560.120 5.240 569.280 5.560 ;
                RECT 571.000 5.240 580.160 5.560 ;
                RECT 581.880 5.240 591.040 5.560 ;
                RECT 592.760 5.240 601.920 5.560 ;
                RECT 603.640 5.240 612.800 5.560 ;
                RECT 614.520 5.240 624.360 5.560 ;
                RECT 625.400 5.240 635.240 5.560 ;
                RECT 636.280 5.240 646.120 5.560 ;
                RECT 647.160 5.240 657.000 5.560 ;
                RECT 658.040 5.240 667.880 5.560 ;
                RECT 668.920 5.240 678.760 5.560 ;
                RECT 679.800 5.240 689.640 5.560 ;
                RECT 690.680 5.240 700.520 5.560 ;
                RECT 701.560 5.240 711.400 5.560 ;
                RECT 712.440 5.240 722.280 5.560 ;
                RECT 724.000 5.240 733.160 5.560 ;
                RECT 734.880 5.240 744.040 5.560 ;
                RECT 745.760 5.240 754.920 5.560 ;
                RECT 756.640 5.240 765.800 5.560 ;
                RECT 767.520 5.240 776.680 5.560 ;
                RECT 778.400 5.240 787.560 5.560 ;
                RECT 789.280 5.240 798.440 5.560 ;
                RECT 800.160 5.240 809.320 5.560 ;
                RECT 811.040 5.240 820.200 5.560 ;
                RECT 821.920 5.240 831.080 5.560 ;
                RECT 832.800 5.240 841.960 5.560 ;
                RECT 843.680 5.240 852.840 5.560 ;
                RECT 854.560 5.240 863.720 5.560 ;
                RECT 865.440 5.240 874.600 5.560 ;
                RECT 876.320 5.240 885.480 5.560 ;
                RECT 887.200 5.240 896.360 5.560 ;
                RECT 898.080 5.240 907.240 5.560 ;
                RECT 908.960 5.240 918.120 5.560 ;
                RECT 919.840 5.240 929.000 5.560 ;
                RECT 930.720 5.240 939.880 5.560 ;
                RECT 941.600 5.240 950.760 5.560 ;
                RECT 952.480 5.240 961.640 5.560 ;
                RECT 963.360 5.240 972.520 5.560 ;
                RECT 974.240 5.240 983.400 5.560 ;
                RECT 985.120 5.240 994.960 5.560 ;
                RECT 996.000 5.240 1005.840 5.560 ;
                RECT 1006.880 5.240 1016.720 5.560 ;
                RECT 1017.760 5.240 1027.600 5.560 ;
                RECT 1028.640 5.240 1038.480 5.560 ;
                RECT 1039.520 5.240 1049.360 5.560 ;
                RECT 1050.400 5.240 1060.240 5.560 ;
                RECT 1061.280 5.240 1071.120 5.560 ;
                RECT 1072.160 5.240 1082.000 5.560 ;
                RECT 1083.040 5.240 1092.880 5.560 ;
                RECT 1094.600 5.240 1103.760 5.560 ;
                RECT 1105.480 5.240 1123.120 5.560 ;
                RECT 2.880 6.600 1123.120 6.920 ;
                RECT 2.880 7.960 1123.120 8.280 ;
                RECT 2.880 9.320 351.000 9.640 ;
                RECT 409.840 9.320 1123.120 9.640 ;
                RECT 2.880 10.680 1123.120 11.000 ;
                RECT 2.880 12.040 1123.120 12.360 ;
                RECT 2.880 13.400 270.080 13.720 ;
                RECT 352.040 13.400 404.040 13.720 ;
                RECT 1116.360 13.400 1123.120 13.720 ;
                RECT 2.880 14.760 404.040 15.080 ;
                RECT 1116.360 14.760 1123.120 15.080 ;
                RECT 2.880 16.120 404.040 16.440 ;
                RECT 1116.360 16.120 1123.120 16.440 ;
                RECT 2.880 17.480 270.080 17.800 ;
                RECT 351.360 17.480 404.040 17.800 ;
                RECT 1116.360 17.480 1123.120 17.800 ;
                RECT 2.880 18.840 404.040 19.160 ;
                RECT 1116.360 18.840 1123.120 19.160 ;
                RECT 2.880 20.200 404.040 20.520 ;
                RECT 1116.360 20.200 1123.120 20.520 ;
                RECT 2.880 21.560 404.040 21.880 ;
                RECT 1116.360 21.560 1123.120 21.880 ;
                RECT 2.880 22.920 404.040 23.240 ;
                RECT 1116.360 22.920 1123.120 23.240 ;
                RECT 2.880 24.280 404.040 24.600 ;
                RECT 1116.360 24.280 1123.120 24.600 ;
                RECT 2.880 25.640 404.040 25.960 ;
                RECT 1116.360 25.640 1123.120 25.960 ;
                RECT 2.880 27.000 404.040 27.320 ;
                RECT 1116.360 27.000 1123.120 27.320 ;
                RECT 2.880 28.360 404.040 28.680 ;
                RECT 1116.360 28.360 1123.120 28.680 ;
                RECT 2.880 29.720 404.040 30.040 ;
                RECT 1116.360 29.720 1123.120 30.040 ;
                RECT 2.880 31.080 403.360 31.400 ;
                RECT 1116.360 31.080 1123.120 31.400 ;
                RECT 2.880 32.440 404.040 32.760 ;
                RECT 1116.360 32.440 1123.120 32.760 ;
                RECT 2.880 33.800 404.040 34.120 ;
                RECT 1116.360 33.800 1123.120 34.120 ;
                RECT 2.880 35.160 404.040 35.480 ;
                RECT 1116.360 35.160 1123.120 35.480 ;
                RECT 2.880 36.520 113.680 36.840 ;
                RECT 324.160 36.520 404.040 36.840 ;
                RECT 1116.360 36.520 1123.120 36.840 ;
                RECT 2.880 37.880 112.320 38.200 ;
                RECT 330.280 37.880 404.040 38.200 ;
                RECT 1116.360 37.880 1123.120 38.200 ;
                RECT 2.880 39.240 110.960 39.560 ;
                RECT 336.400 39.240 404.040 39.560 ;
                RECT 1116.360 39.240 1123.120 39.560 ;
                RECT 2.880 40.600 87.840 40.920 ;
                RECT 351.360 40.600 404.040 40.920 ;
                RECT 1116.360 40.600 1123.120 40.920 ;
                RECT 2.880 41.960 89.200 42.280 ;
                RECT 341.840 41.960 404.040 42.280 ;
                RECT 1116.360 41.960 1123.120 42.280 ;
                RECT 2.880 43.320 404.040 43.640 ;
                RECT 1116.360 43.320 1123.120 43.640 ;
                RECT 2.880 44.680 404.040 45.000 ;
                RECT 1116.360 44.680 1123.120 45.000 ;
                RECT 2.880 46.040 344.200 46.360 ;
                RECT 350.000 46.040 404.040 46.360 ;
                RECT 1116.360 46.040 1123.120 46.360 ;
                RECT 2.880 47.400 344.200 47.720 ;
                RECT 1116.360 47.400 1123.120 47.720 ;
                RECT 2.880 48.760 344.200 49.080 ;
                RECT 1116.360 48.760 1123.120 49.080 ;
                RECT 2.880 50.120 344.200 50.440 ;
                RECT 350.000 50.120 404.040 50.440 ;
                RECT 1116.360 50.120 1123.120 50.440 ;
                RECT 2.880 51.480 344.200 51.800 ;
                RECT 350.000 51.480 404.040 51.800 ;
                RECT 1116.360 51.480 1123.120 51.800 ;
                RECT 2.880 52.840 404.040 53.160 ;
                RECT 1116.360 52.840 1123.120 53.160 ;
                RECT 2.880 54.200 404.040 54.520 ;
                RECT 1116.360 54.200 1123.120 54.520 ;
                RECT 2.880 55.560 404.040 55.880 ;
                RECT 1116.360 55.560 1123.120 55.880 ;
                RECT 2.880 56.920 125.240 57.240 ;
                RECT 348.640 56.920 404.040 57.240 ;
                RECT 1116.360 56.920 1123.120 57.240 ;
                RECT 2.880 58.280 110.960 58.600 ;
                RECT 118.120 58.280 125.240 58.600 ;
                RECT 348.640 58.280 404.040 58.600 ;
                RECT 1116.360 58.280 1123.120 58.600 ;
                RECT 2.880 59.640 112.320 59.960 ;
                RECT 117.440 59.640 125.240 59.960 ;
                RECT 362.920 59.640 404.040 59.960 ;
                RECT 1116.360 59.640 1123.120 59.960 ;
                RECT 2.880 61.000 113.680 61.320 ;
                RECT 116.080 61.000 125.240 61.320 ;
                RECT 365.640 61.000 404.040 61.320 ;
                RECT 1116.360 61.000 1123.120 61.320 ;
                RECT 2.880 62.360 125.240 62.680 ;
                RECT 365.640 62.360 404.040 62.680 ;
                RECT 1116.360 62.360 1123.120 62.680 ;
                RECT 2.880 63.720 125.240 64.040 ;
                RECT 362.920 63.720 404.040 64.040 ;
                RECT 1116.360 63.720 1123.120 64.040 ;
                RECT 2.880 65.080 125.240 65.400 ;
                RECT 365.640 65.080 404.040 65.400 ;
                RECT 1116.360 65.080 1123.120 65.400 ;
                RECT 2.880 66.440 125.240 66.760 ;
                RECT 348.640 66.440 404.040 66.760 ;
                RECT 1116.360 66.440 1123.120 66.760 ;
                RECT 2.880 67.800 125.240 68.120 ;
                RECT 371.080 67.800 404.040 68.120 ;
                RECT 1116.360 67.800 1123.120 68.120 ;
                RECT 2.880 69.160 125.240 69.480 ;
                RECT 371.080 69.160 404.040 69.480 ;
                RECT 1116.360 69.160 1123.120 69.480 ;
                RECT 2.880 70.520 125.240 70.840 ;
                RECT 368.360 70.520 404.040 70.840 ;
                RECT 1116.360 70.520 1123.120 70.840 ;
                RECT 2.880 71.880 125.240 72.200 ;
                RECT 371.080 71.880 404.040 72.200 ;
                RECT 1116.360 71.880 1123.120 72.200 ;
                RECT 2.880 73.240 125.240 73.560 ;
                RECT 371.080 73.240 404.040 73.560 ;
                RECT 1116.360 73.240 1123.120 73.560 ;
                RECT 2.880 74.600 125.240 74.920 ;
                RECT 348.640 74.600 404.040 74.920 ;
                RECT 1116.360 74.600 1123.120 74.920 ;
                RECT 2.880 75.960 125.240 76.280 ;
                RECT 376.520 75.960 404.040 76.280 ;
                RECT 1116.360 75.960 1123.120 76.280 ;
                RECT 2.880 77.320 125.240 77.640 ;
                RECT 373.800 77.320 404.040 77.640 ;
                RECT 1116.360 77.320 1123.120 77.640 ;
                RECT 2.880 78.680 125.240 79.000 ;
                RECT 376.520 78.680 404.040 79.000 ;
                RECT 1116.360 78.680 1123.120 79.000 ;
                RECT 2.880 80.040 125.240 80.360 ;
                RECT 376.520 80.040 404.040 80.360 ;
                RECT 1116.360 80.040 1123.120 80.360 ;
                RECT 2.880 81.400 125.240 81.720 ;
                RECT 376.520 81.400 404.040 81.720 ;
                RECT 1116.360 81.400 1123.120 81.720 ;
                RECT 2.880 82.760 125.240 83.080 ;
                RECT 373.800 82.760 404.040 83.080 ;
                RECT 1116.360 82.760 1123.120 83.080 ;
                RECT 2.880 84.120 125.240 84.440 ;
                RECT 348.640 84.120 404.040 84.440 ;
                RECT 1116.360 84.120 1123.120 84.440 ;
                RECT 2.880 85.480 125.240 85.800 ;
                RECT 379.240 85.480 404.040 85.800 ;
                RECT 1116.360 85.480 1123.120 85.800 ;
                RECT 2.880 86.840 125.240 87.160 ;
                RECT 381.960 86.840 404.040 87.160 ;
                RECT 1116.360 86.840 1123.120 87.160 ;
                RECT 2.880 88.200 125.240 88.520 ;
                RECT 381.960 88.200 404.040 88.520 ;
                RECT 1116.360 88.200 1123.120 88.520 ;
                RECT 2.880 89.560 125.240 89.880 ;
                RECT 379.240 89.560 404.040 89.880 ;
                RECT 1116.360 89.560 1123.120 89.880 ;
                RECT 2.880 90.920 125.240 91.240 ;
                RECT 381.960 90.920 404.040 91.240 ;
                RECT 1116.360 90.920 1123.120 91.240 ;
                RECT 2.880 92.280 125.240 92.600 ;
                RECT 348.640 92.280 404.040 92.600 ;
                RECT 1116.360 92.280 1123.120 92.600 ;
                RECT 2.880 93.640 125.240 93.960 ;
                RECT 387.400 93.640 404.040 93.960 ;
                RECT 1116.360 93.640 1123.120 93.960 ;
                RECT 2.880 95.000 125.240 95.320 ;
                RECT 387.400 95.000 404.040 95.320 ;
                RECT 1116.360 95.000 1123.120 95.320 ;
                RECT 2.880 96.360 125.240 96.680 ;
                RECT 384.680 96.360 404.040 96.680 ;
                RECT 1116.360 96.360 1123.120 96.680 ;
                RECT 2.880 97.720 125.240 98.040 ;
                RECT 387.400 97.720 404.040 98.040 ;
                RECT 1116.360 97.720 1123.120 98.040 ;
                RECT 2.880 99.080 125.240 99.400 ;
                RECT 387.400 99.080 404.040 99.400 ;
                RECT 1116.360 99.080 1123.120 99.400 ;
                RECT 2.880 100.440 125.240 100.760 ;
                RECT 348.640 100.440 404.040 100.760 ;
                RECT 1116.360 100.440 1123.120 100.760 ;
                RECT 2.880 101.800 125.240 102.120 ;
                RECT 392.840 101.800 404.040 102.120 ;
                RECT 1116.360 101.800 1123.120 102.120 ;
                RECT 2.880 103.160 125.240 103.480 ;
                RECT 390.120 103.160 404.040 103.480 ;
                RECT 1116.360 103.160 1123.120 103.480 ;
                RECT 2.880 104.520 125.240 104.840 ;
                RECT 392.840 104.520 404.040 104.840 ;
                RECT 1116.360 104.520 1123.120 104.840 ;
                RECT 2.880 105.880 125.240 106.200 ;
                RECT 392.840 105.880 404.040 106.200 ;
                RECT 1116.360 105.880 1123.120 106.200 ;
                RECT 2.880 107.240 125.240 107.560 ;
                RECT 392.840 107.240 404.040 107.560 ;
                RECT 1116.360 107.240 1123.120 107.560 ;
                RECT 2.880 108.600 125.240 108.920 ;
                RECT 390.120 108.600 404.040 108.920 ;
                RECT 1116.360 108.600 1123.120 108.920 ;
                RECT 2.880 109.960 125.240 110.280 ;
                RECT 348.640 109.960 404.040 110.280 ;
                RECT 1116.360 109.960 1123.120 110.280 ;
                RECT 2.880 111.320 125.240 111.640 ;
                RECT 395.560 111.320 404.040 111.640 ;
                RECT 1116.360 111.320 1123.120 111.640 ;
                RECT 2.880 112.680 125.240 113.000 ;
                RECT 398.280 112.680 404.040 113.000 ;
                RECT 1116.360 112.680 1123.120 113.000 ;
                RECT 2.880 114.040 125.240 114.360 ;
                RECT 398.280 114.040 404.040 114.360 ;
                RECT 1116.360 114.040 1123.120 114.360 ;
                RECT 2.880 115.400 125.240 115.720 ;
                RECT 395.560 115.400 404.040 115.720 ;
                RECT 1116.360 115.400 1123.120 115.720 ;
                RECT 2.880 116.760 125.240 117.080 ;
                RECT 398.280 116.760 404.040 117.080 ;
                RECT 1116.360 116.760 1123.120 117.080 ;
                RECT 2.880 118.120 125.240 118.440 ;
                RECT 348.640 118.120 404.040 118.440 ;
                RECT 1116.360 118.120 1123.120 118.440 ;
                RECT 2.880 119.480 125.240 119.800 ;
                RECT 1116.360 119.480 1123.120 119.800 ;
                RECT 2.880 120.840 125.240 121.160 ;
                RECT 1116.360 120.840 1123.120 121.160 ;
                RECT 2.880 122.200 125.240 122.520 ;
                RECT 401.000 122.200 404.040 122.520 ;
                RECT 1116.360 122.200 1123.120 122.520 ;
                RECT 2.880 123.560 125.240 123.880 ;
                RECT 1116.360 123.560 1123.120 123.880 ;
                RECT 2.880 124.920 125.240 125.240 ;
                RECT 1116.360 124.920 1123.120 125.240 ;
                RECT 2.880 126.280 125.240 126.600 ;
                RECT 348.640 126.280 404.040 126.600 ;
                RECT 1116.360 126.280 1123.120 126.600 ;
                RECT 2.880 127.640 404.040 127.960 ;
                RECT 1116.360 127.640 1123.120 127.960 ;
                RECT 2.880 129.000 404.040 129.320 ;
                RECT 1116.360 129.000 1123.120 129.320 ;
                RECT 2.880 130.360 357.120 130.680 ;
                RECT 1116.360 130.360 1123.120 130.680 ;
                RECT 2.880 131.720 397.920 132.040 ;
                RECT 1116.360 131.720 1123.120 132.040 ;
                RECT 2.880 133.080 397.920 133.400 ;
                RECT 1116.360 133.080 1123.120 133.400 ;
                RECT 2.880 134.440 392.480 134.760 ;
                RECT 1116.360 134.440 1123.120 134.760 ;
                RECT 2.880 135.800 392.480 136.120 ;
                RECT 1116.360 135.800 1123.120 136.120 ;
                RECT 2.880 137.160 387.040 137.480 ;
                RECT 1116.360 137.160 1123.120 137.480 ;
                RECT 2.880 138.520 387.040 138.840 ;
                RECT 1116.360 138.520 1123.120 138.840 ;
                RECT 2.880 139.880 381.600 140.200 ;
                RECT 1116.360 139.880 1123.120 140.200 ;
                RECT 2.880 141.240 381.600 141.560 ;
                RECT 1116.360 141.240 1123.120 141.560 ;
                RECT 2.880 142.600 376.160 142.920 ;
                RECT 1116.360 142.600 1123.120 142.920 ;
                RECT 2.880 143.960 376.160 144.280 ;
                RECT 1116.360 143.960 1123.120 144.280 ;
                RECT 2.880 145.320 376.160 145.640 ;
                RECT 1116.360 145.320 1123.120 145.640 ;
                RECT 2.880 146.680 370.720 147.000 ;
                RECT 1116.360 146.680 1123.120 147.000 ;
                RECT 2.880 148.040 86.480 148.360 ;
                RECT 97.040 148.040 370.720 148.360 ;
                RECT 1116.360 148.040 1123.120 148.360 ;
                RECT 2.880 149.400 87.840 149.720 ;
                RECT 90.920 149.400 365.280 149.720 ;
                RECT 1116.360 149.400 1123.120 149.720 ;
                RECT 2.880 150.760 89.200 151.080 ;
                RECT 93.640 150.760 100.760 151.080 ;
                RECT 103.840 150.760 365.280 151.080 ;
                RECT 1116.360 150.760 1123.120 151.080 ;
                RECT 2.880 152.120 359.840 152.440 ;
                RECT 1116.360 152.120 1123.120 152.440 ;
                RECT 2.880 153.480 95.320 153.800 ;
                RECT 103.840 153.480 359.840 153.800 ;
                RECT 1116.360 153.480 1123.120 153.800 ;
                RECT 2.880 154.840 87.840 155.160 ;
                RECT 97.040 154.840 404.040 155.160 ;
                RECT 1116.360 154.840 1123.120 155.160 ;
                RECT 2.880 156.200 91.920 156.520 ;
                RECT 97.040 156.200 404.040 156.520 ;
                RECT 1116.360 156.200 1123.120 156.520 ;
                RECT 2.880 157.560 404.040 157.880 ;
                RECT 1116.360 157.560 1123.120 157.880 ;
                RECT 2.880 158.920 87.840 159.240 ;
                RECT 97.040 158.920 404.040 159.240 ;
                RECT 1116.360 158.920 1123.120 159.240 ;
                RECT 2.880 160.280 95.320 160.600 ;
                RECT 103.160 160.280 404.040 160.600 ;
                RECT 1116.360 160.280 1123.120 160.600 ;
                RECT 2.880 161.640 94.640 161.960 ;
                RECT 97.040 161.640 404.040 161.960 ;
                RECT 1116.360 161.640 1123.120 161.960 ;
                RECT 2.880 163.000 404.040 163.320 ;
                RECT 1116.360 163.000 1123.120 163.320 ;
                RECT 2.880 164.360 95.320 164.680 ;
                RECT 103.840 164.360 404.040 164.680 ;
                RECT 1116.360 164.360 1123.120 164.680 ;
                RECT 2.880 165.720 92.600 166.040 ;
                RECT 97.040 165.720 404.040 166.040 ;
                RECT 1116.360 165.720 1123.120 166.040 ;
                RECT 2.880 167.080 94.640 167.400 ;
                RECT 97.040 167.080 404.040 167.400 ;
                RECT 1116.360 167.080 1123.120 167.400 ;
                RECT 2.880 168.440 98.040 168.760 ;
                RECT 108.600 168.440 404.040 168.760 ;
                RECT 1116.360 168.440 1123.120 168.760 ;
                RECT 2.880 169.800 85.800 170.120 ;
                RECT 103.840 169.800 404.040 170.120 ;
                RECT 1116.360 169.800 1123.120 170.120 ;
                RECT 2.880 171.160 94.640 171.480 ;
                RECT 97.040 171.160 102.800 171.480 ;
                RECT 109.960 171.160 404.040 171.480 ;
                RECT 1116.360 171.160 1123.120 171.480 ;
                RECT 2.880 172.520 106.880 172.840 ;
                RECT 110.640 172.520 404.040 172.840 ;
                RECT 1116.360 172.520 1123.120 172.840 ;
                RECT 2.880 173.880 86.480 174.200 ;
                RECT 99.760 173.880 404.040 174.200 ;
                RECT 1116.360 173.880 1123.120 174.200 ;
                RECT 2.880 175.240 95.320 175.560 ;
                RECT 103.840 175.240 404.040 175.560 ;
                RECT 1116.360 175.240 1123.120 175.560 ;
                RECT 2.880 176.600 92.600 176.920 ;
                RECT 103.840 176.600 404.040 176.920 ;
                RECT 1116.360 176.600 1123.120 176.920 ;
                RECT 2.880 177.960 64.720 178.280 ;
                RECT 82.760 177.960 404.040 178.280 ;
                RECT 1116.360 177.960 1123.120 178.280 ;
                RECT 2.880 179.320 64.720 179.640 ;
                RECT 82.760 179.320 88.520 179.640 ;
                RECT 90.920 179.320 404.040 179.640 ;
                RECT 1116.360 179.320 1123.120 179.640 ;
                RECT 2.880 180.680 64.720 181.000 ;
                RECT 82.760 180.680 92.600 181.000 ;
                RECT 97.040 180.680 404.040 181.000 ;
                RECT 1116.360 180.680 1123.120 181.000 ;
                RECT 2.880 182.040 64.720 182.360 ;
                RECT 82.760 182.040 404.040 182.360 ;
                RECT 1116.360 182.040 1123.120 182.360 ;
                RECT 2.880 183.400 64.720 183.720 ;
                RECT 82.760 183.400 404.040 183.720 ;
                RECT 1116.360 183.400 1123.120 183.720 ;
                RECT 2.880 184.760 64.720 185.080 ;
                RECT 82.760 184.760 94.640 185.080 ;
                RECT 97.040 184.760 404.040 185.080 ;
                RECT 1116.360 184.760 1123.120 185.080 ;
                RECT 2.880 186.120 64.720 186.440 ;
                RECT 82.760 186.120 95.320 186.440 ;
                RECT 97.720 186.120 404.040 186.440 ;
                RECT 1116.360 186.120 1123.120 186.440 ;
                RECT 2.880 187.480 64.720 187.800 ;
                RECT 82.760 187.480 94.640 187.800 ;
                RECT 97.040 187.480 404.040 187.800 ;
                RECT 1116.360 187.480 1123.120 187.800 ;
                RECT 2.880 188.840 64.720 189.160 ;
                RECT 82.760 188.840 404.040 189.160 ;
                RECT 1116.360 188.840 1123.120 189.160 ;
                RECT 2.880 190.200 64.720 190.520 ;
                RECT 82.760 190.200 85.120 190.520 ;
                RECT 97.040 190.200 404.040 190.520 ;
                RECT 1116.360 190.200 1123.120 190.520 ;
                RECT 2.880 191.560 64.720 191.880 ;
                RECT 82.760 191.560 95.320 191.880 ;
                RECT 97.720 191.560 404.040 191.880 ;
                RECT 1116.360 191.560 1123.120 191.880 ;
                RECT 2.880 192.920 64.720 193.240 ;
                RECT 82.760 192.920 404.040 193.240 ;
                RECT 1116.360 192.920 1123.120 193.240 ;
                RECT 2.880 194.280 64.720 194.600 ;
                RECT 82.760 194.280 404.040 194.600 ;
                RECT 1116.360 194.280 1123.120 194.600 ;
                RECT 2.880 195.640 64.720 195.960 ;
                RECT 96.360 195.640 404.040 195.960 ;
                RECT 1116.360 195.640 1123.120 195.960 ;
                RECT 2.880 197.000 64.720 197.320 ;
                RECT 82.760 197.000 92.600 197.320 ;
                RECT 99.760 197.000 404.040 197.320 ;
                RECT 1116.360 197.000 1123.120 197.320 ;
                RECT 2.880 198.360 64.720 198.680 ;
                RECT 82.760 198.360 109.600 198.680 ;
                RECT 347.960 198.360 404.040 198.680 ;
                RECT 1116.360 198.360 1123.120 198.680 ;
                RECT 2.880 199.720 64.720 200.040 ;
                RECT 82.760 199.720 87.840 200.040 ;
                RECT 93.640 199.720 274.160 200.040 ;
                RECT 347.960 199.720 404.040 200.040 ;
                RECT 1116.360 199.720 1123.120 200.040 ;
                RECT 2.880 201.080 64.720 201.400 ;
                RECT 82.760 201.080 87.840 201.400 ;
                RECT 104.520 201.080 274.160 201.400 ;
                RECT 347.960 201.080 404.040 201.400 ;
                RECT 1116.360 201.080 1123.120 201.400 ;
                RECT 2.880 202.440 64.720 202.760 ;
                RECT 82.760 202.440 274.160 202.760 ;
                RECT 347.960 202.440 362.560 202.760 ;
                RECT 1116.360 202.440 1123.120 202.760 ;
                RECT 2.880 203.800 64.720 204.120 ;
                RECT 82.760 203.800 89.200 204.120 ;
                RECT 103.840 203.800 362.560 204.120 ;
                RECT 1116.360 203.800 1123.120 204.120 ;
                RECT 2.880 205.160 64.720 205.480 ;
                RECT 82.760 205.160 91.920 205.480 ;
                RECT 103.840 205.160 362.560 205.480 ;
                RECT 1116.360 205.160 1123.120 205.480 ;
                RECT 2.880 206.520 64.720 206.840 ;
                RECT 82.760 206.520 85.800 206.840 ;
                RECT 89.560 206.520 368.000 206.840 ;
                RECT 1116.360 206.520 1123.120 206.840 ;
                RECT 2.880 207.880 64.720 208.200 ;
                RECT 82.760 207.880 368.000 208.200 ;
                RECT 1116.360 207.880 1123.120 208.200 ;
                RECT 2.880 209.240 64.720 209.560 ;
                RECT 82.760 209.240 219.080 209.560 ;
                RECT 349.320 209.240 373.440 209.560 ;
                RECT 1116.360 209.240 1123.120 209.560 ;
                RECT 2.880 210.600 64.720 210.920 ;
                RECT 82.760 210.600 86.480 210.920 ;
                RECT 93.640 210.600 219.080 210.920 ;
                RECT 349.320 210.600 373.440 210.920 ;
                RECT 1116.360 210.600 1123.120 210.920 ;
                RECT 2.880 211.960 64.720 212.280 ;
                RECT 82.760 211.960 91.920 212.280 ;
                RECT 96.360 211.960 219.080 212.280 ;
                RECT 349.320 211.960 378.880 212.280 ;
                RECT 1116.360 211.960 1123.120 212.280 ;
                RECT 2.880 213.320 64.720 213.640 ;
                RECT 82.760 213.320 219.080 213.640 ;
                RECT 349.320 213.320 378.880 213.640 ;
                RECT 1116.360 213.320 1123.120 213.640 ;
                RECT 2.880 214.680 64.720 215.000 ;
                RECT 83.440 214.680 87.840 215.000 ;
                RECT 92.960 214.680 219.080 215.000 ;
                RECT 349.320 214.680 384.320 215.000 ;
                RECT 1116.360 214.680 1123.120 215.000 ;
                RECT 2.880 216.040 64.720 216.360 ;
                RECT 82.760 216.040 91.240 216.360 ;
                RECT 103.840 216.040 219.080 216.360 ;
                RECT 349.320 216.040 384.320 216.360 ;
                RECT 1116.360 216.040 1123.120 216.360 ;
                RECT 2.880 217.400 64.720 217.720 ;
                RECT 82.760 217.400 219.080 217.720 ;
                RECT 349.320 217.400 384.320 217.720 ;
                RECT 1116.360 217.400 1123.120 217.720 ;
                RECT 2.880 218.760 64.720 219.080 ;
                RECT 82.760 218.760 219.080 219.080 ;
                RECT 349.320 218.760 389.760 219.080 ;
                RECT 1116.360 218.760 1123.120 219.080 ;
                RECT 2.880 220.120 64.720 220.440 ;
                RECT 82.760 220.120 219.080 220.440 ;
                RECT 349.320 220.120 389.760 220.440 ;
                RECT 1116.360 220.120 1123.120 220.440 ;
                RECT 2.880 221.480 64.720 221.800 ;
                RECT 82.760 221.480 89.200 221.800 ;
                RECT 90.920 221.480 219.080 221.800 ;
                RECT 349.320 221.480 395.200 221.800 ;
                RECT 1116.360 221.480 1123.120 221.800 ;
                RECT 2.880 222.840 64.720 223.160 ;
                RECT 82.760 222.840 219.080 223.160 ;
                RECT 349.320 222.840 395.200 223.160 ;
                RECT 1116.360 222.840 1123.120 223.160 ;
                RECT 2.880 224.200 64.720 224.520 ;
                RECT 82.760 224.200 219.080 224.520 ;
                RECT 349.320 224.200 400.640 224.520 ;
                RECT 1116.360 224.200 1123.120 224.520 ;
                RECT 2.880 225.560 64.720 225.880 ;
                RECT 82.760 225.560 101.440 225.880 ;
                RECT 103.840 225.560 219.080 225.880 ;
                RECT 349.320 225.560 400.640 225.880 ;
                RECT 1116.360 225.560 1123.120 225.880 ;
                RECT 2.880 226.920 64.720 227.240 ;
                RECT 82.760 226.920 219.080 227.240 ;
                RECT 349.320 226.920 404.040 227.240 ;
                RECT 1116.360 226.920 1123.120 227.240 ;
                RECT 2.880 228.280 64.720 228.600 ;
                RECT 82.760 228.280 219.080 228.600 ;
                RECT 1116.360 228.280 1123.120 228.600 ;
                RECT 2.880 229.640 64.720 229.960 ;
                RECT 82.760 229.640 219.080 229.960 ;
                RECT 1116.360 229.640 1123.120 229.960 ;
                RECT 2.880 231.000 64.720 231.320 ;
                RECT 82.760 231.000 219.080 231.320 ;
                RECT 1116.360 231.000 1123.120 231.320 ;
                RECT 2.880 232.360 64.720 232.680 ;
                RECT 82.760 232.360 219.080 232.680 ;
                RECT 1116.360 232.360 1123.120 232.680 ;
                RECT 2.880 233.720 64.720 234.040 ;
                RECT 82.760 233.720 94.640 234.040 ;
                RECT 103.160 233.720 219.080 234.040 ;
                RECT 349.320 233.720 404.040 234.040 ;
                RECT 1116.360 233.720 1123.120 234.040 ;
                RECT 2.880 235.080 64.720 235.400 ;
                RECT 82.760 235.080 219.080 235.400 ;
                RECT 349.320 235.080 404.040 235.400 ;
                RECT 1116.360 235.080 1123.120 235.400 ;
                RECT 2.880 236.440 64.720 236.760 ;
                RECT 82.760 236.440 219.080 236.760 ;
                RECT 349.320 236.440 404.040 236.760 ;
                RECT 1116.360 236.440 1123.120 236.760 ;
                RECT 2.880 237.800 64.720 238.120 ;
                RECT 82.760 237.800 219.080 238.120 ;
                RECT 349.320 237.800 404.040 238.120 ;
                RECT 1116.360 237.800 1123.120 238.120 ;
                RECT 2.880 239.160 64.720 239.480 ;
                RECT 82.760 239.160 219.080 239.480 ;
                RECT 349.320 239.160 404.040 239.480 ;
                RECT 1116.360 239.160 1123.120 239.480 ;
                RECT 2.880 240.520 64.720 240.840 ;
                RECT 82.760 240.520 219.080 240.840 ;
                RECT 349.320 240.520 404.040 240.840 ;
                RECT 1116.360 240.520 1123.120 240.840 ;
                RECT 2.880 241.880 64.720 242.200 ;
                RECT 82.760 241.880 219.080 242.200 ;
                RECT 349.320 241.880 404.040 242.200 ;
                RECT 1116.360 241.880 1123.120 242.200 ;
                RECT 2.880 243.240 64.720 243.560 ;
                RECT 82.760 243.240 219.080 243.560 ;
                RECT 349.320 243.240 404.040 243.560 ;
                RECT 1116.360 243.240 1123.120 243.560 ;
                RECT 2.880 244.600 64.720 244.920 ;
                RECT 82.760 244.600 90.560 244.920 ;
                RECT 93.640 244.600 219.080 244.920 ;
                RECT 349.320 244.600 404.040 244.920 ;
                RECT 1116.360 244.600 1123.120 244.920 ;
                RECT 2.880 245.960 64.720 246.280 ;
                RECT 82.760 245.960 219.080 246.280 ;
                RECT 349.320 245.960 404.040 246.280 ;
                RECT 1116.360 245.960 1123.120 246.280 ;
                RECT 2.880 247.320 64.720 247.640 ;
                RECT 82.760 247.320 219.080 247.640 ;
                RECT 349.320 247.320 404.040 247.640 ;
                RECT 1116.360 247.320 1123.120 247.640 ;
                RECT 2.880 248.680 64.720 249.000 ;
                RECT 82.760 248.680 219.080 249.000 ;
                RECT 349.320 248.680 404.040 249.000 ;
                RECT 1116.360 248.680 1123.120 249.000 ;
                RECT 2.880 250.040 64.720 250.360 ;
                RECT 82.760 250.040 219.080 250.360 ;
                RECT 349.320 250.040 404.040 250.360 ;
                RECT 1116.360 250.040 1123.120 250.360 ;
                RECT 2.880 251.400 64.720 251.720 ;
                RECT 82.760 251.400 219.080 251.720 ;
                RECT 349.320 251.400 404.040 251.720 ;
                RECT 1116.360 251.400 1123.120 251.720 ;
                RECT 2.880 252.760 219.080 253.080 ;
                RECT 349.320 252.760 404.040 253.080 ;
                RECT 1116.360 252.760 1123.120 253.080 ;
                RECT 2.880 254.120 219.080 254.440 ;
                RECT 349.320 254.120 404.040 254.440 ;
                RECT 1116.360 254.120 1123.120 254.440 ;
                RECT 2.880 255.480 87.840 255.800 ;
                RECT 93.640 255.480 219.080 255.800 ;
                RECT 349.320 255.480 404.040 255.800 ;
                RECT 1116.360 255.480 1123.120 255.800 ;
                RECT 2.880 256.840 43.640 257.160 ;
                RECT 64.400 256.840 219.080 257.160 ;
                RECT 349.320 256.840 404.040 257.160 ;
                RECT 1116.360 256.840 1123.120 257.160 ;
                RECT 2.880 258.200 43.640 258.520 ;
                RECT 64.400 258.200 219.080 258.520 ;
                RECT 349.320 258.200 404.040 258.520 ;
                RECT 1116.360 258.200 1123.120 258.520 ;
                RECT 2.880 259.560 43.640 259.880 ;
                RECT 64.400 259.560 70.840 259.880 ;
                RECT 78.000 259.560 219.080 259.880 ;
                RECT 349.320 259.560 404.040 259.880 ;
                RECT 1116.360 259.560 1123.120 259.880 ;
                RECT 2.880 260.920 91.920 261.240 ;
                RECT 97.720 260.920 219.080 261.240 ;
                RECT 1116.360 260.920 1123.120 261.240 ;
                RECT 2.880 262.280 43.640 262.600 ;
                RECT 64.400 262.280 65.400 262.600 ;
                RECT 82.760 262.280 219.080 262.600 ;
                RECT 1116.360 262.280 1123.120 262.600 ;
                RECT 2.880 263.640 43.640 263.960 ;
                RECT 64.400 263.640 65.400 263.960 ;
                RECT 82.760 263.640 219.080 263.960 ;
                RECT 1116.360 263.640 1123.120 263.960 ;
                RECT 2.880 265.000 43.640 265.320 ;
                RECT 64.400 265.000 219.080 265.320 ;
                RECT 1116.360 265.000 1123.120 265.320 ;
                RECT 2.880 266.360 21.880 266.680 ;
                RECT 78.000 266.360 85.120 266.680 ;
                RECT 96.360 266.360 219.080 266.680 ;
                RECT 349.320 266.360 404.040 266.680 ;
                RECT 1116.360 266.360 1123.120 266.680 ;
                RECT 2.880 267.720 70.840 268.040 ;
                RECT 90.920 267.720 1123.120 268.040 ;
                RECT 2.880 269.080 87.840 269.400 ;
                RECT 131.720 269.080 1123.120 269.400 ;
                RECT 2.880 270.440 401.320 270.760 ;
                RECT 1118.400 270.440 1123.120 270.760 ;
                RECT 2.880 271.800 401.320 272.120 ;
                RECT 1118.400 271.800 1123.120 272.120 ;
                RECT 2.880 273.160 125.920 273.480 ;
                RECT 132.400 273.160 202.760 273.480 ;
                RECT 1118.400 273.160 1123.120 273.480 ;
                RECT 2.880 274.520 123.880 274.840 ;
                RECT 148.040 274.520 202.760 274.840 ;
                RECT 1118.400 274.520 1123.120 274.840 ;
                RECT 2.880 275.880 123.880 276.200 ;
                RECT 147.360 275.880 159.920 276.200 ;
                RECT 161.640 275.880 174.880 276.200 ;
                RECT 192.240 275.880 202.760 276.200 ;
                RECT 1118.400 275.880 1123.120 276.200 ;
                RECT 2.880 277.240 159.920 277.560 ;
                RECT 161.640 277.240 174.880 277.560 ;
                RECT 192.240 277.240 202.760 277.560 ;
                RECT 1118.400 277.240 1123.120 277.560 ;
                RECT 2.880 278.600 123.880 278.920 ;
                RECT 134.440 278.600 159.920 278.920 ;
                RECT 164.360 278.600 174.880 278.920 ;
                RECT 192.240 278.600 202.760 278.920 ;
                RECT 1118.400 278.600 1123.120 278.920 ;
                RECT 2.880 279.960 159.920 280.280 ;
                RECT 165.040 279.960 174.880 280.280 ;
                RECT 192.240 279.960 202.760 280.280 ;
                RECT 1118.400 279.960 1123.120 280.280 ;
                RECT 2.880 281.320 123.880 281.640 ;
                RECT 134.440 281.320 159.920 281.640 ;
                RECT 165.720 281.320 174.880 281.640 ;
                RECT 192.240 281.320 202.760 281.640 ;
                RECT 1118.400 281.320 1123.120 281.640 ;
                RECT 2.880 282.680 123.880 283.000 ;
                RECT 134.440 282.680 202.760 283.000 ;
                RECT 1118.400 282.680 1123.120 283.000 ;
                RECT 2.880 284.040 174.880 284.360 ;
                RECT 192.240 284.040 202.760 284.360 ;
                RECT 1118.400 284.040 1123.120 284.360 ;
                RECT 2.880 285.400 174.880 285.720 ;
                RECT 192.240 285.400 202.760 285.720 ;
                RECT 1118.400 285.400 1123.120 285.720 ;
                RECT 2.880 286.760 174.880 287.080 ;
                RECT 192.240 286.760 202.760 287.080 ;
                RECT 1118.400 286.760 1123.120 287.080 ;
                RECT 2.880 288.120 21.200 288.440 ;
                RECT 119.480 288.120 132.720 288.440 ;
                RECT 135.120 288.120 174.880 288.440 ;
                RECT 192.240 288.120 202.760 288.440 ;
                RECT 1118.400 288.120 1123.120 288.440 ;
                RECT 2.880 289.480 20.520 289.800 ;
                RECT 119.480 289.480 136.800 289.800 ;
                RECT 148.720 289.480 174.880 289.800 ;
                RECT 185.440 289.480 202.760 289.800 ;
                RECT 1118.400 289.480 1123.120 289.800 ;
                RECT 2.880 290.840 19.840 291.160 ;
                RECT 119.480 290.840 138.160 291.160 ;
                RECT 147.360 290.840 187.120 291.160 ;
                RECT 192.240 290.840 202.760 291.160 ;
                RECT 1118.400 290.840 1123.120 291.160 ;
                RECT 2.880 292.200 19.160 292.520 ;
                RECT 119.480 292.200 159.920 292.520 ;
                RECT 162.320 292.200 174.880 292.520 ;
                RECT 192.240 292.200 202.760 292.520 ;
                RECT 1118.400 292.200 1123.120 292.520 ;
                RECT 2.880 293.560 159.920 293.880 ;
                RECT 162.320 293.560 174.880 293.880 ;
                RECT 192.240 293.560 202.760 293.880 ;
                RECT 1118.400 293.560 1123.120 293.880 ;
                RECT 2.880 294.920 18.480 295.240 ;
                RECT 119.480 294.920 159.920 295.240 ;
                RECT 163.000 294.920 174.880 295.240 ;
                RECT 192.240 294.920 202.760 295.240 ;
                RECT 1118.400 294.920 1123.120 295.240 ;
                RECT 2.880 296.280 17.800 296.600 ;
                RECT 119.480 296.280 159.920 296.600 ;
                RECT 161.640 296.280 174.880 296.600 ;
                RECT 192.240 296.280 202.760 296.600 ;
                RECT 1118.400 296.280 1123.120 296.600 ;
                RECT 2.880 297.640 159.920 297.960 ;
                RECT 163.680 297.640 174.880 297.960 ;
                RECT 186.120 297.640 202.760 297.960 ;
                RECT 1118.400 297.640 1123.120 297.960 ;
                RECT 2.880 299.000 17.120 299.320 ;
                RECT 119.480 299.000 132.720 299.320 ;
                RECT 139.200 299.000 174.880 299.320 ;
                RECT 192.240 299.000 202.760 299.320 ;
                RECT 1118.400 299.000 1123.120 299.320 ;
                RECT 2.880 300.360 16.440 300.680 ;
                RECT 119.480 300.360 132.720 300.680 ;
                RECT 139.880 300.360 174.880 300.680 ;
                RECT 192.240 300.360 202.760 300.680 ;
                RECT 1118.400 300.360 1123.120 300.680 ;
                RECT 2.880 301.720 174.880 302.040 ;
                RECT 192.240 301.720 202.760 302.040 ;
                RECT 1118.400 301.720 1123.120 302.040 ;
                RECT 2.880 303.080 15.760 303.400 ;
                RECT 119.480 303.080 132.720 303.400 ;
                RECT 139.880 303.080 174.880 303.400 ;
                RECT 192.240 303.080 202.760 303.400 ;
                RECT 1118.400 303.080 1123.120 303.400 ;
                RECT 2.880 304.440 15.080 304.760 ;
                RECT 119.480 304.440 132.720 304.760 ;
                RECT 139.200 304.440 174.880 304.760 ;
                RECT 192.240 304.440 202.760 304.760 ;
                RECT 1118.400 304.440 1123.120 304.760 ;
                RECT 2.880 305.800 14.400 306.120 ;
                RECT 119.480 305.800 202.760 306.120 ;
                RECT 1118.400 305.800 1123.120 306.120 ;
                RECT 2.880 307.160 13.720 307.480 ;
                RECT 119.480 307.160 174.880 307.480 ;
                RECT 192.240 307.160 202.760 307.480 ;
                RECT 1118.400 307.160 1123.120 307.480 ;
                RECT 2.880 308.520 174.880 308.840 ;
                RECT 192.240 308.520 202.760 308.840 ;
                RECT 1118.400 308.520 1123.120 308.840 ;
                RECT 2.880 309.880 13.040 310.200 ;
                RECT 119.480 309.880 174.880 310.200 ;
                RECT 192.240 309.880 202.760 310.200 ;
                RECT 1118.400 309.880 1123.120 310.200 ;
                RECT 2.880 311.240 12.360 311.560 ;
                RECT 119.480 311.240 174.880 311.560 ;
                RECT 192.240 311.240 202.760 311.560 ;
                RECT 1118.400 311.240 1123.120 311.560 ;
                RECT 2.880 312.600 11.680 312.920 ;
                RECT 119.480 312.600 174.880 312.920 ;
                RECT 192.240 312.600 202.760 312.920 ;
                RECT 1118.400 312.600 1123.120 312.920 ;
                RECT 2.880 313.960 202.760 314.280 ;
                RECT 1118.400 313.960 1123.120 314.280 ;
                RECT 2.880 315.320 11.000 315.640 ;
                RECT 119.480 315.320 132.720 315.640 ;
                RECT 135.120 315.320 174.880 315.640 ;
                RECT 192.240 315.320 202.760 315.640 ;
                RECT 1118.400 315.320 1123.120 315.640 ;
                RECT 2.880 316.680 174.880 317.000 ;
                RECT 192.240 316.680 202.760 317.000 ;
                RECT 1118.400 316.680 1123.120 317.000 ;
                RECT 2.880 318.040 174.880 318.360 ;
                RECT 192.240 318.040 202.760 318.360 ;
                RECT 1118.400 318.040 1123.120 318.360 ;
                RECT 2.880 319.400 174.880 319.720 ;
                RECT 192.240 319.400 202.760 319.720 ;
                RECT 1118.400 319.400 1123.120 319.720 ;
                RECT 2.880 320.760 174.880 321.080 ;
                RECT 192.240 320.760 202.760 321.080 ;
                RECT 1118.400 320.760 1123.120 321.080 ;
                RECT 2.880 322.120 202.760 322.440 ;
                RECT 1118.400 322.120 1123.120 322.440 ;
                RECT 2.880 323.480 174.880 323.800 ;
                RECT 192.240 323.480 202.760 323.800 ;
                RECT 1118.400 323.480 1123.120 323.800 ;
                RECT 2.880 324.840 174.880 325.160 ;
                RECT 192.240 324.840 202.760 325.160 ;
                RECT 1118.400 324.840 1123.120 325.160 ;
                RECT 2.880 326.200 174.880 326.520 ;
                RECT 192.240 326.200 202.760 326.520 ;
                RECT 1118.400 326.200 1123.120 326.520 ;
                RECT 2.880 327.560 174.880 327.880 ;
                RECT 192.240 327.560 202.760 327.880 ;
                RECT 1118.400 327.560 1123.120 327.880 ;
                RECT 2.880 328.920 174.880 329.240 ;
                RECT 188.840 328.920 202.760 329.240 ;
                RECT 1118.400 328.920 1123.120 329.240 ;
                RECT 2.880 330.280 188.480 330.600 ;
                RECT 192.240 330.280 202.760 330.600 ;
                RECT 1118.400 330.280 1123.120 330.600 ;
                RECT 2.880 331.640 174.880 331.960 ;
                RECT 192.240 331.640 202.760 331.960 ;
                RECT 1118.400 331.640 1123.120 331.960 ;
                RECT 2.880 333.000 174.880 333.320 ;
                RECT 192.240 333.000 202.760 333.320 ;
                RECT 1118.400 333.000 1123.120 333.320 ;
                RECT 2.880 334.360 174.880 334.680 ;
                RECT 192.240 334.360 202.760 334.680 ;
                RECT 1118.400 334.360 1123.120 334.680 ;
                RECT 2.880 335.720 174.880 336.040 ;
                RECT 192.240 335.720 202.760 336.040 ;
                RECT 1118.400 335.720 1123.120 336.040 ;
                RECT 2.880 337.080 174.880 337.400 ;
                RECT 189.520 337.080 202.760 337.400 ;
                RECT 1118.400 337.080 1123.120 337.400 ;
                RECT 2.880 338.440 174.880 338.760 ;
                RECT 192.240 338.440 202.760 338.760 ;
                RECT 1118.400 338.440 1123.120 338.760 ;
                RECT 2.880 339.800 174.880 340.120 ;
                RECT 192.240 339.800 202.760 340.120 ;
                RECT 1118.400 339.800 1123.120 340.120 ;
                RECT 2.880 341.160 174.880 341.480 ;
                RECT 192.240 341.160 202.760 341.480 ;
                RECT 1118.400 341.160 1123.120 341.480 ;
                RECT 2.880 342.520 174.880 342.840 ;
                RECT 192.240 342.520 202.760 342.840 ;
                RECT 1118.400 342.520 1123.120 342.840 ;
                RECT 2.880 343.880 174.880 344.200 ;
                RECT 192.240 343.880 202.760 344.200 ;
                RECT 1118.400 343.880 1123.120 344.200 ;
                RECT 2.880 345.240 202.760 345.560 ;
                RECT 1118.400 345.240 1123.120 345.560 ;
                RECT 2.880 346.600 174.880 346.920 ;
                RECT 192.240 346.600 202.760 346.920 ;
                RECT 1118.400 346.600 1123.120 346.920 ;
                RECT 2.880 347.960 174.880 348.280 ;
                RECT 192.240 347.960 202.760 348.280 ;
                RECT 1118.400 347.960 1123.120 348.280 ;
                RECT 2.880 349.320 174.880 349.640 ;
                RECT 192.240 349.320 202.760 349.640 ;
                RECT 1118.400 349.320 1123.120 349.640 ;
                RECT 2.880 350.680 174.880 351.000 ;
                RECT 192.240 350.680 202.760 351.000 ;
                RECT 1118.400 350.680 1123.120 351.000 ;
                RECT 2.880 352.040 174.880 352.360 ;
                RECT 192.240 352.040 202.760 352.360 ;
                RECT 1118.400 352.040 1123.120 352.360 ;
                RECT 2.880 353.400 202.760 353.720 ;
                RECT 1118.400 353.400 1123.120 353.720 ;
                RECT 2.880 354.760 174.880 355.080 ;
                RECT 192.240 354.760 202.760 355.080 ;
                RECT 1118.400 354.760 1123.120 355.080 ;
                RECT 2.880 356.120 174.880 356.440 ;
                RECT 192.240 356.120 202.760 356.440 ;
                RECT 1118.400 356.120 1123.120 356.440 ;
                RECT 2.880 357.480 174.880 357.800 ;
                RECT 192.240 357.480 202.760 357.800 ;
                RECT 1118.400 357.480 1123.120 357.800 ;
                RECT 2.880 358.840 174.880 359.160 ;
                RECT 192.240 358.840 202.760 359.160 ;
                RECT 1118.400 358.840 1123.120 359.160 ;
                RECT 2.880 360.200 174.880 360.520 ;
                RECT 192.240 360.200 202.760 360.520 ;
                RECT 1118.400 360.200 1123.120 360.520 ;
                RECT 2.880 361.560 202.760 361.880 ;
                RECT 1118.400 361.560 1123.120 361.880 ;
                RECT 2.880 362.920 174.880 363.240 ;
                RECT 192.240 362.920 202.760 363.240 ;
                RECT 1118.400 362.920 1123.120 363.240 ;
                RECT 2.880 364.280 174.880 364.600 ;
                RECT 192.240 364.280 202.760 364.600 ;
                RECT 1118.400 364.280 1123.120 364.600 ;
                RECT 2.880 365.640 174.880 365.960 ;
                RECT 192.240 365.640 202.760 365.960 ;
                RECT 1118.400 365.640 1123.120 365.960 ;
                RECT 2.880 367.000 174.880 367.320 ;
                RECT 192.240 367.000 202.760 367.320 ;
                RECT 1118.400 367.000 1123.120 367.320 ;
                RECT 2.880 368.360 174.880 368.680 ;
                RECT 192.240 368.360 202.760 368.680 ;
                RECT 1118.400 368.360 1123.120 368.680 ;
                RECT 2.880 369.720 183.040 370.040 ;
                RECT 192.240 369.720 202.760 370.040 ;
                RECT 1118.400 369.720 1123.120 370.040 ;
                RECT 2.880 371.080 176.920 371.400 ;
                RECT 192.240 371.080 202.760 371.400 ;
                RECT 1118.400 371.080 1123.120 371.400 ;
                RECT 2.880 372.440 176.920 372.760 ;
                RECT 192.240 372.440 202.760 372.760 ;
                RECT 1118.400 372.440 1123.120 372.760 ;
                RECT 2.880 373.800 176.920 374.120 ;
                RECT 192.240 373.800 202.760 374.120 ;
                RECT 1118.400 373.800 1123.120 374.120 ;
                RECT 2.880 375.160 176.920 375.480 ;
                RECT 192.240 375.160 202.760 375.480 ;
                RECT 1118.400 375.160 1123.120 375.480 ;
                RECT 2.880 376.520 138.840 376.840 ;
                RECT 148.720 376.520 202.760 376.840 ;
                RECT 1118.400 376.520 1123.120 376.840 ;
                RECT 2.880 377.880 137.480 378.200 ;
                RECT 147.360 377.880 159.920 378.200 ;
                RECT 161.640 377.880 174.880 378.200 ;
                RECT 192.240 377.880 202.760 378.200 ;
                RECT 1118.400 377.880 1123.120 378.200 ;
                RECT 2.880 379.240 159.920 379.560 ;
                RECT 163.680 379.240 174.880 379.560 ;
                RECT 192.240 379.240 202.760 379.560 ;
                RECT 1118.400 379.240 1123.120 379.560 ;
                RECT 2.880 380.600 159.920 380.920 ;
                RECT 164.360 380.600 174.880 380.920 ;
                RECT 192.240 380.600 202.760 380.920 ;
                RECT 1118.400 380.600 1123.120 380.920 ;
                RECT 2.880 381.960 159.920 382.280 ;
                RECT 165.040 381.960 174.880 382.280 ;
                RECT 192.240 381.960 202.760 382.280 ;
                RECT 1118.400 381.960 1123.120 382.280 ;
                RECT 2.880 383.320 159.920 383.640 ;
                RECT 161.640 383.320 174.880 383.640 ;
                RECT 192.240 383.320 202.760 383.640 ;
                RECT 1118.400 383.320 1123.120 383.640 ;
                RECT 2.880 384.680 202.760 385.000 ;
                RECT 1118.400 384.680 1123.120 385.000 ;
                RECT 2.880 386.040 174.880 386.360 ;
                RECT 192.240 386.040 202.760 386.360 ;
                RECT 1118.400 386.040 1123.120 386.360 ;
                RECT 2.880 387.400 174.880 387.720 ;
                RECT 192.240 387.400 202.760 387.720 ;
                RECT 1118.400 387.400 1123.120 387.720 ;
                RECT 2.880 388.760 174.880 389.080 ;
                RECT 192.240 388.760 202.760 389.080 ;
                RECT 1118.400 388.760 1123.120 389.080 ;
                RECT 2.880 390.120 174.880 390.440 ;
                RECT 192.240 390.120 202.760 390.440 ;
                RECT 1118.400 390.120 1123.120 390.440 ;
                RECT 2.880 391.480 174.880 391.800 ;
                RECT 192.240 391.480 202.760 391.800 ;
                RECT 1118.400 391.480 1123.120 391.800 ;
                RECT 2.880 392.840 135.440 393.160 ;
                RECT 148.040 392.840 202.760 393.160 ;
                RECT 1118.400 392.840 1123.120 393.160 ;
                RECT 2.880 394.200 134.080 394.520 ;
                RECT 147.360 394.200 159.920 394.520 ;
                RECT 161.640 394.200 174.880 394.520 ;
                RECT 192.240 394.200 202.760 394.520 ;
                RECT 1118.400 394.200 1123.120 394.520 ;
                RECT 2.880 395.560 159.920 395.880 ;
                RECT 162.320 395.560 174.880 395.880 ;
                RECT 192.240 395.560 202.760 395.880 ;
                RECT 1118.400 395.560 1123.120 395.880 ;
                RECT 2.880 396.920 159.920 397.240 ;
                RECT 162.320 396.920 174.880 397.240 ;
                RECT 192.240 396.920 202.760 397.240 ;
                RECT 1118.400 396.920 1123.120 397.240 ;
                RECT 2.880 398.280 159.920 398.600 ;
                RECT 163.000 398.280 174.880 398.600 ;
                RECT 192.240 398.280 202.760 398.600 ;
                RECT 1118.400 398.280 1123.120 398.600 ;
                RECT 2.880 399.640 159.920 399.960 ;
                RECT 163.680 399.640 174.880 399.960 ;
                RECT 192.240 399.640 202.760 399.960 ;
                RECT 1118.400 399.640 1123.120 399.960 ;
                RECT 2.880 401.000 202.760 401.320 ;
                RECT 1118.400 401.000 1123.120 401.320 ;
                RECT 2.880 402.360 174.880 402.680 ;
                RECT 192.240 402.360 202.760 402.680 ;
                RECT 1118.400 402.360 1123.120 402.680 ;
                RECT 2.880 403.720 174.880 404.040 ;
                RECT 192.240 403.720 202.760 404.040 ;
                RECT 1118.400 403.720 1123.120 404.040 ;
                RECT 2.880 405.080 174.880 405.400 ;
                RECT 192.240 405.080 202.760 405.400 ;
                RECT 1118.400 405.080 1123.120 405.400 ;
                RECT 2.880 406.440 174.880 406.760 ;
                RECT 192.240 406.440 202.760 406.760 ;
                RECT 1118.400 406.440 1123.120 406.760 ;
                RECT 2.880 407.800 174.880 408.120 ;
                RECT 179.320 407.800 202.760 408.120 ;
                RECT 1118.400 407.800 1123.120 408.120 ;
                RECT 2.880 409.160 202.760 409.480 ;
                RECT 1118.400 409.160 1123.120 409.480 ;
                RECT 2.880 410.520 174.880 410.840 ;
                RECT 192.240 410.520 202.760 410.840 ;
                RECT 1118.400 410.520 1123.120 410.840 ;
                RECT 2.880 411.880 174.880 412.200 ;
                RECT 192.240 411.880 202.760 412.200 ;
                RECT 1118.400 411.880 1123.120 412.200 ;
                RECT 2.880 413.240 174.880 413.560 ;
                RECT 192.240 413.240 202.760 413.560 ;
                RECT 1118.400 413.240 1123.120 413.560 ;
                RECT 2.880 414.600 174.880 414.920 ;
                RECT 192.240 414.600 202.760 414.920 ;
                RECT 1118.400 414.600 1123.120 414.920 ;
                RECT 2.880 415.960 174.880 416.280 ;
                RECT 180.000 415.960 202.760 416.280 ;
                RECT 1118.400 415.960 1123.120 416.280 ;
                RECT 2.880 417.320 174.880 417.640 ;
                RECT 192.240 417.320 202.760 417.640 ;
                RECT 1118.400 417.320 1123.120 417.640 ;
                RECT 2.880 418.680 174.880 419.000 ;
                RECT 192.240 418.680 202.760 419.000 ;
                RECT 1118.400 418.680 1123.120 419.000 ;
                RECT 2.880 420.040 174.880 420.360 ;
                RECT 192.240 420.040 202.760 420.360 ;
                RECT 1118.400 420.040 1123.120 420.360 ;
                RECT 2.880 421.400 174.880 421.720 ;
                RECT 192.240 421.400 202.760 421.720 ;
                RECT 1118.400 421.400 1123.120 421.720 ;
                RECT 2.880 422.760 174.880 423.080 ;
                RECT 192.240 422.760 202.760 423.080 ;
                RECT 1118.400 422.760 1123.120 423.080 ;
                RECT 2.880 424.120 174.880 424.440 ;
                RECT 180.680 424.120 202.760 424.440 ;
                RECT 1118.400 424.120 1123.120 424.440 ;
                RECT 2.880 425.480 174.880 425.800 ;
                RECT 192.240 425.480 202.760 425.800 ;
                RECT 1118.400 425.480 1123.120 425.800 ;
                RECT 2.880 426.840 174.880 427.160 ;
                RECT 192.240 426.840 202.760 427.160 ;
                RECT 1118.400 426.840 1123.120 427.160 ;
                RECT 2.880 428.200 174.880 428.520 ;
                RECT 192.240 428.200 202.760 428.520 ;
                RECT 1118.400 428.200 1123.120 428.520 ;
                RECT 2.880 429.560 174.880 429.880 ;
                RECT 192.240 429.560 202.760 429.880 ;
                RECT 1118.400 429.560 1123.120 429.880 ;
                RECT 2.880 430.920 174.880 431.240 ;
                RECT 192.240 430.920 202.760 431.240 ;
                RECT 1118.400 430.920 1123.120 431.240 ;
                RECT 2.880 432.280 202.760 432.600 ;
                RECT 1118.400 432.280 1123.120 432.600 ;
                RECT 2.880 433.640 174.880 433.960 ;
                RECT 192.240 433.640 202.760 433.960 ;
                RECT 1118.400 433.640 1123.120 433.960 ;
                RECT 2.880 435.000 174.880 435.320 ;
                RECT 192.240 435.000 202.760 435.320 ;
                RECT 1118.400 435.000 1123.120 435.320 ;
                RECT 2.880 436.360 174.880 436.680 ;
                RECT 192.240 436.360 202.760 436.680 ;
                RECT 1118.400 436.360 1123.120 436.680 ;
                RECT 2.880 437.720 174.880 438.040 ;
                RECT 192.240 437.720 202.760 438.040 ;
                RECT 1118.400 437.720 1123.120 438.040 ;
                RECT 2.880 439.080 174.880 439.400 ;
                RECT 192.240 439.080 202.760 439.400 ;
                RECT 1118.400 439.080 1123.120 439.400 ;
                RECT 2.880 440.440 202.760 440.760 ;
                RECT 1118.400 440.440 1123.120 440.760 ;
                RECT 2.880 441.800 174.880 442.120 ;
                RECT 192.240 441.800 202.760 442.120 ;
                RECT 1118.400 441.800 1123.120 442.120 ;
                RECT 2.880 443.160 174.880 443.480 ;
                RECT 192.240 443.160 202.760 443.480 ;
                RECT 1118.400 443.160 1123.120 443.480 ;
                RECT 2.880 444.520 174.880 444.840 ;
                RECT 192.240 444.520 202.760 444.840 ;
                RECT 1118.400 444.520 1123.120 444.840 ;
                RECT 2.880 445.880 174.880 446.200 ;
                RECT 192.240 445.880 202.760 446.200 ;
                RECT 1118.400 445.880 1123.120 446.200 ;
                RECT 2.880 447.240 174.880 447.560 ;
                RECT 192.240 447.240 202.760 447.560 ;
                RECT 1118.400 447.240 1123.120 447.560 ;
                RECT 2.880 448.600 202.760 448.920 ;
                RECT 1118.400 448.600 1123.120 448.920 ;
                RECT 2.880 449.960 174.880 450.280 ;
                RECT 192.240 449.960 202.760 450.280 ;
                RECT 1118.400 449.960 1123.120 450.280 ;
                RECT 2.880 451.320 174.880 451.640 ;
                RECT 192.240 451.320 202.760 451.640 ;
                RECT 1118.400 451.320 1123.120 451.640 ;
                RECT 2.880 452.680 174.880 453.000 ;
                RECT 192.240 452.680 202.760 453.000 ;
                RECT 1118.400 452.680 1123.120 453.000 ;
                RECT 2.880 454.040 174.880 454.360 ;
                RECT 192.240 454.040 202.760 454.360 ;
                RECT 1118.400 454.040 1123.120 454.360 ;
                RECT 2.880 455.400 174.880 455.720 ;
                RECT 183.400 455.400 202.760 455.720 ;
                RECT 1118.400 455.400 1123.120 455.720 ;
                RECT 2.880 456.760 188.480 457.080 ;
                RECT 192.240 456.760 202.760 457.080 ;
                RECT 1118.400 456.760 1123.120 457.080 ;
                RECT 2.880 458.120 174.880 458.440 ;
                RECT 192.240 458.120 202.760 458.440 ;
                RECT 1118.400 458.120 1123.120 458.440 ;
                RECT 2.880 459.480 174.880 459.800 ;
                RECT 192.240 459.480 202.760 459.800 ;
                RECT 1118.400 459.480 1123.120 459.800 ;
                RECT 2.880 460.840 174.880 461.160 ;
                RECT 192.240 460.840 202.760 461.160 ;
                RECT 1118.400 460.840 1123.120 461.160 ;
                RECT 2.880 462.200 174.880 462.520 ;
                RECT 192.240 462.200 202.760 462.520 ;
                RECT 1118.400 462.200 1123.120 462.520 ;
                RECT 2.880 463.560 174.880 463.880 ;
                RECT 184.080 463.560 202.760 463.880 ;
                RECT 1118.400 463.560 1123.120 463.880 ;
                RECT 2.880 464.920 174.880 465.240 ;
                RECT 192.240 464.920 202.760 465.240 ;
                RECT 1118.400 464.920 1123.120 465.240 ;
                RECT 2.880 466.280 174.880 466.600 ;
                RECT 192.240 466.280 202.760 466.600 ;
                RECT 1118.400 466.280 1123.120 466.600 ;
                RECT 2.880 467.640 174.880 467.960 ;
                RECT 192.240 467.640 202.760 467.960 ;
                RECT 1118.400 467.640 1123.120 467.960 ;
                RECT 2.880 469.000 174.880 469.320 ;
                RECT 192.240 469.000 202.760 469.320 ;
                RECT 1118.400 469.000 1123.120 469.320 ;
                RECT 2.880 470.360 174.880 470.680 ;
                RECT 192.240 470.360 202.760 470.680 ;
                RECT 1118.400 470.360 1123.120 470.680 ;
                RECT 2.880 471.720 202.760 472.040 ;
                RECT 1118.400 471.720 1123.120 472.040 ;
                RECT 2.880 473.080 178.280 473.400 ;
                RECT 192.240 473.080 202.760 473.400 ;
                RECT 1118.400 473.080 1123.120 473.400 ;
                RECT 2.880 474.440 178.280 474.760 ;
                RECT 192.240 474.440 202.760 474.760 ;
                RECT 1118.400 474.440 1123.120 474.760 ;
                RECT 2.880 475.800 185.760 476.120 ;
                RECT 192.240 475.800 202.760 476.120 ;
                RECT 1118.400 475.800 1123.120 476.120 ;
                RECT 2.880 477.160 178.280 477.480 ;
                RECT 192.240 477.160 202.760 477.480 ;
                RECT 1118.400 477.160 1123.120 477.480 ;
                RECT 2.880 478.520 178.280 478.840 ;
                RECT 192.240 478.520 202.760 478.840 ;
                RECT 1118.400 478.520 1123.120 478.840 ;
                RECT 2.880 479.880 202.760 480.200 ;
                RECT 1118.400 479.880 1123.120 480.200 ;
                RECT 2.880 481.240 178.280 481.560 ;
                RECT 192.240 481.240 202.760 481.560 ;
                RECT 1118.400 481.240 1123.120 481.560 ;
                RECT 2.880 482.600 178.280 482.920 ;
                RECT 192.240 482.600 202.760 482.920 ;
                RECT 1118.400 482.600 1123.120 482.920 ;
                RECT 2.880 483.960 178.280 484.280 ;
                RECT 192.240 483.960 202.760 484.280 ;
                RECT 1118.400 483.960 1123.120 484.280 ;
                RECT 2.880 485.320 188.480 485.640 ;
                RECT 192.240 485.320 202.760 485.640 ;
                RECT 1118.400 485.320 1123.120 485.640 ;
                RECT 2.880 486.680 178.280 487.000 ;
                RECT 192.240 486.680 202.760 487.000 ;
                RECT 1118.400 486.680 1123.120 487.000 ;
                RECT 2.880 488.040 202.760 488.360 ;
                RECT 1118.400 488.040 1123.120 488.360 ;
                RECT 2.880 489.400 178.280 489.720 ;
                RECT 192.240 489.400 202.760 489.720 ;
                RECT 1118.400 489.400 1123.120 489.720 ;
                RECT 2.880 490.760 178.280 491.080 ;
                RECT 192.240 490.760 202.760 491.080 ;
                RECT 1118.400 490.760 1123.120 491.080 ;
                RECT 2.880 492.120 178.280 492.440 ;
                RECT 192.240 492.120 202.760 492.440 ;
                RECT 1118.400 492.120 1123.120 492.440 ;
                RECT 2.880 493.480 178.280 493.800 ;
                RECT 192.240 493.480 202.760 493.800 ;
                RECT 1118.400 493.480 1123.120 493.800 ;
                RECT 2.880 494.840 202.760 495.160 ;
                RECT 1118.400 494.840 1123.120 495.160 ;
                RECT 2.880 496.200 183.040 496.520 ;
                RECT 192.240 496.200 202.760 496.520 ;
                RECT 1118.400 496.200 1123.120 496.520 ;
                RECT 2.880 497.560 178.960 497.880 ;
                RECT 192.240 497.560 202.760 497.880 ;
                RECT 1118.400 497.560 1123.120 497.880 ;
                RECT 2.880 498.920 178.960 499.240 ;
                RECT 192.240 498.920 202.760 499.240 ;
                RECT 1118.400 498.920 1123.120 499.240 ;
                RECT 2.880 500.280 178.960 500.600 ;
                RECT 192.240 500.280 202.760 500.600 ;
                RECT 1118.400 500.280 1123.120 500.600 ;
                RECT 2.880 501.640 178.960 501.960 ;
                RECT 192.240 501.640 202.760 501.960 ;
                RECT 1118.400 501.640 1123.120 501.960 ;
                RECT 2.880 503.000 202.760 503.320 ;
                RECT 1118.400 503.000 1123.120 503.320 ;
                RECT 2.880 504.360 185.080 504.680 ;
                RECT 192.240 504.360 202.760 504.680 ;
                RECT 1118.400 504.360 1123.120 504.680 ;
                RECT 2.880 505.720 178.960 506.040 ;
                RECT 192.240 505.720 202.760 506.040 ;
                RECT 1118.400 505.720 1123.120 506.040 ;
                RECT 2.880 507.080 178.960 507.400 ;
                RECT 192.240 507.080 202.760 507.400 ;
                RECT 1118.400 507.080 1123.120 507.400 ;
                RECT 2.880 508.440 178.960 508.760 ;
                RECT 192.240 508.440 202.760 508.760 ;
                RECT 1118.400 508.440 1123.120 508.760 ;
                RECT 2.880 509.800 178.960 510.120 ;
                RECT 192.240 509.800 202.760 510.120 ;
                RECT 1118.400 509.800 1123.120 510.120 ;
                RECT 2.880 511.160 202.760 511.480 ;
                RECT 1118.400 511.160 1123.120 511.480 ;
                RECT 2.880 512.520 178.960 512.840 ;
                RECT 192.240 512.520 202.760 512.840 ;
                RECT 1118.400 512.520 1123.120 512.840 ;
                RECT 2.880 513.880 187.120 514.200 ;
                RECT 192.240 513.880 202.760 514.200 ;
                RECT 1118.400 513.880 1123.120 514.200 ;
                RECT 2.880 515.240 187.800 515.560 ;
                RECT 192.240 515.240 202.760 515.560 ;
                RECT 1118.400 515.240 1123.120 515.560 ;
                RECT 2.880 516.600 178.960 516.920 ;
                RECT 192.240 516.600 202.760 516.920 ;
                RECT 1118.400 516.600 1123.120 516.920 ;
                RECT 2.880 517.960 178.960 518.280 ;
                RECT 192.240 517.960 202.760 518.280 ;
                RECT 1118.400 517.960 1123.120 518.280 ;
                RECT 2.880 519.320 202.760 519.640 ;
                RECT 1118.400 519.320 1123.120 519.640 ;
                RECT 2.880 520.680 178.960 521.000 ;
                RECT 192.240 520.680 202.760 521.000 ;
                RECT 1118.400 520.680 1123.120 521.000 ;
                RECT 2.880 522.040 178.960 522.360 ;
                RECT 192.240 522.040 202.760 522.360 ;
                RECT 1118.400 522.040 1123.120 522.360 ;
                RECT 2.880 523.400 189.840 523.720 ;
                RECT 192.240 523.400 202.760 523.720 ;
                RECT 1118.400 523.400 1123.120 523.720 ;
                RECT 2.880 524.760 190.520 525.080 ;
                RECT 192.240 524.760 202.760 525.080 ;
                RECT 1118.400 524.760 1123.120 525.080 ;
                RECT 2.880 526.120 178.960 526.440 ;
                RECT 192.240 526.120 202.760 526.440 ;
                RECT 1118.400 526.120 1123.120 526.440 ;
                RECT 2.880 527.480 202.760 527.800 ;
                RECT 1118.400 527.480 1123.120 527.800 ;
                RECT 2.880 528.840 178.960 529.160 ;
                RECT 192.240 528.840 202.760 529.160 ;
                RECT 1118.400 528.840 1123.120 529.160 ;
                RECT 2.880 530.200 178.960 530.520 ;
                RECT 192.240 530.200 202.760 530.520 ;
                RECT 1118.400 530.200 1123.120 530.520 ;
                RECT 2.880 531.560 178.960 531.880 ;
                RECT 192.240 531.560 202.760 531.880 ;
                RECT 1118.400 531.560 1123.120 531.880 ;
                RECT 2.880 532.920 178.960 533.240 ;
                RECT 192.240 532.920 202.760 533.240 ;
                RECT 1118.400 532.920 1123.120 533.240 ;
                RECT 2.880 534.280 202.760 534.600 ;
                RECT 1118.400 534.280 1123.120 534.600 ;
                RECT 2.880 535.640 185.080 535.960 ;
                RECT 192.240 535.640 202.760 535.960 ;
                RECT 1118.400 535.640 1123.120 535.960 ;
                RECT 2.880 537.000 178.960 537.320 ;
                RECT 192.240 537.000 202.760 537.320 ;
                RECT 1118.400 537.000 1123.120 537.320 ;
                RECT 2.880 538.360 178.960 538.680 ;
                RECT 192.240 538.360 202.760 538.680 ;
                RECT 1118.400 538.360 1123.120 538.680 ;
                RECT 2.880 539.720 178.960 540.040 ;
                RECT 192.240 539.720 202.760 540.040 ;
                RECT 1118.400 539.720 1123.120 540.040 ;
                RECT 2.880 541.080 178.960 541.400 ;
                RECT 192.240 541.080 202.760 541.400 ;
                RECT 1118.400 541.080 1123.120 541.400 ;
                RECT 2.880 542.440 202.760 542.760 ;
                RECT 1118.400 542.440 1123.120 542.760 ;
                RECT 2.880 543.800 187.120 544.120 ;
                RECT 192.240 543.800 202.760 544.120 ;
                RECT 1118.400 543.800 1123.120 544.120 ;
                RECT 2.880 545.160 178.960 545.480 ;
                RECT 192.240 545.160 202.760 545.480 ;
                RECT 1118.400 545.160 1123.120 545.480 ;
                RECT 2.880 546.520 178.960 546.840 ;
                RECT 192.240 546.520 202.760 546.840 ;
                RECT 1118.400 546.520 1123.120 546.840 ;
                RECT 2.880 547.880 178.960 548.200 ;
                RECT 192.240 547.880 202.760 548.200 ;
                RECT 1118.400 547.880 1123.120 548.200 ;
                RECT 2.880 549.240 178.960 549.560 ;
                RECT 192.240 549.240 202.760 549.560 ;
                RECT 1118.400 549.240 1123.120 549.560 ;
                RECT 2.880 550.600 202.760 550.920 ;
                RECT 1118.400 550.600 1123.120 550.920 ;
                RECT 2.880 551.960 178.960 552.280 ;
                RECT 192.240 551.960 202.760 552.280 ;
                RECT 1118.400 551.960 1123.120 552.280 ;
                RECT 2.880 553.320 189.160 553.640 ;
                RECT 192.240 553.320 202.760 553.640 ;
                RECT 1118.400 553.320 1123.120 553.640 ;
                RECT 2.880 554.680 178.960 555.000 ;
                RECT 192.240 554.680 202.760 555.000 ;
                RECT 1118.400 554.680 1123.120 555.000 ;
                RECT 2.880 556.040 178.960 556.360 ;
                RECT 192.240 556.040 202.760 556.360 ;
                RECT 1118.400 556.040 1123.120 556.360 ;
                RECT 2.880 557.400 178.960 557.720 ;
                RECT 192.240 557.400 202.760 557.720 ;
                RECT 1118.400 557.400 1123.120 557.720 ;
                RECT 2.880 558.760 202.760 559.080 ;
                RECT 1118.400 558.760 1123.120 559.080 ;
                RECT 2.880 560.120 179.640 560.440 ;
                RECT 192.240 560.120 202.760 560.440 ;
                RECT 1118.400 560.120 1123.120 560.440 ;
                RECT 2.880 561.480 179.640 561.800 ;
                RECT 192.240 561.480 202.760 561.800 ;
                RECT 1118.400 561.480 1123.120 561.800 ;
                RECT 2.880 562.840 183.720 563.160 ;
                RECT 192.240 562.840 202.760 563.160 ;
                RECT 1118.400 562.840 1123.120 563.160 ;
                RECT 2.880 564.200 179.640 564.520 ;
                RECT 192.240 564.200 202.760 564.520 ;
                RECT 1118.400 564.200 1123.120 564.520 ;
                RECT 2.880 565.560 179.640 565.880 ;
                RECT 192.240 565.560 202.760 565.880 ;
                RECT 1118.400 565.560 1123.120 565.880 ;
                RECT 2.880 566.920 202.760 567.240 ;
                RECT 1118.400 566.920 1123.120 567.240 ;
                RECT 2.880 568.280 179.640 568.600 ;
                RECT 192.240 568.280 202.760 568.600 ;
                RECT 1118.400 568.280 1123.120 568.600 ;
                RECT 2.880 569.640 179.640 569.960 ;
                RECT 192.240 569.640 202.760 569.960 ;
                RECT 1118.400 569.640 1123.120 569.960 ;
                RECT 2.880 571.000 179.640 571.320 ;
                RECT 192.240 571.000 202.760 571.320 ;
                RECT 1118.400 571.000 1123.120 571.320 ;
                RECT 2.880 572.360 186.440 572.680 ;
                RECT 192.240 572.360 202.760 572.680 ;
                RECT 1118.400 572.360 1123.120 572.680 ;
                RECT 2.880 573.720 202.760 574.040 ;
                RECT 1118.400 573.720 1123.120 574.040 ;
                RECT 2.880 575.080 187.120 575.400 ;
                RECT 192.240 575.080 202.760 575.400 ;
                RECT 1118.400 575.080 1123.120 575.400 ;
                RECT 2.880 576.440 179.640 576.760 ;
                RECT 192.240 576.440 202.760 576.760 ;
                RECT 1118.400 576.440 1123.120 576.760 ;
                RECT 2.880 577.800 179.640 578.120 ;
                RECT 192.240 577.800 202.760 578.120 ;
                RECT 1118.400 577.800 1123.120 578.120 ;
                RECT 2.880 579.160 179.640 579.480 ;
                RECT 192.240 579.160 202.760 579.480 ;
                RECT 1118.400 579.160 1123.120 579.480 ;
                RECT 2.880 580.520 179.640 580.840 ;
                RECT 192.240 580.520 202.760 580.840 ;
                RECT 1118.400 580.520 1123.120 580.840 ;
                RECT 2.880 581.880 202.760 582.200 ;
                RECT 1118.400 581.880 1123.120 582.200 ;
                RECT 2.880 583.240 188.480 583.560 ;
                RECT 192.240 583.240 202.760 583.560 ;
                RECT 1118.400 583.240 1123.120 583.560 ;
                RECT 2.880 584.600 179.640 584.920 ;
                RECT 192.240 584.600 202.760 584.920 ;
                RECT 1118.400 584.600 1123.120 584.920 ;
                RECT 2.880 585.960 179.640 586.280 ;
                RECT 192.240 585.960 202.760 586.280 ;
                RECT 1118.400 585.960 1123.120 586.280 ;
                RECT 2.880 587.320 179.640 587.640 ;
                RECT 192.240 587.320 202.760 587.640 ;
                RECT 1118.400 587.320 1123.120 587.640 ;
                RECT 2.880 588.680 179.640 589.000 ;
                RECT 192.240 588.680 202.760 589.000 ;
                RECT 1118.400 588.680 1123.120 589.000 ;
                RECT 2.880 590.040 202.760 590.360 ;
                RECT 1118.400 590.040 1123.120 590.360 ;
                RECT 2.880 591.400 180.320 591.720 ;
                RECT 192.240 591.400 202.760 591.720 ;
                RECT 1118.400 591.400 1123.120 591.720 ;
                RECT 2.880 592.760 183.720 593.080 ;
                RECT 192.240 592.760 202.760 593.080 ;
                RECT 1118.400 592.760 1123.120 593.080 ;
                RECT 2.880 594.120 180.320 594.440 ;
                RECT 192.240 594.120 202.760 594.440 ;
                RECT 1118.400 594.120 1123.120 594.440 ;
                RECT 2.880 595.480 180.320 595.800 ;
                RECT 192.240 595.480 202.760 595.800 ;
                RECT 1118.400 595.480 1123.120 595.800 ;
                RECT 2.880 596.840 180.320 597.160 ;
                RECT 192.240 596.840 202.760 597.160 ;
                RECT 1118.400 596.840 1123.120 597.160 ;
                RECT 2.880 598.200 202.760 598.520 ;
                RECT 1118.400 598.200 1123.120 598.520 ;
                RECT 2.880 599.560 180.320 599.880 ;
                RECT 192.240 599.560 202.760 599.880 ;
                RECT 1118.400 599.560 1123.120 599.880 ;
                RECT 2.880 600.920 180.320 601.240 ;
                RECT 192.240 600.920 202.760 601.240 ;
                RECT 1118.400 600.920 1123.120 601.240 ;
                RECT 2.880 602.280 185.760 602.600 ;
                RECT 192.240 602.280 202.760 602.600 ;
                RECT 1118.400 602.280 1123.120 602.600 ;
                RECT 2.880 603.640 180.320 603.960 ;
                RECT 192.240 603.640 202.760 603.960 ;
                RECT 1118.400 603.640 1123.120 603.960 ;
                RECT 2.880 605.000 180.320 605.320 ;
                RECT 192.240 605.000 202.760 605.320 ;
                RECT 1118.400 605.000 1123.120 605.320 ;
                RECT 2.880 606.360 202.760 606.680 ;
                RECT 1118.400 606.360 1123.120 606.680 ;
                RECT 2.880 607.720 180.320 608.040 ;
                RECT 192.240 607.720 202.760 608.040 ;
                RECT 1118.400 607.720 1123.120 608.040 ;
                RECT 2.880 609.080 180.320 609.400 ;
                RECT 192.240 609.080 202.760 609.400 ;
                RECT 1118.400 609.080 1123.120 609.400 ;
                RECT 2.880 610.440 180.320 610.760 ;
                RECT 192.240 610.440 202.760 610.760 ;
                RECT 1118.400 610.440 1123.120 610.760 ;
                RECT 2.880 611.800 188.480 612.120 ;
                RECT 192.240 611.800 202.760 612.120 ;
                RECT 1118.400 611.800 1123.120 612.120 ;
                RECT 2.880 613.160 180.320 613.480 ;
                RECT 192.240 613.160 202.760 613.480 ;
                RECT 1118.400 613.160 1123.120 613.480 ;
                RECT 2.880 614.520 202.760 614.840 ;
                RECT 1118.400 614.520 1123.120 614.840 ;
                RECT 2.880 615.880 180.320 616.200 ;
                RECT 192.240 615.880 202.760 616.200 ;
                RECT 1118.400 615.880 1123.120 616.200 ;
                RECT 2.880 617.240 180.320 617.560 ;
                RECT 192.240 617.240 202.760 617.560 ;
                RECT 1118.400 617.240 1123.120 617.560 ;
                RECT 2.880 618.600 180.320 618.920 ;
                RECT 192.240 618.600 202.760 618.920 ;
                RECT 1118.400 618.600 1123.120 618.920 ;
                RECT 2.880 619.960 180.320 620.280 ;
                RECT 192.240 619.960 202.760 620.280 ;
                RECT 1118.400 619.960 1123.120 620.280 ;
                RECT 2.880 621.320 202.760 621.640 ;
                RECT 1118.400 621.320 1123.120 621.640 ;
                RECT 2.880 622.680 183.040 623.000 ;
                RECT 192.240 622.680 202.760 623.000 ;
                RECT 1118.400 622.680 1123.120 623.000 ;
                RECT 2.880 624.040 180.320 624.360 ;
                RECT 192.240 624.040 202.760 624.360 ;
                RECT 1118.400 624.040 1123.120 624.360 ;
                RECT 2.880 625.400 180.320 625.720 ;
                RECT 192.240 625.400 202.760 625.720 ;
                RECT 1118.400 625.400 1123.120 625.720 ;
                RECT 2.880 626.760 180.320 627.080 ;
                RECT 192.240 626.760 202.760 627.080 ;
                RECT 1118.400 626.760 1123.120 627.080 ;
                RECT 2.880 628.120 180.320 628.440 ;
                RECT 192.240 628.120 202.760 628.440 ;
                RECT 1118.400 628.120 1123.120 628.440 ;
                RECT 2.880 629.480 202.760 629.800 ;
                RECT 1118.400 629.480 1123.120 629.800 ;
                RECT 2.880 630.840 185.080 631.160 ;
                RECT 192.240 630.840 202.760 631.160 ;
                RECT 1118.400 630.840 1123.120 631.160 ;
                RECT 2.880 632.200 185.080 632.520 ;
                RECT 192.240 632.200 202.760 632.520 ;
                RECT 1118.400 632.200 1123.120 632.520 ;
                RECT 2.880 633.560 180.320 633.880 ;
                RECT 192.240 633.560 202.760 633.880 ;
                RECT 1118.400 633.560 1123.120 633.880 ;
                RECT 2.880 634.920 180.320 635.240 ;
                RECT 192.240 634.920 202.760 635.240 ;
                RECT 1118.400 634.920 1123.120 635.240 ;
                RECT 2.880 636.280 180.320 636.600 ;
                RECT 192.240 636.280 202.760 636.600 ;
                RECT 1118.400 636.280 1123.120 636.600 ;
                RECT 2.880 637.640 202.760 637.960 ;
                RECT 1118.400 637.640 1123.120 637.960 ;
                RECT 2.880 639.000 180.320 639.320 ;
                RECT 192.240 639.000 202.760 639.320 ;
                RECT 1118.400 639.000 1123.120 639.320 ;
                RECT 2.880 640.360 180.320 640.680 ;
                RECT 192.240 640.360 202.760 640.680 ;
                RECT 1118.400 640.360 1123.120 640.680 ;
                RECT 2.880 641.720 187.800 642.040 ;
                RECT 192.240 641.720 202.760 642.040 ;
                RECT 1118.400 641.720 1123.120 642.040 ;
                RECT 2.880 643.080 180.320 643.400 ;
                RECT 192.240 643.080 202.760 643.400 ;
                RECT 1118.400 643.080 1123.120 643.400 ;
                RECT 2.880 644.440 180.320 644.760 ;
                RECT 192.240 644.440 202.760 644.760 ;
                RECT 1118.400 644.440 1123.120 644.760 ;
                RECT 2.880 645.800 202.760 646.120 ;
                RECT 1118.400 645.800 1123.120 646.120 ;
                RECT 2.880 647.160 180.320 647.480 ;
                RECT 192.240 647.160 202.760 647.480 ;
                RECT 1118.400 647.160 1123.120 647.480 ;
                RECT 2.880 648.520 180.320 648.840 ;
                RECT 192.240 648.520 202.760 648.840 ;
                RECT 1118.400 648.520 1123.120 648.840 ;
                RECT 2.880 649.880 180.320 650.200 ;
                RECT 192.240 649.880 202.760 650.200 ;
                RECT 1118.400 649.880 1123.120 650.200 ;
                RECT 2.880 651.240 190.520 651.560 ;
                RECT 192.240 651.240 202.760 651.560 ;
                RECT 1118.400 651.240 1123.120 651.560 ;
                RECT 2.880 652.600 180.320 652.920 ;
                RECT 192.240 652.600 202.760 652.920 ;
                RECT 1118.400 652.600 1123.120 652.920 ;
                RECT 2.880 653.960 202.760 654.280 ;
                RECT 1118.400 653.960 1123.120 654.280 ;
                RECT 2.880 655.320 181.000 655.640 ;
                RECT 192.240 655.320 202.760 655.640 ;
                RECT 1118.400 655.320 1123.120 655.640 ;
                RECT 2.880 656.680 181.000 657.000 ;
                RECT 192.240 656.680 202.760 657.000 ;
                RECT 1118.400 656.680 1123.120 657.000 ;
                RECT 2.880 658.040 181.000 658.360 ;
                RECT 192.240 658.040 202.760 658.360 ;
                RECT 1118.400 658.040 1123.120 658.360 ;
                RECT 2.880 659.400 181.000 659.720 ;
                RECT 192.240 659.400 202.760 659.720 ;
                RECT 1118.400 659.400 1123.120 659.720 ;
                RECT 2.880 660.760 202.760 661.080 ;
                RECT 1118.400 660.760 1123.120 661.080 ;
                RECT 2.880 662.120 185.080 662.440 ;
                RECT 192.240 662.120 202.760 662.440 ;
                RECT 1118.400 662.120 1123.120 662.440 ;
                RECT 2.880 663.480 181.000 663.800 ;
                RECT 192.240 663.480 202.760 663.800 ;
                RECT 1118.400 663.480 1123.120 663.800 ;
                RECT 2.880 664.840 181.000 665.160 ;
                RECT 192.240 664.840 202.760 665.160 ;
                RECT 1118.400 664.840 1123.120 665.160 ;
                RECT 2.880 666.200 181.000 666.520 ;
                RECT 192.240 666.200 202.760 666.520 ;
                RECT 1118.400 666.200 1123.120 666.520 ;
                RECT 2.880 667.560 181.000 667.880 ;
                RECT 192.240 667.560 202.760 667.880 ;
                RECT 1118.400 667.560 1123.120 667.880 ;
                RECT 2.880 668.920 202.760 669.240 ;
                RECT 1118.400 668.920 1123.120 669.240 ;
                RECT 2.880 670.280 187.120 670.600 ;
                RECT 192.240 670.280 202.760 670.600 ;
                RECT 1118.400 670.280 1123.120 670.600 ;
                RECT 2.880 671.640 181.000 671.960 ;
                RECT 192.240 671.640 202.760 671.960 ;
                RECT 1118.400 671.640 1123.120 671.960 ;
                RECT 2.880 673.000 181.000 673.320 ;
                RECT 192.240 673.000 202.760 673.320 ;
                RECT 1118.400 673.000 1123.120 673.320 ;
                RECT 2.880 674.360 181.000 674.680 ;
                RECT 192.240 674.360 202.760 674.680 ;
                RECT 1118.400 674.360 1123.120 674.680 ;
                RECT 2.880 675.720 181.000 676.040 ;
                RECT 192.240 675.720 202.760 676.040 ;
                RECT 1118.400 675.720 1123.120 676.040 ;
                RECT 2.880 677.080 202.760 677.400 ;
                RECT 1118.400 677.080 1123.120 677.400 ;
                RECT 2.880 678.440 181.000 678.760 ;
                RECT 192.240 678.440 202.760 678.760 ;
                RECT 1118.400 678.440 1123.120 678.760 ;
                RECT 2.880 679.800 189.160 680.120 ;
                RECT 192.240 679.800 202.760 680.120 ;
                RECT 1118.400 679.800 1123.120 680.120 ;
                RECT 2.880 681.160 189.840 681.480 ;
                RECT 192.240 681.160 202.760 681.480 ;
                RECT 1118.400 681.160 1123.120 681.480 ;
                RECT 2.880 682.520 181.000 682.840 ;
                RECT 192.240 682.520 202.760 682.840 ;
                RECT 1118.400 682.520 1123.120 682.840 ;
                RECT 2.880 683.880 181.000 684.200 ;
                RECT 192.240 683.880 202.760 684.200 ;
                RECT 1118.400 683.880 1123.120 684.200 ;
                RECT 2.880 685.240 202.760 685.560 ;
                RECT 1118.400 685.240 1123.120 685.560 ;
                RECT 2.880 686.600 181.680 686.920 ;
                RECT 192.240 686.600 202.760 686.920 ;
                RECT 1118.400 686.600 1123.120 686.920 ;
                RECT 2.880 687.960 181.680 688.280 ;
                RECT 192.240 687.960 202.760 688.280 ;
                RECT 1118.400 687.960 1123.120 688.280 ;
                RECT 2.880 689.320 181.680 689.640 ;
                RECT 192.240 689.320 202.760 689.640 ;
                RECT 1118.400 689.320 1123.120 689.640 ;
                RECT 2.880 690.680 184.400 691.000 ;
                RECT 192.240 690.680 202.760 691.000 ;
                RECT 1118.400 690.680 1123.120 691.000 ;
                RECT 2.880 692.040 181.680 692.360 ;
                RECT 192.240 692.040 202.760 692.360 ;
                RECT 1118.400 692.040 1123.120 692.360 ;
                RECT 2.880 693.400 202.760 693.720 ;
                RECT 1118.400 693.400 1123.120 693.720 ;
                RECT 2.880 694.760 181.680 695.080 ;
                RECT 192.240 694.760 202.760 695.080 ;
                RECT 1118.400 694.760 1123.120 695.080 ;
                RECT 2.880 696.120 181.680 696.440 ;
                RECT 192.240 696.120 202.760 696.440 ;
                RECT 1118.400 696.120 1123.120 696.440 ;
                RECT 2.880 697.480 181.680 697.800 ;
                RECT 192.240 697.480 202.760 697.800 ;
                RECT 1118.400 697.480 1123.120 697.800 ;
                RECT 2.880 698.840 181.680 699.160 ;
                RECT 192.240 698.840 202.760 699.160 ;
                RECT 1118.400 698.840 1123.120 699.160 ;
                RECT 2.880 700.200 202.760 700.520 ;
                RECT 1118.400 700.200 1123.120 700.520 ;
                RECT 2.880 701.560 187.120 701.880 ;
                RECT 192.240 701.560 202.760 701.880 ;
                RECT 1118.400 701.560 1123.120 701.880 ;
                RECT 2.880 702.920 181.680 703.240 ;
                RECT 192.240 702.920 202.760 703.240 ;
                RECT 1118.400 702.920 1123.120 703.240 ;
                RECT 2.880 704.280 181.680 704.600 ;
                RECT 192.240 704.280 202.760 704.600 ;
                RECT 1118.400 704.280 1123.120 704.600 ;
                RECT 2.880 705.640 181.680 705.960 ;
                RECT 192.240 705.640 202.760 705.960 ;
                RECT 1118.400 705.640 1123.120 705.960 ;
                RECT 2.880 707.000 181.680 707.320 ;
                RECT 192.240 707.000 202.760 707.320 ;
                RECT 1118.400 707.000 1123.120 707.320 ;
                RECT 2.880 708.360 202.760 708.680 ;
                RECT 1118.400 708.360 1123.120 708.680 ;
                RECT 2.880 709.720 188.480 710.040 ;
                RECT 192.240 709.720 202.760 710.040 ;
                RECT 1118.400 709.720 1123.120 710.040 ;
                RECT 2.880 711.080 181.680 711.400 ;
                RECT 192.240 711.080 202.760 711.400 ;
                RECT 1118.400 711.080 1123.120 711.400 ;
                RECT 2.880 712.440 181.680 712.760 ;
                RECT 192.240 712.440 202.760 712.760 ;
                RECT 1118.400 712.440 1123.120 712.760 ;
                RECT 2.880 713.800 181.680 714.120 ;
                RECT 192.240 713.800 202.760 714.120 ;
                RECT 1118.400 713.800 1123.120 714.120 ;
                RECT 2.880 715.160 181.680 715.480 ;
                RECT 192.240 715.160 202.760 715.480 ;
                RECT 1118.400 715.160 1123.120 715.480 ;
                RECT 2.880 716.520 202.760 716.840 ;
                RECT 1118.400 716.520 1123.120 716.840 ;
                RECT 2.880 717.880 182.360 718.200 ;
                RECT 192.240 717.880 202.760 718.200 ;
                RECT 1118.400 717.880 1123.120 718.200 ;
                RECT 2.880 719.240 183.720 719.560 ;
                RECT 192.240 719.240 202.760 719.560 ;
                RECT 1118.400 719.240 1123.120 719.560 ;
                RECT 2.880 720.600 182.360 720.920 ;
                RECT 192.240 720.600 202.760 720.920 ;
                RECT 1118.400 720.600 1123.120 720.920 ;
                RECT 2.880 721.960 182.360 722.280 ;
                RECT 192.240 721.960 202.760 722.280 ;
                RECT 1118.400 721.960 1123.120 722.280 ;
                RECT 2.880 723.320 182.360 723.640 ;
                RECT 192.240 723.320 202.760 723.640 ;
                RECT 1118.400 723.320 1123.120 723.640 ;
                RECT 2.880 724.680 202.760 725.000 ;
                RECT 1118.400 724.680 1123.120 725.000 ;
                RECT 2.880 726.040 182.360 726.360 ;
                RECT 192.240 726.040 202.760 726.360 ;
                RECT 1118.400 726.040 1123.120 726.360 ;
                RECT 2.880 727.400 182.360 727.720 ;
                RECT 192.240 727.400 202.760 727.720 ;
                RECT 1118.400 727.400 1123.120 727.720 ;
                RECT 2.880 728.760 185.760 729.080 ;
                RECT 192.240 728.760 202.760 729.080 ;
                RECT 1118.400 728.760 1123.120 729.080 ;
                RECT 2.880 730.120 186.440 730.440 ;
                RECT 192.240 730.120 202.760 730.440 ;
                RECT 1118.400 730.120 1123.120 730.440 ;
                RECT 2.880 731.480 182.360 731.800 ;
                RECT 192.240 731.480 202.760 731.800 ;
                RECT 1118.400 731.480 1123.120 731.800 ;
                RECT 2.880 732.840 202.760 733.160 ;
                RECT 1118.400 732.840 1123.120 733.160 ;
                RECT 2.880 734.200 182.360 734.520 ;
                RECT 192.240 734.200 202.760 734.520 ;
                RECT 1118.400 734.200 1123.120 734.520 ;
                RECT 2.880 735.560 182.360 735.880 ;
                RECT 192.240 735.560 202.760 735.880 ;
                RECT 1118.400 735.560 1123.120 735.880 ;
                RECT 2.880 736.920 182.360 737.240 ;
                RECT 192.240 736.920 202.760 737.240 ;
                RECT 1118.400 736.920 1123.120 737.240 ;
                RECT 2.880 738.280 188.480 738.600 ;
                RECT 192.240 738.280 202.760 738.600 ;
                RECT 1118.400 738.280 1123.120 738.600 ;
                RECT 2.880 739.640 202.760 739.960 ;
                RECT 1118.400 739.640 1123.120 739.960 ;
                RECT 2.880 741.000 188.480 741.320 ;
                RECT 192.240 741.000 202.760 741.320 ;
                RECT 1118.400 741.000 1123.120 741.320 ;
                RECT 2.880 742.360 182.360 742.680 ;
                RECT 192.240 742.360 202.760 742.680 ;
                RECT 1118.400 742.360 1123.120 742.680 ;
                RECT 2.880 743.720 182.360 744.040 ;
                RECT 192.240 743.720 202.760 744.040 ;
                RECT 1118.400 743.720 1123.120 744.040 ;
                RECT 2.880 745.080 182.360 745.400 ;
                RECT 192.240 745.080 202.760 745.400 ;
                RECT 1118.400 745.080 1123.120 745.400 ;
                RECT 2.880 746.440 182.360 746.760 ;
                RECT 192.240 746.440 202.760 746.760 ;
                RECT 1118.400 746.440 1123.120 746.760 ;
                RECT 2.880 747.800 202.760 748.120 ;
                RECT 1118.400 747.800 1123.120 748.120 ;
                RECT 2.880 749.160 183.040 749.480 ;
                RECT 192.240 749.160 202.760 749.480 ;
                RECT 1118.400 749.160 1123.120 749.480 ;
                RECT 2.880 750.520 182.360 750.840 ;
                RECT 192.240 750.520 202.760 750.840 ;
                RECT 1118.400 750.520 1123.120 750.840 ;
                RECT 2.880 751.880 182.360 752.200 ;
                RECT 192.240 751.880 202.760 752.200 ;
                RECT 1118.400 751.880 1123.120 752.200 ;
                RECT 2.880 753.240 182.360 753.560 ;
                RECT 192.240 753.240 202.760 753.560 ;
                RECT 1118.400 753.240 1123.120 753.560 ;
                RECT 2.880 754.600 182.360 754.920 ;
                RECT 192.240 754.600 202.760 754.920 ;
                RECT 1118.400 754.600 1123.120 754.920 ;
                RECT 2.880 755.960 202.760 756.280 ;
                RECT 1118.400 755.960 1123.120 756.280 ;
                RECT 2.880 757.320 182.360 757.640 ;
                RECT 192.240 757.320 202.760 757.640 ;
                RECT 1118.400 757.320 1123.120 757.640 ;
                RECT 2.880 758.680 185.080 759.000 ;
                RECT 192.240 758.680 202.760 759.000 ;
                RECT 1118.400 758.680 1123.120 759.000 ;
                RECT 2.880 760.040 182.360 760.360 ;
                RECT 192.240 760.040 202.760 760.360 ;
                RECT 1118.400 760.040 1123.120 760.360 ;
                RECT 2.880 761.400 182.360 761.720 ;
                RECT 192.240 761.400 202.760 761.720 ;
                RECT 1118.400 761.400 1123.120 761.720 ;
                RECT 2.880 762.760 182.360 763.080 ;
                RECT 192.240 762.760 202.760 763.080 ;
                RECT 1118.400 762.760 1123.120 763.080 ;
                RECT 2.880 764.120 202.760 764.440 ;
                RECT 1118.400 764.120 1123.120 764.440 ;
                RECT 2.880 765.480 182.360 765.800 ;
                RECT 192.240 765.480 202.760 765.800 ;
                RECT 1118.400 765.480 1123.120 765.800 ;
                RECT 2.880 766.840 182.360 767.160 ;
                RECT 192.240 766.840 202.760 767.160 ;
                RECT 1118.400 766.840 1123.120 767.160 ;
                RECT 2.880 768.200 187.800 768.520 ;
                RECT 192.240 768.200 202.760 768.520 ;
                RECT 1118.400 768.200 1123.120 768.520 ;
                RECT 2.880 769.560 182.360 769.880 ;
                RECT 192.240 769.560 202.760 769.880 ;
                RECT 1118.400 769.560 1123.120 769.880 ;
                RECT 2.880 770.920 182.360 771.240 ;
                RECT 192.240 770.920 202.760 771.240 ;
                RECT 1118.400 770.920 1123.120 771.240 ;
                RECT 2.880 772.280 202.760 772.600 ;
                RECT 1118.400 772.280 1123.120 772.600 ;
                RECT 2.880 773.640 182.360 773.960 ;
                RECT 192.240 773.640 202.760 773.960 ;
                RECT 1118.400 773.640 1123.120 773.960 ;
                RECT 2.880 775.000 182.360 775.320 ;
                RECT 192.240 775.000 202.760 775.320 ;
                RECT 1118.400 775.000 1123.120 775.320 ;
                RECT 2.880 776.360 182.360 776.680 ;
                RECT 192.240 776.360 202.760 776.680 ;
                RECT 1118.400 776.360 1123.120 776.680 ;
                RECT 2.880 777.720 190.520 778.040 ;
                RECT 192.240 777.720 202.760 778.040 ;
                RECT 1118.400 777.720 1123.120 778.040 ;
                RECT 2.880 779.080 182.360 779.400 ;
                RECT 192.240 779.080 202.760 779.400 ;
                RECT 1118.400 779.080 1123.120 779.400 ;
                RECT 2.880 780.440 202.760 780.760 ;
                RECT 1118.400 780.440 1123.120 780.760 ;
                RECT 2.880 781.800 401.320 782.120 ;
                RECT 1118.400 781.800 1123.120 782.120 ;
                RECT 2.880 783.160 401.320 783.480 ;
                RECT 1118.400 783.160 1123.120 783.480 ;
                RECT 2.880 784.520 401.320 784.840 ;
                RECT 1118.400 784.520 1123.120 784.840 ;
                RECT 2.880 785.880 1123.120 786.200 ;
                RECT 2.880 787.240 1123.120 787.560 ;
                RECT 2.880 788.600 1123.120 788.920 ;
                RECT 2.880 789.960 1123.120 790.280 ;
                RECT 2.880 2.880 1123.120 4.240 ;
                RECT 2.880 791.960 1123.120 793.320 ;
                RECT 405.460 32.185 411.260 33.305 ;
                RECT 1108.560 32.185 1114.360 33.305 ;
                RECT 405.460 38.005 411.260 38.695 ;
                RECT 1108.560 38.005 1114.360 38.695 ;
                RECT 405.460 43.580 411.260 44.370 ;
                RECT 1108.560 43.580 1114.360 44.370 ;
                RECT 405.460 49.700 411.260 50.280 ;
                RECT 1108.560 49.700 1114.360 50.280 ;
                RECT 405.460 54.420 411.260 55.010 ;
                RECT 1108.560 54.420 1114.360 55.010 ;
                RECT 405.460 59.240 411.260 59.830 ;
                RECT 1108.560 59.240 1114.360 59.830 ;
                RECT 405.460 192.230 1114.360 194.030 ;
                RECT 405.460 84.800 1114.360 85.600 ;
                RECT 405.460 95.800 1114.360 99.400 ;
                RECT 405.460 128.535 1114.360 128.825 ;
                RECT 405.460 81.790 1114.360 82.590 ;
                RECT 405.460 86.480 1114.360 87.280 ;
                RECT 405.460 72.740 1114.360 74.540 ;
                RECT 405.460 89.690 1114.360 90.490 ;
                RECT 405.460 22.815 1114.360 24.615 ;
                RECT 203.730 273.555 205.480 780.735 ;
                RECT 217.715 273.555 219.635 780.735 ;
                RECT 242.135 273.555 244.055 780.735 ;
                RECT 245.975 273.555 247.895 780.735 ;
                RECT 249.815 273.555 251.735 780.735 ;
                RECT 292.400 273.555 294.320 780.735 ;
                RECT 296.240 273.555 298.160 780.735 ;
                RECT 300.080 273.555 302.000 780.735 ;
                RECT 303.920 273.555 305.840 780.735 ;
                RECT 307.760 273.555 309.680 780.735 ;
                RECT 311.600 273.555 313.520 780.735 ;
                RECT 315.440 273.555 317.360 780.735 ;
                RECT 319.280 273.555 321.200 780.735 ;
                RECT 125.770 57.175 126.660 126.975 ;
                RECT 132.100 57.175 132.990 126.975 ;
                RECT 138.860 57.175 139.750 126.975 ;
                RECT 146.050 57.175 147.800 126.975 ;
                RECT 160.465 57.175 162.385 126.975 ;
                RECT 185.315 57.175 187.235 126.975 ;
                RECT 189.155 57.175 191.075 126.975 ;
                RECT 192.995 57.175 194.915 126.975 ;
                RECT 236.440 57.175 238.360 126.975 ;
                RECT 240.280 57.175 242.200 126.975 ;
                RECT 244.120 57.175 246.040 126.975 ;
                RECT 247.960 57.175 249.880 126.975 ;
                RECT 251.800 57.175 253.720 126.975 ;
                RECT 255.640 57.175 257.560 126.975 ;
                RECT 259.480 57.175 261.400 126.975 ;
                RECT 263.320 57.175 265.240 126.975 ;
                RECT 220.025 208.940 221.135 266.920 ;
                RECT 227.970 208.940 228.860 266.920 ;
                RECT 234.730 208.940 235.620 266.920 ;
                RECT 241.060 208.940 241.950 266.920 ;
                RECT 247.710 208.940 249.250 266.920 ;
                RECT 260.730 208.940 262.650 266.920 ;
                RECT 286.885 208.940 288.805 266.920 ;
                RECT 290.725 208.940 292.645 266.920 ;
                RECT 294.565 208.940 296.485 266.920 ;
                RECT 298.405 208.940 300.325 266.920 ;
                RECT 274.910 197.780 275.800 202.940 ;
                RECT 282.015 197.780 283.935 202.940 ;
                RECT 299.770 197.780 301.690 202.940 ;
                RECT 303.610 197.780 305.530 202.940 ;
                RECT 307.450 197.780 309.370 202.940 ;
                RECT 344.760 46.015 345.650 51.175 ;
                RECT 124.420 274.620 133.580 274.990 ;
                RECT 124.420 278.060 133.580 279.170 ;
                RECT 44.180 256.280 63.820 256.950 ;
                RECT 44.180 257.510 63.820 260.560 ;
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 1126.000 796.200 ;
        LAYER met2 ;
            RECT 0.000 0.000 1126.000 796.200 ;
    END 
END sram22_2048x64m8w8 
END LIBRARY 

