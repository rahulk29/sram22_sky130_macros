VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_256x8m8w1
    CLASS BLOCK  ;
    FOREIGN sram22_256x8m8w1   ;
    SIZE 261.720 BY 225.680 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.684800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 163.990 0.000 164.130 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.684800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 174.890 0.000 175.030 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.684800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 185.790 0.000 185.930 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.684800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 196.690 0.000 196.830 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.684800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 207.590 0.000 207.730 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.684800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 218.490 0.000 218.630 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.684800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 229.390 0.000 229.530 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.684800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 240.290 0.000 240.430 0.140 ; 
        END 
    END dout[7] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.636500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.406400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 163.570 0.000 163.710 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.636500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.406400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 174.470 0.000 174.610 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.636500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.406400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 185.370 0.000 185.510 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.636500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.406400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 196.270 0.000 196.410 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.636500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.406400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 207.170 0.000 207.310 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.636500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.406400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 218.070 0.000 218.210 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.636500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.406400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 228.970 0.000 229.110 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 4.636500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 5.406400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 239.870 0.000 240.010 0.140 ; 
        END 
    END din[7] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.446900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 163.220 0.000 163.360 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.446900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 174.120 0.000 174.260 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.446900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 185.020 0.000 185.160 0.140 ; 
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.446900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 195.920 0.000 196.060 0.140 ; 
        END 
    END wmask[3] 
    PIN wmask[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.446900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 206.820 0.000 206.960 0.140 ; 
        END 
    END wmask[4] 
    PIN wmask[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.446900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 217.720 0.000 217.860 0.140 ; 
        END 
    END wmask[5] 
    PIN wmask[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.446900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 228.620 0.000 228.760 0.140 ; 
        END 
    END wmask[6] 
    PIN wmask[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.446900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 239.520 0.000 239.660 0.140 ; 
        END 
    END wmask[7] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.855100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 107.920 0.000 108.240 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.855100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 101.800 0.000 102.120 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.855100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 95.680 0.000 96.000 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.855100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 89.560 0.000 89.880 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.855100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 84.120 0.000 84.440 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.855100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 78.000 0.000 78.320 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.855100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 71.880 0.000 72.200 0.320 ; 
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.855100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 65.760 0.000 66.080 0.320 ; 
        END 
    END addr[7] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.855100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 120.160 0.000 120.480 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.855100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 114.040 0.000 114.360 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 10.044000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 123.560 0.000 123.880 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 13.950000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 124.240 0.000 124.560 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 163.320 6.240 ; 
                RECT 165.040 5.920 174.200 6.240 ; 
                RECT 175.920 5.920 185.080 6.240 ; 
                RECT 186.800 5.920 195.960 6.240 ; 
                RECT 197.680 5.920 206.840 6.240 ; 
                RECT 208.560 5.920 217.720 6.240 ; 
                RECT 219.440 5.920 228.600 6.240 ; 
                RECT 230.320 5.920 239.480 6.240 ; 
                RECT 241.200 5.920 261.560 6.240 ; 
                RECT 0.160 7.280 261.560 7.600 ; 
                RECT 0.160 8.640 261.560 8.960 ; 
                RECT 0.160 10.000 123.200 10.320 ; 
                RECT 156.880 10.000 261.560 10.320 ; 
                RECT 0.160 11.360 261.560 11.680 ; 
                RECT 0.160 12.720 261.560 13.040 ; 
                RECT 0.160 14.080 61.320 14.400 ; 
                RECT 124.920 14.080 261.560 14.400 ; 
                RECT 0.160 15.440 162.640 15.760 ; 
                RECT 240.520 15.440 261.560 15.760 ; 
                RECT 0.160 16.800 150.400 17.120 ; 
                RECT 252.080 16.800 261.560 17.120 ; 
                RECT 0.160 18.160 61.320 18.480 ; 
                RECT 124.240 18.160 150.400 18.480 ; 
                RECT 252.080 18.160 261.560 18.480 ; 
                RECT 0.160 19.520 150.400 19.840 ; 
                RECT 252.080 19.520 261.560 19.840 ; 
                RECT 0.160 20.880 150.400 21.200 ; 
                RECT 252.080 20.880 261.560 21.200 ; 
                RECT 0.160 22.240 150.400 22.560 ; 
                RECT 252.080 22.240 261.560 22.560 ; 
                RECT 0.160 23.600 150.400 23.920 ; 
                RECT 252.080 23.600 261.560 23.920 ; 
                RECT 0.160 24.960 150.400 25.280 ; 
                RECT 252.080 24.960 261.560 25.280 ; 
                RECT 0.160 26.320 150.400 26.640 ; 
                RECT 252.080 26.320 261.560 26.640 ; 
                RECT 0.160 27.680 150.400 28.000 ; 
                RECT 252.080 27.680 261.560 28.000 ; 
                RECT 0.160 29.040 150.400 29.360 ; 
                RECT 252.080 29.040 261.560 29.360 ; 
                RECT 0.160 30.400 150.400 30.720 ; 
                RECT 252.080 30.400 261.560 30.720 ; 
                RECT 0.160 31.760 150.400 32.080 ; 
                RECT 252.080 31.760 261.560 32.080 ; 
                RECT 0.160 33.120 87.840 33.440 ; 
                RECT 95.680 33.120 150.400 33.440 ; 
                RECT 252.080 33.120 261.560 33.440 ; 
                RECT 0.160 34.480 86.480 34.800 ; 
                RECT 101.800 34.480 149.720 34.800 ; 
                RECT 252.080 34.480 261.560 34.800 ; 
                RECT 0.160 35.840 85.120 36.160 ; 
                RECT 107.920 35.840 150.400 36.160 ; 
                RECT 252.080 35.840 261.560 36.160 ; 
                RECT 0.160 37.200 65.400 37.520 ; 
                RECT 124.920 37.200 150.400 37.520 ; 
                RECT 252.080 37.200 261.560 37.520 ; 
                RECT 0.160 38.560 64.720 38.880 ; 
                RECT 120.840 38.560 150.400 38.880 ; 
                RECT 252.080 38.560 261.560 38.880 ; 
                RECT 0.160 39.920 150.400 40.240 ; 
                RECT 252.080 39.920 261.560 40.240 ; 
                RECT 0.160 41.280 150.400 41.600 ; 
                RECT 252.080 41.280 261.560 41.600 ; 
                RECT 0.160 42.640 150.400 42.960 ; 
                RECT 252.080 42.640 261.560 42.960 ; 
                RECT 0.160 44.000 150.400 44.320 ; 
                RECT 252.080 44.000 261.560 44.320 ; 
                RECT 0.160 45.360 60.640 45.680 ; 
                RECT 71.880 45.360 150.400 45.680 ; 
                RECT 252.080 45.360 261.560 45.680 ; 
                RECT 0.160 46.720 62.000 47.040 ; 
                RECT 67.800 46.720 75.600 47.040 ; 
                RECT 78.000 46.720 150.400 47.040 ; 
                RECT 252.080 46.720 261.560 47.040 ; 
                RECT 0.160 48.080 63.360 48.400 ; 
                RECT 67.120 48.080 150.400 48.400 ; 
                RECT 252.080 48.080 261.560 48.400 ; 
                RECT 0.160 49.440 150.400 49.760 ; 
                RECT 252.080 49.440 261.560 49.760 ; 
                RECT 0.160 50.800 70.160 51.120 ; 
                RECT 78.680 50.800 117.080 51.120 ; 
                RECT 122.880 50.800 150.400 51.120 ; 
                RECT 252.080 50.800 261.560 51.120 ; 
                RECT 0.160 52.160 62.680 52.480 ; 
                RECT 71.880 52.160 117.080 52.480 ; 
                RECT 252.080 52.160 261.560 52.480 ; 
                RECT 0.160 53.520 66.080 53.840 ; 
                RECT 71.200 53.520 117.080 53.840 ; 
                RECT 252.080 53.520 261.560 53.840 ; 
                RECT 0.160 54.880 117.080 55.200 ; 
                RECT 122.880 54.880 150.400 55.200 ; 
                RECT 252.080 54.880 261.560 55.200 ; 
                RECT 0.160 56.240 62.000 56.560 ; 
                RECT 71.880 56.240 117.080 56.560 ; 
                RECT 122.880 56.240 150.400 56.560 ; 
                RECT 252.080 56.240 261.560 56.560 ; 
                RECT 0.160 57.600 69.480 57.920 ; 
                RECT 78.000 57.600 150.400 57.920 ; 
                RECT 252.080 57.600 261.560 57.920 ; 
                RECT 0.160 58.960 150.400 59.280 ; 
                RECT 252.080 58.960 261.560 59.280 ; 
                RECT 0.160 60.320 70.160 60.640 ; 
                RECT 75.960 60.320 150.400 60.640 ; 
                RECT 252.080 60.320 261.560 60.640 ; 
                RECT 0.160 61.680 72.880 62.000 ; 
                RECT 78.000 61.680 99.400 62.000 ; 
                RECT 122.200 61.680 150.400 62.000 ; 
                RECT 252.080 61.680 261.560 62.000 ; 
                RECT 0.160 63.040 66.760 63.360 ; 
                RECT 71.880 63.040 85.800 63.360 ; 
                RECT 92.960 63.040 99.400 63.360 ; 
                RECT 122.200 63.040 150.400 63.360 ; 
                RECT 252.080 63.040 261.560 63.360 ; 
                RECT 0.160 64.400 87.160 64.720 ; 
                RECT 91.600 64.400 99.400 64.720 ; 
                RECT 131.720 64.400 150.400 64.720 ; 
                RECT 252.080 64.400 261.560 64.720 ; 
                RECT 0.160 65.760 60.640 66.080 ; 
                RECT 83.440 65.760 88.520 66.080 ; 
                RECT 90.920 65.760 99.400 66.080 ; 
                RECT 131.720 65.760 150.400 66.080 ; 
                RECT 252.080 65.760 261.560 66.080 ; 
                RECT 0.160 67.120 70.160 67.440 ; 
                RECT 78.000 67.120 99.400 67.440 ; 
                RECT 134.440 67.120 150.400 67.440 ; 
                RECT 252.080 67.120 261.560 67.440 ; 
                RECT 0.160 68.480 69.480 68.800 ; 
                RECT 71.880 68.480 79.000 68.800 ; 
                RECT 85.480 68.480 99.400 68.800 ; 
                RECT 133.080 68.480 150.400 68.800 ; 
                RECT 252.080 68.480 261.560 68.800 ; 
                RECT 0.160 69.840 60.640 70.160 ; 
                RECT 74.600 69.840 99.400 70.160 ; 
                RECT 134.440 69.840 150.400 70.160 ; 
                RECT 252.080 69.840 261.560 70.160 ; 
                RECT 0.160 71.200 69.480 71.520 ; 
                RECT 78.000 71.200 99.400 71.520 ; 
                RECT 122.200 71.200 150.400 71.520 ; 
                RECT 252.080 71.200 261.560 71.520 ; 
                RECT 0.160 72.560 67.440 72.880 ; 
                RECT 71.200 72.560 99.400 72.880 ; 
                RECT 137.160 72.560 150.400 72.880 ; 
                RECT 252.080 72.560 261.560 72.880 ; 
                RECT 0.160 73.920 62.680 74.240 ; 
                RECT 67.120 73.920 70.160 74.240 ; 
                RECT 78.680 73.920 99.400 74.240 ; 
                RECT 137.160 73.920 150.400 74.240 ; 
                RECT 252.080 73.920 261.560 74.240 ; 
                RECT 0.160 75.280 65.400 75.600 ; 
                RECT 69.160 75.280 99.400 75.600 ; 
                RECT 135.800 75.280 150.400 75.600 ; 
                RECT 252.080 75.280 261.560 75.600 ; 
                RECT 0.160 76.640 62.000 76.960 ; 
                RECT 65.760 76.640 99.400 76.960 ; 
                RECT 139.880 76.640 150.400 76.960 ; 
                RECT 252.080 76.640 261.560 76.960 ; 
                RECT 0.160 78.000 66.080 78.320 ; 
                RECT 71.880 78.000 99.400 78.320 ; 
                RECT 139.880 78.000 150.400 78.320 ; 
                RECT 252.080 78.000 261.560 78.320 ; 
                RECT 0.160 79.360 62.000 79.680 ; 
                RECT 77.320 79.360 99.400 79.680 ; 
                RECT 122.200 79.360 150.400 79.680 ; 
                RECT 252.080 79.360 261.560 79.680 ; 
                RECT 0.160 80.720 99.400 81.040 ; 
                RECT 142.600 80.720 150.400 81.040 ; 
                RECT 252.080 80.720 261.560 81.040 ; 
                RECT 0.160 82.080 69.480 82.400 ; 
                RECT 71.200 82.080 99.400 82.400 ; 
                RECT 141.240 82.080 150.400 82.400 ; 
                RECT 252.080 82.080 261.560 82.400 ; 
                RECT 0.160 83.440 70.160 83.760 ; 
                RECT 72.560 83.440 99.400 83.760 ; 
                RECT 142.600 83.440 150.400 83.760 ; 
                RECT 252.080 83.440 261.560 83.760 ; 
                RECT 0.160 84.800 60.640 85.120 ; 
                RECT 67.800 84.800 69.480 85.120 ; 
                RECT 71.200 84.800 99.400 85.120 ; 
                RECT 145.320 84.800 150.400 85.120 ; 
                RECT 252.080 84.800 261.560 85.120 ; 
                RECT 0.160 86.160 66.080 86.480 ; 
                RECT 78.000 86.160 99.400 86.480 ; 
                RECT 145.320 86.160 150.400 86.480 ; 
                RECT 252.080 86.160 261.560 86.480 ; 
                RECT 0.160 87.520 60.640 87.840 ; 
                RECT 71.880 87.520 99.400 87.840 ; 
                RECT 143.960 87.520 150.400 87.840 ; 
                RECT 252.080 87.520 261.560 87.840 ; 
                RECT 0.160 88.880 69.480 89.200 ; 
                RECT 72.560 88.880 99.400 89.200 ; 
                RECT 122.200 88.880 150.400 89.200 ; 
                RECT 252.080 88.880 261.560 89.200 ; 
                RECT 0.160 90.240 99.400 90.560 ; 
                RECT 146.680 90.240 150.400 90.560 ; 
                RECT 252.080 90.240 261.560 90.560 ; 
                RECT 0.160 91.600 99.400 91.920 ; 
                RECT 148.040 91.600 150.400 91.920 ; 
                RECT 252.080 91.600 261.560 91.920 ; 
                RECT 0.160 92.960 57.240 93.280 ; 
                RECT 74.600 92.960 99.400 93.280 ; 
                RECT 252.080 92.960 261.560 93.280 ; 
                RECT 0.160 94.320 99.400 94.640 ; 
                RECT 252.080 94.320 261.560 94.640 ; 
                RECT 0.160 95.680 99.400 96.000 ; 
                RECT 252.080 95.680 261.560 96.000 ; 
                RECT 0.160 97.040 66.080 97.360 ; 
                RECT 78.000 97.040 99.400 97.360 ; 
                RECT 122.200 97.040 150.400 97.360 ; 
                RECT 252.080 97.040 261.560 97.360 ; 
                RECT 0.160 98.400 72.880 98.720 ; 
                RECT 80.720 98.400 150.400 98.720 ; 
                RECT 252.080 98.400 261.560 98.720 ; 
                RECT 0.160 99.760 125.920 100.080 ; 
                RECT 252.080 99.760 261.560 100.080 ; 
                RECT 0.160 101.120 150.400 101.440 ; 
                RECT 252.080 101.120 261.560 101.440 ; 
                RECT 0.160 102.480 60.640 102.800 ; 
                RECT 65.760 102.480 144.960 102.800 ; 
                RECT 252.080 102.480 261.560 102.800 ; 
                RECT 0.160 103.840 142.240 104.160 ; 
                RECT 252.080 103.840 261.560 104.160 ; 
                RECT 0.160 105.200 139.520 105.520 ; 
                RECT 252.080 105.200 261.560 105.520 ; 
                RECT 0.160 106.560 76.280 106.880 ; 
                RECT 78.680 106.560 136.800 106.880 ; 
                RECT 252.080 106.560 261.560 106.880 ; 
                RECT 0.160 107.920 134.080 108.240 ; 
                RECT 252.080 107.920 261.560 108.240 ; 
                RECT 0.160 109.280 131.360 109.600 ; 
                RECT 252.080 109.280 261.560 109.600 ; 
                RECT 0.160 110.640 128.640 110.960 ; 
                RECT 252.080 110.640 261.560 110.960 ; 
                RECT 0.160 112.000 38.880 112.320 ; 
                RECT 57.600 112.000 62.680 112.320 ; 
                RECT 67.800 112.000 116.400 112.320 ; 
                RECT 122.200 112.000 150.400 112.320 ; 
                RECT 252.080 112.000 261.560 112.320 ; 
                RECT 0.160 113.360 38.880 113.680 ; 
                RECT 57.600 113.360 116.400 113.680 ; 
                RECT 122.200 113.360 150.400 113.680 ; 
                RECT 252.080 113.360 261.560 113.680 ; 
                RECT 0.160 114.720 38.880 115.040 ; 
                RECT 57.600 114.720 69.480 115.040 ; 
                RECT 78.000 114.720 116.400 115.040 ; 
                RECT 122.200 114.720 150.400 115.040 ; 
                RECT 252.080 114.720 261.560 115.040 ; 
                RECT 0.160 116.080 38.880 116.400 ; 
                RECT 57.600 116.080 116.400 116.400 ; 
                RECT 122.200 116.080 150.400 116.400 ; 
                RECT 252.080 116.080 261.560 116.400 ; 
                RECT 0.160 117.440 38.880 117.760 ; 
                RECT 57.600 117.440 65.400 117.760 ; 
                RECT 67.800 117.440 116.400 117.760 ; 
                RECT 122.200 117.440 150.400 117.760 ; 
                RECT 252.080 117.440 261.560 117.760 ; 
                RECT 0.160 118.800 38.880 119.120 ; 
                RECT 57.600 118.800 62.000 119.120 ; 
                RECT 65.080 118.800 150.400 119.120 ; 
                RECT 252.080 118.800 261.560 119.120 ; 
                RECT 0.160 120.160 38.880 120.480 ; 
                RECT 57.600 120.160 130.000 120.480 ; 
                RECT 252.080 120.160 261.560 120.480 ; 
                RECT 0.160 121.520 38.880 121.840 ; 
                RECT 57.600 121.520 130.000 121.840 ; 
                RECT 252.080 121.520 261.560 121.840 ; 
                RECT 0.160 122.880 38.880 123.200 ; 
                RECT 57.600 122.880 102.120 123.200 ; 
                RECT 122.200 122.880 132.720 123.200 ; 
                RECT 252.080 122.880 261.560 123.200 ; 
                RECT 0.160 124.240 38.880 124.560 ; 
                RECT 57.600 124.240 102.120 124.560 ; 
                RECT 122.200 124.240 138.160 124.560 ; 
                RECT 252.080 124.240 261.560 124.560 ; 
                RECT 0.160 125.600 38.880 125.920 ; 
                RECT 57.600 125.600 102.120 125.920 ; 
                RECT 122.200 125.600 140.880 125.920 ; 
                RECT 252.080 125.600 261.560 125.920 ; 
                RECT 0.160 126.960 102.120 127.280 ; 
                RECT 122.200 126.960 143.600 127.280 ; 
                RECT 252.080 126.960 261.560 127.280 ; 
                RECT 0.160 128.320 64.040 128.640 ; 
                RECT 67.800 128.320 102.120 128.640 ; 
                RECT 122.200 128.320 146.320 128.640 ; 
                RECT 252.080 128.320 261.560 128.640 ; 
                RECT 0.160 129.680 102.120 130.000 ; 
                RECT 122.200 129.680 149.040 130.000 ; 
                RECT 252.080 129.680 261.560 130.000 ; 
                RECT 0.160 131.040 22.560 131.360 ; 
                RECT 39.240 131.040 102.120 131.360 ; 
                RECT 252.080 131.040 261.560 131.360 ; 
                RECT 0.160 132.400 22.560 132.720 ; 
                RECT 39.240 132.400 66.080 132.720 ; 
                RECT 72.560 132.400 102.120 132.720 ; 
                RECT 122.200 132.400 150.400 132.720 ; 
                RECT 252.080 132.400 261.560 132.720 ; 
                RECT 0.160 133.760 22.560 134.080 ; 
                RECT 39.240 133.760 45.000 134.080 ; 
                RECT 52.840 133.760 102.120 134.080 ; 
                RECT 122.200 133.760 150.400 134.080 ; 
                RECT 252.080 133.760 261.560 134.080 ; 
                RECT 0.160 135.120 22.560 135.440 ; 
                RECT 56.920 135.120 102.120 135.440 ; 
                RECT 122.200 135.120 150.400 135.440 ; 
                RECT 252.080 135.120 261.560 135.440 ; 
                RECT 0.160 136.480 22.560 136.800 ; 
                RECT 56.920 136.480 102.120 136.800 ; 
                RECT 252.080 136.480 261.560 136.800 ; 
                RECT 0.160 137.840 22.560 138.160 ; 
                RECT 39.240 137.840 45.000 138.160 ; 
                RECT 52.840 137.840 60.640 138.160 ; 
                RECT 70.520 137.840 102.120 138.160 ; 
                RECT 252.080 137.840 261.560 138.160 ; 
                RECT 0.160 139.200 17.120 139.520 ; 
                RECT 52.160 139.200 102.120 139.520 ; 
                RECT 122.200 139.200 261.560 139.520 ; 
                RECT 0.160 140.560 51.800 140.880 ; 
                RECT 99.760 140.560 261.560 140.880 ; 
                RECT 0.160 141.920 147.680 142.240 ; 
                RECT 254.800 141.920 261.560 142.240 ; 
                RECT 0.160 143.280 147.680 143.600 ; 
                RECT 254.800 143.280 261.560 143.600 ; 
                RECT 0.160 144.640 147.680 144.960 ; 
                RECT 254.800 144.640 261.560 144.960 ; 
                RECT 0.160 146.000 56.560 146.320 ; 
                RECT 63.040 146.000 64.720 146.320 ; 
                RECT 75.960 146.000 106.200 146.320 ; 
                RECT 254.800 146.000 261.560 146.320 ; 
                RECT 0.160 147.360 54.520 147.680 ; 
                RECT 75.280 147.360 89.200 147.680 ; 
                RECT 95.000 147.360 106.200 147.680 ; 
                RECT 254.800 147.360 261.560 147.680 ; 
                RECT 0.160 148.720 54.520 149.040 ; 
                RECT 74.600 148.720 87.160 149.040 ; 
                RECT 95.000 148.720 106.200 149.040 ; 
                RECT 254.800 148.720 261.560 149.040 ; 
                RECT 0.160 150.080 54.520 150.400 ; 
                RECT 65.080 150.080 87.160 150.400 ; 
                RECT 90.920 150.080 106.200 150.400 ; 
                RECT 254.800 150.080 261.560 150.400 ; 
                RECT 0.160 151.440 87.160 151.760 ; 
                RECT 95.000 151.440 106.200 151.760 ; 
                RECT 254.800 151.440 261.560 151.760 ; 
                RECT 0.160 152.800 54.520 153.120 ; 
                RECT 65.080 152.800 87.160 153.120 ; 
                RECT 95.000 152.800 106.200 153.120 ; 
                RECT 254.800 152.800 261.560 153.120 ; 
                RECT 0.160 154.160 54.520 154.480 ; 
                RECT 65.080 154.160 106.200 154.480 ; 
                RECT 254.800 154.160 261.560 154.480 ; 
                RECT 0.160 155.520 91.240 155.840 ; 
                RECT 95.000 155.520 106.200 155.840 ; 
                RECT 254.800 155.520 261.560 155.840 ; 
                RECT 0.160 156.880 87.160 157.200 ; 
                RECT 95.000 156.880 106.200 157.200 ; 
                RECT 254.800 156.880 261.560 157.200 ; 
                RECT 0.160 158.240 87.160 158.560 ; 
                RECT 95.000 158.240 106.200 158.560 ; 
                RECT 254.800 158.240 261.560 158.560 ; 
                RECT 0.160 159.600 17.120 159.920 ; 
                RECT 50.120 159.600 63.360 159.920 ; 
                RECT 65.760 159.600 87.160 159.920 ; 
                RECT 88.880 159.600 106.200 159.920 ; 
                RECT 254.800 159.600 261.560 159.920 ; 
                RECT 0.160 160.960 16.440 161.280 ; 
                RECT 50.120 160.960 63.360 161.280 ; 
                RECT 66.440 160.960 87.160 161.280 ; 
                RECT 95.000 160.960 106.200 161.280 ; 
                RECT 254.800 160.960 261.560 161.280 ; 
                RECT 0.160 162.320 15.760 162.640 ; 
                RECT 50.120 162.320 106.200 162.640 ; 
                RECT 254.800 162.320 261.560 162.640 ; 
                RECT 0.160 163.680 15.080 164.000 ; 
                RECT 50.120 163.680 89.200 164.000 ; 
                RECT 95.000 163.680 106.200 164.000 ; 
                RECT 254.800 163.680 261.560 164.000 ; 
                RECT 0.160 165.040 87.160 165.360 ; 
                RECT 95.000 165.040 106.200 165.360 ; 
                RECT 254.800 165.040 261.560 165.360 ; 
                RECT 0.160 166.400 14.400 166.720 ; 
                RECT 50.120 166.400 87.160 166.720 ; 
                RECT 95.000 166.400 106.200 166.720 ; 
                RECT 254.800 166.400 261.560 166.720 ; 
                RECT 0.160 167.760 13.720 168.080 ; 
                RECT 50.120 167.760 87.160 168.080 ; 
                RECT 95.000 167.760 106.200 168.080 ; 
                RECT 254.800 167.760 261.560 168.080 ; 
                RECT 0.160 169.120 87.160 169.440 ; 
                RECT 93.640 169.120 106.200 169.440 ; 
                RECT 254.800 169.120 261.560 169.440 ; 
                RECT 0.160 170.480 13.040 170.800 ; 
                RECT 50.120 170.480 106.200 170.800 ; 
                RECT 254.800 170.480 261.560 170.800 ; 
                RECT 0.160 171.840 12.360 172.160 ; 
                RECT 50.120 171.840 63.360 172.160 ; 
                RECT 67.120 171.840 87.160 172.160 ; 
                RECT 95.000 171.840 106.200 172.160 ; 
                RECT 254.800 171.840 261.560 172.160 ; 
                RECT 0.160 173.200 87.160 173.520 ; 
                RECT 95.000 173.200 106.200 173.520 ; 
                RECT 254.800 173.200 261.560 173.520 ; 
                RECT 0.160 174.560 11.680 174.880 ; 
                RECT 50.120 174.560 63.360 174.880 ; 
                RECT 66.440 174.560 87.160 174.880 ; 
                RECT 95.000 174.560 106.200 174.880 ; 
                RECT 254.800 174.560 261.560 174.880 ; 
                RECT 0.160 175.920 11.000 176.240 ; 
                RECT 50.120 175.920 63.360 176.240 ; 
                RECT 65.760 175.920 87.160 176.240 ; 
                RECT 95.000 175.920 106.200 176.240 ; 
                RECT 254.800 175.920 261.560 176.240 ; 
                RECT 0.160 177.280 87.160 177.600 ; 
                RECT 94.320 177.280 106.200 177.600 ; 
                RECT 254.800 177.280 261.560 177.600 ; 
                RECT 0.160 178.640 89.200 178.960 ; 
                RECT 95.000 178.640 106.200 178.960 ; 
                RECT 254.800 178.640 261.560 178.960 ; 
                RECT 0.160 180.000 106.200 180.320 ; 
                RECT 254.800 180.000 261.560 180.320 ; 
                RECT 0.160 181.360 89.880 181.680 ; 
                RECT 95.000 181.360 106.200 181.680 ; 
                RECT 254.800 181.360 261.560 181.680 ; 
                RECT 0.160 182.720 90.560 183.040 ; 
                RECT 95.000 182.720 106.200 183.040 ; 
                RECT 254.800 182.720 261.560 183.040 ; 
                RECT 0.160 184.080 90.560 184.400 ; 
                RECT 95.000 184.080 106.200 184.400 ; 
                RECT 254.800 184.080 261.560 184.400 ; 
                RECT 0.160 185.440 66.760 185.760 ; 
                RECT 75.280 185.440 106.200 185.760 ; 
                RECT 254.800 185.440 261.560 185.760 ; 
                RECT 0.160 186.800 65.400 187.120 ; 
                RECT 74.600 186.800 87.160 187.120 ; 
                RECT 95.000 186.800 106.200 187.120 ; 
                RECT 254.800 186.800 261.560 187.120 ; 
                RECT 0.160 188.160 87.160 188.480 ; 
                RECT 95.000 188.160 106.200 188.480 ; 
                RECT 254.800 188.160 261.560 188.480 ; 
                RECT 0.160 189.520 87.160 189.840 ; 
                RECT 89.560 189.520 106.200 189.840 ; 
                RECT 254.800 189.520 261.560 189.840 ; 
                RECT 0.160 190.880 87.160 191.200 ; 
                RECT 95.000 190.880 106.200 191.200 ; 
                RECT 254.800 190.880 261.560 191.200 ; 
                RECT 0.160 192.240 87.160 192.560 ; 
                RECT 95.000 192.240 106.200 192.560 ; 
                RECT 254.800 192.240 261.560 192.560 ; 
                RECT 0.160 193.600 87.160 193.920 ; 
                RECT 90.240 193.600 106.200 193.920 ; 
                RECT 254.800 193.600 261.560 193.920 ; 
                RECT 0.160 194.960 89.200 195.280 ; 
                RECT 95.000 194.960 106.200 195.280 ; 
                RECT 254.800 194.960 261.560 195.280 ; 
                RECT 0.160 196.320 89.880 196.640 ; 
                RECT 95.000 196.320 106.200 196.640 ; 
                RECT 254.800 196.320 261.560 196.640 ; 
                RECT 0.160 197.680 90.560 198.000 ; 
                RECT 95.000 197.680 106.200 198.000 ; 
                RECT 254.800 197.680 261.560 198.000 ; 
                RECT 0.160 199.040 106.200 199.360 ; 
                RECT 254.800 199.040 261.560 199.360 ; 
                RECT 0.160 200.400 90.560 200.720 ; 
                RECT 95.000 200.400 106.200 200.720 ; 
                RECT 254.800 200.400 261.560 200.720 ; 
                RECT 0.160 201.760 106.200 202.080 ; 
                RECT 254.800 201.760 261.560 202.080 ; 
                RECT 0.160 203.120 91.240 203.440 ; 
                RECT 95.000 203.120 106.200 203.440 ; 
                RECT 254.800 203.120 261.560 203.440 ; 
                RECT 0.160 204.480 91.920 204.800 ; 
                RECT 95.000 204.480 106.200 204.800 ; 
                RECT 254.800 204.480 261.560 204.800 ; 
                RECT 0.160 205.840 91.920 206.160 ; 
                RECT 95.000 205.840 106.200 206.160 ; 
                RECT 254.800 205.840 261.560 206.160 ; 
                RECT 0.160 207.200 92.600 207.520 ; 
                RECT 95.000 207.200 106.200 207.520 ; 
                RECT 254.800 207.200 261.560 207.520 ; 
                RECT 0.160 208.560 106.200 208.880 ; 
                RECT 254.800 208.560 261.560 208.880 ; 
                RECT 0.160 209.920 106.200 210.240 ; 
                RECT 254.800 209.920 261.560 210.240 ; 
                RECT 0.160 211.280 147.680 211.600 ; 
                RECT 254.800 211.280 261.560 211.600 ; 
                RECT 0.160 212.640 147.680 212.960 ; 
                RECT 254.800 212.640 261.560 212.960 ; 
                RECT 0.160 214.000 147.680 214.320 ; 
                RECT 254.800 214.000 261.560 214.320 ; 
                RECT 0.160 215.360 261.560 215.680 ; 
                RECT 0.160 216.720 261.560 217.040 ; 
                RECT 0.160 218.080 261.560 218.400 ; 
                RECT 0.160 219.440 261.560 219.760 ; 
                RECT 0.160 0.160 261.560 1.520 ; 
                RECT 0.160 224.160 261.560 225.520 ; 
                RECT 151.820 37.975 157.620 39.345 ; 
                RECT 244.520 37.975 250.320 39.345 ; 
                RECT 151.820 42.245 157.620 43.015 ; 
                RECT 244.520 42.245 250.320 43.015 ; 
                RECT 151.820 45.660 157.620 46.480 ; 
                RECT 244.520 45.660 250.320 46.480 ; 
                RECT 151.820 49.150 157.620 49.970 ; 
                RECT 244.520 49.150 250.320 49.970 ; 
                RECT 151.820 86.365 250.320 86.655 ; 
                RECT 151.820 70.870 250.320 71.670 ; 
                RECT 151.820 82.075 250.320 83.145 ; 
                RECT 151.820 113.670 250.320 114.640 ; 
                RECT 151.820 75.760 250.320 76.560 ; 
                RECT 151.820 67.860 250.320 68.660 ; 
                RECT 151.820 133.920 250.320 135.270 ; 
                RECT 151.820 56.390 250.320 58.190 ; 
                RECT 151.820 22.220 250.320 24.020 ; 
                RECT 111.590 145.715 113.510 210.495 ; 
                RECT 115.430 145.715 117.350 210.495 ; 
                RECT 128.715 145.715 130.635 210.495 ; 
                RECT 132.555 145.715 134.475 210.495 ; 
                RECT 136.395 145.715 138.315 210.495 ; 
                RECT 140.235 145.715 142.155 210.495 ; 
                RECT 144.075 145.715 145.995 210.495 ; 
                RECT 102.735 61.965 104.275 97.365 ; 
                RECT 110.595 61.965 112.515 97.365 ; 
                RECT 119.290 61.965 121.210 97.365 ; 
                RECT 106.180 123.440 108.100 139.080 ; 
                RECT 113.155 123.440 115.075 139.080 ; 
                RECT 119.915 123.440 121.835 139.080 ; 
                RECT 119.915 112.280 121.835 117.440 ; 
                RECT 120.215 50.805 121.965 55.965 ; 
                RECT 55.210 147.985 64.370 148.735 ; 
                RECT 55.210 152.740 64.370 154.660 ; 
                RECT 40.360 135.770 56.400 136.570 ; 
                RECT 23.560 135.125 38.400 138.175 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 163.320 5.560 ; 
                RECT 165.040 5.240 174.200 5.560 ; 
                RECT 175.920 5.240 185.080 5.560 ; 
                RECT 186.800 5.240 195.960 5.560 ; 
                RECT 197.680 5.240 206.840 5.560 ; 
                RECT 208.560 5.240 217.720 5.560 ; 
                RECT 219.440 5.240 228.600 5.560 ; 
                RECT 230.320 5.240 239.480 5.560 ; 
                RECT 241.200 5.240 258.840 5.560 ; 
                RECT 2.880 6.600 258.840 6.920 ; 
                RECT 2.880 7.960 258.840 8.280 ; 
                RECT 2.880 9.320 123.880 9.640 ; 
                RECT 156.200 9.320 258.840 9.640 ; 
                RECT 2.880 10.680 258.840 11.000 ; 
                RECT 2.880 12.040 258.840 12.360 ; 
                RECT 2.880 13.400 61.320 13.720 ; 
                RECT 124.920 13.400 258.840 13.720 ; 
                RECT 2.880 14.760 258.840 15.080 ; 
                RECT 2.880 16.120 150.400 16.440 ; 
                RECT 252.080 16.120 258.840 16.440 ; 
                RECT 2.880 17.480 61.320 17.800 ; 
                RECT 124.240 17.480 150.400 17.800 ; 
                RECT 252.080 17.480 258.840 17.800 ; 
                RECT 2.880 18.840 150.400 19.160 ; 
                RECT 252.080 18.840 258.840 19.160 ; 
                RECT 2.880 20.200 150.400 20.520 ; 
                RECT 252.080 20.200 258.840 20.520 ; 
                RECT 2.880 21.560 150.400 21.880 ; 
                RECT 252.080 21.560 258.840 21.880 ; 
                RECT 2.880 22.920 150.400 23.240 ; 
                RECT 252.080 22.920 258.840 23.240 ; 
                RECT 2.880 24.280 150.400 24.600 ; 
                RECT 252.080 24.280 258.840 24.600 ; 
                RECT 2.880 25.640 150.400 25.960 ; 
                RECT 252.080 25.640 258.840 25.960 ; 
                RECT 2.880 27.000 150.400 27.320 ; 
                RECT 252.080 27.000 258.840 27.320 ; 
                RECT 2.880 28.360 150.400 28.680 ; 
                RECT 252.080 28.360 258.840 28.680 ; 
                RECT 2.880 29.720 150.400 30.040 ; 
                RECT 252.080 29.720 258.840 30.040 ; 
                RECT 2.880 31.080 150.400 31.400 ; 
                RECT 252.080 31.080 258.840 31.400 ; 
                RECT 2.880 32.440 88.520 32.760 ; 
                RECT 97.040 32.440 150.400 32.760 ; 
                RECT 252.080 32.440 258.840 32.760 ; 
                RECT 2.880 33.800 87.160 34.120 ; 
                RECT 103.160 33.800 149.720 34.120 ; 
                RECT 252.080 33.800 258.840 34.120 ; 
                RECT 2.880 35.160 85.800 35.480 ; 
                RECT 109.280 35.160 150.400 35.480 ; 
                RECT 252.080 35.160 258.840 35.480 ; 
                RECT 2.880 36.520 62.680 36.840 ; 
                RECT 124.240 36.520 150.400 36.840 ; 
                RECT 252.080 36.520 258.840 36.840 ; 
                RECT 2.880 37.880 63.360 38.200 ; 
                RECT 114.720 37.880 150.400 38.200 ; 
                RECT 252.080 37.880 258.840 38.200 ; 
                RECT 2.880 39.240 150.400 39.560 ; 
                RECT 252.080 39.240 258.840 39.560 ; 
                RECT 2.880 40.600 150.400 40.920 ; 
                RECT 252.080 40.600 258.840 40.920 ; 
                RECT 2.880 41.960 150.400 42.280 ; 
                RECT 252.080 41.960 258.840 42.280 ; 
                RECT 2.880 43.320 150.400 43.640 ; 
                RECT 252.080 43.320 258.840 43.640 ; 
                RECT 2.880 44.680 60.640 45.000 ; 
                RECT 71.880 44.680 150.400 45.000 ; 
                RECT 252.080 44.680 258.840 45.000 ; 
                RECT 2.880 46.040 62.000 46.360 ; 
                RECT 64.400 46.040 150.400 46.360 ; 
                RECT 252.080 46.040 258.840 46.360 ; 
                RECT 2.880 47.400 63.360 47.720 ; 
                RECT 67.800 47.400 75.600 47.720 ; 
                RECT 78.000 47.400 150.400 47.720 ; 
                RECT 252.080 47.400 258.840 47.720 ; 
                RECT 2.880 48.760 63.360 49.080 ; 
                RECT 67.120 48.760 150.400 49.080 ; 
                RECT 252.080 48.760 258.840 49.080 ; 
                RECT 2.880 50.120 70.160 50.440 ; 
                RECT 78.680 50.120 150.400 50.440 ; 
                RECT 252.080 50.120 258.840 50.440 ; 
                RECT 2.880 51.480 65.400 51.800 ; 
                RECT 71.880 51.480 117.080 51.800 ; 
                RECT 122.880 51.480 150.400 51.800 ; 
                RECT 252.080 51.480 258.840 51.800 ; 
                RECT 2.880 52.840 62.680 53.160 ; 
                RECT 71.880 52.840 117.080 53.160 ; 
                RECT 252.080 52.840 258.840 53.160 ; 
                RECT 2.880 54.200 117.080 54.520 ; 
                RECT 252.080 54.200 258.840 54.520 ; 
                RECT 2.880 55.560 62.000 55.880 ; 
                RECT 71.880 55.560 83.760 55.880 ; 
                RECT 114.040 55.560 117.080 55.880 ; 
                RECT 122.880 55.560 150.400 55.880 ; 
                RECT 252.080 55.560 258.840 55.880 ; 
                RECT 2.880 56.920 70.160 57.240 ; 
                RECT 78.000 56.920 150.400 57.240 ; 
                RECT 252.080 56.920 258.840 57.240 ; 
                RECT 2.880 58.280 69.480 58.600 ; 
                RECT 71.880 58.280 150.400 58.600 ; 
                RECT 252.080 58.280 258.840 58.600 ; 
                RECT 2.880 59.640 150.400 59.960 ; 
                RECT 252.080 59.640 258.840 59.960 ; 
                RECT 2.880 61.000 70.160 61.320 ; 
                RECT 78.000 61.000 150.400 61.320 ; 
                RECT 252.080 61.000 258.840 61.320 ; 
                RECT 2.880 62.360 66.760 62.680 ; 
                RECT 71.880 62.360 85.120 62.680 ; 
                RECT 92.960 62.360 99.400 62.680 ; 
                RECT 122.200 62.360 150.400 62.680 ; 
                RECT 252.080 62.360 258.840 62.680 ; 
                RECT 2.880 63.720 69.480 64.040 ; 
                RECT 71.880 63.720 86.480 64.040 ; 
                RECT 92.280 63.720 99.400 64.040 ; 
                RECT 131.720 63.720 150.400 64.040 ; 
                RECT 252.080 63.720 258.840 64.040 ; 
                RECT 2.880 65.080 87.840 65.400 ; 
                RECT 91.600 65.080 99.400 65.400 ; 
                RECT 131.720 65.080 150.400 65.400 ; 
                RECT 252.080 65.080 258.840 65.400 ; 
                RECT 2.880 66.440 60.640 66.760 ; 
                RECT 83.440 66.440 99.400 66.760 ; 
                RECT 130.360 66.440 150.400 66.760 ; 
                RECT 252.080 66.440 258.840 66.760 ; 
                RECT 2.880 67.800 79.000 68.120 ; 
                RECT 84.800 67.800 99.400 68.120 ; 
                RECT 134.440 67.800 150.400 68.120 ; 
                RECT 252.080 67.800 258.840 68.120 ; 
                RECT 2.880 69.160 69.480 69.480 ; 
                RECT 71.880 69.160 81.720 69.480 ; 
                RECT 85.480 69.160 99.400 69.480 ; 
                RECT 134.440 69.160 150.400 69.480 ; 
                RECT 252.080 69.160 258.840 69.480 ; 
                RECT 2.880 70.520 60.640 70.840 ; 
                RECT 74.600 70.520 99.400 70.840 ; 
                RECT 133.080 70.520 150.400 70.840 ; 
                RECT 252.080 70.520 258.840 70.840 ; 
                RECT 2.880 71.880 69.480 72.200 ; 
                RECT 78.000 71.880 99.400 72.200 ; 
                RECT 137.160 71.880 150.400 72.200 ; 
                RECT 252.080 71.880 258.840 72.200 ; 
                RECT 2.880 73.240 67.440 73.560 ; 
                RECT 78.680 73.240 99.400 73.560 ; 
                RECT 135.800 73.240 150.400 73.560 ; 
                RECT 252.080 73.240 258.840 73.560 ; 
                RECT 2.880 74.600 62.680 74.920 ; 
                RECT 69.160 74.600 99.400 74.920 ; 
                RECT 137.160 74.600 150.400 74.920 ; 
                RECT 252.080 74.600 258.840 74.920 ; 
                RECT 2.880 75.960 99.400 76.280 ; 
                RECT 139.880 75.960 150.400 76.280 ; 
                RECT 252.080 75.960 258.840 76.280 ; 
                RECT 2.880 77.320 62.000 77.640 ; 
                RECT 65.760 77.320 99.400 77.640 ; 
                RECT 138.520 77.320 150.400 77.640 ; 
                RECT 252.080 77.320 258.840 77.640 ; 
                RECT 2.880 78.680 62.000 79.000 ; 
                RECT 71.880 78.680 99.400 79.000 ; 
                RECT 139.880 78.680 150.400 79.000 ; 
                RECT 252.080 78.680 258.840 79.000 ; 
                RECT 2.880 80.040 66.080 80.360 ; 
                RECT 77.320 80.040 99.400 80.360 ; 
                RECT 122.200 80.040 150.400 80.360 ; 
                RECT 252.080 80.040 258.840 80.360 ; 
                RECT 2.880 81.400 69.480 81.720 ; 
                RECT 71.200 81.400 99.400 81.720 ; 
                RECT 142.600 81.400 150.400 81.720 ; 
                RECT 252.080 81.400 258.840 81.720 ; 
                RECT 2.880 82.760 70.160 83.080 ; 
                RECT 72.560 82.760 99.400 83.080 ; 
                RECT 142.600 82.760 150.400 83.080 ; 
                RECT 252.080 82.760 258.840 83.080 ; 
                RECT 2.880 84.120 99.400 84.440 ; 
                RECT 122.200 84.120 150.400 84.440 ; 
                RECT 252.080 84.120 258.840 84.440 ; 
                RECT 2.880 85.480 60.640 85.800 ; 
                RECT 78.000 85.480 99.400 85.800 ; 
                RECT 143.960 85.480 150.400 85.800 ; 
                RECT 252.080 85.480 258.840 85.800 ; 
                RECT 2.880 86.840 60.640 87.160 ; 
                RECT 71.880 86.840 76.280 87.160 ; 
                RECT 78.000 86.840 99.400 87.160 ; 
                RECT 145.320 86.840 150.400 87.160 ; 
                RECT 252.080 86.840 258.840 87.160 ; 
                RECT 2.880 88.200 69.480 88.520 ; 
                RECT 72.560 88.200 99.400 88.520 ; 
                RECT 122.200 88.200 150.400 88.520 ; 
                RECT 252.080 88.200 258.840 88.520 ; 
                RECT 2.880 89.560 99.400 89.880 ; 
                RECT 148.040 89.560 150.400 89.880 ; 
                RECT 252.080 89.560 258.840 89.880 ; 
                RECT 2.880 90.920 99.400 91.240 ; 
                RECT 148.040 90.920 150.400 91.240 ; 
                RECT 252.080 90.920 258.840 91.240 ; 
                RECT 2.880 92.280 57.240 92.600 ; 
                RECT 70.520 92.280 99.400 92.600 ; 
                RECT 146.680 92.280 150.400 92.600 ; 
                RECT 252.080 92.280 258.840 92.600 ; 
                RECT 2.880 93.640 67.440 93.960 ; 
                RECT 74.600 93.640 99.400 93.960 ; 
                RECT 252.080 93.640 258.840 93.960 ; 
                RECT 2.880 95.000 99.400 95.320 ; 
                RECT 252.080 95.000 258.840 95.320 ; 
                RECT 2.880 96.360 99.400 96.680 ; 
                RECT 252.080 96.360 258.840 96.680 ; 
                RECT 2.880 97.720 66.080 98.040 ; 
                RECT 80.720 97.720 99.400 98.040 ; 
                RECT 122.200 97.720 150.400 98.040 ; 
                RECT 252.080 97.720 258.840 98.040 ; 
                RECT 2.880 99.080 150.400 99.400 ; 
                RECT 252.080 99.080 258.840 99.400 ; 
                RECT 2.880 100.440 125.920 100.760 ; 
                RECT 252.080 100.440 258.840 100.760 ; 
                RECT 2.880 101.800 62.680 102.120 ; 
                RECT 65.760 101.800 147.680 102.120 ; 
                RECT 252.080 101.800 258.840 102.120 ; 
                RECT 2.880 103.160 60.640 103.480 ; 
                RECT 64.400 103.160 144.960 103.480 ; 
                RECT 252.080 103.160 258.840 103.480 ; 
                RECT 2.880 104.520 142.240 104.840 ; 
                RECT 252.080 104.520 258.840 104.840 ; 
                RECT 2.880 105.880 76.280 106.200 ; 
                RECT 78.680 105.880 139.520 106.200 ; 
                RECT 252.080 105.880 258.840 106.200 ; 
                RECT 2.880 107.240 136.800 107.560 ; 
                RECT 252.080 107.240 258.840 107.560 ; 
                RECT 2.880 108.600 134.080 108.920 ; 
                RECT 252.080 108.600 258.840 108.920 ; 
                RECT 2.880 109.960 128.640 110.280 ; 
                RECT 252.080 109.960 258.840 110.280 ; 
                RECT 2.880 111.320 62.680 111.640 ; 
                RECT 67.800 111.320 128.640 111.640 ; 
                RECT 252.080 111.320 258.840 111.640 ; 
                RECT 2.880 112.680 38.880 113.000 ; 
                RECT 57.600 112.680 84.440 113.000 ; 
                RECT 122.200 112.680 150.400 113.000 ; 
                RECT 252.080 112.680 258.840 113.000 ; 
                RECT 2.880 114.040 38.880 114.360 ; 
                RECT 57.600 114.040 69.480 114.360 ; 
                RECT 78.000 114.040 116.400 114.360 ; 
                RECT 122.200 114.040 150.400 114.360 ; 
                RECT 252.080 114.040 258.840 114.360 ; 
                RECT 2.880 115.400 38.880 115.720 ; 
                RECT 57.600 115.400 116.400 115.720 ; 
                RECT 122.200 115.400 150.400 115.720 ; 
                RECT 252.080 115.400 258.840 115.720 ; 
                RECT 2.880 116.760 38.880 117.080 ; 
                RECT 57.600 116.760 65.400 117.080 ; 
                RECT 67.800 116.760 116.400 117.080 ; 
                RECT 122.200 116.760 150.400 117.080 ; 
                RECT 252.080 116.760 258.840 117.080 ; 
                RECT 2.880 118.120 38.880 118.440 ; 
                RECT 58.280 118.120 62.000 118.440 ; 
                RECT 65.080 118.120 150.400 118.440 ; 
                RECT 252.080 118.120 258.840 118.440 ; 
                RECT 2.880 119.480 38.880 119.800 ; 
                RECT 57.600 119.480 150.400 119.800 ; 
                RECT 252.080 119.480 258.840 119.800 ; 
                RECT 2.880 120.840 38.880 121.160 ; 
                RECT 57.600 120.840 130.000 121.160 ; 
                RECT 252.080 120.840 258.840 121.160 ; 
                RECT 2.880 122.200 38.880 122.520 ; 
                RECT 57.600 122.200 132.720 122.520 ; 
                RECT 252.080 122.200 258.840 122.520 ; 
                RECT 2.880 123.560 38.880 123.880 ; 
                RECT 57.600 123.560 102.120 123.880 ; 
                RECT 122.200 123.560 135.440 123.880 ; 
                RECT 252.080 123.560 258.840 123.880 ; 
                RECT 2.880 124.920 38.880 125.240 ; 
                RECT 57.600 124.920 102.120 125.240 ; 
                RECT 122.200 124.920 138.160 125.240 ; 
                RECT 252.080 124.920 258.840 125.240 ; 
                RECT 2.880 126.280 38.880 126.600 ; 
                RECT 57.600 126.280 102.120 126.600 ; 
                RECT 122.200 126.280 140.880 126.600 ; 
                RECT 252.080 126.280 258.840 126.600 ; 
                RECT 2.880 127.640 64.040 127.960 ; 
                RECT 67.800 127.640 102.120 127.960 ; 
                RECT 122.200 127.640 143.600 127.960 ; 
                RECT 252.080 127.640 258.840 127.960 ; 
                RECT 2.880 129.000 102.120 129.320 ; 
                RECT 122.200 129.000 146.320 129.320 ; 
                RECT 252.080 129.000 258.840 129.320 ; 
                RECT 2.880 130.360 22.560 130.680 ; 
                RECT 39.240 130.360 102.120 130.680 ; 
                RECT 252.080 130.360 258.840 130.680 ; 
                RECT 2.880 131.720 22.560 132.040 ; 
                RECT 39.240 131.720 102.120 132.040 ; 
                RECT 252.080 131.720 258.840 132.040 ; 
                RECT 2.880 133.080 22.560 133.400 ; 
                RECT 39.240 133.080 66.080 133.400 ; 
                RECT 72.560 133.080 102.120 133.400 ; 
                RECT 122.200 133.080 150.400 133.400 ; 
                RECT 252.080 133.080 258.840 133.400 ; 
                RECT 2.880 134.440 22.560 134.760 ; 
                RECT 39.240 134.440 45.000 134.760 ; 
                RECT 52.840 134.440 102.120 134.760 ; 
                RECT 122.200 134.440 150.400 134.760 ; 
                RECT 252.080 134.440 258.840 134.760 ; 
                RECT 2.880 135.800 22.560 136.120 ; 
                RECT 56.920 135.800 102.120 136.120 ; 
                RECT 122.200 135.800 150.400 136.120 ; 
                RECT 252.080 135.800 258.840 136.120 ; 
                RECT 2.880 137.160 22.560 137.480 ; 
                RECT 39.240 137.160 102.120 137.480 ; 
                RECT 252.080 137.160 258.840 137.480 ; 
                RECT 2.880 138.520 17.120 138.840 ; 
                RECT 52.840 138.520 60.640 138.840 ; 
                RECT 70.520 138.520 102.120 138.840 ; 
                RECT 122.200 138.520 150.400 138.840 ; 
                RECT 252.080 138.520 258.840 138.840 ; 
                RECT 2.880 139.880 45.000 140.200 ; 
                RECT 65.080 139.880 258.840 140.200 ; 
                RECT 2.880 141.240 61.320 141.560 ; 
                RECT 64.400 141.240 258.840 141.560 ; 
                RECT 2.880 142.600 147.680 142.920 ; 
                RECT 254.800 142.600 258.840 142.920 ; 
                RECT 2.880 143.960 147.680 144.280 ; 
                RECT 254.800 143.960 258.840 144.280 ; 
                RECT 2.880 145.320 56.560 145.640 ; 
                RECT 63.040 145.320 106.200 145.640 ; 
                RECT 254.800 145.320 258.840 145.640 ; 
                RECT 2.880 146.680 54.520 147.000 ; 
                RECT 75.960 146.680 106.200 147.000 ; 
                RECT 254.800 146.680 258.840 147.000 ; 
                RECT 2.880 148.040 54.520 148.360 ; 
                RECT 74.600 148.040 87.160 148.360 ; 
                RECT 95.000 148.040 106.200 148.360 ; 
                RECT 254.800 148.040 258.840 148.360 ; 
                RECT 2.880 149.400 68.120 149.720 ; 
                RECT 73.920 149.400 87.160 149.720 ; 
                RECT 95.000 149.400 106.200 149.720 ; 
                RECT 254.800 149.400 258.840 149.720 ; 
                RECT 2.880 150.760 54.520 151.080 ; 
                RECT 65.080 150.760 87.160 151.080 ; 
                RECT 95.000 150.760 106.200 151.080 ; 
                RECT 254.800 150.760 258.840 151.080 ; 
                RECT 2.880 152.120 54.520 152.440 ; 
                RECT 65.080 152.120 87.160 152.440 ; 
                RECT 95.000 152.120 106.200 152.440 ; 
                RECT 254.800 152.120 258.840 152.440 ; 
                RECT 2.880 153.480 54.520 153.800 ; 
                RECT 65.080 153.480 87.160 153.800 ; 
                RECT 91.600 153.480 106.200 153.800 ; 
                RECT 254.800 153.480 258.840 153.800 ; 
                RECT 2.880 154.840 54.520 155.160 ; 
                RECT 65.080 154.840 106.200 155.160 ; 
                RECT 254.800 154.840 258.840 155.160 ; 
                RECT 2.880 156.200 87.160 156.520 ; 
                RECT 95.000 156.200 106.200 156.520 ; 
                RECT 254.800 156.200 258.840 156.520 ; 
                RECT 2.880 157.560 87.160 157.880 ; 
                RECT 95.000 157.560 106.200 157.880 ; 
                RECT 254.800 157.560 258.840 157.880 ; 
                RECT 2.880 158.920 17.120 159.240 ; 
                RECT 50.120 158.920 91.920 159.240 ; 
                RECT 95.000 158.920 106.200 159.240 ; 
                RECT 254.800 158.920 258.840 159.240 ; 
                RECT 2.880 160.280 16.440 160.600 ; 
                RECT 50.120 160.280 87.160 160.600 ; 
                RECT 95.000 160.280 106.200 160.600 ; 
                RECT 254.800 160.280 258.840 160.600 ; 
                RECT 2.880 161.640 87.160 161.960 ; 
                RECT 92.280 161.640 106.200 161.960 ; 
                RECT 254.800 161.640 258.840 161.960 ; 
                RECT 2.880 163.000 15.760 163.320 ; 
                RECT 50.120 163.000 63.360 163.320 ; 
                RECT 67.120 163.000 89.200 163.320 ; 
                RECT 95.000 163.000 106.200 163.320 ; 
                RECT 254.800 163.000 258.840 163.320 ; 
                RECT 2.880 164.360 15.080 164.680 ; 
                RECT 50.120 164.360 63.360 164.680 ; 
                RECT 67.800 164.360 87.160 164.680 ; 
                RECT 88.880 164.360 106.200 164.680 ; 
                RECT 254.800 164.360 258.840 164.680 ; 
                RECT 2.880 165.720 87.160 166.040 ; 
                RECT 92.960 165.720 106.200 166.040 ; 
                RECT 254.800 165.720 258.840 166.040 ; 
                RECT 2.880 167.080 14.400 167.400 ; 
                RECT 50.120 167.080 63.360 167.400 ; 
                RECT 68.480 167.080 87.160 167.400 ; 
                RECT 95.000 167.080 106.200 167.400 ; 
                RECT 254.800 167.080 258.840 167.400 ; 
                RECT 2.880 168.440 13.720 168.760 ; 
                RECT 50.120 168.440 63.360 168.760 ; 
                RECT 69.160 168.440 87.160 168.760 ; 
                RECT 95.000 168.440 106.200 168.760 ; 
                RECT 254.800 168.440 258.840 168.760 ; 
                RECT 2.880 169.800 13.040 170.120 ; 
                RECT 50.120 169.800 63.360 170.120 ; 
                RECT 67.800 169.800 87.160 170.120 ; 
                RECT 93.640 169.800 106.200 170.120 ; 
                RECT 254.800 169.800 258.840 170.120 ; 
                RECT 2.880 171.160 12.360 171.480 ; 
                RECT 50.120 171.160 91.240 171.480 ; 
                RECT 95.000 171.160 106.200 171.480 ; 
                RECT 254.800 171.160 258.840 171.480 ; 
                RECT 2.880 172.520 87.160 172.840 ; 
                RECT 95.000 172.520 106.200 172.840 ; 
                RECT 254.800 172.520 258.840 172.840 ; 
                RECT 2.880 173.880 11.680 174.200 ; 
                RECT 50.120 173.880 87.160 174.200 ; 
                RECT 93.640 173.880 106.200 174.200 ; 
                RECT 254.800 173.880 258.840 174.200 ; 
                RECT 2.880 175.240 11.000 175.560 ; 
                RECT 50.120 175.240 87.160 175.560 ; 
                RECT 88.880 175.240 106.200 175.560 ; 
                RECT 254.800 175.240 258.840 175.560 ; 
                RECT 2.880 176.600 87.160 176.920 ; 
                RECT 95.000 176.600 106.200 176.920 ; 
                RECT 254.800 176.600 258.840 176.920 ; 
                RECT 2.880 177.960 106.200 178.280 ; 
                RECT 254.800 177.960 258.840 178.280 ; 
                RECT 2.880 179.320 89.200 179.640 ; 
                RECT 95.000 179.320 106.200 179.640 ; 
                RECT 254.800 179.320 258.840 179.640 ; 
                RECT 2.880 180.680 89.880 181.000 ; 
                RECT 95.000 180.680 106.200 181.000 ; 
                RECT 254.800 180.680 258.840 181.000 ; 
                RECT 2.880 182.040 90.560 182.360 ; 
                RECT 95.000 182.040 106.200 182.360 ; 
                RECT 254.800 182.040 258.840 182.360 ; 
                RECT 2.880 183.400 90.560 183.720 ; 
                RECT 95.000 183.400 106.200 183.720 ; 
                RECT 254.800 183.400 258.840 183.720 ; 
                RECT 2.880 184.760 106.200 185.080 ; 
                RECT 254.800 184.760 258.840 185.080 ; 
                RECT 2.880 186.120 66.080 186.440 ; 
                RECT 75.280 186.120 106.200 186.440 ; 
                RECT 254.800 186.120 258.840 186.440 ; 
                RECT 2.880 187.480 64.720 187.800 ; 
                RECT 73.920 187.480 87.160 187.800 ; 
                RECT 95.000 187.480 106.200 187.800 ; 
                RECT 254.800 187.480 258.840 187.800 ; 
                RECT 2.880 188.840 87.160 189.160 ; 
                RECT 95.000 188.840 106.200 189.160 ; 
                RECT 254.800 188.840 258.840 189.160 ; 
                RECT 2.880 190.200 87.160 190.520 ; 
                RECT 95.000 190.200 106.200 190.520 ; 
                RECT 254.800 190.200 258.840 190.520 ; 
                RECT 2.880 191.560 87.160 191.880 ; 
                RECT 95.000 191.560 106.200 191.880 ; 
                RECT 254.800 191.560 258.840 191.880 ; 
                RECT 2.880 192.920 87.160 193.240 ; 
                RECT 90.240 192.920 106.200 193.240 ; 
                RECT 254.800 192.920 258.840 193.240 ; 
                RECT 2.880 194.280 106.200 194.600 ; 
                RECT 254.800 194.280 258.840 194.600 ; 
                RECT 2.880 195.640 89.200 195.960 ; 
                RECT 95.000 195.640 106.200 195.960 ; 
                RECT 254.800 195.640 258.840 195.960 ; 
                RECT 2.880 197.000 89.880 197.320 ; 
                RECT 95.000 197.000 106.200 197.320 ; 
                RECT 254.800 197.000 258.840 197.320 ; 
                RECT 2.880 198.360 90.560 198.680 ; 
                RECT 95.000 198.360 106.200 198.680 ; 
                RECT 254.800 198.360 258.840 198.680 ; 
                RECT 2.880 199.720 90.560 200.040 ; 
                RECT 95.000 199.720 106.200 200.040 ; 
                RECT 254.800 199.720 258.840 200.040 ; 
                RECT 2.880 201.080 106.200 201.400 ; 
                RECT 254.800 201.080 258.840 201.400 ; 
                RECT 2.880 202.440 91.240 202.760 ; 
                RECT 95.000 202.440 106.200 202.760 ; 
                RECT 254.800 202.440 258.840 202.760 ; 
                RECT 2.880 203.800 106.200 204.120 ; 
                RECT 254.800 203.800 258.840 204.120 ; 
                RECT 2.880 205.160 91.920 205.480 ; 
                RECT 95.000 205.160 106.200 205.480 ; 
                RECT 254.800 205.160 258.840 205.480 ; 
                RECT 2.880 206.520 91.920 206.840 ; 
                RECT 95.000 206.520 106.200 206.840 ; 
                RECT 254.800 206.520 258.840 206.840 ; 
                RECT 2.880 207.880 92.600 208.200 ; 
                RECT 95.000 207.880 106.200 208.200 ; 
                RECT 254.800 207.880 258.840 208.200 ; 
                RECT 2.880 209.240 106.200 209.560 ; 
                RECT 254.800 209.240 258.840 209.560 ; 
                RECT 2.880 210.600 106.200 210.920 ; 
                RECT 254.800 210.600 258.840 210.920 ; 
                RECT 2.880 211.960 147.680 212.280 ; 
                RECT 254.800 211.960 258.840 212.280 ; 
                RECT 2.880 213.320 147.680 213.640 ; 
                RECT 254.800 213.320 258.840 213.640 ; 
                RECT 2.880 214.680 258.840 215.000 ; 
                RECT 2.880 216.040 258.840 216.360 ; 
                RECT 2.880 217.400 258.840 217.720 ; 
                RECT 2.880 218.760 258.840 219.080 ; 
                RECT 2.880 220.120 258.840 220.440 ; 
                RECT 2.880 2.880 258.840 4.240 ; 
                RECT 2.880 221.440 258.840 222.800 ; 
                RECT 151.820 35.330 157.620 36.450 ; 
                RECT 244.520 35.330 250.320 36.450 ; 
                RECT 151.820 41.000 157.620 41.390 ; 
                RECT 244.520 41.000 250.320 41.390 ; 
                RECT 151.820 44.375 157.620 44.775 ; 
                RECT 244.520 44.375 250.320 44.775 ; 
                RECT 151.820 47.865 157.620 48.265 ; 
                RECT 244.520 47.865 250.320 48.265 ; 
                RECT 151.820 80.205 250.320 81.275 ; 
                RECT 151.820 118.150 250.320 118.520 ; 
                RECT 151.820 98.925 250.320 99.215 ; 
                RECT 151.820 72.190 250.320 72.990 ; 
                RECT 151.820 77.080 250.320 77.880 ; 
                RECT 151.820 73.870 250.320 74.670 ; 
                RECT 151.820 69.180 250.320 69.980 ; 
                RECT 151.820 60.130 250.320 61.930 ; 
                RECT 151.820 25.960 250.320 27.760 ; 
                RECT 106.930 145.715 108.850 210.495 ; 
                RECT 120.585 145.715 122.505 210.495 ; 
                RECT 124.425 145.715 126.345 210.495 ; 
                RECT 100.350 61.965 101.240 97.365 ; 
                RECT 106.465 61.965 107.785 97.365 ; 
                RECT 115.695 61.965 116.805 97.365 ; 
                RECT 103.015 123.440 104.125 139.080 ; 
                RECT 110.530 123.440 111.420 139.080 ; 
                RECT 117.290 123.440 118.180 139.080 ; 
                RECT 117.290 112.280 118.180 117.440 ; 
                RECT 117.720 50.805 118.610 55.965 ; 
                RECT 55.210 146.780 64.370 147.150 ; 
                RECT 55.210 150.115 64.370 151.005 ; 
                RECT 23.560 130.840 38.400 131.510 ; 
                RECT 23.560 132.105 38.400 134.135 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 261.720 225.680 ; 
        LAYER met2 ;
            RECT 0.000 0.000 261.720 225.680 ; 
    END 
END sram22_256x8m8w1 
END LIBRARY 

