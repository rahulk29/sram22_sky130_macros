VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_256x128m4w8
    CLASS BLOCK  ;
    FOREIGN sram22_256x128m4w8   ;
    SIZE 1085.880 BY 313.400 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 292.150 0.000 292.290 0.140 ;
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 298.250 0.000 298.390 0.140 ;
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 304.350 0.000 304.490 0.140 ;
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 310.450 0.000 310.590 0.140 ;
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 316.550 0.000 316.690 0.140 ;
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 322.650 0.000 322.790 0.140 ;
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 328.750 0.000 328.890 0.140 ;
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 334.850 0.000 334.990 0.140 ;
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 340.950 0.000 341.090 0.140 ;
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 347.050 0.000 347.190 0.140 ;
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 353.150 0.000 353.290 0.140 ;
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 359.250 0.000 359.390 0.140 ;
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 365.350 0.000 365.490 0.140 ;
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 371.450 0.000 371.590 0.140 ;
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 377.550 0.000 377.690 0.140 ;
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 383.650 0.000 383.790 0.140 ;
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 389.750 0.000 389.890 0.140 ;
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 395.850 0.000 395.990 0.140 ;
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 401.950 0.000 402.090 0.140 ;
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 408.050 0.000 408.190 0.140 ;
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 414.150 0.000 414.290 0.140 ;
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 420.250 0.000 420.390 0.140 ;
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 426.350 0.000 426.490 0.140 ;
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 432.450 0.000 432.590 0.140 ;
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 438.550 0.000 438.690 0.140 ;
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 444.650 0.000 444.790 0.140 ;
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 450.750 0.000 450.890 0.140 ;
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 456.850 0.000 456.990 0.140 ;
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 462.950 0.000 463.090 0.140 ;
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 469.050 0.000 469.190 0.140 ;
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 475.150 0.000 475.290 0.140 ;
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 481.250 0.000 481.390 0.140 ;
        END 
    END dout[31] 
    PIN dout[32] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 487.350 0.000 487.490 0.140 ;
        END 
    END dout[32] 
    PIN dout[33] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 493.450 0.000 493.590 0.140 ;
        END 
    END dout[33] 
    PIN dout[34] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 499.550 0.000 499.690 0.140 ;
        END 
    END dout[34] 
    PIN dout[35] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 505.650 0.000 505.790 0.140 ;
        END 
    END dout[35] 
    PIN dout[36] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 511.750 0.000 511.890 0.140 ;
        END 
    END dout[36] 
    PIN dout[37] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 517.850 0.000 517.990 0.140 ;
        END 
    END dout[37] 
    PIN dout[38] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 523.950 0.000 524.090 0.140 ;
        END 
    END dout[38] 
    PIN dout[39] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 530.050 0.000 530.190 0.140 ;
        END 
    END dout[39] 
    PIN dout[40] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 536.150 0.000 536.290 0.140 ;
        END 
    END dout[40] 
    PIN dout[41] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 542.250 0.000 542.390 0.140 ;
        END 
    END dout[41] 
    PIN dout[42] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 548.350 0.000 548.490 0.140 ;
        END 
    END dout[42] 
    PIN dout[43] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 554.450 0.000 554.590 0.140 ;
        END 
    END dout[43] 
    PIN dout[44] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 560.550 0.000 560.690 0.140 ;
        END 
    END dout[44] 
    PIN dout[45] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 566.650 0.000 566.790 0.140 ;
        END 
    END dout[45] 
    PIN dout[46] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 572.750 0.000 572.890 0.140 ;
        END 
    END dout[46] 
    PIN dout[47] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 578.850 0.000 578.990 0.140 ;
        END 
    END dout[47] 
    PIN dout[48] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 584.950 0.000 585.090 0.140 ;
        END 
    END dout[48] 
    PIN dout[49] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 591.050 0.000 591.190 0.140 ;
        END 
    END dout[49] 
    PIN dout[50] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 597.150 0.000 597.290 0.140 ;
        END 
    END dout[50] 
    PIN dout[51] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 603.250 0.000 603.390 0.140 ;
        END 
    END dout[51] 
    PIN dout[52] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 609.350 0.000 609.490 0.140 ;
        END 
    END dout[52] 
    PIN dout[53] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 615.450 0.000 615.590 0.140 ;
        END 
    END dout[53] 
    PIN dout[54] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 621.550 0.000 621.690 0.140 ;
        END 
    END dout[54] 
    PIN dout[55] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 627.650 0.000 627.790 0.140 ;
        END 
    END dout[55] 
    PIN dout[56] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 633.750 0.000 633.890 0.140 ;
        END 
    END dout[56] 
    PIN dout[57] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 639.850 0.000 639.990 0.140 ;
        END 
    END dout[57] 
    PIN dout[58] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 645.950 0.000 646.090 0.140 ;
        END 
    END dout[58] 
    PIN dout[59] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 652.050 0.000 652.190 0.140 ;
        END 
    END dout[59] 
    PIN dout[60] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 658.150 0.000 658.290 0.140 ;
        END 
    END dout[60] 
    PIN dout[61] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 664.250 0.000 664.390 0.140 ;
        END 
    END dout[61] 
    PIN dout[62] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 670.350 0.000 670.490 0.140 ;
        END 
    END dout[62] 
    PIN dout[63] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 676.450 0.000 676.590 0.140 ;
        END 
    END dout[63] 
    PIN dout[64] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 682.550 0.000 682.690 0.140 ;
        END 
    END dout[64] 
    PIN dout[65] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 688.650 0.000 688.790 0.140 ;
        END 
    END dout[65] 
    PIN dout[66] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 694.750 0.000 694.890 0.140 ;
        END 
    END dout[66] 
    PIN dout[67] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 700.850 0.000 700.990 0.140 ;
        END 
    END dout[67] 
    PIN dout[68] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 706.950 0.000 707.090 0.140 ;
        END 
    END dout[68] 
    PIN dout[69] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 713.050 0.000 713.190 0.140 ;
        END 
    END dout[69] 
    PIN dout[70] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 719.150 0.000 719.290 0.140 ;
        END 
    END dout[70] 
    PIN dout[71] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 725.250 0.000 725.390 0.140 ;
        END 
    END dout[71] 
    PIN dout[72] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 731.350 0.000 731.490 0.140 ;
        END 
    END dout[72] 
    PIN dout[73] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 737.450 0.000 737.590 0.140 ;
        END 
    END dout[73] 
    PIN dout[74] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 743.550 0.000 743.690 0.140 ;
        END 
    END dout[74] 
    PIN dout[75] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 749.650 0.000 749.790 0.140 ;
        END 
    END dout[75] 
    PIN dout[76] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 755.750 0.000 755.890 0.140 ;
        END 
    END dout[76] 
    PIN dout[77] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 761.850 0.000 761.990 0.140 ;
        END 
    END dout[77] 
    PIN dout[78] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 767.950 0.000 768.090 0.140 ;
        END 
    END dout[78] 
    PIN dout[79] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 774.050 0.000 774.190 0.140 ;
        END 
    END dout[79] 
    PIN dout[80] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 780.150 0.000 780.290 0.140 ;
        END 
    END dout[80] 
    PIN dout[81] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 786.250 0.000 786.390 0.140 ;
        END 
    END dout[81] 
    PIN dout[82] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 792.350 0.000 792.490 0.140 ;
        END 
    END dout[82] 
    PIN dout[83] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 798.450 0.000 798.590 0.140 ;
        END 
    END dout[83] 
    PIN dout[84] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 804.550 0.000 804.690 0.140 ;
        END 
    END dout[84] 
    PIN dout[85] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 810.650 0.000 810.790 0.140 ;
        END 
    END dout[85] 
    PIN dout[86] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 816.750 0.000 816.890 0.140 ;
        END 
    END dout[86] 
    PIN dout[87] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 822.850 0.000 822.990 0.140 ;
        END 
    END dout[87] 
    PIN dout[88] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 828.950 0.000 829.090 0.140 ;
        END 
    END dout[88] 
    PIN dout[89] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 835.050 0.000 835.190 0.140 ;
        END 
    END dout[89] 
    PIN dout[90] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 841.150 0.000 841.290 0.140 ;
        END 
    END dout[90] 
    PIN dout[91] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 847.250 0.000 847.390 0.140 ;
        END 
    END dout[91] 
    PIN dout[92] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 853.350 0.000 853.490 0.140 ;
        END 
    END dout[92] 
    PIN dout[93] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 859.450 0.000 859.590 0.140 ;
        END 
    END dout[93] 
    PIN dout[94] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 865.550 0.000 865.690 0.140 ;
        END 
    END dout[94] 
    PIN dout[95] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 871.650 0.000 871.790 0.140 ;
        END 
    END dout[95] 
    PIN dout[96] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 877.750 0.000 877.890 0.140 ;
        END 
    END dout[96] 
    PIN dout[97] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 883.850 0.000 883.990 0.140 ;
        END 
    END dout[97] 
    PIN dout[98] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 889.950 0.000 890.090 0.140 ;
        END 
    END dout[98] 
    PIN dout[99] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 896.050 0.000 896.190 0.140 ;
        END 
    END dout[99] 
    PIN dout[100] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 902.150 0.000 902.290 0.140 ;
        END 
    END dout[100] 
    PIN dout[101] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 908.250 0.000 908.390 0.140 ;
        END 
    END dout[101] 
    PIN dout[102] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 914.350 0.000 914.490 0.140 ;
        END 
    END dout[102] 
    PIN dout[103] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 920.450 0.000 920.590 0.140 ;
        END 
    END dout[103] 
    PIN dout[104] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 926.550 0.000 926.690 0.140 ;
        END 
    END dout[104] 
    PIN dout[105] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 932.650 0.000 932.790 0.140 ;
        END 
    END dout[105] 
    PIN dout[106] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 938.750 0.000 938.890 0.140 ;
        END 
    END dout[106] 
    PIN dout[107] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 944.850 0.000 944.990 0.140 ;
        END 
    END dout[107] 
    PIN dout[108] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 950.950 0.000 951.090 0.140 ;
        END 
    END dout[108] 
    PIN dout[109] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 957.050 0.000 957.190 0.140 ;
        END 
    END dout[109] 
    PIN dout[110] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 963.150 0.000 963.290 0.140 ;
        END 
    END dout[110] 
    PIN dout[111] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 969.250 0.000 969.390 0.140 ;
        END 
    END dout[111] 
    PIN dout[112] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 975.350 0.000 975.490 0.140 ;
        END 
    END dout[112] 
    PIN dout[113] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 981.450 0.000 981.590 0.140 ;
        END 
    END dout[113] 
    PIN dout[114] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 987.550 0.000 987.690 0.140 ;
        END 
    END dout[114] 
    PIN dout[115] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 993.650 0.000 993.790 0.140 ;
        END 
    END dout[115] 
    PIN dout[116] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 999.750 0.000 999.890 0.140 ;
        END 
    END dout[116] 
    PIN dout[117] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1005.850 0.000 1005.990 0.140 ;
        END 
    END dout[117] 
    PIN dout[118] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1011.950 0.000 1012.090 0.140 ;
        END 
    END dout[118] 
    PIN dout[119] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1018.050 0.000 1018.190 0.140 ;
        END 
    END dout[119] 
    PIN dout[120] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1024.150 0.000 1024.290 0.140 ;
        END 
    END dout[120] 
    PIN dout[121] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1030.250 0.000 1030.390 0.140 ;
        END 
    END dout[121] 
    PIN dout[122] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1036.350 0.000 1036.490 0.140 ;
        END 
    END dout[122] 
    PIN dout[123] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1042.450 0.000 1042.590 0.140 ;
        END 
    END dout[123] 
    PIN dout[124] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1048.550 0.000 1048.690 0.140 ;
        END 
    END dout[124] 
    PIN dout[125] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1054.650 0.000 1054.790 0.140 ;
        END 
    END dout[125] 
    PIN dout[126] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1060.750 0.000 1060.890 0.140 ;
        END 
    END dout[126] 
    PIN dout[127] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.636400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1066.850 0.000 1066.990 0.140 ;
        END 
    END dout[127] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 291.730 0.000 291.870 0.140 ;
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 297.830 0.000 297.970 0.140 ;
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 303.930 0.000 304.070 0.140 ;
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 310.030 0.000 310.170 0.140 ;
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 316.130 0.000 316.270 0.140 ;
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 322.230 0.000 322.370 0.140 ;
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 328.330 0.000 328.470 0.140 ;
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 334.430 0.000 334.570 0.140 ;
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 340.530 0.000 340.670 0.140 ;
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 346.630 0.000 346.770 0.140 ;
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 352.730 0.000 352.870 0.140 ;
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 358.830 0.000 358.970 0.140 ;
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 364.930 0.000 365.070 0.140 ;
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 371.030 0.000 371.170 0.140 ;
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 377.130 0.000 377.270 0.140 ;
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 383.230 0.000 383.370 0.140 ;
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 389.330 0.000 389.470 0.140 ;
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 395.430 0.000 395.570 0.140 ;
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 401.530 0.000 401.670 0.140 ;
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 407.630 0.000 407.770 0.140 ;
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 413.730 0.000 413.870 0.140 ;
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 419.830 0.000 419.970 0.140 ;
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 425.930 0.000 426.070 0.140 ;
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 432.030 0.000 432.170 0.140 ;
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 438.130 0.000 438.270 0.140 ;
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 444.230 0.000 444.370 0.140 ;
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 450.330 0.000 450.470 0.140 ;
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 456.430 0.000 456.570 0.140 ;
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 462.530 0.000 462.670 0.140 ;
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 468.630 0.000 468.770 0.140 ;
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 474.730 0.000 474.870 0.140 ;
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 480.830 0.000 480.970 0.140 ;
        END 
    END din[31] 
    PIN din[32] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 486.930 0.000 487.070 0.140 ;
        END 
    END din[32] 
    PIN din[33] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 493.030 0.000 493.170 0.140 ;
        END 
    END din[33] 
    PIN din[34] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 499.130 0.000 499.270 0.140 ;
        END 
    END din[34] 
    PIN din[35] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 505.230 0.000 505.370 0.140 ;
        END 
    END din[35] 
    PIN din[36] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 511.330 0.000 511.470 0.140 ;
        END 
    END din[36] 
    PIN din[37] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 517.430 0.000 517.570 0.140 ;
        END 
    END din[37] 
    PIN din[38] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 523.530 0.000 523.670 0.140 ;
        END 
    END din[38] 
    PIN din[39] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 529.630 0.000 529.770 0.140 ;
        END 
    END din[39] 
    PIN din[40] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 535.730 0.000 535.870 0.140 ;
        END 
    END din[40] 
    PIN din[41] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 541.830 0.000 541.970 0.140 ;
        END 
    END din[41] 
    PIN din[42] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 547.930 0.000 548.070 0.140 ;
        END 
    END din[42] 
    PIN din[43] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 554.030 0.000 554.170 0.140 ;
        END 
    END din[43] 
    PIN din[44] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 560.130 0.000 560.270 0.140 ;
        END 
    END din[44] 
    PIN din[45] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 566.230 0.000 566.370 0.140 ;
        END 
    END din[45] 
    PIN din[46] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 572.330 0.000 572.470 0.140 ;
        END 
    END din[46] 
    PIN din[47] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 578.430 0.000 578.570 0.140 ;
        END 
    END din[47] 
    PIN din[48] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 584.530 0.000 584.670 0.140 ;
        END 
    END din[48] 
    PIN din[49] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 590.630 0.000 590.770 0.140 ;
        END 
    END din[49] 
    PIN din[50] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 596.730 0.000 596.870 0.140 ;
        END 
    END din[50] 
    PIN din[51] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 602.830 0.000 602.970 0.140 ;
        END 
    END din[51] 
    PIN din[52] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 608.930 0.000 609.070 0.140 ;
        END 
    END din[52] 
    PIN din[53] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 615.030 0.000 615.170 0.140 ;
        END 
    END din[53] 
    PIN din[54] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 621.130 0.000 621.270 0.140 ;
        END 
    END din[54] 
    PIN din[55] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 627.230 0.000 627.370 0.140 ;
        END 
    END din[55] 
    PIN din[56] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 633.330 0.000 633.470 0.140 ;
        END 
    END din[56] 
    PIN din[57] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 639.430 0.000 639.570 0.140 ;
        END 
    END din[57] 
    PIN din[58] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 645.530 0.000 645.670 0.140 ;
        END 
    END din[58] 
    PIN din[59] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 651.630 0.000 651.770 0.140 ;
        END 
    END din[59] 
    PIN din[60] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 657.730 0.000 657.870 0.140 ;
        END 
    END din[60] 
    PIN din[61] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 663.830 0.000 663.970 0.140 ;
        END 
    END din[61] 
    PIN din[62] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 669.930 0.000 670.070 0.140 ;
        END 
    END din[62] 
    PIN din[63] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 676.030 0.000 676.170 0.140 ;
        END 
    END din[63] 
    PIN din[64] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 682.130 0.000 682.270 0.140 ;
        END 
    END din[64] 
    PIN din[65] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 688.230 0.000 688.370 0.140 ;
        END 
    END din[65] 
    PIN din[66] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 694.330 0.000 694.470 0.140 ;
        END 
    END din[66] 
    PIN din[67] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 700.430 0.000 700.570 0.140 ;
        END 
    END din[67] 
    PIN din[68] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 706.530 0.000 706.670 0.140 ;
        END 
    END din[68] 
    PIN din[69] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 712.630 0.000 712.770 0.140 ;
        END 
    END din[69] 
    PIN din[70] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 718.730 0.000 718.870 0.140 ;
        END 
    END din[70] 
    PIN din[71] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 724.830 0.000 724.970 0.140 ;
        END 
    END din[71] 
    PIN din[72] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 730.930 0.000 731.070 0.140 ;
        END 
    END din[72] 
    PIN din[73] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 737.030 0.000 737.170 0.140 ;
        END 
    END din[73] 
    PIN din[74] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 743.130 0.000 743.270 0.140 ;
        END 
    END din[74] 
    PIN din[75] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 749.230 0.000 749.370 0.140 ;
        END 
    END din[75] 
    PIN din[76] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 755.330 0.000 755.470 0.140 ;
        END 
    END din[76] 
    PIN din[77] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 761.430 0.000 761.570 0.140 ;
        END 
    END din[77] 
    PIN din[78] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 767.530 0.000 767.670 0.140 ;
        END 
    END din[78] 
    PIN din[79] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 773.630 0.000 773.770 0.140 ;
        END 
    END din[79] 
    PIN din[80] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 779.730 0.000 779.870 0.140 ;
        END 
    END din[80] 
    PIN din[81] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 785.830 0.000 785.970 0.140 ;
        END 
    END din[81] 
    PIN din[82] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 791.930 0.000 792.070 0.140 ;
        END 
    END din[82] 
    PIN din[83] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 798.030 0.000 798.170 0.140 ;
        END 
    END din[83] 
    PIN din[84] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 804.130 0.000 804.270 0.140 ;
        END 
    END din[84] 
    PIN din[85] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 810.230 0.000 810.370 0.140 ;
        END 
    END din[85] 
    PIN din[86] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 816.330 0.000 816.470 0.140 ;
        END 
    END din[86] 
    PIN din[87] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 822.430 0.000 822.570 0.140 ;
        END 
    END din[87] 
    PIN din[88] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 828.530 0.000 828.670 0.140 ;
        END 
    END din[88] 
    PIN din[89] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 834.630 0.000 834.770 0.140 ;
        END 
    END din[89] 
    PIN din[90] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 840.730 0.000 840.870 0.140 ;
        END 
    END din[90] 
    PIN din[91] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 846.830 0.000 846.970 0.140 ;
        END 
    END din[91] 
    PIN din[92] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 852.930 0.000 853.070 0.140 ;
        END 
    END din[92] 
    PIN din[93] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 859.030 0.000 859.170 0.140 ;
        END 
    END din[93] 
    PIN din[94] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 865.130 0.000 865.270 0.140 ;
        END 
    END din[94] 
    PIN din[95] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 871.230 0.000 871.370 0.140 ;
        END 
    END din[95] 
    PIN din[96] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 877.330 0.000 877.470 0.140 ;
        END 
    END din[96] 
    PIN din[97] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 883.430 0.000 883.570 0.140 ;
        END 
    END din[97] 
    PIN din[98] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 889.530 0.000 889.670 0.140 ;
        END 
    END din[98] 
    PIN din[99] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 895.630 0.000 895.770 0.140 ;
        END 
    END din[99] 
    PIN din[100] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 901.730 0.000 901.870 0.140 ;
        END 
    END din[100] 
    PIN din[101] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 907.830 0.000 907.970 0.140 ;
        END 
    END din[101] 
    PIN din[102] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 913.930 0.000 914.070 0.140 ;
        END 
    END din[102] 
    PIN din[103] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 920.030 0.000 920.170 0.140 ;
        END 
    END din[103] 
    PIN din[104] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 926.130 0.000 926.270 0.140 ;
        END 
    END din[104] 
    PIN din[105] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 932.230 0.000 932.370 0.140 ;
        END 
    END din[105] 
    PIN din[106] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 938.330 0.000 938.470 0.140 ;
        END 
    END din[106] 
    PIN din[107] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 944.430 0.000 944.570 0.140 ;
        END 
    END din[107] 
    PIN din[108] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 950.530 0.000 950.670 0.140 ;
        END 
    END din[108] 
    PIN din[109] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 956.630 0.000 956.770 0.140 ;
        END 
    END din[109] 
    PIN din[110] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 962.730 0.000 962.870 0.140 ;
        END 
    END din[110] 
    PIN din[111] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 968.830 0.000 968.970 0.140 ;
        END 
    END din[111] 
    PIN din[112] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 974.930 0.000 975.070 0.140 ;
        END 
    END din[112] 
    PIN din[113] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 981.030 0.000 981.170 0.140 ;
        END 
    END din[113] 
    PIN din[114] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 987.130 0.000 987.270 0.140 ;
        END 
    END din[114] 
    PIN din[115] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 993.230 0.000 993.370 0.140 ;
        END 
    END din[115] 
    PIN din[116] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 999.330 0.000 999.470 0.140 ;
        END 
    END din[116] 
    PIN din[117] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1005.430 0.000 1005.570 0.140 ;
        END 
    END din[117] 
    PIN din[118] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1011.530 0.000 1011.670 0.140 ;
        END 
    END din[118] 
    PIN din[119] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1017.630 0.000 1017.770 0.140 ;
        END 
    END din[119] 
    PIN din[120] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1023.730 0.000 1023.870 0.140 ;
        END 
    END din[120] 
    PIN din[121] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1029.830 0.000 1029.970 0.140 ;
        END 
    END din[121] 
    PIN din[122] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1035.930 0.000 1036.070 0.140 ;
        END 
    END din[122] 
    PIN din[123] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1042.030 0.000 1042.170 0.140 ;
        END 
    END din[123] 
    PIN din[124] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1048.130 0.000 1048.270 0.140 ;
        END 
    END din[124] 
    PIN din[125] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1054.230 0.000 1054.370 0.140 ;
        END 
    END din[125] 
    PIN din[126] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1060.330 0.000 1060.470 0.140 ;
        END 
    END din[126] 
    PIN din[127] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.745300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.358000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1066.430 0.000 1066.570 0.140 ;
        END 
    END din[127] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 291.380 0.000 291.520 0.140 ;
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 340.180 0.000 340.320 0.140 ;
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 388.980 0.000 389.120 0.140 ;
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 437.780 0.000 437.920 0.140 ;
        END 
    END wmask[3] 
    PIN wmask[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 486.580 0.000 486.720 0.140 ;
        END 
    END wmask[4] 
    PIN wmask[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 535.380 0.000 535.520 0.140 ;
        END 
    END wmask[5] 
    PIN wmask[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 584.180 0.000 584.320 0.140 ;
        END 
    END wmask[6] 
    PIN wmask[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 632.980 0.000 633.120 0.140 ;
        END 
    END wmask[7] 
    PIN wmask[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 681.780 0.000 681.920 0.140 ;
        END 
    END wmask[8] 
    PIN wmask[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 730.580 0.000 730.720 0.140 ;
        END 
    END wmask[9] 
    PIN wmask[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 779.380 0.000 779.520 0.140 ;
        END 
    END wmask[10] 
    PIN wmask[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 828.180 0.000 828.320 0.140 ;
        END 
    END wmask[11] 
    PIN wmask[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 876.980 0.000 877.120 0.140 ;
        END 
    END wmask[12] 
    PIN wmask[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 925.780 0.000 925.920 0.140 ;
        END 
    END wmask[13] 
    PIN wmask[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 974.580 0.000 974.720 0.140 ;
        END 
    END wmask[14] 
    PIN wmask[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.555700 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 1023.380 0.000 1023.520 0.140 ;
        END 
    END wmask[15] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.739900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 242.560 0.000 242.880 0.320 ;
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.739900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 236.440 0.000 236.760 0.320 ;
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.739900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 230.320 0.000 230.640 0.320 ;
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.739900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 224.200 0.000 224.520 0.320 ;
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.739900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 218.080 0.000 218.400 0.320 ;
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.739900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 211.960 0.000 212.280 0.320 ;
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.739900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 205.840 0.000 206.160 0.320 ;
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.739900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 199.720 0.000 200.040 0.320 ;
        END 
    END addr[7] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.739900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 254.120 0.000 254.440 0.320 ;
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.739900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 248.680 0.000 249.000 0.320 ;
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 79.236000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 257.520 0.000 257.840 0.320 ;
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 83.142000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 258.200 0.000 258.520 0.320 ;
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 291.160 6.240 ;
                RECT 292.880 5.920 297.280 6.240 ;
                RECT 299.000 5.920 303.400 6.240 ;
                RECT 305.120 5.920 309.520 6.240 ;
                RECT 311.240 5.920 315.640 6.240 ;
                RECT 317.360 5.920 321.760 6.240 ;
                RECT 323.480 5.920 327.880 6.240 ;
                RECT 329.600 5.920 334.000 6.240 ;
                RECT 335.720 5.920 340.120 6.240 ;
                RECT 341.840 5.920 346.240 6.240 ;
                RECT 347.960 5.920 352.360 6.240 ;
                RECT 354.080 5.920 358.480 6.240 ;
                RECT 360.200 5.920 364.600 6.240 ;
                RECT 366.320 5.920 370.720 6.240 ;
                RECT 372.440 5.920 376.840 6.240 ;
                RECT 378.560 5.920 382.960 6.240 ;
                RECT 384.680 5.920 389.080 6.240 ;
                RECT 390.800 5.920 395.200 6.240 ;
                RECT 396.920 5.920 401.320 6.240 ;
                RECT 403.040 5.920 407.440 6.240 ;
                RECT 409.160 5.920 413.560 6.240 ;
                RECT 415.280 5.920 419.680 6.240 ;
                RECT 421.400 5.920 425.800 6.240 ;
                RECT 427.520 5.920 431.920 6.240 ;
                RECT 432.960 5.920 438.040 6.240 ;
                RECT 439.080 5.920 444.160 6.240 ;
                RECT 445.200 5.920 450.280 6.240 ;
                RECT 451.320 5.920 456.400 6.240 ;
                RECT 457.440 5.920 462.520 6.240 ;
                RECT 463.560 5.920 468.640 6.240 ;
                RECT 469.680 5.920 474.760 6.240 ;
                RECT 475.800 5.920 480.880 6.240 ;
                RECT 481.920 5.920 486.320 6.240 ;
                RECT 488.040 5.920 492.440 6.240 ;
                RECT 494.160 5.920 498.560 6.240 ;
                RECT 500.280 5.920 504.680 6.240 ;
                RECT 506.400 5.920 510.800 6.240 ;
                RECT 512.520 5.920 516.920 6.240 ;
                RECT 518.640 5.920 523.040 6.240 ;
                RECT 524.760 5.920 529.160 6.240 ;
                RECT 530.880 5.920 535.280 6.240 ;
                RECT 537.000 5.920 541.400 6.240 ;
                RECT 543.120 5.920 547.520 6.240 ;
                RECT 549.240 5.920 553.640 6.240 ;
                RECT 555.360 5.920 559.760 6.240 ;
                RECT 561.480 5.920 565.880 6.240 ;
                RECT 567.600 5.920 572.000 6.240 ;
                RECT 573.720 5.920 578.120 6.240 ;
                RECT 579.840 5.920 584.240 6.240 ;
                RECT 585.960 5.920 590.360 6.240 ;
                RECT 592.080 5.920 596.480 6.240 ;
                RECT 598.200 5.920 602.600 6.240 ;
                RECT 604.320 5.920 608.720 6.240 ;
                RECT 610.440 5.920 614.840 6.240 ;
                RECT 616.560 5.920 620.960 6.240 ;
                RECT 622.680 5.920 627.080 6.240 ;
                RECT 628.800 5.920 633.200 6.240 ;
                RECT 634.920 5.920 639.320 6.240 ;
                RECT 640.360 5.920 645.440 6.240 ;
                RECT 646.480 5.920 651.560 6.240 ;
                RECT 652.600 5.920 657.680 6.240 ;
                RECT 658.720 5.920 663.800 6.240 ;
                RECT 664.840 5.920 669.920 6.240 ;
                RECT 670.960 5.920 676.040 6.240 ;
                RECT 677.080 5.920 682.160 6.240 ;
                RECT 683.200 5.920 688.280 6.240 ;
                RECT 689.320 5.920 693.720 6.240 ;
                RECT 695.440 5.920 699.840 6.240 ;
                RECT 701.560 5.920 705.960 6.240 ;
                RECT 707.680 5.920 712.080 6.240 ;
                RECT 713.800 5.920 718.200 6.240 ;
                RECT 719.920 5.920 724.320 6.240 ;
                RECT 726.040 5.920 730.440 6.240 ;
                RECT 732.160 5.920 736.560 6.240 ;
                RECT 738.280 5.920 742.680 6.240 ;
                RECT 744.400 5.920 748.800 6.240 ;
                RECT 750.520 5.920 754.920 6.240 ;
                RECT 756.640 5.920 761.040 6.240 ;
                RECT 762.760 5.920 767.160 6.240 ;
                RECT 768.880 5.920 773.280 6.240 ;
                RECT 775.000 5.920 779.400 6.240 ;
                RECT 781.120 5.920 785.520 6.240 ;
                RECT 787.240 5.920 791.640 6.240 ;
                RECT 793.360 5.920 797.760 6.240 ;
                RECT 799.480 5.920 803.880 6.240 ;
                RECT 805.600 5.920 810.000 6.240 ;
                RECT 811.720 5.920 816.120 6.240 ;
                RECT 817.840 5.920 822.240 6.240 ;
                RECT 823.960 5.920 828.360 6.240 ;
                RECT 830.080 5.920 834.480 6.240 ;
                RECT 836.200 5.920 840.600 6.240 ;
                RECT 842.320 5.920 846.720 6.240 ;
                RECT 847.760 5.920 852.840 6.240 ;
                RECT 853.880 5.920 858.960 6.240 ;
                RECT 860.000 5.920 865.080 6.240 ;
                RECT 866.120 5.920 871.200 6.240 ;
                RECT 872.240 5.920 877.320 6.240 ;
                RECT 878.360 5.920 883.440 6.240 ;
                RECT 884.480 5.920 889.560 6.240 ;
                RECT 890.600 5.920 895.680 6.240 ;
                RECT 896.720 5.920 901.120 6.240 ;
                RECT 902.840 5.920 907.240 6.240 ;
                RECT 908.960 5.920 913.360 6.240 ;
                RECT 915.080 5.920 919.480 6.240 ;
                RECT 921.200 5.920 925.600 6.240 ;
                RECT 927.320 5.920 931.720 6.240 ;
                RECT 933.440 5.920 937.840 6.240 ;
                RECT 939.560 5.920 943.960 6.240 ;
                RECT 945.680 5.920 950.080 6.240 ;
                RECT 951.800 5.920 956.200 6.240 ;
                RECT 957.920 5.920 962.320 6.240 ;
                RECT 964.040 5.920 968.440 6.240 ;
                RECT 970.160 5.920 974.560 6.240 ;
                RECT 976.280 5.920 980.680 6.240 ;
                RECT 982.400 5.920 986.800 6.240 ;
                RECT 988.520 5.920 992.920 6.240 ;
                RECT 994.640 5.920 999.040 6.240 ;
                RECT 1000.760 5.920 1005.160 6.240 ;
                RECT 1006.880 5.920 1011.280 6.240 ;
                RECT 1013.000 5.920 1017.400 6.240 ;
                RECT 1019.120 5.920 1023.520 6.240 ;
                RECT 1025.240 5.920 1029.640 6.240 ;
                RECT 1031.360 5.920 1035.760 6.240 ;
                RECT 1037.480 5.920 1041.880 6.240 ;
                RECT 1043.600 5.920 1048.000 6.240 ;
                RECT 1049.720 5.920 1054.120 6.240 ;
                RECT 1055.160 5.920 1060.240 6.240 ;
                RECT 1061.280 5.920 1066.360 6.240 ;
                RECT 1067.400 5.920 1085.720 6.240 ;
                RECT 0.160 7.280 1085.720 7.600 ;
                RECT 0.160 8.640 1085.720 8.960 ;
                RECT 0.160 10.000 257.160 10.320 ;
                RECT 287.440 10.000 1085.720 10.320 ;
                RECT 0.160 11.360 1085.720 11.680 ;
                RECT 0.160 12.720 195.280 13.040 ;
                RECT 258.880 12.720 1085.720 13.040 ;
                RECT 0.160 14.080 1085.720 14.400 ;
                RECT 0.160 15.440 1085.720 15.760 ;
                RECT 0.160 16.800 195.280 17.120 ;
                RECT 258.200 16.800 1085.720 17.120 ;
                RECT 0.160 18.160 1085.720 18.480 ;
                RECT 0.160 19.520 1085.720 19.840 ;
                RECT 0.160 20.880 1085.720 21.200 ;
                RECT 0.160 22.240 1085.720 22.560 ;
                RECT 0.160 23.600 290.480 23.920 ;
                RECT 1023.880 23.600 1085.720 23.920 ;
                RECT 0.160 24.960 280.960 25.280 ;
                RECT 1076.240 24.960 1085.720 25.280 ;
                RECT 0.160 26.320 280.960 26.640 ;
                RECT 1076.240 26.320 1085.720 26.640 ;
                RECT 0.160 27.680 280.960 28.000 ;
                RECT 1076.240 27.680 1085.720 28.000 ;
                RECT 0.160 29.040 280.960 29.360 ;
                RECT 1076.240 29.040 1085.720 29.360 ;
                RECT 0.160 30.400 280.960 30.720 ;
                RECT 1076.240 30.400 1085.720 30.720 ;
                RECT 0.160 31.760 280.960 32.080 ;
                RECT 1076.240 31.760 1085.720 32.080 ;
                RECT 0.160 33.120 144.960 33.440 ;
                RECT 237.120 33.120 280.960 33.440 ;
                RECT 1076.240 33.120 1085.720 33.440 ;
                RECT 0.160 34.480 143.600 34.800 ;
                RECT 243.240 34.480 280.960 34.800 ;
                RECT 1076.240 34.480 1085.720 34.800 ;
                RECT 0.160 35.840 120.480 36.160 ;
                RECT 258.200 35.840 280.960 36.160 ;
                RECT 1076.240 35.840 1085.720 36.160 ;
                RECT 0.160 37.200 121.160 37.520 ;
                RECT 248.680 37.200 280.960 37.520 ;
                RECT 1076.240 37.200 1085.720 37.520 ;
                RECT 0.160 38.560 280.960 38.880 ;
                RECT 1076.240 38.560 1085.720 38.880 ;
                RECT 0.160 39.920 280.960 40.240 ;
                RECT 1076.240 39.920 1085.720 40.240 ;
                RECT 0.160 41.280 280.280 41.600 ;
                RECT 1076.240 41.280 1085.720 41.600 ;
                RECT 0.160 42.640 280.960 42.960 ;
                RECT 1076.240 42.640 1085.720 42.960 ;
                RECT 0.160 44.000 280.960 44.320 ;
                RECT 1076.240 44.000 1085.720 44.320 ;
                RECT 0.160 45.360 118.440 45.680 ;
                RECT 129.680 45.360 280.960 45.680 ;
                RECT 1076.240 45.360 1085.720 45.680 ;
                RECT 0.160 46.720 119.800 47.040 ;
                RECT 125.600 46.720 133.400 47.040 ;
                RECT 135.800 46.720 280.960 47.040 ;
                RECT 1076.240 46.720 1085.720 47.040 ;
                RECT 0.160 48.080 121.160 48.400 ;
                RECT 124.920 48.080 280.960 48.400 ;
                RECT 1076.240 48.080 1085.720 48.400 ;
                RECT 0.160 49.440 127.960 49.760 ;
                RECT 135.120 49.440 225.200 49.760 ;
                RECT 254.800 49.440 280.960 49.760 ;
                RECT 1076.240 49.440 1085.720 49.760 ;
                RECT 0.160 50.800 123.200 51.120 ;
                RECT 136.480 50.800 225.200 51.120 ;
                RECT 1076.240 50.800 1085.720 51.120 ;
                RECT 0.160 52.160 120.480 52.480 ;
                RECT 129.680 52.160 225.200 52.480 ;
                RECT 1076.240 52.160 1085.720 52.480 ;
                RECT 0.160 53.520 225.200 53.840 ;
                RECT 254.800 53.520 280.960 53.840 ;
                RECT 1076.240 53.520 1085.720 53.840 ;
                RECT 0.160 54.880 119.800 55.200 ;
                RECT 122.880 54.880 225.200 55.200 ;
                RECT 254.800 54.880 280.960 55.200 ;
                RECT 1076.240 54.880 1085.720 55.200 ;
                RECT 0.160 56.240 120.480 56.560 ;
                RECT 135.120 56.240 280.960 56.560 ;
                RECT 1076.240 56.240 1085.720 56.560 ;
                RECT 0.160 57.600 126.600 57.920 ;
                RECT 129.680 57.600 280.960 57.920 ;
                RECT 1076.240 57.600 1085.720 57.920 ;
                RECT 0.160 58.960 280.960 59.280 ;
                RECT 1076.240 58.960 1085.720 59.280 ;
                RECT 0.160 60.320 127.960 60.640 ;
                RECT 135.800 60.320 153.800 60.640 ;
                RECT 256.160 60.320 280.960 60.640 ;
                RECT 1076.240 60.320 1085.720 60.640 ;
                RECT 0.160 61.680 124.560 62.000 ;
                RECT 129.680 61.680 143.600 62.000 ;
                RECT 148.040 61.680 153.800 62.000 ;
                RECT 256.160 61.680 280.960 62.000 ;
                RECT 1076.240 61.680 1085.720 62.000 ;
                RECT 0.160 63.040 126.600 63.360 ;
                RECT 129.680 63.040 144.960 63.360 ;
                RECT 147.360 63.040 153.800 63.360 ;
                RECT 269.080 63.040 280.960 63.360 ;
                RECT 1076.240 63.040 1085.720 63.360 ;
                RECT 0.160 64.400 153.800 64.720 ;
                RECT 269.080 64.400 280.960 64.720 ;
                RECT 1076.240 64.400 1085.720 64.720 ;
                RECT 0.160 65.760 117.760 66.080 ;
                RECT 141.240 65.760 153.800 66.080 ;
                RECT 269.080 65.760 280.960 66.080 ;
                RECT 1076.240 65.760 1085.720 66.080 ;
                RECT 0.160 67.120 136.800 67.440 ;
                RECT 142.600 67.120 153.800 67.440 ;
                RECT 267.040 67.120 280.960 67.440 ;
                RECT 1076.240 67.120 1085.720 67.440 ;
                RECT 0.160 68.480 126.600 68.800 ;
                RECT 129.680 68.480 139.520 68.800 ;
                RECT 143.280 68.480 153.800 68.800 ;
                RECT 269.080 68.480 280.960 68.800 ;
                RECT 1076.240 68.480 1085.720 68.800 ;
                RECT 0.160 69.840 118.440 70.160 ;
                RECT 132.400 69.840 153.800 70.160 ;
                RECT 256.160 69.840 280.960 70.160 ;
                RECT 1076.240 69.840 1085.720 70.160 ;
                RECT 0.160 71.200 127.280 71.520 ;
                RECT 135.800 71.200 153.800 71.520 ;
                RECT 269.080 71.200 280.960 71.520 ;
                RECT 1076.240 71.200 1085.720 71.520 ;
                RECT 0.160 72.560 125.240 72.880 ;
                RECT 129.000 72.560 153.800 72.880 ;
                RECT 273.160 72.560 280.960 72.880 ;
                RECT 1076.240 72.560 1085.720 72.880 ;
                RECT 0.160 73.920 127.960 74.240 ;
                RECT 136.480 73.920 153.800 74.240 ;
                RECT 271.120 73.920 280.960 74.240 ;
                RECT 1076.240 73.920 1085.720 74.240 ;
                RECT 0.160 75.280 153.800 75.600 ;
                RECT 273.160 75.280 280.960 75.600 ;
                RECT 1076.240 75.280 1085.720 75.600 ;
                RECT 0.160 76.640 119.800 76.960 ;
                RECT 124.920 76.640 153.800 76.960 ;
                RECT 273.160 76.640 280.960 76.960 ;
                RECT 1076.240 76.640 1085.720 76.960 ;
                RECT 0.160 78.000 123.200 78.320 ;
                RECT 129.680 78.000 153.800 78.320 ;
                RECT 256.160 78.000 280.960 78.320 ;
                RECT 1076.240 78.000 1085.720 78.320 ;
                RECT 0.160 79.360 153.800 79.680 ;
                RECT 273.160 79.360 280.960 79.680 ;
                RECT 1076.240 79.360 1085.720 79.680 ;
                RECT 0.160 80.720 126.600 81.040 ;
                RECT 129.000 80.720 153.800 81.040 ;
                RECT 271.120 80.720 280.960 81.040 ;
                RECT 1076.240 80.720 1085.720 81.040 ;
                RECT 0.160 82.080 127.960 82.400 ;
                RECT 129.680 82.080 153.800 82.400 ;
                RECT 273.160 82.080 280.960 82.400 ;
                RECT 1076.240 82.080 1085.720 82.400 ;
                RECT 0.160 83.440 153.800 83.760 ;
                RECT 277.240 83.440 280.960 83.760 ;
                RECT 1076.240 83.440 1085.720 83.760 ;
                RECT 0.160 84.800 125.240 85.120 ;
                RECT 135.800 84.800 153.800 85.120 ;
                RECT 277.240 84.800 280.960 85.120 ;
                RECT 1076.240 84.800 1085.720 85.120 ;
                RECT 0.160 86.160 117.760 86.480 ;
                RECT 135.800 86.160 153.800 86.480 ;
                RECT 275.200 86.160 280.960 86.480 ;
                RECT 1076.240 86.160 1085.720 86.480 ;
                RECT 0.160 87.520 127.280 87.840 ;
                RECT 129.680 87.520 153.800 87.840 ;
                RECT 256.160 87.520 280.960 87.840 ;
                RECT 1076.240 87.520 1085.720 87.840 ;
                RECT 0.160 88.880 153.800 89.200 ;
                RECT 277.240 88.880 280.960 89.200 ;
                RECT 1076.240 88.880 1085.720 89.200 ;
                RECT 0.160 90.240 153.800 90.560 ;
                RECT 277.240 90.240 280.960 90.560 ;
                RECT 1076.240 90.240 1085.720 90.560 ;
                RECT 0.160 91.600 115.040 91.920 ;
                RECT 128.320 91.600 153.800 91.920 ;
                RECT 277.240 91.600 280.960 91.920 ;
                RECT 1076.240 91.600 1085.720 91.920 ;
                RECT 0.160 92.960 124.560 93.280 ;
                RECT 132.400 92.960 153.800 93.280 ;
                RECT 275.200 92.960 280.960 93.280 ;
                RECT 1076.240 92.960 1085.720 93.280 ;
                RECT 0.160 94.320 153.800 94.640 ;
                RECT 1076.240 94.320 1085.720 94.640 ;
                RECT 0.160 95.680 121.840 96.000 ;
                RECT 124.920 95.680 153.800 96.000 ;
                RECT 256.160 95.680 280.960 96.000 ;
                RECT 1076.240 95.680 1085.720 96.000 ;
                RECT 0.160 97.040 120.480 97.360 ;
                RECT 138.520 97.040 153.800 97.360 ;
                RECT 1076.240 97.040 1085.720 97.360 ;
                RECT 0.160 98.400 153.800 98.720 ;
                RECT 1076.240 98.400 1085.720 98.720 ;
                RECT 0.160 99.760 153.800 100.080 ;
                RECT 1076.240 99.760 1085.720 100.080 ;
                RECT 0.160 101.120 121.840 101.440 ;
                RECT 135.120 101.120 153.800 101.440 ;
                RECT 1076.240 101.120 1085.720 101.440 ;
                RECT 0.160 102.480 117.760 102.800 ;
                RECT 122.200 102.480 153.800 102.800 ;
                RECT 1076.240 102.480 1085.720 102.800 ;
                RECT 0.160 103.840 153.800 104.160 ;
                RECT 256.160 103.840 280.960 104.160 ;
                RECT 1076.240 103.840 1085.720 104.160 ;
                RECT 0.160 105.200 280.960 105.520 ;
                RECT 1076.240 105.200 1085.720 105.520 ;
                RECT 0.160 106.560 118.440 106.880 ;
                RECT 125.600 106.560 133.400 106.880 ;
                RECT 136.480 106.560 280.960 106.880 ;
                RECT 1076.240 106.560 1085.720 106.880 ;
                RECT 0.160 107.920 280.960 108.240 ;
                RECT 1076.240 107.920 1085.720 108.240 ;
                RECT 0.160 109.280 123.880 109.600 ;
                RECT 128.320 109.280 280.960 109.600 ;
                RECT 1076.240 109.280 1085.720 109.600 ;
                RECT 0.160 110.640 142.240 110.960 ;
                RECT 186.120 110.640 189.160 110.960 ;
                RECT 254.800 110.640 280.960 110.960 ;
                RECT 1076.240 110.640 1085.720 110.960 ;
                RECT 0.160 112.000 120.480 112.320 ;
                RECT 125.600 112.000 189.160 112.320 ;
                RECT 254.800 112.000 280.960 112.320 ;
                RECT 1076.240 112.000 1085.720 112.320 ;
                RECT 0.160 113.360 189.160 113.680 ;
                RECT 254.800 113.360 280.960 113.680 ;
                RECT 1076.240 113.360 1085.720 113.680 ;
                RECT 0.160 114.720 126.600 115.040 ;
                RECT 135.120 114.720 189.160 115.040 ;
                RECT 254.800 114.720 280.960 115.040 ;
                RECT 1076.240 114.720 1085.720 115.040 ;
                RECT 0.160 116.080 189.160 116.400 ;
                RECT 254.800 116.080 280.960 116.400 ;
                RECT 1076.240 116.080 1085.720 116.400 ;
                RECT 0.160 117.440 189.160 117.760 ;
                RECT 1076.240 117.440 1085.720 117.760 ;
                RECT 0.160 118.800 121.160 119.120 ;
                RECT 123.560 118.800 189.160 119.120 ;
                RECT 254.800 118.800 276.880 119.120 ;
                RECT 1076.240 118.800 1085.720 119.120 ;
                RECT 0.160 120.160 96.680 120.480 ;
                RECT 115.400 120.160 189.160 120.480 ;
                RECT 254.800 120.160 276.880 120.480 ;
                RECT 1076.240 120.160 1085.720 120.480 ;
                RECT 0.160 121.520 96.680 121.840 ;
                RECT 115.400 121.520 189.160 121.840 ;
                RECT 254.800 121.520 272.800 121.840 ;
                RECT 1076.240 121.520 1085.720 121.840 ;
                RECT 0.160 122.880 96.680 123.200 ;
                RECT 115.400 122.880 189.160 123.200 ;
                RECT 254.800 122.880 268.720 123.200 ;
                RECT 1076.240 122.880 1085.720 123.200 ;
                RECT 0.160 124.240 96.680 124.560 ;
                RECT 115.400 124.240 189.160 124.560 ;
                RECT 254.800 124.240 268.720 124.560 ;
                RECT 1076.240 124.240 1085.720 124.560 ;
                RECT 0.160 125.600 96.680 125.920 ;
                RECT 115.400 125.600 189.160 125.920 ;
                RECT 254.800 125.600 264.640 125.920 ;
                RECT 1076.240 125.600 1085.720 125.920 ;
                RECT 0.160 126.960 96.680 127.280 ;
                RECT 115.400 126.960 189.160 127.280 ;
                RECT 254.800 126.960 264.640 127.280 ;
                RECT 1076.240 126.960 1085.720 127.280 ;
                RECT 0.160 128.320 96.680 128.640 ;
                RECT 115.400 128.320 189.160 128.640 ;
                RECT 254.800 128.320 280.960 128.640 ;
                RECT 1076.240 128.320 1085.720 128.640 ;
                RECT 0.160 129.680 96.680 130.000 ;
                RECT 115.400 129.680 280.960 130.000 ;
                RECT 1076.240 129.680 1085.720 130.000 ;
                RECT 0.160 131.040 96.680 131.360 ;
                RECT 115.400 131.040 280.960 131.360 ;
                RECT 1076.240 131.040 1085.720 131.360 ;
                RECT 0.160 132.400 96.680 132.720 ;
                RECT 115.400 132.400 280.960 132.720 ;
                RECT 1076.240 132.400 1085.720 132.720 ;
                RECT 0.160 133.760 96.680 134.080 ;
                RECT 115.400 133.760 280.960 134.080 ;
                RECT 1076.240 133.760 1085.720 134.080 ;
                RECT 0.160 135.120 96.680 135.440 ;
                RECT 116.080 135.120 187.800 135.440 ;
                RECT 256.160 135.120 280.960 135.440 ;
                RECT 1076.240 135.120 1085.720 135.440 ;
                RECT 0.160 136.480 96.680 136.800 ;
                RECT 115.400 136.480 187.800 136.800 ;
                RECT 256.160 136.480 280.960 136.800 ;
                RECT 1076.240 136.480 1085.720 136.800 ;
                RECT 0.160 137.840 96.680 138.160 ;
                RECT 115.400 137.840 187.800 138.160 ;
                RECT 256.160 137.840 280.960 138.160 ;
                RECT 1076.240 137.840 1085.720 138.160 ;
                RECT 0.160 139.200 96.680 139.520 ;
                RECT 115.400 139.200 187.800 139.520 ;
                RECT 256.160 139.200 280.960 139.520 ;
                RECT 1076.240 139.200 1085.720 139.520 ;
                RECT 0.160 140.560 96.680 140.880 ;
                RECT 115.400 140.560 187.800 140.880 ;
                RECT 256.160 140.560 280.960 140.880 ;
                RECT 1076.240 140.560 1085.720 140.880 ;
                RECT 0.160 141.920 96.680 142.240 ;
                RECT 115.400 141.920 123.200 142.240 ;
                RECT 125.600 141.920 187.800 142.240 ;
                RECT 256.160 141.920 266.680 142.240 ;
                RECT 1076.240 141.920 1085.720 142.240 ;
                RECT 0.160 143.280 96.680 143.600 ;
                RECT 115.400 143.280 187.800 143.600 ;
                RECT 256.160 143.280 266.680 143.600 ;
                RECT 1076.240 143.280 1085.720 143.600 ;
                RECT 0.160 144.640 96.680 144.960 ;
                RECT 115.400 144.640 187.800 144.960 ;
                RECT 256.160 144.640 270.760 144.960 ;
                RECT 1076.240 144.640 1085.720 144.960 ;
                RECT 0.160 146.000 96.680 146.320 ;
                RECT 115.400 146.000 187.800 146.320 ;
                RECT 256.160 146.000 274.840 146.320 ;
                RECT 1076.240 146.000 1085.720 146.320 ;
                RECT 0.160 147.360 96.680 147.680 ;
                RECT 115.400 147.360 187.800 147.680 ;
                RECT 256.160 147.360 274.840 147.680 ;
                RECT 1076.240 147.360 1085.720 147.680 ;
                RECT 0.160 148.720 96.680 149.040 ;
                RECT 115.400 148.720 187.800 149.040 ;
                RECT 256.160 148.720 278.920 149.040 ;
                RECT 1076.240 148.720 1085.720 149.040 ;
                RECT 0.160 150.080 96.680 150.400 ;
                RECT 115.400 150.080 187.800 150.400 ;
                RECT 1076.240 150.080 1085.720 150.400 ;
                RECT 0.160 151.440 96.680 151.760 ;
                RECT 115.400 151.440 187.800 151.760 ;
                RECT 1076.240 151.440 1085.720 151.760 ;
                RECT 0.160 152.800 96.680 153.120 ;
                RECT 115.400 152.800 119.800 153.120 ;
                RECT 125.600 152.800 187.800 153.120 ;
                RECT 256.160 152.800 280.960 153.120 ;
                RECT 1076.240 152.800 1085.720 153.120 ;
                RECT 0.160 154.160 187.800 154.480 ;
                RECT 256.160 154.160 280.960 154.480 ;
                RECT 1076.240 154.160 1085.720 154.480 ;
                RECT 0.160 155.520 187.800 155.840 ;
                RECT 256.160 155.520 280.960 155.840 ;
                RECT 1076.240 155.520 1085.720 155.840 ;
                RECT 0.160 156.880 123.880 157.200 ;
                RECT 129.680 156.880 187.800 157.200 ;
                RECT 256.160 156.880 280.960 157.200 ;
                RECT 1076.240 156.880 1085.720 157.200 ;
                RECT 0.160 158.240 78.320 158.560 ;
                RECT 97.040 158.240 102.800 158.560 ;
                RECT 109.960 158.240 187.800 158.560 ;
                RECT 256.160 158.240 280.960 158.560 ;
                RECT 1076.240 158.240 1085.720 158.560 ;
                RECT 0.160 159.600 78.320 159.920 ;
                RECT 114.720 159.600 187.800 159.920 ;
                RECT 256.160 159.600 280.960 159.920 ;
                RECT 1076.240 159.600 1085.720 159.920 ;
                RECT 0.160 160.960 78.320 161.280 ;
                RECT 114.720 160.960 187.800 161.280 ;
                RECT 1076.240 160.960 1085.720 161.280 ;
                RECT 0.160 162.320 78.320 162.640 ;
                RECT 97.040 162.320 102.800 162.640 ;
                RECT 109.960 162.320 117.760 162.640 ;
                RECT 128.320 162.320 187.800 162.640 ;
                RECT 256.160 162.320 261.240 162.640 ;
                RECT 1076.240 162.320 1085.720 162.640 ;
                RECT 0.160 163.680 75.600 164.000 ;
                RECT 109.280 163.680 187.800 164.000 ;
                RECT 256.160 163.680 1085.720 164.000 ;
                RECT 0.160 165.040 108.920 165.360 ;
                RECT 185.440 165.040 1085.720 165.360 ;
                RECT 0.160 166.400 278.240 166.720 ;
                RECT 1078.960 166.400 1085.720 166.720 ;
                RECT 0.160 167.760 278.240 168.080 ;
                RECT 1078.960 167.760 1085.720 168.080 ;
                RECT 0.160 169.120 278.240 169.440 ;
                RECT 1078.960 169.120 1085.720 169.440 ;
                RECT 0.160 170.480 25.960 170.800 ;
                RECT 32.440 170.480 34.800 170.800 ;
                RECT 47.400 170.480 79.680 170.800 ;
                RECT 1078.960 170.480 1085.720 170.800 ;
                RECT 0.160 171.840 23.920 172.160 ;
                RECT 34.480 171.840 36.160 172.160 ;
                RECT 46.040 171.840 64.040 172.160 ;
                RECT 69.160 171.840 79.680 172.160 ;
                RECT 1078.960 171.840 1085.720 172.160 ;
                RECT 0.160 173.200 23.920 173.520 ;
                RECT 34.480 173.200 37.520 173.520 ;
                RECT 45.360 173.200 59.280 173.520 ;
                RECT 69.160 173.200 79.680 173.520 ;
                RECT 1078.960 173.200 1085.720 173.520 ;
                RECT 0.160 174.560 23.920 174.880 ;
                RECT 34.480 174.560 59.280 174.880 ;
                RECT 69.160 174.560 79.680 174.880 ;
                RECT 1078.960 174.560 1085.720 174.880 ;
                RECT 0.160 175.920 59.280 176.240 ;
                RECT 69.160 175.920 79.680 176.240 ;
                RECT 1078.960 175.920 1085.720 176.240 ;
                RECT 0.160 177.280 23.920 177.600 ;
                RECT 34.480 177.280 59.280 177.600 ;
                RECT 69.160 177.280 79.680 177.600 ;
                RECT 1078.960 177.280 1085.720 177.600 ;
                RECT 0.160 178.640 23.920 178.960 ;
                RECT 34.480 178.640 79.680 178.960 ;
                RECT 1078.960 178.640 1085.720 178.960 ;
                RECT 0.160 180.000 59.960 180.320 ;
                RECT 69.160 180.000 79.680 180.320 ;
                RECT 1078.960 180.000 1085.720 180.320 ;
                RECT 0.160 181.360 59.280 181.680 ;
                RECT 69.160 181.360 79.680 181.680 ;
                RECT 1078.960 181.360 1085.720 181.680 ;
                RECT 0.160 182.720 59.280 183.040 ;
                RECT 69.160 182.720 79.680 183.040 ;
                RECT 1078.960 182.720 1085.720 183.040 ;
                RECT 0.160 184.080 17.120 184.400 ;
                RECT 19.520 184.080 32.760 184.400 ;
                RECT 35.840 184.080 59.280 184.400 ;
                RECT 69.160 184.080 79.680 184.400 ;
                RECT 1078.960 184.080 1085.720 184.400 ;
                RECT 0.160 185.440 16.440 185.760 ;
                RECT 19.520 185.440 32.760 185.760 ;
                RECT 36.520 185.440 59.280 185.760 ;
                RECT 69.160 185.440 79.680 185.760 ;
                RECT 1078.960 185.440 1085.720 185.760 ;
                RECT 0.160 186.800 15.760 187.120 ;
                RECT 19.520 186.800 79.680 187.120 ;
                RECT 1078.960 186.800 1085.720 187.120 ;
                RECT 0.160 188.160 15.080 188.480 ;
                RECT 19.520 188.160 60.640 188.480 ;
                RECT 69.160 188.160 79.680 188.480 ;
                RECT 1078.960 188.160 1085.720 188.480 ;
                RECT 0.160 189.520 59.280 189.840 ;
                RECT 69.160 189.520 79.680 189.840 ;
                RECT 1078.960 189.520 1085.720 189.840 ;
                RECT 0.160 190.880 14.400 191.200 ;
                RECT 19.520 190.880 59.280 191.200 ;
                RECT 69.160 190.880 79.680 191.200 ;
                RECT 1078.960 190.880 1085.720 191.200 ;
                RECT 0.160 192.240 13.720 192.560 ;
                RECT 19.520 192.240 59.280 192.560 ;
                RECT 69.160 192.240 79.680 192.560 ;
                RECT 1078.960 192.240 1085.720 192.560 ;
                RECT 0.160 193.600 59.280 193.920 ;
                RECT 69.160 193.600 79.680 193.920 ;
                RECT 1078.960 193.600 1085.720 193.920 ;
                RECT 0.160 194.960 13.040 195.280 ;
                RECT 19.520 194.960 79.680 195.280 ;
                RECT 1078.960 194.960 1085.720 195.280 ;
                RECT 0.160 196.320 12.360 196.640 ;
                RECT 19.520 196.320 32.760 196.640 ;
                RECT 38.560 196.320 59.280 196.640 ;
                RECT 69.160 196.320 79.680 196.640 ;
                RECT 1078.960 196.320 1085.720 196.640 ;
                RECT 0.160 197.680 59.280 198.000 ;
                RECT 69.160 197.680 79.680 198.000 ;
                RECT 1078.960 197.680 1085.720 198.000 ;
                RECT 0.160 199.040 11.680 199.360 ;
                RECT 19.520 199.040 32.760 199.360 ;
                RECT 37.880 199.040 59.280 199.360 ;
                RECT 69.160 199.040 79.680 199.360 ;
                RECT 1078.960 199.040 1085.720 199.360 ;
                RECT 0.160 200.400 11.000 200.720 ;
                RECT 19.520 200.400 32.760 200.720 ;
                RECT 37.200 200.400 59.280 200.720 ;
                RECT 69.160 200.400 79.680 200.720 ;
                RECT 1078.960 200.400 1085.720 200.720 ;
                RECT 0.160 201.760 10.320 202.080 ;
                RECT 19.520 201.760 32.760 202.080 ;
                RECT 36.520 201.760 59.280 202.080 ;
                RECT 69.160 201.760 79.680 202.080 ;
                RECT 1078.960 201.760 1085.720 202.080 ;
                RECT 0.160 203.120 9.640 203.440 ;
                RECT 19.520 203.120 64.040 203.440 ;
                RECT 69.160 203.120 79.680 203.440 ;
                RECT 1078.960 203.120 1085.720 203.440 ;
                RECT 0.160 204.480 60.640 204.800 ;
                RECT 69.160 204.480 79.680 204.800 ;
                RECT 1078.960 204.480 1085.720 204.800 ;
                RECT 0.160 205.840 60.640 206.160 ;
                RECT 69.160 205.840 79.680 206.160 ;
                RECT 1078.960 205.840 1085.720 206.160 ;
                RECT 0.160 207.200 60.640 207.520 ;
                RECT 69.160 207.200 79.680 207.520 ;
                RECT 1078.960 207.200 1085.720 207.520 ;
                RECT 0.160 208.560 60.640 208.880 ;
                RECT 69.160 208.560 79.680 208.880 ;
                RECT 1078.960 208.560 1085.720 208.880 ;
                RECT 0.160 209.920 38.200 210.240 ;
                RECT 47.400 209.920 79.680 210.240 ;
                RECT 1078.960 209.920 1085.720 210.240 ;
                RECT 0.160 211.280 36.840 211.600 ;
                RECT 46.040 211.280 65.400 211.600 ;
                RECT 69.160 211.280 79.680 211.600 ;
                RECT 1078.960 211.280 1085.720 211.600 ;
                RECT 0.160 212.640 35.480 212.960 ;
                RECT 45.360 212.640 59.280 212.960 ;
                RECT 69.160 212.640 79.680 212.960 ;
                RECT 1078.960 212.640 1085.720 212.960 ;
                RECT 0.160 214.000 59.280 214.320 ;
                RECT 69.160 214.000 79.680 214.320 ;
                RECT 1078.960 214.000 1085.720 214.320 ;
                RECT 0.160 215.360 59.280 215.680 ;
                RECT 69.160 215.360 79.680 215.680 ;
                RECT 1078.960 215.360 1085.720 215.680 ;
                RECT 0.160 216.720 59.280 217.040 ;
                RECT 69.160 216.720 79.680 217.040 ;
                RECT 1078.960 216.720 1085.720 217.040 ;
                RECT 0.160 218.080 59.280 218.400 ;
                RECT 62.360 218.080 79.680 218.400 ;
                RECT 1078.960 218.080 1085.720 218.400 ;
                RECT 0.160 219.440 61.320 219.760 ;
                RECT 69.160 219.440 79.680 219.760 ;
                RECT 1078.960 219.440 1085.720 219.760 ;
                RECT 0.160 220.800 59.280 221.120 ;
                RECT 69.160 220.800 79.680 221.120 ;
                RECT 1078.960 220.800 1085.720 221.120 ;
                RECT 0.160 222.160 59.280 222.480 ;
                RECT 69.160 222.160 79.680 222.480 ;
                RECT 1078.960 222.160 1085.720 222.480 ;
                RECT 0.160 223.520 59.280 223.840 ;
                RECT 69.160 223.520 79.680 223.840 ;
                RECT 1078.960 223.520 1085.720 223.840 ;
                RECT 0.160 224.880 59.280 225.200 ;
                RECT 69.160 224.880 79.680 225.200 ;
                RECT 1078.960 224.880 1085.720 225.200 ;
                RECT 0.160 226.240 79.680 226.560 ;
                RECT 1078.960 226.240 1085.720 226.560 ;
                RECT 0.160 227.600 61.320 227.920 ;
                RECT 69.160 227.600 79.680 227.920 ;
                RECT 1078.960 227.600 1085.720 227.920 ;
                RECT 0.160 228.960 59.280 229.280 ;
                RECT 69.160 228.960 79.680 229.280 ;
                RECT 1078.960 228.960 1085.720 229.280 ;
                RECT 0.160 230.320 59.280 230.640 ;
                RECT 69.160 230.320 79.680 230.640 ;
                RECT 1078.960 230.320 1085.720 230.640 ;
                RECT 0.160 231.680 59.280 232.000 ;
                RECT 69.160 231.680 79.680 232.000 ;
                RECT 1078.960 231.680 1085.720 232.000 ;
                RECT 0.160 233.040 59.280 233.360 ;
                RECT 69.160 233.040 79.680 233.360 ;
                RECT 1078.960 233.040 1085.720 233.360 ;
                RECT 0.160 234.400 79.680 234.720 ;
                RECT 1078.960 234.400 1085.720 234.720 ;
                RECT 0.160 235.760 59.280 236.080 ;
                RECT 69.160 235.760 79.680 236.080 ;
                RECT 1078.960 235.760 1085.720 236.080 ;
                RECT 0.160 237.120 59.280 237.440 ;
                RECT 69.160 237.120 79.680 237.440 ;
                RECT 1078.960 237.120 1085.720 237.440 ;
                RECT 0.160 238.480 59.280 238.800 ;
                RECT 69.160 238.480 79.680 238.800 ;
                RECT 1078.960 238.480 1085.720 238.800 ;
                RECT 0.160 239.840 59.280 240.160 ;
                RECT 69.160 239.840 79.680 240.160 ;
                RECT 1078.960 239.840 1085.720 240.160 ;
                RECT 0.160 241.200 59.280 241.520 ;
                RECT 69.160 241.200 79.680 241.520 ;
                RECT 1078.960 241.200 1085.720 241.520 ;
                RECT 0.160 242.560 79.680 242.880 ;
                RECT 1078.960 242.560 1085.720 242.880 ;
                RECT 0.160 243.920 62.000 244.240 ;
                RECT 69.160 243.920 79.680 244.240 ;
                RECT 1078.960 243.920 1085.720 244.240 ;
                RECT 0.160 245.280 62.000 245.600 ;
                RECT 69.160 245.280 79.680 245.600 ;
                RECT 1078.960 245.280 1085.720 245.600 ;
                RECT 0.160 246.640 62.000 246.960 ;
                RECT 69.160 246.640 79.680 246.960 ;
                RECT 1078.960 246.640 1085.720 246.960 ;
                RECT 0.160 248.000 62.000 248.320 ;
                RECT 69.160 248.000 79.680 248.320 ;
                RECT 1078.960 248.000 1085.720 248.320 ;
                RECT 0.160 249.360 79.680 249.680 ;
                RECT 1078.960 249.360 1085.720 249.680 ;
                RECT 0.160 250.720 64.040 251.040 ;
                RECT 69.160 250.720 79.680 251.040 ;
                RECT 1078.960 250.720 1085.720 251.040 ;
                RECT 0.160 252.080 62.000 252.400 ;
                RECT 69.160 252.080 79.680 252.400 ;
                RECT 1078.960 252.080 1085.720 252.400 ;
                RECT 0.160 253.440 62.000 253.760 ;
                RECT 69.160 253.440 79.680 253.760 ;
                RECT 1078.960 253.440 1085.720 253.760 ;
                RECT 0.160 254.800 62.000 255.120 ;
                RECT 69.160 254.800 79.680 255.120 ;
                RECT 1078.960 254.800 1085.720 255.120 ;
                RECT 0.160 256.160 62.000 256.480 ;
                RECT 69.160 256.160 79.680 256.480 ;
                RECT 1078.960 256.160 1085.720 256.480 ;
                RECT 0.160 257.520 79.680 257.840 ;
                RECT 1078.960 257.520 1085.720 257.840 ;
                RECT 0.160 258.880 65.400 259.200 ;
                RECT 69.160 258.880 79.680 259.200 ;
                RECT 1078.960 258.880 1085.720 259.200 ;
                RECT 0.160 260.240 66.080 260.560 ;
                RECT 69.160 260.240 79.680 260.560 ;
                RECT 1078.960 260.240 1085.720 260.560 ;
                RECT 0.160 261.600 62.000 261.920 ;
                RECT 69.160 261.600 79.680 261.920 ;
                RECT 1078.960 261.600 1085.720 261.920 ;
                RECT 0.160 262.960 62.000 263.280 ;
                RECT 69.160 262.960 79.680 263.280 ;
                RECT 1078.960 262.960 1085.720 263.280 ;
                RECT 0.160 264.320 62.000 264.640 ;
                RECT 69.160 264.320 79.680 264.640 ;
                RECT 1078.960 264.320 1085.720 264.640 ;
                RECT 0.160 265.680 79.680 266.000 ;
                RECT 1078.960 265.680 1085.720 266.000 ;
                RECT 0.160 267.040 62.680 267.360 ;
                RECT 69.160 267.040 79.680 267.360 ;
                RECT 1078.960 267.040 1085.720 267.360 ;
                RECT 0.160 268.400 62.680 268.720 ;
                RECT 69.160 268.400 79.680 268.720 ;
                RECT 1078.960 268.400 1085.720 268.720 ;
                RECT 0.160 269.760 64.720 270.080 ;
                RECT 69.160 269.760 79.680 270.080 ;
                RECT 1078.960 269.760 1085.720 270.080 ;
                RECT 0.160 271.120 62.680 271.440 ;
                RECT 69.160 271.120 79.680 271.440 ;
                RECT 1078.960 271.120 1085.720 271.440 ;
                RECT 0.160 272.480 62.680 272.800 ;
                RECT 69.160 272.480 79.680 272.800 ;
                RECT 1078.960 272.480 1085.720 272.800 ;
                RECT 0.160 273.840 79.680 274.160 ;
                RECT 1078.960 273.840 1085.720 274.160 ;
                RECT 0.160 275.200 62.680 275.520 ;
                RECT 69.160 275.200 79.680 275.520 ;
                RECT 1078.960 275.200 1085.720 275.520 ;
                RECT 0.160 276.560 62.680 276.880 ;
                RECT 69.160 276.560 79.680 276.880 ;
                RECT 1078.960 276.560 1085.720 276.880 ;
                RECT 0.160 277.920 62.680 278.240 ;
                RECT 69.160 277.920 79.680 278.240 ;
                RECT 1078.960 277.920 1085.720 278.240 ;
                RECT 0.160 279.280 67.440 279.600 ;
                RECT 69.160 279.280 79.680 279.600 ;
                RECT 1078.960 279.280 1085.720 279.600 ;
                RECT 0.160 280.640 62.680 280.960 ;
                RECT 69.160 280.640 79.680 280.960 ;
                RECT 1078.960 280.640 1085.720 280.960 ;
                RECT 0.160 282.000 79.680 282.320 ;
                RECT 1078.960 282.000 1085.720 282.320 ;
                RECT 0.160 283.360 63.360 283.680 ;
                RECT 69.160 283.360 79.680 283.680 ;
                RECT 1078.960 283.360 1085.720 283.680 ;
                RECT 0.160 284.720 63.360 285.040 ;
                RECT 69.160 284.720 79.680 285.040 ;
                RECT 1078.960 284.720 1085.720 285.040 ;
                RECT 0.160 286.080 63.360 286.400 ;
                RECT 69.160 286.080 79.680 286.400 ;
                RECT 1078.960 286.080 1085.720 286.400 ;
                RECT 0.160 287.440 63.360 287.760 ;
                RECT 69.160 287.440 79.680 287.760 ;
                RECT 1078.960 287.440 1085.720 287.760 ;
                RECT 0.160 288.800 79.680 289.120 ;
                RECT 1078.960 288.800 1085.720 289.120 ;
                RECT 0.160 290.160 65.400 290.480 ;
                RECT 69.160 290.160 79.680 290.480 ;
                RECT 1078.960 290.160 1085.720 290.480 ;
                RECT 0.160 291.520 63.360 291.840 ;
                RECT 69.160 291.520 79.680 291.840 ;
                RECT 1078.960 291.520 1085.720 291.840 ;
                RECT 0.160 292.880 63.360 293.200 ;
                RECT 69.160 292.880 79.680 293.200 ;
                RECT 1078.960 292.880 1085.720 293.200 ;
                RECT 0.160 294.240 63.360 294.560 ;
                RECT 69.160 294.240 79.680 294.560 ;
                RECT 1078.960 294.240 1085.720 294.560 ;
                RECT 0.160 295.600 63.360 295.920 ;
                RECT 69.160 295.600 79.680 295.920 ;
                RECT 1078.960 295.600 1085.720 295.920 ;
                RECT 0.160 296.960 79.680 297.280 ;
                RECT 1078.960 296.960 1085.720 297.280 ;
                RECT 0.160 298.320 79.680 298.640 ;
                RECT 1078.960 298.320 1085.720 298.640 ;
                RECT 0.160 299.680 278.240 300.000 ;
                RECT 1078.960 299.680 1085.720 300.000 ;
                RECT 0.160 301.040 278.240 301.360 ;
                RECT 1078.960 301.040 1085.720 301.360 ;
                RECT 0.160 302.400 1085.720 302.720 ;
                RECT 0.160 303.760 1085.720 304.080 ;
                RECT 0.160 305.120 1085.720 305.440 ;
                RECT 0.160 306.480 1085.720 306.800 ;
                RECT 0.160 307.840 1085.720 308.160 ;
                RECT 0.160 0.160 1085.720 1.520 ;
                RECT 0.160 311.880 1085.720 313.240 ;
                RECT 282.380 45.895 288.180 47.265 ;
                RECT 1068.680 45.895 1074.480 47.265 ;
                RECT 282.380 51.415 288.180 53.155 ;
                RECT 1068.680 51.415 1074.480 53.155 ;
                RECT 282.380 57.260 288.180 58.830 ;
                RECT 1068.680 57.260 1074.480 58.830 ;
                RECT 282.380 62.850 288.180 64.420 ;
                RECT 1068.680 62.850 1074.480 64.420 ;
                RECT 282.380 90.650 1074.480 91.450 ;
                RECT 282.380 98.330 1074.480 100.420 ;
                RECT 282.380 130.625 1074.480 132.425 ;
                RECT 282.380 85.760 1074.480 86.560 ;
                RECT 282.380 82.750 1074.480 83.550 ;
                RECT 282.380 71.280 1074.480 73.080 ;
                RECT 282.380 155.865 1074.480 158.465 ;
                RECT 282.380 103.755 1074.480 104.045 ;
                RECT 282.380 30.140 1074.480 31.940 ;
                RECT 84.580 170.195 86.500 298.175 ;
                RECT 88.420 170.195 90.340 298.175 ;
                RECT 100.830 170.195 102.750 298.175 ;
                RECT 104.670 170.195 106.590 298.175 ;
                RECT 108.510 170.195 110.430 298.175 ;
                RECT 112.350 170.195 114.270 298.175 ;
                RECT 133.035 170.195 134.955 298.175 ;
                RECT 136.875 170.195 138.795 298.175 ;
                RECT 140.715 170.195 142.635 298.175 ;
                RECT 144.555 170.195 146.475 298.175 ;
                RECT 148.395 170.195 150.315 298.175 ;
                RECT 152.235 170.195 154.155 298.175 ;
                RECT 156.075 170.195 157.995 298.175 ;
                RECT 159.915 170.195 161.835 298.175 ;
                RECT 163.755 170.195 165.675 298.175 ;
                RECT 201.235 170.195 203.155 298.175 ;
                RECT 205.075 170.195 206.995 298.175 ;
                RECT 208.915 170.195 210.835 298.175 ;
                RECT 212.755 170.195 214.675 298.175 ;
                RECT 216.595 170.195 218.515 298.175 ;
                RECT 220.435 170.195 222.355 298.175 ;
                RECT 224.275 170.195 226.195 298.175 ;
                RECT 228.115 170.195 230.035 298.175 ;
                RECT 231.955 170.195 233.875 298.175 ;
                RECT 235.795 170.195 237.715 298.175 ;
                RECT 239.635 170.195 241.555 298.175 ;
                RECT 243.475 170.195 245.395 298.175 ;
                RECT 247.315 170.195 249.235 298.175 ;
                RECT 251.155 170.195 253.075 298.175 ;
                RECT 254.995 170.195 256.915 298.175 ;
                RECT 258.835 170.195 260.755 298.175 ;
                RECT 262.675 170.195 264.595 298.175 ;
                RECT 266.515 170.195 268.435 298.175 ;
                RECT 270.355 170.195 272.275 298.175 ;
                RECT 274.195 170.195 276.115 298.175 ;
                RECT 157.940 60.640 159.860 104.640 ;
                RECT 164.915 60.640 166.835 104.640 ;
                RECT 173.610 60.640 175.530 104.640 ;
                RECT 187.925 60.640 189.845 104.640 ;
                RECT 191.765 60.640 193.685 104.640 ;
                RECT 195.605 60.640 197.525 104.640 ;
                RECT 218.870 60.640 220.790 104.640 ;
                RECT 222.710 60.640 224.630 104.640 ;
                RECT 226.550 60.640 228.470 104.640 ;
                RECT 230.390 60.640 232.310 104.640 ;
                RECT 234.230 60.640 236.150 104.640 ;
                RECT 238.070 60.640 239.990 104.640 ;
                RECT 241.910 60.640 243.830 104.640 ;
                RECT 245.750 60.640 247.670 104.640 ;
                RECT 249.590 60.640 251.510 104.640 ;
                RECT 253.430 60.640 255.350 104.640 ;
                RECT 192.320 134.860 194.240 163.560 ;
                RECT 199.725 134.860 201.645 163.560 ;
                RECT 206.355 134.860 208.105 163.560 ;
                RECT 214.765 134.860 216.685 163.560 ;
                RECT 218.605 134.860 220.525 163.560 ;
                RECT 234.270 134.860 236.190 163.560 ;
                RECT 238.110 134.860 240.030 163.560 ;
                RECT 241.950 134.860 243.870 163.560 ;
                RECT 245.790 134.860 247.710 163.560 ;
                RECT 249.630 134.860 251.550 163.560 ;
                RECT 253.470 134.860 255.390 163.560 ;
                RECT 192.965 110.640 194.885 128.860 ;
                RECT 200.155 110.640 202.075 128.860 ;
                RECT 206.785 110.640 208.535 128.860 ;
                RECT 216.055 110.640 217.975 128.860 ;
                RECT 219.895 110.640 221.815 128.860 ;
                RECT 236.835 110.640 238.755 128.860 ;
                RECT 240.675 110.640 242.595 128.860 ;
                RECT 244.515 110.640 246.435 128.860 ;
                RECT 248.355 110.640 250.275 128.860 ;
                RECT 252.195 110.640 254.115 128.860 ;
                RECT 229.060 49.480 230.980 54.640 ;
                RECT 236.895 49.480 238.815 54.640 ;
                RECT 248.615 49.480 250.535 54.640 ;
                RECT 252.455 49.480 254.375 54.640 ;
                RECT 24.860 172.465 34.020 173.215 ;
                RECT 24.860 177.220 34.020 179.140 ;
                RECT 98.040 160.250 114.080 161.050 ;
                RECT 78.840 160.960 96.080 162.650 ;
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 291.160 5.560 ;
                RECT 292.880 5.240 297.280 5.560 ;
                RECT 299.000 5.240 303.400 5.560 ;
                RECT 305.120 5.240 309.520 5.560 ;
                RECT 311.240 5.240 315.640 5.560 ;
                RECT 317.360 5.240 321.760 5.560 ;
                RECT 323.480 5.240 327.880 5.560 ;
                RECT 329.600 5.240 334.000 5.560 ;
                RECT 335.720 5.240 340.120 5.560 ;
                RECT 341.840 5.240 346.240 5.560 ;
                RECT 347.960 5.240 352.360 5.560 ;
                RECT 354.080 5.240 358.480 5.560 ;
                RECT 360.200 5.240 364.600 5.560 ;
                RECT 366.320 5.240 370.720 5.560 ;
                RECT 372.440 5.240 376.840 5.560 ;
                RECT 378.560 5.240 382.960 5.560 ;
                RECT 384.680 5.240 389.080 5.560 ;
                RECT 390.800 5.240 395.200 5.560 ;
                RECT 396.920 5.240 401.320 5.560 ;
                RECT 403.040 5.240 407.440 5.560 ;
                RECT 409.160 5.240 413.560 5.560 ;
                RECT 415.280 5.240 419.680 5.560 ;
                RECT 421.400 5.240 425.800 5.560 ;
                RECT 427.520 5.240 431.920 5.560 ;
                RECT 432.960 5.240 438.040 5.560 ;
                RECT 439.080 5.240 444.160 5.560 ;
                RECT 445.200 5.240 450.280 5.560 ;
                RECT 451.320 5.240 456.400 5.560 ;
                RECT 457.440 5.240 462.520 5.560 ;
                RECT 463.560 5.240 468.640 5.560 ;
                RECT 469.680 5.240 474.760 5.560 ;
                RECT 475.800 5.240 480.880 5.560 ;
                RECT 481.920 5.240 486.320 5.560 ;
                RECT 488.040 5.240 492.440 5.560 ;
                RECT 494.160 5.240 498.560 5.560 ;
                RECT 500.280 5.240 504.680 5.560 ;
                RECT 506.400 5.240 510.800 5.560 ;
                RECT 512.520 5.240 516.920 5.560 ;
                RECT 518.640 5.240 523.040 5.560 ;
                RECT 524.760 5.240 529.160 5.560 ;
                RECT 530.880 5.240 535.280 5.560 ;
                RECT 537.000 5.240 541.400 5.560 ;
                RECT 543.120 5.240 547.520 5.560 ;
                RECT 549.240 5.240 553.640 5.560 ;
                RECT 555.360 5.240 559.760 5.560 ;
                RECT 561.480 5.240 565.880 5.560 ;
                RECT 567.600 5.240 572.000 5.560 ;
                RECT 573.720 5.240 578.120 5.560 ;
                RECT 579.840 5.240 584.240 5.560 ;
                RECT 585.960 5.240 590.360 5.560 ;
                RECT 592.080 5.240 596.480 5.560 ;
                RECT 598.200 5.240 602.600 5.560 ;
                RECT 604.320 5.240 608.720 5.560 ;
                RECT 610.440 5.240 614.840 5.560 ;
                RECT 616.560 5.240 620.960 5.560 ;
                RECT 622.680 5.240 627.080 5.560 ;
                RECT 628.800 5.240 633.200 5.560 ;
                RECT 634.920 5.240 639.320 5.560 ;
                RECT 640.360 5.240 645.440 5.560 ;
                RECT 646.480 5.240 651.560 5.560 ;
                RECT 652.600 5.240 657.680 5.560 ;
                RECT 658.720 5.240 663.800 5.560 ;
                RECT 664.840 5.240 669.920 5.560 ;
                RECT 670.960 5.240 676.040 5.560 ;
                RECT 677.080 5.240 682.160 5.560 ;
                RECT 683.200 5.240 688.280 5.560 ;
                RECT 689.320 5.240 693.720 5.560 ;
                RECT 695.440 5.240 699.840 5.560 ;
                RECT 701.560 5.240 705.960 5.560 ;
                RECT 707.680 5.240 712.080 5.560 ;
                RECT 713.800 5.240 718.200 5.560 ;
                RECT 719.920 5.240 724.320 5.560 ;
                RECT 726.040 5.240 730.440 5.560 ;
                RECT 732.160 5.240 736.560 5.560 ;
                RECT 738.280 5.240 742.680 5.560 ;
                RECT 744.400 5.240 748.800 5.560 ;
                RECT 750.520 5.240 754.920 5.560 ;
                RECT 756.640 5.240 761.040 5.560 ;
                RECT 762.760 5.240 767.160 5.560 ;
                RECT 768.880 5.240 773.280 5.560 ;
                RECT 775.000 5.240 779.400 5.560 ;
                RECT 781.120 5.240 785.520 5.560 ;
                RECT 787.240 5.240 791.640 5.560 ;
                RECT 793.360 5.240 797.760 5.560 ;
                RECT 799.480 5.240 803.880 5.560 ;
                RECT 805.600 5.240 810.000 5.560 ;
                RECT 811.720 5.240 816.120 5.560 ;
                RECT 817.840 5.240 822.240 5.560 ;
                RECT 823.960 5.240 828.360 5.560 ;
                RECT 830.080 5.240 834.480 5.560 ;
                RECT 836.200 5.240 840.600 5.560 ;
                RECT 842.320 5.240 846.720 5.560 ;
                RECT 847.760 5.240 852.840 5.560 ;
                RECT 853.880 5.240 858.960 5.560 ;
                RECT 860.000 5.240 865.080 5.560 ;
                RECT 866.120 5.240 871.200 5.560 ;
                RECT 872.240 5.240 877.320 5.560 ;
                RECT 878.360 5.240 883.440 5.560 ;
                RECT 884.480 5.240 889.560 5.560 ;
                RECT 890.600 5.240 895.680 5.560 ;
                RECT 896.720 5.240 901.120 5.560 ;
                RECT 902.840 5.240 907.240 5.560 ;
                RECT 908.960 5.240 913.360 5.560 ;
                RECT 915.080 5.240 919.480 5.560 ;
                RECT 921.200 5.240 925.600 5.560 ;
                RECT 927.320 5.240 931.720 5.560 ;
                RECT 933.440 5.240 937.840 5.560 ;
                RECT 939.560 5.240 943.960 5.560 ;
                RECT 945.680 5.240 950.080 5.560 ;
                RECT 951.800 5.240 956.200 5.560 ;
                RECT 957.920 5.240 962.320 5.560 ;
                RECT 964.040 5.240 968.440 5.560 ;
                RECT 970.160 5.240 974.560 5.560 ;
                RECT 976.280 5.240 980.680 5.560 ;
                RECT 982.400 5.240 986.800 5.560 ;
                RECT 988.520 5.240 992.920 5.560 ;
                RECT 994.640 5.240 999.040 5.560 ;
                RECT 1000.760 5.240 1005.160 5.560 ;
                RECT 1006.880 5.240 1011.280 5.560 ;
                RECT 1013.000 5.240 1017.400 5.560 ;
                RECT 1019.120 5.240 1023.520 5.560 ;
                RECT 1025.240 5.240 1029.640 5.560 ;
                RECT 1031.360 5.240 1035.760 5.560 ;
                RECT 1037.480 5.240 1041.880 5.560 ;
                RECT 1043.600 5.240 1048.000 5.560 ;
                RECT 1049.720 5.240 1054.120 5.560 ;
                RECT 1055.160 5.240 1060.240 5.560 ;
                RECT 1061.280 5.240 1066.360 5.560 ;
                RECT 1067.400 5.240 1083.000 5.560 ;
                RECT 2.880 6.600 1083.000 6.920 ;
                RECT 2.880 7.960 1083.000 8.280 ;
                RECT 2.880 9.320 257.840 9.640 ;
                RECT 286.760 9.320 1083.000 9.640 ;
                RECT 2.880 10.680 1083.000 11.000 ;
                RECT 2.880 12.040 1083.000 12.360 ;
                RECT 2.880 13.400 195.280 13.720 ;
                RECT 258.880 13.400 1083.000 13.720 ;
                RECT 2.880 14.760 1083.000 15.080 ;
                RECT 2.880 16.120 1083.000 16.440 ;
                RECT 2.880 17.480 195.280 17.800 ;
                RECT 258.200 17.480 1083.000 17.800 ;
                RECT 2.880 18.840 1083.000 19.160 ;
                RECT 2.880 20.200 1083.000 20.520 ;
                RECT 2.880 21.560 1083.000 21.880 ;
                RECT 2.880 22.920 1083.000 23.240 ;
                RECT 2.880 24.280 280.960 24.600 ;
                RECT 1076.240 24.280 1083.000 24.600 ;
                RECT 2.880 25.640 280.960 25.960 ;
                RECT 1076.240 25.640 1083.000 25.960 ;
                RECT 2.880 27.000 280.960 27.320 ;
                RECT 1076.240 27.000 1083.000 27.320 ;
                RECT 2.880 28.360 280.960 28.680 ;
                RECT 1076.240 28.360 1083.000 28.680 ;
                RECT 2.880 29.720 280.960 30.040 ;
                RECT 1076.240 29.720 1083.000 30.040 ;
                RECT 2.880 31.080 280.960 31.400 ;
                RECT 1076.240 31.080 1083.000 31.400 ;
                RECT 2.880 32.440 280.960 32.760 ;
                RECT 1076.240 32.440 1083.000 32.760 ;
                RECT 2.880 33.800 144.280 34.120 ;
                RECT 235.760 33.800 280.960 34.120 ;
                RECT 1076.240 33.800 1083.000 34.120 ;
                RECT 2.880 35.160 142.920 35.480 ;
                RECT 241.880 35.160 280.960 35.480 ;
                RECT 1076.240 35.160 1083.000 35.480 ;
                RECT 2.880 36.520 123.200 36.840 ;
                RECT 258.880 36.520 280.960 36.840 ;
                RECT 1076.240 36.520 1083.000 36.840 ;
                RECT 2.880 37.880 122.520 38.200 ;
                RECT 254.800 37.880 280.960 38.200 ;
                RECT 1076.240 37.880 1083.000 38.200 ;
                RECT 2.880 39.240 280.960 39.560 ;
                RECT 1076.240 39.240 1083.000 39.560 ;
                RECT 2.880 40.600 280.960 40.920 ;
                RECT 1076.240 40.600 1083.000 40.920 ;
                RECT 2.880 41.960 280.280 42.280 ;
                RECT 1076.240 41.960 1083.000 42.280 ;
                RECT 2.880 43.320 280.960 43.640 ;
                RECT 1076.240 43.320 1083.000 43.640 ;
                RECT 2.880 44.680 118.440 45.000 ;
                RECT 129.680 44.680 280.960 45.000 ;
                RECT 1076.240 44.680 1083.000 45.000 ;
                RECT 2.880 46.040 119.800 46.360 ;
                RECT 123.560 46.040 280.960 46.360 ;
                RECT 1076.240 46.040 1083.000 46.360 ;
                RECT 2.880 47.400 121.160 47.720 ;
                RECT 125.600 47.400 133.400 47.720 ;
                RECT 135.800 47.400 280.960 47.720 ;
                RECT 1076.240 47.400 1083.000 47.720 ;
                RECT 2.880 48.760 280.960 49.080 ;
                RECT 1076.240 48.760 1083.000 49.080 ;
                RECT 2.880 50.120 127.960 50.440 ;
                RECT 136.480 50.120 225.200 50.440 ;
                RECT 254.800 50.120 280.960 50.440 ;
                RECT 1076.240 50.120 1083.000 50.440 ;
                RECT 2.880 51.480 120.480 51.800 ;
                RECT 129.680 51.480 225.200 51.800 ;
                RECT 1076.240 51.480 1083.000 51.800 ;
                RECT 2.880 52.840 123.880 53.160 ;
                RECT 129.000 52.840 225.200 53.160 ;
                RECT 1076.240 52.840 1083.000 53.160 ;
                RECT 2.880 54.200 141.560 54.520 ;
                RECT 222.840 54.200 225.200 54.520 ;
                RECT 254.800 54.200 280.960 54.520 ;
                RECT 1076.240 54.200 1083.000 54.520 ;
                RECT 2.880 55.560 119.800 55.880 ;
                RECT 129.680 55.560 280.960 55.880 ;
                RECT 1076.240 55.560 1083.000 55.880 ;
                RECT 2.880 56.920 127.960 57.240 ;
                RECT 135.120 56.920 280.960 57.240 ;
                RECT 1076.240 56.920 1083.000 57.240 ;
                RECT 2.880 58.280 126.600 58.600 ;
                RECT 129.680 58.280 280.960 58.600 ;
                RECT 1076.240 58.280 1083.000 58.600 ;
                RECT 2.880 59.640 280.960 59.960 ;
                RECT 1076.240 59.640 1083.000 59.960 ;
                RECT 2.880 61.000 127.960 61.320 ;
                RECT 135.800 61.000 142.920 61.320 ;
                RECT 148.720 61.000 153.800 61.320 ;
                RECT 256.160 61.000 280.960 61.320 ;
                RECT 1076.240 61.000 1083.000 61.320 ;
                RECT 2.880 62.360 124.560 62.680 ;
                RECT 129.680 62.360 144.280 62.680 ;
                RECT 147.360 62.360 153.800 62.680 ;
                RECT 269.080 62.360 280.960 62.680 ;
                RECT 1076.240 62.360 1083.000 62.680 ;
                RECT 2.880 63.720 126.600 64.040 ;
                RECT 129.680 63.720 153.800 64.040 ;
                RECT 256.160 63.720 280.960 64.040 ;
                RECT 1076.240 63.720 1083.000 64.040 ;
                RECT 2.880 65.080 130.680 65.400 ;
                RECT 141.240 65.080 153.800 65.400 ;
                RECT 267.040 65.080 280.960 65.400 ;
                RECT 1076.240 65.080 1083.000 65.400 ;
                RECT 2.880 66.440 117.760 66.760 ;
                RECT 135.800 66.440 153.800 66.760 ;
                RECT 269.080 66.440 280.960 66.760 ;
                RECT 1076.240 66.440 1083.000 66.760 ;
                RECT 2.880 67.800 126.600 68.120 ;
                RECT 129.680 67.800 136.800 68.120 ;
                RECT 142.600 67.800 153.800 68.120 ;
                RECT 269.080 67.800 280.960 68.120 ;
                RECT 1076.240 67.800 1083.000 68.120 ;
                RECT 2.880 69.160 139.520 69.480 ;
                RECT 143.280 69.160 153.800 69.480 ;
                RECT 267.040 69.160 280.960 69.480 ;
                RECT 1076.240 69.160 1083.000 69.480 ;
                RECT 2.880 70.520 118.440 70.840 ;
                RECT 132.400 70.520 153.800 70.840 ;
                RECT 269.080 70.520 280.960 70.840 ;
                RECT 1076.240 70.520 1083.000 70.840 ;
                RECT 2.880 71.880 127.280 72.200 ;
                RECT 135.800 71.880 153.800 72.200 ;
                RECT 267.040 71.880 280.960 72.200 ;
                RECT 1076.240 71.880 1083.000 72.200 ;
                RECT 2.880 73.240 125.240 73.560 ;
                RECT 136.480 73.240 153.800 73.560 ;
                RECT 273.160 73.240 280.960 73.560 ;
                RECT 1076.240 73.240 1083.000 73.560 ;
                RECT 2.880 74.600 153.800 74.920 ;
                RECT 273.160 74.600 280.960 74.920 ;
                RECT 1076.240 74.600 1083.000 74.920 ;
                RECT 2.880 75.960 121.160 76.280 ;
                RECT 123.560 75.960 153.800 76.280 ;
                RECT 271.120 75.960 280.960 76.280 ;
                RECT 1076.240 75.960 1083.000 76.280 ;
                RECT 2.880 77.320 119.800 77.640 ;
                RECT 129.680 77.320 153.800 77.640 ;
                RECT 273.160 77.320 280.960 77.640 ;
                RECT 1076.240 77.320 1083.000 77.640 ;
                RECT 2.880 78.680 153.800 79.000 ;
                RECT 256.160 78.680 280.960 79.000 ;
                RECT 1076.240 78.680 1083.000 79.000 ;
                RECT 2.880 80.040 153.800 80.360 ;
                RECT 273.160 80.040 280.960 80.360 ;
                RECT 1076.240 80.040 1083.000 80.360 ;
                RECT 2.880 81.400 126.600 81.720 ;
                RECT 129.000 81.400 153.800 81.720 ;
                RECT 273.160 81.400 280.960 81.720 ;
                RECT 1076.240 81.400 1083.000 81.720 ;
                RECT 2.880 82.760 127.960 83.080 ;
                RECT 129.680 82.760 153.800 83.080 ;
                RECT 256.160 82.760 280.960 83.080 ;
                RECT 1076.240 82.760 1083.000 83.080 ;
                RECT 2.880 84.120 126.600 84.440 ;
                RECT 129.000 84.120 153.800 84.440 ;
                RECT 275.200 84.120 280.960 84.440 ;
                RECT 1076.240 84.120 1083.000 84.440 ;
                RECT 2.880 85.480 125.240 85.800 ;
                RECT 135.800 85.480 153.800 85.800 ;
                RECT 277.240 85.480 280.960 85.800 ;
                RECT 1076.240 85.480 1083.000 85.800 ;
                RECT 2.880 86.840 117.760 87.160 ;
                RECT 129.680 86.840 153.800 87.160 ;
                RECT 256.160 86.840 280.960 87.160 ;
                RECT 1076.240 86.840 1083.000 87.160 ;
                RECT 2.880 88.200 127.280 88.520 ;
                RECT 129.680 88.200 153.800 88.520 ;
                RECT 277.240 88.200 280.960 88.520 ;
                RECT 1076.240 88.200 1083.000 88.520 ;
                RECT 2.880 89.560 153.800 89.880 ;
                RECT 277.240 89.560 280.960 89.880 ;
                RECT 1076.240 89.560 1083.000 89.880 ;
                RECT 2.880 90.920 153.800 91.240 ;
                RECT 275.200 90.920 280.960 91.240 ;
                RECT 1076.240 90.920 1083.000 91.240 ;
                RECT 2.880 92.280 115.040 92.600 ;
                RECT 128.320 92.280 153.800 92.600 ;
                RECT 277.240 92.280 280.960 92.600 ;
                RECT 1076.240 92.280 1083.000 92.600 ;
                RECT 2.880 93.640 124.560 93.960 ;
                RECT 132.400 93.640 153.800 93.960 ;
                RECT 1076.240 93.640 1083.000 93.960 ;
                RECT 2.880 95.000 153.800 95.320 ;
                RECT 1076.240 95.000 1083.000 95.320 ;
                RECT 2.880 96.360 121.840 96.680 ;
                RECT 125.600 96.360 153.800 96.680 ;
                RECT 1076.240 96.360 1083.000 96.680 ;
                RECT 2.880 97.720 120.480 98.040 ;
                RECT 138.520 97.720 153.800 98.040 ;
                RECT 1076.240 97.720 1083.000 98.040 ;
                RECT 2.880 99.080 153.800 99.400 ;
                RECT 1076.240 99.080 1083.000 99.400 ;
                RECT 2.880 100.440 121.840 100.760 ;
                RECT 125.600 100.440 153.800 100.760 ;
                RECT 1076.240 100.440 1083.000 100.760 ;
                RECT 2.880 101.800 123.880 102.120 ;
                RECT 135.120 101.800 153.800 102.120 ;
                RECT 1076.240 101.800 1083.000 102.120 ;
                RECT 2.880 103.160 117.760 103.480 ;
                RECT 122.200 103.160 153.800 103.480 ;
                RECT 1076.240 103.160 1083.000 103.480 ;
                RECT 2.880 104.520 153.800 104.840 ;
                RECT 256.160 104.520 280.960 104.840 ;
                RECT 1076.240 104.520 1083.000 104.840 ;
                RECT 2.880 105.880 133.400 106.200 ;
                RECT 136.480 105.880 280.960 106.200 ;
                RECT 1076.240 105.880 1083.000 106.200 ;
                RECT 2.880 107.240 118.440 107.560 ;
                RECT 125.600 107.240 280.960 107.560 ;
                RECT 1076.240 107.240 1083.000 107.560 ;
                RECT 2.880 108.600 123.880 108.920 ;
                RECT 128.320 108.600 280.960 108.920 ;
                RECT 1076.240 108.600 1083.000 108.920 ;
                RECT 2.880 109.960 280.960 110.280 ;
                RECT 1076.240 109.960 1083.000 110.280 ;
                RECT 2.880 111.320 120.480 111.640 ;
                RECT 125.600 111.320 189.160 111.640 ;
                RECT 254.800 111.320 280.960 111.640 ;
                RECT 1076.240 111.320 1083.000 111.640 ;
                RECT 2.880 112.680 189.160 113.000 ;
                RECT 254.800 112.680 280.960 113.000 ;
                RECT 1076.240 112.680 1083.000 113.000 ;
                RECT 2.880 114.040 126.600 114.360 ;
                RECT 135.120 114.040 189.160 114.360 ;
                RECT 254.800 114.040 280.960 114.360 ;
                RECT 1076.240 114.040 1083.000 114.360 ;
                RECT 2.880 115.400 189.160 115.720 ;
                RECT 254.800 115.400 280.960 115.720 ;
                RECT 1076.240 115.400 1083.000 115.720 ;
                RECT 2.880 116.760 189.160 117.080 ;
                RECT 254.800 116.760 280.960 117.080 ;
                RECT 1076.240 116.760 1083.000 117.080 ;
                RECT 2.880 118.120 121.160 118.440 ;
                RECT 123.560 118.120 189.160 118.440 ;
                RECT 1076.240 118.120 1083.000 118.440 ;
                RECT 2.880 119.480 189.160 119.800 ;
                RECT 254.800 119.480 276.880 119.800 ;
                RECT 1076.240 119.480 1083.000 119.800 ;
                RECT 2.880 120.840 96.680 121.160 ;
                RECT 115.400 120.840 189.160 121.160 ;
                RECT 254.800 120.840 272.800 121.160 ;
                RECT 1076.240 120.840 1083.000 121.160 ;
                RECT 2.880 122.200 96.680 122.520 ;
                RECT 115.400 122.200 189.160 122.520 ;
                RECT 254.800 122.200 272.800 122.520 ;
                RECT 1076.240 122.200 1083.000 122.520 ;
                RECT 2.880 123.560 96.680 123.880 ;
                RECT 115.400 123.560 189.160 123.880 ;
                RECT 254.800 123.560 268.720 123.880 ;
                RECT 1076.240 123.560 1083.000 123.880 ;
                RECT 2.880 124.920 96.680 125.240 ;
                RECT 115.400 124.920 189.160 125.240 ;
                RECT 254.800 124.920 264.640 125.240 ;
                RECT 1076.240 124.920 1083.000 125.240 ;
                RECT 2.880 126.280 96.680 126.600 ;
                RECT 115.400 126.280 189.160 126.600 ;
                RECT 254.800 126.280 264.640 126.600 ;
                RECT 1076.240 126.280 1083.000 126.600 ;
                RECT 2.880 127.640 96.680 127.960 ;
                RECT 115.400 127.640 189.160 127.960 ;
                RECT 254.800 127.640 280.960 127.960 ;
                RECT 1076.240 127.640 1083.000 127.960 ;
                RECT 2.880 129.000 96.680 129.320 ;
                RECT 115.400 129.000 189.160 129.320 ;
                RECT 254.800 129.000 280.960 129.320 ;
                RECT 1076.240 129.000 1083.000 129.320 ;
                RECT 2.880 130.360 96.680 130.680 ;
                RECT 115.400 130.360 280.960 130.680 ;
                RECT 1076.240 130.360 1083.000 130.680 ;
                RECT 2.880 131.720 96.680 132.040 ;
                RECT 115.400 131.720 280.960 132.040 ;
                RECT 1076.240 131.720 1083.000 132.040 ;
                RECT 2.880 133.080 96.680 133.400 ;
                RECT 115.400 133.080 280.960 133.400 ;
                RECT 1076.240 133.080 1083.000 133.400 ;
                RECT 2.880 134.440 96.680 134.760 ;
                RECT 115.400 134.440 187.800 134.760 ;
                RECT 256.160 134.440 280.960 134.760 ;
                RECT 1076.240 134.440 1083.000 134.760 ;
                RECT 2.880 135.800 96.680 136.120 ;
                RECT 116.080 135.800 187.800 136.120 ;
                RECT 256.160 135.800 280.960 136.120 ;
                RECT 1076.240 135.800 1083.000 136.120 ;
                RECT 2.880 137.160 96.680 137.480 ;
                RECT 115.400 137.160 187.800 137.480 ;
                RECT 256.160 137.160 280.960 137.480 ;
                RECT 1076.240 137.160 1083.000 137.480 ;
                RECT 2.880 138.520 96.680 138.840 ;
                RECT 115.400 138.520 187.800 138.840 ;
                RECT 256.160 138.520 280.960 138.840 ;
                RECT 1076.240 138.520 1083.000 138.840 ;
                RECT 2.880 139.880 96.680 140.200 ;
                RECT 115.400 139.880 187.800 140.200 ;
                RECT 256.160 139.880 280.960 140.200 ;
                RECT 1076.240 139.880 1083.000 140.200 ;
                RECT 2.880 141.240 96.680 141.560 ;
                RECT 115.400 141.240 123.200 141.560 ;
                RECT 125.600 141.240 187.800 141.560 ;
                RECT 256.160 141.240 266.680 141.560 ;
                RECT 1076.240 141.240 1083.000 141.560 ;
                RECT 2.880 142.600 96.680 142.920 ;
                RECT 115.400 142.600 187.800 142.920 ;
                RECT 256.160 142.600 266.680 142.920 ;
                RECT 1076.240 142.600 1083.000 142.920 ;
                RECT 2.880 143.960 96.680 144.280 ;
                RECT 115.400 143.960 187.800 144.280 ;
                RECT 256.160 143.960 270.760 144.280 ;
                RECT 1076.240 143.960 1083.000 144.280 ;
                RECT 2.880 145.320 96.680 145.640 ;
                RECT 115.400 145.320 187.800 145.640 ;
                RECT 256.160 145.320 270.760 145.640 ;
                RECT 1076.240 145.320 1083.000 145.640 ;
                RECT 2.880 146.680 96.680 147.000 ;
                RECT 115.400 146.680 187.800 147.000 ;
                RECT 256.160 146.680 274.840 147.000 ;
                RECT 1076.240 146.680 1083.000 147.000 ;
                RECT 2.880 148.040 96.680 148.360 ;
                RECT 115.400 148.040 187.800 148.360 ;
                RECT 256.160 148.040 278.920 148.360 ;
                RECT 1076.240 148.040 1083.000 148.360 ;
                RECT 2.880 149.400 96.680 149.720 ;
                RECT 115.400 149.400 187.800 149.720 ;
                RECT 256.160 149.400 278.920 149.720 ;
                RECT 1076.240 149.400 1083.000 149.720 ;
                RECT 2.880 150.760 96.680 151.080 ;
                RECT 115.400 150.760 187.800 151.080 ;
                RECT 1076.240 150.760 1083.000 151.080 ;
                RECT 2.880 152.120 96.680 152.440 ;
                RECT 115.400 152.120 119.800 152.440 ;
                RECT 125.600 152.120 187.800 152.440 ;
                RECT 1076.240 152.120 1083.000 152.440 ;
                RECT 2.880 153.480 96.680 153.800 ;
                RECT 115.400 153.480 187.800 153.800 ;
                RECT 256.160 153.480 280.960 153.800 ;
                RECT 1076.240 153.480 1083.000 153.800 ;
                RECT 2.880 154.840 187.800 155.160 ;
                RECT 256.160 154.840 280.960 155.160 ;
                RECT 1076.240 154.840 1083.000 155.160 ;
                RECT 2.880 156.200 187.800 156.520 ;
                RECT 256.160 156.200 280.960 156.520 ;
                RECT 1076.240 156.200 1083.000 156.520 ;
                RECT 2.880 157.560 78.320 157.880 ;
                RECT 97.040 157.560 123.880 157.880 ;
                RECT 129.680 157.560 187.800 157.880 ;
                RECT 256.160 157.560 280.960 157.880 ;
                RECT 1076.240 157.560 1083.000 157.880 ;
                RECT 2.880 158.920 78.320 159.240 ;
                RECT 97.040 158.920 102.800 159.240 ;
                RECT 109.960 158.920 187.800 159.240 ;
                RECT 256.160 158.920 280.960 159.240 ;
                RECT 1076.240 158.920 1083.000 159.240 ;
                RECT 2.880 160.280 78.320 160.600 ;
                RECT 114.720 160.280 187.800 160.600 ;
                RECT 1076.240 160.280 1083.000 160.600 ;
                RECT 2.880 161.640 78.320 161.960 ;
                RECT 97.040 161.640 187.800 161.960 ;
                RECT 1076.240 161.640 1083.000 161.960 ;
                RECT 2.880 163.000 75.600 163.320 ;
                RECT 109.960 163.000 117.760 163.320 ;
                RECT 128.320 163.000 187.800 163.320 ;
                RECT 256.160 163.000 280.960 163.320 ;
                RECT 1076.240 163.000 1083.000 163.320 ;
                RECT 2.880 164.360 102.800 164.680 ;
                RECT 122.880 164.360 1083.000 164.680 ;
                RECT 2.880 165.720 30.720 166.040 ;
                RECT 122.200 165.720 1083.000 166.040 ;
                RECT 2.880 167.080 278.240 167.400 ;
                RECT 1078.960 167.080 1083.000 167.400 ;
                RECT 2.880 168.440 278.240 168.760 ;
                RECT 1078.960 168.440 1083.000 168.760 ;
                RECT 2.880 169.800 25.960 170.120 ;
                RECT 32.440 169.800 79.680 170.120 ;
                RECT 1078.960 169.800 1083.000 170.120 ;
                RECT 2.880 171.160 23.920 171.480 ;
                RECT 46.720 171.160 79.680 171.480 ;
                RECT 1078.960 171.160 1083.000 171.480 ;
                RECT 2.880 172.520 23.920 172.840 ;
                RECT 46.040 172.520 59.280 172.840 ;
                RECT 69.160 172.520 79.680 172.840 ;
                RECT 1078.960 172.520 1083.000 172.840 ;
                RECT 2.880 173.880 38.200 174.200 ;
                RECT 44.680 173.880 59.280 174.200 ;
                RECT 69.160 173.880 79.680 174.200 ;
                RECT 1078.960 173.880 1083.000 174.200 ;
                RECT 2.880 175.240 23.920 175.560 ;
                RECT 34.480 175.240 59.280 175.560 ;
                RECT 69.160 175.240 79.680 175.560 ;
                RECT 1078.960 175.240 1083.000 175.560 ;
                RECT 2.880 176.600 23.920 176.920 ;
                RECT 34.480 176.600 59.280 176.920 ;
                RECT 69.160 176.600 79.680 176.920 ;
                RECT 1078.960 176.600 1083.000 176.920 ;
                RECT 2.880 177.960 23.920 178.280 ;
                RECT 34.480 177.960 59.280 178.280 ;
                RECT 69.160 177.960 79.680 178.280 ;
                RECT 1078.960 177.960 1083.000 178.280 ;
                RECT 2.880 179.320 23.920 179.640 ;
                RECT 34.480 179.320 79.680 179.640 ;
                RECT 1078.960 179.320 1083.000 179.640 ;
                RECT 2.880 180.680 59.280 181.000 ;
                RECT 69.160 180.680 79.680 181.000 ;
                RECT 1078.960 180.680 1083.000 181.000 ;
                RECT 2.880 182.040 59.280 182.360 ;
                RECT 69.160 182.040 79.680 182.360 ;
                RECT 1078.960 182.040 1083.000 182.360 ;
                RECT 2.880 183.400 17.120 183.720 ;
                RECT 19.520 183.400 59.960 183.720 ;
                RECT 69.160 183.400 79.680 183.720 ;
                RECT 1078.960 183.400 1083.000 183.720 ;
                RECT 2.880 184.760 16.440 185.080 ;
                RECT 19.520 184.760 59.280 185.080 ;
                RECT 69.160 184.760 79.680 185.080 ;
                RECT 1078.960 184.760 1083.000 185.080 ;
                RECT 2.880 186.120 59.280 186.440 ;
                RECT 67.120 186.120 79.680 186.440 ;
                RECT 1078.960 186.120 1083.000 186.440 ;
                RECT 2.880 187.480 15.760 187.800 ;
                RECT 19.520 187.480 32.760 187.800 ;
                RECT 37.200 187.480 64.040 187.800 ;
                RECT 69.160 187.480 79.680 187.800 ;
                RECT 1078.960 187.480 1083.000 187.800 ;
                RECT 2.880 188.840 15.080 189.160 ;
                RECT 19.520 188.840 32.760 189.160 ;
                RECT 37.880 188.840 59.280 189.160 ;
                RECT 69.160 188.840 79.680 189.160 ;
                RECT 1078.960 188.840 1083.000 189.160 ;
                RECT 2.880 190.200 59.280 190.520 ;
                RECT 69.160 190.200 79.680 190.520 ;
                RECT 1078.960 190.200 1083.000 190.520 ;
                RECT 2.880 191.560 14.400 191.880 ;
                RECT 19.520 191.560 32.760 191.880 ;
                RECT 38.560 191.560 59.280 191.880 ;
                RECT 69.160 191.560 79.680 191.880 ;
                RECT 1078.960 191.560 1083.000 191.880 ;
                RECT 2.880 192.920 13.720 193.240 ;
                RECT 19.520 192.920 32.760 193.240 ;
                RECT 39.240 192.920 59.280 193.240 ;
                RECT 69.160 192.920 79.680 193.240 ;
                RECT 1078.960 192.920 1083.000 193.240 ;
                RECT 2.880 194.280 13.040 194.600 ;
                RECT 19.520 194.280 32.760 194.600 ;
                RECT 39.240 194.280 59.280 194.600 ;
                RECT 67.800 194.280 79.680 194.600 ;
                RECT 1078.960 194.280 1083.000 194.600 ;
                RECT 2.880 195.640 12.360 195.960 ;
                RECT 19.520 195.640 65.400 195.960 ;
                RECT 69.160 195.640 79.680 195.960 ;
                RECT 1078.960 195.640 1083.000 195.960 ;
                RECT 2.880 197.000 59.280 197.320 ;
                RECT 69.160 197.000 79.680 197.320 ;
                RECT 1078.960 197.000 1083.000 197.320 ;
                RECT 2.880 198.360 11.680 198.680 ;
                RECT 19.520 198.360 59.280 198.680 ;
                RECT 69.160 198.360 79.680 198.680 ;
                RECT 1078.960 198.360 1083.000 198.680 ;
                RECT 2.880 199.720 11.000 200.040 ;
                RECT 19.520 199.720 59.280 200.040 ;
                RECT 69.160 199.720 79.680 200.040 ;
                RECT 1078.960 199.720 1083.000 200.040 ;
                RECT 2.880 201.080 10.320 201.400 ;
                RECT 19.520 201.080 59.280 201.400 ;
                RECT 69.160 201.080 79.680 201.400 ;
                RECT 1078.960 201.080 1083.000 201.400 ;
                RECT 2.880 202.440 79.680 202.760 ;
                RECT 1078.960 202.440 1083.000 202.760 ;
                RECT 2.880 203.800 9.640 204.120 ;
                RECT 19.520 203.800 32.760 204.120 ;
                RECT 35.840 203.800 60.640 204.120 ;
                RECT 69.160 203.800 79.680 204.120 ;
                RECT 1078.960 203.800 1083.000 204.120 ;
                RECT 2.880 205.160 64.040 205.480 ;
                RECT 69.160 205.160 79.680 205.480 ;
                RECT 1078.960 205.160 1083.000 205.480 ;
                RECT 2.880 206.520 64.720 206.840 ;
                RECT 69.160 206.520 79.680 206.840 ;
                RECT 1078.960 206.520 1083.000 206.840 ;
                RECT 2.880 207.880 60.640 208.200 ;
                RECT 69.160 207.880 79.680 208.200 ;
                RECT 1078.960 207.880 1083.000 208.200 ;
                RECT 2.880 209.240 60.640 209.560 ;
                RECT 69.160 209.240 79.680 209.560 ;
                RECT 1078.960 209.240 1083.000 209.560 ;
                RECT 2.880 210.600 37.520 210.920 ;
                RECT 46.720 210.600 79.680 210.920 ;
                RECT 1078.960 210.600 1083.000 210.920 ;
                RECT 2.880 211.960 36.160 212.280 ;
                RECT 46.040 211.960 60.640 212.280 ;
                RECT 69.160 211.960 79.680 212.280 ;
                RECT 1078.960 211.960 1083.000 212.280 ;
                RECT 2.880 213.320 34.800 213.640 ;
                RECT 44.680 213.320 59.280 213.640 ;
                RECT 69.160 213.320 79.680 213.640 ;
                RECT 1078.960 213.320 1083.000 213.640 ;
                RECT 2.880 214.680 59.280 215.000 ;
                RECT 69.160 214.680 79.680 215.000 ;
                RECT 1078.960 214.680 1083.000 215.000 ;
                RECT 2.880 216.040 59.280 216.360 ;
                RECT 69.160 216.040 79.680 216.360 ;
                RECT 1078.960 216.040 1083.000 216.360 ;
                RECT 2.880 217.400 59.280 217.720 ;
                RECT 69.160 217.400 79.680 217.720 ;
                RECT 1078.960 217.400 1083.000 217.720 ;
                RECT 2.880 218.760 79.680 219.080 ;
                RECT 1078.960 218.760 1083.000 219.080 ;
                RECT 2.880 220.120 59.280 220.440 ;
                RECT 69.160 220.120 79.680 220.440 ;
                RECT 1078.960 220.120 1083.000 220.440 ;
                RECT 2.880 221.480 59.280 221.800 ;
                RECT 69.160 221.480 79.680 221.800 ;
                RECT 1078.960 221.480 1083.000 221.800 ;
                RECT 2.880 222.840 59.280 223.160 ;
                RECT 69.160 222.840 79.680 223.160 ;
                RECT 1078.960 222.840 1083.000 223.160 ;
                RECT 2.880 224.200 59.280 224.520 ;
                RECT 69.160 224.200 79.680 224.520 ;
                RECT 1078.960 224.200 1083.000 224.520 ;
                RECT 2.880 225.560 59.280 225.880 ;
                RECT 63.040 225.560 79.680 225.880 ;
                RECT 1078.960 225.560 1083.000 225.880 ;
                RECT 2.880 226.920 65.400 227.240 ;
                RECT 69.160 226.920 79.680 227.240 ;
                RECT 1078.960 226.920 1083.000 227.240 ;
                RECT 2.880 228.280 59.280 228.600 ;
                RECT 69.160 228.280 79.680 228.600 ;
                RECT 1078.960 228.280 1083.000 228.600 ;
                RECT 2.880 229.640 59.280 229.960 ;
                RECT 69.160 229.640 79.680 229.960 ;
                RECT 1078.960 229.640 1083.000 229.960 ;
                RECT 2.880 231.000 59.280 231.320 ;
                RECT 69.160 231.000 79.680 231.320 ;
                RECT 1078.960 231.000 1083.000 231.320 ;
                RECT 2.880 232.360 59.280 232.680 ;
                RECT 69.160 232.360 79.680 232.680 ;
                RECT 1078.960 232.360 1083.000 232.680 ;
                RECT 2.880 233.720 59.280 234.040 ;
                RECT 63.720 233.720 79.680 234.040 ;
                RECT 1078.960 233.720 1083.000 234.040 ;
                RECT 2.880 235.080 64.040 235.400 ;
                RECT 69.160 235.080 79.680 235.400 ;
                RECT 1078.960 235.080 1083.000 235.400 ;
                RECT 2.880 236.440 59.280 236.760 ;
                RECT 69.160 236.440 79.680 236.760 ;
                RECT 1078.960 236.440 1083.000 236.760 ;
                RECT 2.880 237.800 59.280 238.120 ;
                RECT 69.160 237.800 79.680 238.120 ;
                RECT 1078.960 237.800 1083.000 238.120 ;
                RECT 2.880 239.160 59.280 239.480 ;
                RECT 69.160 239.160 79.680 239.480 ;
                RECT 1078.960 239.160 1083.000 239.480 ;
                RECT 2.880 240.520 59.280 240.840 ;
                RECT 69.160 240.520 79.680 240.840 ;
                RECT 1078.960 240.520 1083.000 240.840 ;
                RECT 2.880 241.880 79.680 242.200 ;
                RECT 1078.960 241.880 1083.000 242.200 ;
                RECT 2.880 243.240 62.000 243.560 ;
                RECT 69.160 243.240 79.680 243.560 ;
                RECT 1078.960 243.240 1083.000 243.560 ;
                RECT 2.880 244.600 66.080 244.920 ;
                RECT 69.160 244.600 79.680 244.920 ;
                RECT 1078.960 244.600 1083.000 244.920 ;
                RECT 2.880 245.960 62.000 246.280 ;
                RECT 69.160 245.960 79.680 246.280 ;
                RECT 1078.960 245.960 1083.000 246.280 ;
                RECT 2.880 247.320 62.000 247.640 ;
                RECT 69.160 247.320 79.680 247.640 ;
                RECT 1078.960 247.320 1083.000 247.640 ;
                RECT 2.880 248.680 62.000 249.000 ;
                RECT 69.160 248.680 79.680 249.000 ;
                RECT 1078.960 248.680 1083.000 249.000 ;
                RECT 2.880 250.040 79.680 250.360 ;
                RECT 1078.960 250.040 1083.000 250.360 ;
                RECT 2.880 251.400 62.000 251.720 ;
                RECT 69.160 251.400 79.680 251.720 ;
                RECT 1078.960 251.400 1083.000 251.720 ;
                RECT 2.880 252.760 62.000 253.080 ;
                RECT 69.160 252.760 79.680 253.080 ;
                RECT 1078.960 252.760 1083.000 253.080 ;
                RECT 2.880 254.120 64.720 254.440 ;
                RECT 69.160 254.120 79.680 254.440 ;
                RECT 1078.960 254.120 1083.000 254.440 ;
                RECT 2.880 255.480 65.400 255.800 ;
                RECT 69.160 255.480 79.680 255.800 ;
                RECT 1078.960 255.480 1083.000 255.800 ;
                RECT 2.880 256.840 62.000 257.160 ;
                RECT 69.160 256.840 79.680 257.160 ;
                RECT 1078.960 256.840 1083.000 257.160 ;
                RECT 2.880 258.200 79.680 258.520 ;
                RECT 1078.960 258.200 1083.000 258.520 ;
                RECT 2.880 259.560 62.000 259.880 ;
                RECT 69.160 259.560 79.680 259.880 ;
                RECT 1078.960 259.560 1083.000 259.880 ;
                RECT 2.880 260.920 62.000 261.240 ;
                RECT 69.160 260.920 79.680 261.240 ;
                RECT 1078.960 260.920 1083.000 261.240 ;
                RECT 2.880 262.280 62.000 262.600 ;
                RECT 69.160 262.280 79.680 262.600 ;
                RECT 1078.960 262.280 1083.000 262.600 ;
                RECT 2.880 263.640 62.000 263.960 ;
                RECT 69.160 263.640 79.680 263.960 ;
                RECT 1078.960 263.640 1083.000 263.960 ;
                RECT 2.880 265.000 79.680 265.320 ;
                RECT 1078.960 265.000 1083.000 265.320 ;
                RECT 2.880 266.360 64.040 266.680 ;
                RECT 69.160 266.360 79.680 266.680 ;
                RECT 1078.960 266.360 1083.000 266.680 ;
                RECT 2.880 267.720 62.680 268.040 ;
                RECT 69.160 267.720 79.680 268.040 ;
                RECT 1078.960 267.720 1083.000 268.040 ;
                RECT 2.880 269.080 62.680 269.400 ;
                RECT 69.160 269.080 79.680 269.400 ;
                RECT 1078.960 269.080 1083.000 269.400 ;
                RECT 2.880 270.440 62.680 270.760 ;
                RECT 69.160 270.440 79.680 270.760 ;
                RECT 1078.960 270.440 1083.000 270.760 ;
                RECT 2.880 271.800 62.680 272.120 ;
                RECT 69.160 271.800 79.680 272.120 ;
                RECT 1078.960 271.800 1083.000 272.120 ;
                RECT 2.880 273.160 79.680 273.480 ;
                RECT 1078.960 273.160 1083.000 273.480 ;
                RECT 2.880 274.520 65.400 274.840 ;
                RECT 69.160 274.520 79.680 274.840 ;
                RECT 1078.960 274.520 1083.000 274.840 ;
                RECT 2.880 275.880 62.680 276.200 ;
                RECT 69.160 275.880 79.680 276.200 ;
                RECT 1078.960 275.880 1083.000 276.200 ;
                RECT 2.880 277.240 62.680 277.560 ;
                RECT 69.160 277.240 79.680 277.560 ;
                RECT 1078.960 277.240 1083.000 277.560 ;
                RECT 2.880 278.600 62.680 278.920 ;
                RECT 69.160 278.600 79.680 278.920 ;
                RECT 1078.960 278.600 1083.000 278.920 ;
                RECT 2.880 279.960 62.680 280.280 ;
                RECT 69.160 279.960 79.680 280.280 ;
                RECT 1078.960 279.960 1083.000 280.280 ;
                RECT 2.880 281.320 79.680 281.640 ;
                RECT 1078.960 281.320 1083.000 281.640 ;
                RECT 2.880 282.680 63.360 283.000 ;
                RECT 69.160 282.680 79.680 283.000 ;
                RECT 1078.960 282.680 1083.000 283.000 ;
                RECT 2.880 284.040 64.040 284.360 ;
                RECT 69.160 284.040 79.680 284.360 ;
                RECT 1078.960 284.040 1083.000 284.360 ;
                RECT 2.880 285.400 63.360 285.720 ;
                RECT 69.160 285.400 79.680 285.720 ;
                RECT 1078.960 285.400 1083.000 285.720 ;
                RECT 2.880 286.760 63.360 287.080 ;
                RECT 69.160 286.760 79.680 287.080 ;
                RECT 1078.960 286.760 1083.000 287.080 ;
                RECT 2.880 288.120 63.360 288.440 ;
                RECT 69.160 288.120 79.680 288.440 ;
                RECT 1078.960 288.120 1083.000 288.440 ;
                RECT 2.880 289.480 79.680 289.800 ;
                RECT 1078.960 289.480 1083.000 289.800 ;
                RECT 2.880 290.840 63.360 291.160 ;
                RECT 69.160 290.840 79.680 291.160 ;
                RECT 1078.960 290.840 1083.000 291.160 ;
                RECT 2.880 292.200 63.360 292.520 ;
                RECT 69.160 292.200 79.680 292.520 ;
                RECT 1078.960 292.200 1083.000 292.520 ;
                RECT 2.880 293.560 66.760 293.880 ;
                RECT 69.160 293.560 79.680 293.880 ;
                RECT 1078.960 293.560 1083.000 293.880 ;
                RECT 2.880 294.920 63.360 295.240 ;
                RECT 69.160 294.920 79.680 295.240 ;
                RECT 1078.960 294.920 1083.000 295.240 ;
                RECT 2.880 296.280 63.360 296.600 ;
                RECT 69.160 296.280 79.680 296.600 ;
                RECT 1078.960 296.280 1083.000 296.600 ;
                RECT 2.880 297.640 79.680 297.960 ;
                RECT 1078.960 297.640 1083.000 297.960 ;
                RECT 2.880 299.000 278.240 299.320 ;
                RECT 1078.960 299.000 1083.000 299.320 ;
                RECT 2.880 300.360 278.240 300.680 ;
                RECT 1078.960 300.360 1083.000 300.680 ;
                RECT 2.880 301.720 278.240 302.040 ;
                RECT 1078.960 301.720 1083.000 302.040 ;
                RECT 2.880 303.080 1083.000 303.400 ;
                RECT 2.880 304.440 1083.000 304.760 ;
                RECT 2.880 305.800 1083.000 306.120 ;
                RECT 2.880 307.160 1083.000 307.480 ;
                RECT 2.880 2.880 1083.000 4.240 ;
                RECT 2.880 309.160 1083.000 310.520 ;
                RECT 282.380 43.250 288.180 44.370 ;
                RECT 1068.680 43.250 1074.480 44.370 ;
                RECT 282.380 49.115 288.180 49.885 ;
                RECT 1068.680 49.115 1074.480 49.885 ;
                RECT 282.380 55.150 288.180 55.850 ;
                RECT 1068.680 55.150 1074.480 55.850 ;
                RECT 282.380 60.740 288.180 61.440 ;
                RECT 1068.680 60.740 1074.480 61.440 ;
                RECT 282.380 116.315 1074.480 116.605 ;
                RECT 282.380 137.820 1074.480 139.225 ;
                RECT 282.380 95.210 1074.480 97.300 ;
                RECT 282.380 84.070 1074.480 84.870 ;
                RECT 282.380 91.970 1074.480 92.770 ;
                RECT 282.380 87.080 1074.480 87.880 ;
                RECT 282.380 88.760 1074.480 89.560 ;
                RECT 282.380 75.020 1074.480 76.820 ;
                RECT 282.380 33.880 1074.480 35.680 ;
                RECT 80.650 170.195 82.400 298.175 ;
                RECT 94.635 170.195 96.555 298.175 ;
                RECT 119.055 170.195 120.975 298.175 ;
                RECT 122.895 170.195 124.815 298.175 ;
                RECT 126.735 170.195 128.655 298.175 ;
                RECT 169.320 170.195 171.240 298.175 ;
                RECT 173.160 170.195 175.080 298.175 ;
                RECT 177.000 170.195 178.920 298.175 ;
                RECT 180.840 170.195 182.760 298.175 ;
                RECT 184.680 170.195 186.600 298.175 ;
                RECT 188.520 170.195 190.440 298.175 ;
                RECT 192.360 170.195 194.280 298.175 ;
                RECT 196.200 170.195 198.120 298.175 ;
                RECT 154.775 60.640 155.885 104.640 ;
                RECT 162.290 60.640 163.180 104.640 ;
                RECT 169.265 60.640 170.585 104.640 ;
                RECT 180.670 60.640 182.590 104.640 ;
                RECT 202.310 60.640 204.230 104.640 ;
                RECT 206.150 60.640 208.070 104.640 ;
                RECT 209.990 60.640 211.910 104.640 ;
                RECT 213.830 60.640 215.750 104.640 ;
                RECT 188.725 134.860 189.835 163.560 ;
                RECT 197.100 134.860 197.990 163.560 ;
                RECT 203.860 134.860 204.750 163.560 ;
                RECT 210.620 134.860 212.370 163.560 ;
                RECT 224.620 134.860 226.540 163.560 ;
                RECT 228.460 134.860 230.380 163.560 ;
                RECT 189.585 110.640 190.695 128.860 ;
                RECT 197.530 110.640 198.420 128.860 ;
                RECT 204.290 110.640 205.180 128.860 ;
                RECT 211.180 110.640 213.100 128.860 ;
                RECT 226.125 110.640 228.045 128.860 ;
                RECT 229.965 110.640 231.885 128.860 ;
                RECT 226.220 49.480 227.110 54.640 ;
                RECT 233.515 49.480 234.625 54.640 ;
                RECT 242.450 49.480 244.370 54.640 ;
                RECT 24.860 171.260 34.020 171.630 ;
                RECT 24.860 174.595 34.020 175.485 ;
                RECT 78.840 157.620 96.080 158.290 ;
                RECT 78.840 158.920 96.080 159.930 ;
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 1085.880 313.400 ;
        LAYER met2 ;
            RECT 0.000 0.000 1085.880 313.400 ;
    END 
END sram22_256x128m4w8 
END LIBRARY 

