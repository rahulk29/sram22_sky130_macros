VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_128x32m4w8
    CLASS BLOCK  ;
    FOREIGN sram22_128x32m4w8   ;
    SIZE 416.760 BY 224.320 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 208.510 0.000 208.650 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 214.610 0.000 214.750 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 220.710 0.000 220.850 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 226.810 0.000 226.950 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 232.910 0.000 233.050 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 239.010 0.000 239.150 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 245.110 0.000 245.250 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 251.210 0.000 251.350 0.140 ; 
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 257.310 0.000 257.450 0.140 ; 
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 263.410 0.000 263.550 0.140 ; 
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 269.510 0.000 269.650 0.140 ; 
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 275.610 0.000 275.750 0.140 ; 
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 281.710 0.000 281.850 0.140 ; 
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 287.810 0.000 287.950 0.140 ; 
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 293.910 0.000 294.050 0.140 ; 
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 300.010 0.000 300.150 0.140 ; 
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 306.110 0.000 306.250 0.140 ; 
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 312.210 0.000 312.350 0.140 ; 
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 318.310 0.000 318.450 0.140 ; 
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 324.410 0.000 324.550 0.140 ; 
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 330.510 0.000 330.650 0.140 ; 
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 336.610 0.000 336.750 0.140 ; 
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 342.710 0.000 342.850 0.140 ; 
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 348.810 0.000 348.950 0.140 ; 
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 354.910 0.000 355.050 0.140 ; 
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 361.010 0.000 361.150 0.140 ; 
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 367.110 0.000 367.250 0.140 ; 
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 373.210 0.000 373.350 0.140 ; 
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 379.310 0.000 379.450 0.140 ; 
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 385.410 0.000 385.550 0.140 ; 
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 391.510 0.000 391.650 0.140 ; 
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.335400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 397.610 0.000 397.750 0.140 ; 
        END 
    END dout[31] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 208.090 0.000 208.230 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 214.190 0.000 214.330 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 220.290 0.000 220.430 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 226.390 0.000 226.530 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 232.490 0.000 232.630 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 238.590 0.000 238.730 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 244.690 0.000 244.830 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 250.790 0.000 250.930 0.140 ; 
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 256.890 0.000 257.030 0.140 ; 
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 262.990 0.000 263.130 0.140 ; 
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 269.090 0.000 269.230 0.140 ; 
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 275.190 0.000 275.330 0.140 ; 
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 281.290 0.000 281.430 0.140 ; 
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 287.390 0.000 287.530 0.140 ; 
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 293.490 0.000 293.630 0.140 ; 
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 299.590 0.000 299.730 0.140 ; 
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 305.690 0.000 305.830 0.140 ; 
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 311.790 0.000 311.930 0.140 ; 
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 317.890 0.000 318.030 0.140 ; 
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 323.990 0.000 324.130 0.140 ; 
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 330.090 0.000 330.230 0.140 ; 
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 336.190 0.000 336.330 0.140 ; 
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 342.290 0.000 342.430 0.140 ; 
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 348.390 0.000 348.530 0.140 ; 
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 354.490 0.000 354.630 0.140 ; 
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 360.590 0.000 360.730 0.140 ; 
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 366.690 0.000 366.830 0.140 ; 
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 372.790 0.000 372.930 0.140 ; 
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 378.890 0.000 379.030 0.140 ; 
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 384.990 0.000 385.130 0.140 ; 
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 391.090 0.000 391.230 0.140 ; 
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.020800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.057000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 397.190 0.000 397.330 0.140 ; 
        END 
    END din[31] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.831200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 207.740 0.000 207.880 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.831200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 256.540 0.000 256.680 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.831200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 305.340 0.000 305.480 0.140 ; 
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 2.831200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 354.140 0.000 354.280 0.140 ; 
        END 
    END wmask[3] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 166.400 0.000 166.720 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 160.280 0.000 160.600 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 154.160 0.000 154.480 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 148.040 0.000 148.360 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 141.920 0.000 142.240 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 135.800 0.000 136.120 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 129.680 0.000 130.000 0.320 ; 
        END 
    END addr[6] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 178.640 0.000 178.960 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.867900 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 172.520 0.000 172.840 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 22.041000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 181.360 0.000 181.680 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 25.947000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 182.040 0.000 182.360 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 207.520 6.240 ; 
                RECT 209.240 5.920 213.640 6.240 ; 
                RECT 215.360 5.920 219.760 6.240 ; 
                RECT 221.480 5.920 225.880 6.240 ; 
                RECT 227.600 5.920 232.000 6.240 ; 
                RECT 233.720 5.920 238.120 6.240 ; 
                RECT 239.840 5.920 244.240 6.240 ; 
                RECT 245.960 5.920 250.360 6.240 ; 
                RECT 252.080 5.920 256.480 6.240 ; 
                RECT 258.200 5.920 262.600 6.240 ; 
                RECT 264.320 5.920 268.720 6.240 ; 
                RECT 270.440 5.920 274.840 6.240 ; 
                RECT 276.560 5.920 280.960 6.240 ; 
                RECT 282.680 5.920 287.080 6.240 ; 
                RECT 288.800 5.920 293.200 6.240 ; 
                RECT 294.920 5.920 299.320 6.240 ; 
                RECT 301.040 5.920 305.440 6.240 ; 
                RECT 307.160 5.920 311.560 6.240 ; 
                RECT 313.280 5.920 317.680 6.240 ; 
                RECT 319.400 5.920 323.800 6.240 ; 
                RECT 325.520 5.920 329.920 6.240 ; 
                RECT 331.640 5.920 336.040 6.240 ; 
                RECT 337.760 5.920 342.160 6.240 ; 
                RECT 343.880 5.920 348.280 6.240 ; 
                RECT 349.320 5.920 354.400 6.240 ; 
                RECT 355.440 5.920 360.520 6.240 ; 
                RECT 361.560 5.920 366.640 6.240 ; 
                RECT 367.680 5.920 372.760 6.240 ; 
                RECT 373.800 5.920 378.880 6.240 ; 
                RECT 379.920 5.920 385.000 6.240 ; 
                RECT 386.040 5.920 391.120 6.240 ; 
                RECT 392.160 5.920 397.240 6.240 ; 
                RECT 398.280 5.920 416.600 6.240 ; 
                RECT 0.160 7.280 416.600 7.600 ; 
                RECT 0.160 8.640 416.600 8.960 ; 
                RECT 0.160 10.000 181.000 10.320 ; 
                RECT 203.800 10.000 416.600 10.320 ; 
                RECT 0.160 11.360 416.600 11.680 ; 
                RECT 0.160 12.720 416.600 13.040 ; 
                RECT 0.160 14.080 125.920 14.400 ; 
                RECT 182.720 14.080 416.600 14.400 ; 
                RECT 0.160 15.440 416.600 15.760 ; 
                RECT 0.160 16.800 416.600 17.120 ; 
                RECT 0.160 18.160 125.920 18.480 ; 
                RECT 182.040 18.160 206.840 18.480 ; 
                RECT 354.760 18.160 416.600 18.480 ; 
                RECT 0.160 19.520 197.320 19.840 ; 
                RECT 407.120 19.520 416.600 19.840 ; 
                RECT 0.160 20.880 197.320 21.200 ; 
                RECT 407.120 20.880 416.600 21.200 ; 
                RECT 0.160 22.240 197.320 22.560 ; 
                RECT 407.120 22.240 416.600 22.560 ; 
                RECT 0.160 23.600 197.320 23.920 ; 
                RECT 407.120 23.600 416.600 23.920 ; 
                RECT 0.160 24.960 197.320 25.280 ; 
                RECT 407.120 24.960 416.600 25.280 ; 
                RECT 0.160 26.320 197.320 26.640 ; 
                RECT 407.120 26.320 416.600 26.640 ; 
                RECT 0.160 27.680 197.320 28.000 ; 
                RECT 407.120 27.680 416.600 28.000 ; 
                RECT 0.160 29.040 197.320 29.360 ; 
                RECT 407.120 29.040 416.600 29.360 ; 
                RECT 0.160 30.400 197.320 30.720 ; 
                RECT 407.120 30.400 416.600 30.720 ; 
                RECT 0.160 31.760 197.320 32.080 ; 
                RECT 407.120 31.760 416.600 32.080 ; 
                RECT 0.160 33.120 142.920 33.440 ; 
                RECT 159.600 33.120 197.320 33.440 ; 
                RECT 407.120 33.120 416.600 33.440 ; 
                RECT 0.160 34.480 141.560 34.800 ; 
                RECT 165.720 34.480 197.320 34.800 ; 
                RECT 407.120 34.480 416.600 34.800 ; 
                RECT 0.160 35.840 121.840 36.160 ; 
                RECT 182.720 35.840 197.320 36.160 ; 
                RECT 407.120 35.840 416.600 36.160 ; 
                RECT 0.160 37.200 121.160 37.520 ; 
                RECT 178.640 37.200 196.640 37.520 ; 
                RECT 407.120 37.200 416.600 37.520 ; 
                RECT 0.160 38.560 197.320 38.880 ; 
                RECT 407.120 38.560 416.600 38.880 ; 
                RECT 0.160 39.920 197.320 40.240 ; 
                RECT 407.120 39.920 416.600 40.240 ; 
                RECT 0.160 41.280 197.320 41.600 ; 
                RECT 407.120 41.280 416.600 41.600 ; 
                RECT 0.160 42.640 197.320 42.960 ; 
                RECT 407.120 42.640 416.600 42.960 ; 
                RECT 0.160 44.000 117.080 44.320 ; 
                RECT 128.320 44.000 197.320 44.320 ; 
                RECT 407.120 44.000 416.600 44.320 ; 
                RECT 0.160 45.360 118.440 45.680 ; 
                RECT 124.240 45.360 132.040 45.680 ; 
                RECT 134.440 45.360 197.320 45.680 ; 
                RECT 407.120 45.360 416.600 45.680 ; 
                RECT 0.160 46.720 119.800 47.040 ; 
                RECT 123.560 46.720 197.320 47.040 ; 
                RECT 407.120 46.720 416.600 47.040 ; 
                RECT 0.160 48.080 197.320 48.400 ; 
                RECT 407.120 48.080 416.600 48.400 ; 
                RECT 0.160 49.440 126.600 49.760 ; 
                RECT 135.120 49.440 197.320 49.760 ; 
                RECT 407.120 49.440 416.600 49.760 ; 
                RECT 0.160 50.800 119.120 51.120 ; 
                RECT 128.320 50.800 197.320 51.120 ; 
                RECT 407.120 50.800 416.600 51.120 ; 
                RECT 0.160 52.160 122.520 52.480 ; 
                RECT 127.640 52.160 197.320 52.480 ; 
                RECT 407.120 52.160 416.600 52.480 ; 
                RECT 0.160 53.520 197.320 53.840 ; 
                RECT 407.120 53.520 416.600 53.840 ; 
                RECT 0.160 54.880 118.440 55.200 ; 
                RECT 128.320 54.880 173.520 55.200 ; 
                RECT 180.000 54.880 197.320 55.200 ; 
                RECT 407.120 54.880 416.600 55.200 ; 
                RECT 0.160 56.240 125.240 56.560 ; 
                RECT 133.760 56.240 173.520 56.560 ; 
                RECT 180.000 56.240 197.320 56.560 ; 
                RECT 407.120 56.240 416.600 56.560 ; 
                RECT 0.160 57.600 173.520 57.920 ; 
                RECT 407.120 57.600 416.600 57.920 ; 
                RECT 0.160 58.960 126.600 59.280 ; 
                RECT 132.400 58.960 173.520 59.280 ; 
                RECT 180.000 58.960 197.320 59.280 ; 
                RECT 407.120 58.960 416.600 59.280 ; 
                RECT 0.160 60.320 129.320 60.640 ; 
                RECT 134.440 60.320 197.320 60.640 ; 
                RECT 407.120 60.320 416.600 60.640 ; 
                RECT 0.160 61.680 123.200 62.000 ; 
                RECT 128.320 61.680 197.320 62.000 ; 
                RECT 407.120 61.680 416.600 62.000 ; 
                RECT 0.160 63.040 197.320 63.360 ; 
                RECT 407.120 63.040 416.600 63.360 ; 
                RECT 0.160 64.400 116.400 64.720 ; 
                RECT 180.000 64.400 197.320 64.720 ; 
                RECT 407.120 64.400 416.600 64.720 ; 
                RECT 0.160 65.760 126.600 66.080 ; 
                RECT 134.440 65.760 142.240 66.080 ; 
                RECT 146.680 65.760 152.440 66.080 ; 
                RECT 180.000 65.760 197.320 66.080 ; 
                RECT 407.120 65.760 416.600 66.080 ; 
                RECT 0.160 67.120 125.240 67.440 ; 
                RECT 128.320 67.120 135.440 67.440 ; 
                RECT 141.920 67.120 143.600 67.440 ; 
                RECT 146.000 67.120 152.440 67.440 ; 
                RECT 189.520 67.120 197.320 67.440 ; 
                RECT 407.120 67.120 416.600 67.440 ; 
                RECT 0.160 68.480 117.080 68.800 ; 
                RECT 131.040 68.480 152.440 68.800 ; 
                RECT 189.520 68.480 197.320 68.800 ; 
                RECT 407.120 68.480 416.600 68.800 ; 
                RECT 0.160 69.840 125.920 70.160 ; 
                RECT 134.440 69.840 152.440 70.160 ; 
                RECT 188.160 69.840 197.320 70.160 ; 
                RECT 407.120 69.840 416.600 70.160 ; 
                RECT 0.160 71.200 123.880 71.520 ; 
                RECT 127.640 71.200 152.440 71.520 ; 
                RECT 189.520 71.200 197.320 71.520 ; 
                RECT 407.120 71.200 416.600 71.520 ; 
                RECT 0.160 72.560 119.120 72.880 ; 
                RECT 123.560 72.560 126.600 72.880 ; 
                RECT 135.120 72.560 152.440 72.880 ; 
                RECT 192.240 72.560 197.320 72.880 ; 
                RECT 407.120 72.560 416.600 72.880 ; 
                RECT 0.160 73.920 121.840 74.240 ; 
                RECT 125.600 73.920 152.440 74.240 ; 
                RECT 180.000 73.920 197.320 74.240 ; 
                RECT 407.120 73.920 416.600 74.240 ; 
                RECT 0.160 75.280 118.440 75.600 ; 
                RECT 122.200 75.280 152.440 75.600 ; 
                RECT 192.240 75.280 197.320 75.600 ; 
                RECT 407.120 75.280 416.600 75.600 ; 
                RECT 0.160 76.640 122.520 76.960 ; 
                RECT 128.320 76.640 152.440 76.960 ; 
                RECT 190.880 76.640 197.320 76.960 ; 
                RECT 407.120 76.640 416.600 76.960 ; 
                RECT 0.160 78.000 118.440 78.320 ; 
                RECT 133.760 78.000 152.440 78.320 ; 
                RECT 192.240 78.000 197.320 78.320 ; 
                RECT 407.120 78.000 416.600 78.320 ; 
                RECT 0.160 79.360 152.440 79.680 ; 
                RECT 194.960 79.360 197.320 79.680 ; 
                RECT 407.120 79.360 416.600 79.680 ; 
                RECT 0.160 80.720 125.240 81.040 ; 
                RECT 127.640 80.720 152.440 81.040 ; 
                RECT 194.960 80.720 197.320 81.040 ; 
                RECT 407.120 80.720 416.600 81.040 ; 
                RECT 0.160 82.080 126.600 82.400 ; 
                RECT 128.320 82.080 152.440 82.400 ; 
                RECT 193.600 82.080 197.320 82.400 ; 
                RECT 407.120 82.080 416.600 82.400 ; 
                RECT 0.160 83.440 117.080 83.760 ; 
                RECT 127.640 83.440 152.440 83.760 ; 
                RECT 180.000 83.440 197.320 83.760 ; 
                RECT 407.120 83.440 416.600 83.760 ; 
                RECT 0.160 84.800 122.520 85.120 ; 
                RECT 134.440 84.800 152.440 85.120 ; 
                RECT 193.600 84.800 197.320 85.120 ; 
                RECT 407.120 84.800 416.600 85.120 ; 
                RECT 0.160 86.160 117.080 86.480 ; 
                RECT 128.320 86.160 152.440 86.480 ; 
                RECT 407.120 86.160 416.600 86.480 ; 
                RECT 0.160 87.520 125.920 87.840 ; 
                RECT 128.320 87.520 152.440 87.840 ; 
                RECT 407.120 87.520 416.600 87.840 ; 
                RECT 0.160 88.880 152.440 89.200 ; 
                RECT 407.120 88.880 416.600 89.200 ; 
                RECT 0.160 90.240 152.440 90.560 ; 
                RECT 407.120 90.240 416.600 90.560 ; 
                RECT 0.160 91.600 113.680 91.920 ; 
                RECT 131.040 91.600 152.440 91.920 ; 
                RECT 180.000 91.600 197.320 91.920 ; 
                RECT 407.120 91.600 416.600 91.920 ; 
                RECT 0.160 92.960 197.320 93.280 ; 
                RECT 407.120 92.960 416.600 93.280 ; 
                RECT 0.160 94.320 197.320 94.640 ; 
                RECT 407.120 94.320 416.600 94.640 ; 
                RECT 0.160 95.680 122.520 96.000 ; 
                RECT 134.440 95.680 197.320 96.000 ; 
                RECT 407.120 95.680 416.600 96.000 ; 
                RECT 0.160 97.040 129.320 97.360 ; 
                RECT 137.160 97.040 197.320 97.360 ; 
                RECT 407.120 97.040 416.600 97.360 ; 
                RECT 0.160 98.400 140.880 98.720 ; 
                RECT 154.160 98.400 157.200 98.720 ; 
                RECT 179.320 98.400 197.320 98.720 ; 
                RECT 407.120 98.400 416.600 98.720 ; 
                RECT 0.160 99.760 157.200 100.080 ; 
                RECT 179.320 99.760 197.320 100.080 ; 
                RECT 407.120 99.760 416.600 100.080 ; 
                RECT 0.160 101.120 116.400 101.440 ; 
                RECT 122.200 101.120 157.200 101.440 ; 
                RECT 179.320 101.120 197.320 101.440 ; 
                RECT 407.120 101.120 416.600 101.440 ; 
                RECT 0.160 102.480 157.200 102.800 ; 
                RECT 179.320 102.480 197.320 102.800 ; 
                RECT 407.120 102.480 416.600 102.800 ; 
                RECT 0.160 103.840 157.200 104.160 ; 
                RECT 179.320 103.840 197.320 104.160 ; 
                RECT 407.120 103.840 416.600 104.160 ; 
                RECT 0.160 105.200 132.040 105.520 ; 
                RECT 135.120 105.200 157.200 105.520 ; 
                RECT 179.320 105.200 197.320 105.520 ; 
                RECT 407.120 105.200 416.600 105.520 ; 
                RECT 0.160 106.560 157.200 106.880 ; 
                RECT 179.320 106.560 197.320 106.880 ; 
                RECT 407.120 106.560 416.600 106.880 ; 
                RECT 0.160 107.920 157.200 108.240 ; 
                RECT 179.320 107.920 197.320 108.240 ; 
                RECT 407.120 107.920 416.600 108.240 ; 
                RECT 0.160 109.280 157.200 109.600 ; 
                RECT 407.120 109.280 416.600 109.600 ; 
                RECT 0.160 110.640 119.120 110.960 ; 
                RECT 124.240 110.640 157.200 110.960 ; 
                RECT 179.320 110.640 194.600 110.960 ; 
                RECT 407.120 110.640 416.600 110.960 ; 
                RECT 0.160 112.000 157.200 112.320 ; 
                RECT 179.320 112.000 191.880 112.320 ; 
                RECT 407.120 112.000 416.600 112.320 ; 
                RECT 0.160 113.360 95.320 113.680 ; 
                RECT 114.040 113.360 125.240 113.680 ; 
                RECT 133.760 113.360 157.200 113.680 ; 
                RECT 179.320 113.360 189.160 113.680 ; 
                RECT 407.120 113.360 416.600 113.680 ; 
                RECT 0.160 114.720 95.320 115.040 ; 
                RECT 114.040 114.720 186.440 115.040 ; 
                RECT 407.120 114.720 416.600 115.040 ; 
                RECT 0.160 116.080 95.320 116.400 ; 
                RECT 114.040 116.080 121.840 116.400 ; 
                RECT 124.240 116.080 197.320 116.400 ; 
                RECT 407.120 116.080 416.600 116.400 ; 
                RECT 0.160 117.440 95.320 117.760 ; 
                RECT 114.040 117.440 118.440 117.760 ; 
                RECT 121.520 117.440 197.320 117.760 ; 
                RECT 407.120 117.440 416.600 117.760 ; 
                RECT 0.160 118.800 95.320 119.120 ; 
                RECT 114.720 118.800 197.320 119.120 ; 
                RECT 407.120 118.800 416.600 119.120 ; 
                RECT 0.160 120.160 95.320 120.480 ; 
                RECT 114.040 120.160 157.200 120.480 ; 
                RECT 180.000 120.160 197.320 120.480 ; 
                RECT 407.120 120.160 416.600 120.480 ; 
                RECT 0.160 121.520 95.320 121.840 ; 
                RECT 114.040 121.520 157.200 121.840 ; 
                RECT 180.000 121.520 197.320 121.840 ; 
                RECT 407.120 121.520 416.600 121.840 ; 
                RECT 0.160 122.880 95.320 123.200 ; 
                RECT 114.040 122.880 157.200 123.200 ; 
                RECT 180.000 122.880 197.320 123.200 ; 
                RECT 407.120 122.880 416.600 123.200 ; 
                RECT 0.160 124.240 95.320 124.560 ; 
                RECT 114.040 124.240 157.200 124.560 ; 
                RECT 180.000 124.240 187.800 124.560 ; 
                RECT 407.120 124.240 416.600 124.560 ; 
                RECT 0.160 125.600 95.320 125.920 ; 
                RECT 114.040 125.600 157.200 125.920 ; 
                RECT 180.000 125.600 190.520 125.920 ; 
                RECT 407.120 125.600 416.600 125.920 ; 
                RECT 0.160 126.960 95.320 127.280 ; 
                RECT 114.040 126.960 120.480 127.280 ; 
                RECT 124.240 126.960 157.200 127.280 ; 
                RECT 180.000 126.960 193.240 127.280 ; 
                RECT 407.120 126.960 416.600 127.280 ; 
                RECT 0.160 128.320 157.200 128.640 ; 
                RECT 180.000 128.320 195.960 128.640 ; 
                RECT 407.120 128.320 416.600 128.640 ; 
                RECT 0.160 129.680 157.200 130.000 ; 
                RECT 407.120 129.680 416.600 130.000 ; 
                RECT 0.160 131.040 79.000 131.360 ; 
                RECT 95.680 131.040 122.520 131.360 ; 
                RECT 128.320 131.040 157.200 131.360 ; 
                RECT 180.000 131.040 197.320 131.360 ; 
                RECT 407.120 131.040 416.600 131.360 ; 
                RECT 0.160 132.400 79.000 132.720 ; 
                RECT 95.680 132.400 101.440 132.720 ; 
                RECT 108.600 132.400 157.200 132.720 ; 
                RECT 180.000 132.400 197.320 132.720 ; 
                RECT 407.120 132.400 416.600 132.720 ; 
                RECT 0.160 133.760 79.000 134.080 ; 
                RECT 113.360 133.760 157.200 134.080 ; 
                RECT 180.000 133.760 197.320 134.080 ; 
                RECT 407.120 133.760 416.600 134.080 ; 
                RECT 0.160 135.120 79.000 135.440 ; 
                RECT 113.360 135.120 157.200 135.440 ; 
                RECT 407.120 135.120 416.600 135.440 ; 
                RECT 0.160 136.480 79.000 136.800 ; 
                RECT 95.680 136.480 101.440 136.800 ; 
                RECT 108.600 136.480 117.080 136.800 ; 
                RECT 126.960 136.480 157.200 136.800 ; 
                RECT 407.120 136.480 416.600 136.800 ; 
                RECT 0.160 137.840 79.680 138.160 ; 
                RECT 107.920 137.840 157.200 138.160 ; 
                RECT 180.000 137.840 416.600 138.160 ; 
                RECT 0.160 139.200 107.560 139.520 ; 
                RECT 154.840 139.200 416.600 139.520 ; 
                RECT 0.160 140.560 194.600 140.880 ; 
                RECT 409.160 140.560 416.600 140.880 ; 
                RECT 0.160 141.920 194.600 142.240 ; 
                RECT 409.160 141.920 416.600 142.240 ; 
                RECT 0.160 143.280 194.600 143.600 ; 
                RECT 409.160 143.280 416.600 143.600 ; 
                RECT 0.160 144.640 24.600 144.960 ; 
                RECT 31.080 144.640 33.440 144.960 ; 
                RECT 44.680 144.640 72.880 144.960 ; 
                RECT 409.160 144.640 416.600 144.960 ; 
                RECT 0.160 146.000 22.560 146.320 ; 
                RECT 33.120 146.000 34.800 146.320 ; 
                RECT 43.320 146.000 57.240 146.320 ; 
                RECT 63.040 146.000 72.880 146.320 ; 
                RECT 409.160 146.000 416.600 146.320 ; 
                RECT 0.160 147.360 22.560 147.680 ; 
                RECT 33.120 147.360 36.160 147.680 ; 
                RECT 42.640 147.360 55.200 147.680 ; 
                RECT 63.040 147.360 72.880 147.680 ; 
                RECT 409.160 147.360 416.600 147.680 ; 
                RECT 0.160 148.720 22.560 149.040 ; 
                RECT 33.120 148.720 55.200 149.040 ; 
                RECT 58.960 148.720 72.880 149.040 ; 
                RECT 409.160 148.720 416.600 149.040 ; 
                RECT 0.160 150.080 55.200 150.400 ; 
                RECT 63.040 150.080 72.880 150.400 ; 
                RECT 409.160 150.080 416.600 150.400 ; 
                RECT 0.160 151.440 22.560 151.760 ; 
                RECT 33.120 151.440 55.200 151.760 ; 
                RECT 63.040 151.440 72.880 151.760 ; 
                RECT 409.160 151.440 416.600 151.760 ; 
                RECT 0.160 152.800 22.560 153.120 ; 
                RECT 33.120 152.800 72.880 153.120 ; 
                RECT 409.160 152.800 416.600 153.120 ; 
                RECT 0.160 154.160 59.280 154.480 ; 
                RECT 63.040 154.160 72.880 154.480 ; 
                RECT 409.160 154.160 416.600 154.480 ; 
                RECT 0.160 155.520 55.200 155.840 ; 
                RECT 63.040 155.520 72.880 155.840 ; 
                RECT 409.160 155.520 416.600 155.840 ; 
                RECT 0.160 156.880 15.760 157.200 ; 
                RECT 18.160 156.880 55.200 157.200 ; 
                RECT 63.040 156.880 72.880 157.200 ; 
                RECT 409.160 156.880 416.600 157.200 ; 
                RECT 0.160 158.240 55.200 158.560 ; 
                RECT 56.920 158.240 72.880 158.560 ; 
                RECT 409.160 158.240 416.600 158.560 ; 
                RECT 0.160 159.600 15.080 159.920 ; 
                RECT 18.160 159.600 31.400 159.920 ; 
                RECT 35.160 159.600 55.200 159.920 ; 
                RECT 63.040 159.600 72.880 159.920 ; 
                RECT 409.160 159.600 416.600 159.920 ; 
                RECT 0.160 160.960 14.400 161.280 ; 
                RECT 18.160 160.960 31.400 161.280 ; 
                RECT 35.840 160.960 72.880 161.280 ; 
                RECT 409.160 160.960 416.600 161.280 ; 
                RECT 0.160 162.320 13.720 162.640 ; 
                RECT 18.160 162.320 31.400 162.640 ; 
                RECT 36.520 162.320 57.240 162.640 ; 
                RECT 63.040 162.320 72.880 162.640 ; 
                RECT 409.160 162.320 416.600 162.640 ; 
                RECT 0.160 163.680 55.200 164.000 ; 
                RECT 63.040 163.680 72.880 164.000 ; 
                RECT 409.160 163.680 416.600 164.000 ; 
                RECT 0.160 165.040 13.040 165.360 ; 
                RECT 18.160 165.040 31.400 165.360 ; 
                RECT 37.200 165.040 55.200 165.360 ; 
                RECT 63.040 165.040 72.880 165.360 ; 
                RECT 409.160 165.040 416.600 165.360 ; 
                RECT 0.160 166.400 12.360 166.720 ; 
                RECT 18.160 166.400 55.200 166.720 ; 
                RECT 63.040 166.400 72.880 166.720 ; 
                RECT 409.160 166.400 416.600 166.720 ; 
                RECT 0.160 167.760 11.680 168.080 ; 
                RECT 18.160 167.760 55.200 168.080 ; 
                RECT 61.680 167.760 72.880 168.080 ; 
                RECT 409.160 167.760 416.600 168.080 ; 
                RECT 0.160 169.120 11.000 169.440 ; 
                RECT 18.160 169.120 72.880 169.440 ; 
                RECT 409.160 169.120 416.600 169.440 ; 
                RECT 0.160 170.480 55.200 170.800 ; 
                RECT 63.040 170.480 72.880 170.800 ; 
                RECT 409.160 170.480 416.600 170.800 ; 
                RECT 0.160 171.840 10.320 172.160 ; 
                RECT 18.160 171.840 55.200 172.160 ; 
                RECT 63.040 171.840 72.880 172.160 ; 
                RECT 409.160 171.840 416.600 172.160 ; 
                RECT 0.160 173.200 9.640 173.520 ; 
                RECT 18.160 173.200 55.200 173.520 ; 
                RECT 63.040 173.200 72.880 173.520 ; 
                RECT 409.160 173.200 416.600 173.520 ; 
                RECT 0.160 174.560 55.200 174.880 ; 
                RECT 63.040 174.560 72.880 174.880 ; 
                RECT 409.160 174.560 416.600 174.880 ; 
                RECT 0.160 175.920 55.200 176.240 ; 
                RECT 62.360 175.920 72.880 176.240 ; 
                RECT 409.160 175.920 416.600 176.240 ; 
                RECT 0.160 177.280 57.240 177.600 ; 
                RECT 63.040 177.280 72.880 177.600 ; 
                RECT 409.160 177.280 416.600 177.600 ; 
                RECT 0.160 178.640 72.880 178.960 ; 
                RECT 409.160 178.640 416.600 178.960 ; 
                RECT 0.160 180.000 57.920 180.320 ; 
                RECT 63.040 180.000 72.880 180.320 ; 
                RECT 409.160 180.000 416.600 180.320 ; 
                RECT 0.160 181.360 58.600 181.680 ; 
                RECT 63.040 181.360 72.880 181.680 ; 
                RECT 409.160 181.360 416.600 181.680 ; 
                RECT 0.160 182.720 59.280 183.040 ; 
                RECT 63.040 182.720 72.880 183.040 ; 
                RECT 409.160 182.720 416.600 183.040 ; 
                RECT 0.160 184.080 35.480 184.400 ; 
                RECT 44.000 184.080 72.880 184.400 ; 
                RECT 409.160 184.080 416.600 184.400 ; 
                RECT 0.160 185.440 34.120 185.760 ; 
                RECT 42.640 185.440 55.200 185.760 ; 
                RECT 63.040 185.440 72.880 185.760 ; 
                RECT 409.160 185.440 416.600 185.760 ; 
                RECT 0.160 186.800 55.200 187.120 ; 
                RECT 63.040 186.800 72.880 187.120 ; 
                RECT 409.160 186.800 416.600 187.120 ; 
                RECT 0.160 188.160 55.200 188.480 ; 
                RECT 57.600 188.160 72.880 188.480 ; 
                RECT 409.160 188.160 416.600 188.480 ; 
                RECT 0.160 189.520 55.200 189.840 ; 
                RECT 63.040 189.520 72.880 189.840 ; 
                RECT 409.160 189.520 416.600 189.840 ; 
                RECT 0.160 190.880 55.200 191.200 ; 
                RECT 63.040 190.880 72.880 191.200 ; 
                RECT 409.160 190.880 416.600 191.200 ; 
                RECT 0.160 192.240 55.200 192.560 ; 
                RECT 58.960 192.240 72.880 192.560 ; 
                RECT 409.160 192.240 416.600 192.560 ; 
                RECT 0.160 193.600 57.240 193.920 ; 
                RECT 63.040 193.600 72.880 193.920 ; 
                RECT 409.160 193.600 416.600 193.920 ; 
                RECT 0.160 194.960 57.920 195.280 ; 
                RECT 63.040 194.960 72.880 195.280 ; 
                RECT 409.160 194.960 416.600 195.280 ; 
                RECT 0.160 196.320 58.600 196.640 ; 
                RECT 63.040 196.320 72.880 196.640 ; 
                RECT 409.160 196.320 416.600 196.640 ; 
                RECT 0.160 197.680 72.880 198.000 ; 
                RECT 409.160 197.680 416.600 198.000 ; 
                RECT 0.160 199.040 59.280 199.360 ; 
                RECT 63.040 199.040 72.880 199.360 ; 
                RECT 409.160 199.040 416.600 199.360 ; 
                RECT 0.160 200.400 72.880 200.720 ; 
                RECT 409.160 200.400 416.600 200.720 ; 
                RECT 0.160 201.760 59.280 202.080 ; 
                RECT 63.040 201.760 72.880 202.080 ; 
                RECT 409.160 201.760 416.600 202.080 ; 
                RECT 0.160 203.120 59.960 203.440 ; 
                RECT 63.040 203.120 72.880 203.440 ; 
                RECT 409.160 203.120 416.600 203.440 ; 
                RECT 0.160 204.480 60.640 204.800 ; 
                RECT 63.040 204.480 72.880 204.800 ; 
                RECT 409.160 204.480 416.600 204.800 ; 
                RECT 0.160 205.840 60.640 206.160 ; 
                RECT 63.040 205.840 72.880 206.160 ; 
                RECT 409.160 205.840 416.600 206.160 ; 
                RECT 0.160 207.200 72.880 207.520 ; 
                RECT 409.160 207.200 416.600 207.520 ; 
                RECT 0.160 208.560 72.880 208.880 ; 
                RECT 409.160 208.560 416.600 208.880 ; 
                RECT 0.160 209.920 194.600 210.240 ; 
                RECT 409.160 209.920 416.600 210.240 ; 
                RECT 0.160 211.280 194.600 211.600 ; 
                RECT 409.160 211.280 416.600 211.600 ; 
                RECT 0.160 212.640 194.600 212.960 ; 
                RECT 409.160 212.640 416.600 212.960 ; 
                RECT 0.160 214.000 416.600 214.320 ; 
                RECT 0.160 215.360 416.600 215.680 ; 
                RECT 0.160 216.720 416.600 217.040 ; 
                RECT 0.160 218.080 416.600 218.400 ; 
                RECT 0.160 0.160 416.600 1.520 ; 
                RECT 0.160 222.800 416.600 224.160 ; 
                RECT 198.740 40.720 204.540 42.090 ; 
                RECT 399.440 40.720 405.240 42.090 ; 
                RECT 198.740 45.835 204.540 47.255 ; 
                RECT 399.440 45.835 405.240 47.255 ; 
                RECT 198.740 51.155 204.540 52.675 ; 
                RECT 399.440 51.155 405.240 52.675 ; 
                RECT 198.740 56.625 204.540 58.145 ; 
                RECT 399.440 56.625 405.240 58.145 ; 
                RECT 198.740 95.005 405.240 95.295 ; 
                RECT 198.740 79.510 405.240 80.310 ; 
                RECT 198.740 84.400 405.240 85.200 ; 
                RECT 198.740 76.500 405.240 77.300 ; 
                RECT 198.740 90.715 405.240 91.785 ; 
                RECT 198.740 65.030 405.240 66.830 ; 
                RECT 198.740 117.310 405.240 118.280 ; 
                RECT 198.740 132.560 405.240 133.910 ; 
                RECT 198.740 24.965 405.240 26.765 ; 
                RECT 78.110 144.355 80.030 209.135 ; 
                RECT 88.985 144.355 90.905 209.135 ; 
                RECT 92.825 144.355 94.745 209.135 ; 
                RECT 96.665 144.355 98.585 209.135 ; 
                RECT 112.330 144.355 114.250 209.135 ; 
                RECT 116.170 144.355 118.090 209.135 ; 
                RECT 120.010 144.355 121.930 209.135 ; 
                RECT 123.850 144.355 125.770 209.135 ; 
                RECT 127.690 144.355 129.610 209.135 ; 
                RECT 152.290 144.355 154.210 209.135 ; 
                RECT 156.130 144.355 158.050 209.135 ; 
                RECT 159.970 144.355 161.890 209.135 ; 
                RECT 163.810 144.355 165.730 209.135 ; 
                RECT 167.650 144.355 169.570 209.135 ; 
                RECT 171.490 144.355 173.410 209.135 ; 
                RECT 175.330 144.355 177.250 209.135 ; 
                RECT 179.170 144.355 181.090 209.135 ; 
                RECT 183.010 144.355 184.930 209.135 ; 
                RECT 186.850 144.355 188.770 209.135 ; 
                RECT 190.690 144.355 192.610 209.135 ; 
                RECT 156.580 65.060 158.500 91.860 ; 
                RECT 163.555 65.060 165.475 91.860 ; 
                RECT 173.340 65.060 175.260 91.860 ; 
                RECT 177.180 65.060 179.100 91.860 ; 
                RECT 161.720 119.500 163.640 137.720 ; 
                RECT 168.995 119.500 170.745 137.720 ; 
                RECT 177.175 119.500 179.095 137.720 ; 
                RECT 161.290 97.860 163.210 113.500 ; 
                RECT 168.565 97.860 170.315 113.500 ; 
                RECT 176.960 97.860 178.880 113.500 ; 
                RECT 177.625 55.480 179.545 59.060 ; 
                RECT 23.460 146.625 32.620 147.375 ; 
                RECT 23.460 151.250 32.620 153.000 ; 
                RECT 96.680 134.410 112.720 135.210 ; 
                RECT 79.880 135.070 94.720 136.760 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 207.520 5.560 ; 
                RECT 209.240 5.240 213.640 5.560 ; 
                RECT 215.360 5.240 219.760 5.560 ; 
                RECT 221.480 5.240 225.880 5.560 ; 
                RECT 227.600 5.240 232.000 5.560 ; 
                RECT 233.720 5.240 238.120 5.560 ; 
                RECT 239.840 5.240 244.240 5.560 ; 
                RECT 245.960 5.240 250.360 5.560 ; 
                RECT 252.080 5.240 256.480 5.560 ; 
                RECT 258.200 5.240 262.600 5.560 ; 
                RECT 264.320 5.240 268.720 5.560 ; 
                RECT 270.440 5.240 274.840 5.560 ; 
                RECT 276.560 5.240 280.960 5.560 ; 
                RECT 282.680 5.240 287.080 5.560 ; 
                RECT 288.800 5.240 293.200 5.560 ; 
                RECT 294.920 5.240 299.320 5.560 ; 
                RECT 301.040 5.240 305.440 5.560 ; 
                RECT 307.160 5.240 311.560 5.560 ; 
                RECT 313.280 5.240 317.680 5.560 ; 
                RECT 319.400 5.240 323.800 5.560 ; 
                RECT 325.520 5.240 329.920 5.560 ; 
                RECT 331.640 5.240 336.040 5.560 ; 
                RECT 337.760 5.240 342.160 5.560 ; 
                RECT 343.880 5.240 348.280 5.560 ; 
                RECT 349.320 5.240 354.400 5.560 ; 
                RECT 355.440 5.240 360.520 5.560 ; 
                RECT 361.560 5.240 366.640 5.560 ; 
                RECT 367.680 5.240 372.760 5.560 ; 
                RECT 373.800 5.240 378.880 5.560 ; 
                RECT 379.920 5.240 385.000 5.560 ; 
                RECT 386.040 5.240 391.120 5.560 ; 
                RECT 392.160 5.240 397.240 5.560 ; 
                RECT 398.280 5.240 413.880 5.560 ; 
                RECT 2.880 6.600 413.880 6.920 ; 
                RECT 2.880 7.960 413.880 8.280 ; 
                RECT 2.880 9.320 181.680 9.640 ; 
                RECT 203.120 9.320 413.880 9.640 ; 
                RECT 2.880 10.680 413.880 11.000 ; 
                RECT 2.880 12.040 413.880 12.360 ; 
                RECT 2.880 13.400 125.920 13.720 ; 
                RECT 182.720 13.400 413.880 13.720 ; 
                RECT 2.880 14.760 413.880 15.080 ; 
                RECT 2.880 16.120 413.880 16.440 ; 
                RECT 2.880 17.480 125.920 17.800 ; 
                RECT 182.040 17.480 413.880 17.800 ; 
                RECT 2.880 18.840 197.320 19.160 ; 
                RECT 407.120 18.840 413.880 19.160 ; 
                RECT 2.880 20.200 197.320 20.520 ; 
                RECT 407.120 20.200 413.880 20.520 ; 
                RECT 2.880 21.560 197.320 21.880 ; 
                RECT 407.120 21.560 413.880 21.880 ; 
                RECT 2.880 22.920 197.320 23.240 ; 
                RECT 407.120 22.920 413.880 23.240 ; 
                RECT 2.880 24.280 197.320 24.600 ; 
                RECT 407.120 24.280 413.880 24.600 ; 
                RECT 2.880 25.640 197.320 25.960 ; 
                RECT 407.120 25.640 413.880 25.960 ; 
                RECT 2.880 27.000 197.320 27.320 ; 
                RECT 407.120 27.000 413.880 27.320 ; 
                RECT 2.880 28.360 197.320 28.680 ; 
                RECT 407.120 28.360 413.880 28.680 ; 
                RECT 2.880 29.720 197.320 30.040 ; 
                RECT 407.120 29.720 413.880 30.040 ; 
                RECT 2.880 31.080 197.320 31.400 ; 
                RECT 407.120 31.080 413.880 31.400 ; 
                RECT 2.880 32.440 143.600 32.760 ; 
                RECT 160.960 32.440 197.320 32.760 ; 
                RECT 407.120 32.440 413.880 32.760 ; 
                RECT 2.880 33.800 142.240 34.120 ; 
                RECT 167.080 33.800 197.320 34.120 ; 
                RECT 407.120 33.800 413.880 34.120 ; 
                RECT 2.880 35.160 119.120 35.480 ; 
                RECT 182.040 35.160 197.320 35.480 ; 
                RECT 407.120 35.160 413.880 35.480 ; 
                RECT 2.880 36.520 119.800 36.840 ; 
                RECT 172.520 36.520 196.640 36.840 ; 
                RECT 407.120 36.520 413.880 36.840 ; 
                RECT 2.880 37.880 197.320 38.200 ; 
                RECT 407.120 37.880 413.880 38.200 ; 
                RECT 2.880 39.240 197.320 39.560 ; 
                RECT 407.120 39.240 413.880 39.560 ; 
                RECT 2.880 40.600 197.320 40.920 ; 
                RECT 407.120 40.600 413.880 40.920 ; 
                RECT 2.880 41.960 197.320 42.280 ; 
                RECT 407.120 41.960 413.880 42.280 ; 
                RECT 2.880 43.320 117.080 43.640 ; 
                RECT 128.320 43.320 197.320 43.640 ; 
                RECT 407.120 43.320 413.880 43.640 ; 
                RECT 2.880 44.680 118.440 45.000 ; 
                RECT 120.840 44.680 197.320 45.000 ; 
                RECT 407.120 44.680 413.880 45.000 ; 
                RECT 2.880 46.040 119.800 46.360 ; 
                RECT 124.240 46.040 132.040 46.360 ; 
                RECT 134.440 46.040 197.320 46.360 ; 
                RECT 407.120 46.040 413.880 46.360 ; 
                RECT 2.880 47.400 119.800 47.720 ; 
                RECT 123.560 47.400 197.320 47.720 ; 
                RECT 407.120 47.400 413.880 47.720 ; 
                RECT 2.880 48.760 126.600 49.080 ; 
                RECT 135.120 48.760 197.320 49.080 ; 
                RECT 407.120 48.760 413.880 49.080 ; 
                RECT 2.880 50.120 121.840 50.440 ; 
                RECT 128.320 50.120 197.320 50.440 ; 
                RECT 407.120 50.120 413.880 50.440 ; 
                RECT 2.880 51.480 119.120 51.800 ; 
                RECT 128.320 51.480 197.320 51.800 ; 
                RECT 407.120 51.480 413.880 51.800 ; 
                RECT 2.880 52.840 197.320 53.160 ; 
                RECT 407.120 52.840 413.880 53.160 ; 
                RECT 2.880 54.200 118.440 54.520 ; 
                RECT 128.320 54.200 197.320 54.520 ; 
                RECT 407.120 54.200 413.880 54.520 ; 
                RECT 2.880 55.560 126.600 55.880 ; 
                RECT 133.760 55.560 173.520 55.880 ; 
                RECT 180.000 55.560 197.320 55.880 ; 
                RECT 407.120 55.560 413.880 55.880 ; 
                RECT 2.880 56.920 125.240 57.240 ; 
                RECT 128.320 56.920 173.520 57.240 ; 
                RECT 407.120 56.920 413.880 57.240 ; 
                RECT 2.880 58.280 140.200 58.600 ; 
                RECT 170.480 58.280 173.520 58.600 ; 
                RECT 180.000 58.280 197.320 58.600 ; 
                RECT 407.120 58.280 413.880 58.600 ; 
                RECT 2.880 59.640 126.600 59.960 ; 
                RECT 134.440 59.640 197.320 59.960 ; 
                RECT 407.120 59.640 413.880 59.960 ; 
                RECT 2.880 61.000 123.200 61.320 ; 
                RECT 128.320 61.000 197.320 61.320 ; 
                RECT 407.120 61.000 413.880 61.320 ; 
                RECT 2.880 62.360 125.240 62.680 ; 
                RECT 128.320 62.360 197.320 62.680 ; 
                RECT 407.120 62.360 413.880 62.680 ; 
                RECT 2.880 63.720 197.320 64.040 ; 
                RECT 407.120 63.720 413.880 64.040 ; 
                RECT 2.880 65.080 116.400 65.400 ; 
                RECT 139.880 65.080 141.560 65.400 ; 
                RECT 147.360 65.080 152.440 65.400 ; 
                RECT 180.000 65.080 197.320 65.400 ; 
                RECT 407.120 65.080 413.880 65.400 ; 
                RECT 2.880 66.440 135.440 66.760 ; 
                RECT 141.240 66.440 142.920 66.760 ; 
                RECT 146.000 66.440 152.440 66.760 ; 
                RECT 189.520 66.440 197.320 66.760 ; 
                RECT 407.120 66.440 413.880 66.760 ; 
                RECT 2.880 67.800 125.240 68.120 ; 
                RECT 128.320 67.800 138.160 68.120 ; 
                RECT 141.920 67.800 152.440 68.120 ; 
                RECT 188.160 67.800 197.320 68.120 ; 
                RECT 407.120 67.800 413.880 68.120 ; 
                RECT 2.880 69.160 117.080 69.480 ; 
                RECT 131.040 69.160 152.440 69.480 ; 
                RECT 189.520 69.160 197.320 69.480 ; 
                RECT 407.120 69.160 413.880 69.480 ; 
                RECT 2.880 70.520 125.920 70.840 ; 
                RECT 134.440 70.520 152.440 70.840 ; 
                RECT 189.520 70.520 197.320 70.840 ; 
                RECT 407.120 70.520 413.880 70.840 ; 
                RECT 2.880 71.880 123.880 72.200 ; 
                RECT 135.120 71.880 152.440 72.200 ; 
                RECT 180.000 71.880 197.320 72.200 ; 
                RECT 407.120 71.880 413.880 72.200 ; 
                RECT 2.880 73.240 119.120 73.560 ; 
                RECT 125.600 73.240 152.440 73.560 ; 
                RECT 190.880 73.240 197.320 73.560 ; 
                RECT 407.120 73.240 413.880 73.560 ; 
                RECT 2.880 74.600 152.440 74.920 ; 
                RECT 180.000 74.600 197.320 74.920 ; 
                RECT 407.120 74.600 413.880 74.920 ; 
                RECT 2.880 75.960 118.440 76.280 ; 
                RECT 122.200 75.960 152.440 76.280 ; 
                RECT 192.240 75.960 197.320 76.280 ; 
                RECT 407.120 75.960 413.880 76.280 ; 
                RECT 2.880 77.320 118.440 77.640 ; 
                RECT 128.320 77.320 152.440 77.640 ; 
                RECT 192.240 77.320 197.320 77.640 ; 
                RECT 407.120 77.320 413.880 77.640 ; 
                RECT 2.880 78.680 122.520 79.000 ; 
                RECT 133.760 78.680 152.440 79.000 ; 
                RECT 194.960 78.680 197.320 79.000 ; 
                RECT 407.120 78.680 413.880 79.000 ; 
                RECT 2.880 80.040 125.240 80.360 ; 
                RECT 127.640 80.040 152.440 80.360 ; 
                RECT 193.600 80.040 197.320 80.360 ; 
                RECT 407.120 80.040 413.880 80.360 ; 
                RECT 2.880 81.400 126.600 81.720 ; 
                RECT 128.320 81.400 152.440 81.720 ; 
                RECT 194.960 81.400 197.320 81.720 ; 
                RECT 407.120 81.400 413.880 81.720 ; 
                RECT 2.880 82.760 152.440 83.080 ; 
                RECT 180.000 82.760 197.320 83.080 ; 
                RECT 407.120 82.760 413.880 83.080 ; 
                RECT 2.880 84.120 117.080 84.440 ; 
                RECT 134.440 84.120 152.440 84.440 ; 
                RECT 194.960 84.120 197.320 84.440 ; 
                RECT 407.120 84.120 413.880 84.440 ; 
                RECT 2.880 85.480 117.080 85.800 ; 
                RECT 128.320 85.480 132.040 85.800 ; 
                RECT 134.440 85.480 152.440 85.800 ; 
                RECT 407.120 85.480 413.880 85.800 ; 
                RECT 2.880 86.840 125.920 87.160 ; 
                RECT 128.320 86.840 152.440 87.160 ; 
                RECT 407.120 86.840 413.880 87.160 ; 
                RECT 2.880 88.200 152.440 88.520 ; 
                RECT 407.120 88.200 413.880 88.520 ; 
                RECT 2.880 89.560 152.440 89.880 ; 
                RECT 407.120 89.560 413.880 89.880 ; 
                RECT 2.880 90.920 113.680 91.240 ; 
                RECT 126.960 90.920 152.440 91.240 ; 
                RECT 407.120 90.920 413.880 91.240 ; 
                RECT 2.880 92.280 123.880 92.600 ; 
                RECT 131.040 92.280 197.320 92.600 ; 
                RECT 407.120 92.280 413.880 92.600 ; 
                RECT 2.880 93.640 197.320 93.960 ; 
                RECT 407.120 93.640 413.880 93.960 ; 
                RECT 2.880 95.000 197.320 95.320 ; 
                RECT 407.120 95.000 413.880 95.320 ; 
                RECT 2.880 96.360 122.520 96.680 ; 
                RECT 137.160 96.360 197.320 96.680 ; 
                RECT 407.120 96.360 413.880 96.680 ; 
                RECT 2.880 97.720 157.200 98.040 ; 
                RECT 179.320 97.720 197.320 98.040 ; 
                RECT 407.120 97.720 413.880 98.040 ; 
                RECT 2.880 99.080 157.200 99.400 ; 
                RECT 179.320 99.080 197.320 99.400 ; 
                RECT 407.120 99.080 413.880 99.400 ; 
                RECT 2.880 100.440 119.120 100.760 ; 
                RECT 122.200 100.440 157.200 100.760 ; 
                RECT 179.320 100.440 197.320 100.760 ; 
                RECT 407.120 100.440 413.880 100.760 ; 
                RECT 2.880 101.800 116.400 102.120 ; 
                RECT 120.840 101.800 157.200 102.120 ; 
                RECT 179.320 101.800 197.320 102.120 ; 
                RECT 407.120 101.800 413.880 102.120 ; 
                RECT 2.880 103.160 157.200 103.480 ; 
                RECT 179.320 103.160 197.320 103.480 ; 
                RECT 407.120 103.160 413.880 103.480 ; 
                RECT 2.880 104.520 132.040 104.840 ; 
                RECT 135.120 104.520 157.200 104.840 ; 
                RECT 179.320 104.520 197.320 104.840 ; 
                RECT 407.120 104.520 413.880 104.840 ; 
                RECT 2.880 105.880 157.200 106.200 ; 
                RECT 179.320 105.880 197.320 106.200 ; 
                RECT 407.120 105.880 413.880 106.200 ; 
                RECT 2.880 107.240 157.200 107.560 ; 
                RECT 179.320 107.240 197.320 107.560 ; 
                RECT 407.120 107.240 413.880 107.560 ; 
                RECT 2.880 108.600 157.200 108.920 ; 
                RECT 407.120 108.600 413.880 108.920 ; 
                RECT 2.880 109.960 119.120 110.280 ; 
                RECT 124.240 109.960 157.200 110.280 ; 
                RECT 179.320 109.960 194.600 110.280 ; 
                RECT 407.120 109.960 413.880 110.280 ; 
                RECT 2.880 111.320 157.200 111.640 ; 
                RECT 179.320 111.320 191.880 111.640 ; 
                RECT 407.120 111.320 413.880 111.640 ; 
                RECT 2.880 112.680 95.320 113.000 ; 
                RECT 114.040 112.680 125.240 113.000 ; 
                RECT 133.760 112.680 157.200 113.000 ; 
                RECT 179.320 112.680 189.160 113.000 ; 
                RECT 407.120 112.680 413.880 113.000 ; 
                RECT 2.880 114.040 95.320 114.360 ; 
                RECT 114.040 114.040 186.440 114.360 ; 
                RECT 407.120 114.040 413.880 114.360 ; 
                RECT 2.880 115.400 95.320 115.720 ; 
                RECT 114.040 115.400 121.840 115.720 ; 
                RECT 124.240 115.400 186.440 115.720 ; 
                RECT 407.120 115.400 413.880 115.720 ; 
                RECT 2.880 116.760 95.320 117.080 ; 
                RECT 114.040 116.760 118.440 117.080 ; 
                RECT 121.520 116.760 197.320 117.080 ; 
                RECT 407.120 116.760 413.880 117.080 ; 
                RECT 2.880 118.120 95.320 118.440 ; 
                RECT 114.040 118.120 197.320 118.440 ; 
                RECT 407.120 118.120 413.880 118.440 ; 
                RECT 2.880 119.480 95.320 119.800 ; 
                RECT 114.040 119.480 157.200 119.800 ; 
                RECT 180.000 119.480 197.320 119.800 ; 
                RECT 407.120 119.480 413.880 119.800 ; 
                RECT 2.880 120.840 95.320 121.160 ; 
                RECT 114.040 120.840 157.200 121.160 ; 
                RECT 180.000 120.840 197.320 121.160 ; 
                RECT 407.120 120.840 413.880 121.160 ; 
                RECT 2.880 122.200 95.320 122.520 ; 
                RECT 114.040 122.200 157.200 122.520 ; 
                RECT 180.000 122.200 197.320 122.520 ; 
                RECT 407.120 122.200 413.880 122.520 ; 
                RECT 2.880 123.560 95.320 123.880 ; 
                RECT 114.040 123.560 157.200 123.880 ; 
                RECT 180.000 123.560 187.800 123.880 ; 
                RECT 407.120 123.560 413.880 123.880 ; 
                RECT 2.880 124.920 95.320 125.240 ; 
                RECT 114.040 124.920 157.200 125.240 ; 
                RECT 180.000 124.920 187.800 125.240 ; 
                RECT 407.120 124.920 413.880 125.240 ; 
                RECT 2.880 126.280 95.320 126.600 ; 
                RECT 114.040 126.280 120.480 126.600 ; 
                RECT 124.240 126.280 157.200 126.600 ; 
                RECT 180.000 126.280 190.520 126.600 ; 
                RECT 407.120 126.280 413.880 126.600 ; 
                RECT 2.880 127.640 157.200 127.960 ; 
                RECT 180.000 127.640 193.240 127.960 ; 
                RECT 407.120 127.640 413.880 127.960 ; 
                RECT 2.880 129.000 157.200 129.320 ; 
                RECT 407.120 129.000 413.880 129.320 ; 
                RECT 2.880 130.360 157.200 130.680 ; 
                RECT 407.120 130.360 413.880 130.680 ; 
                RECT 2.880 131.720 79.000 132.040 ; 
                RECT 95.680 131.720 122.520 132.040 ; 
                RECT 128.320 131.720 157.200 132.040 ; 
                RECT 180.000 131.720 197.320 132.040 ; 
                RECT 407.120 131.720 413.880 132.040 ; 
                RECT 2.880 133.080 79.000 133.400 ; 
                RECT 95.680 133.080 101.440 133.400 ; 
                RECT 108.600 133.080 157.200 133.400 ; 
                RECT 180.000 133.080 197.320 133.400 ; 
                RECT 407.120 133.080 413.880 133.400 ; 
                RECT 2.880 134.440 79.000 134.760 ; 
                RECT 113.360 134.440 157.200 134.760 ; 
                RECT 180.000 134.440 197.320 134.760 ; 
                RECT 407.120 134.440 413.880 134.760 ; 
                RECT 2.880 135.800 79.000 136.120 ; 
                RECT 95.680 135.800 157.200 136.120 ; 
                RECT 407.120 135.800 413.880 136.120 ; 
                RECT 2.880 137.160 79.680 137.480 ; 
                RECT 108.600 137.160 117.080 137.480 ; 
                RECT 126.960 137.160 157.200 137.480 ; 
                RECT 180.000 137.160 197.320 137.480 ; 
                RECT 407.120 137.160 413.880 137.480 ; 
                RECT 2.880 138.520 101.440 138.840 ; 
                RECT 121.520 138.520 413.880 138.840 ; 
                RECT 2.880 139.880 29.360 140.200 ; 
                RECT 120.840 139.880 413.880 140.200 ; 
                RECT 2.880 141.240 194.600 141.560 ; 
                RECT 409.160 141.240 413.880 141.560 ; 
                RECT 2.880 142.600 194.600 142.920 ; 
                RECT 409.160 142.600 413.880 142.920 ; 
                RECT 2.880 143.960 24.600 144.280 ; 
                RECT 31.080 143.960 72.880 144.280 ; 
                RECT 409.160 143.960 413.880 144.280 ; 
                RECT 2.880 145.320 22.560 145.640 ; 
                RECT 44.000 145.320 72.880 145.640 ; 
                RECT 409.160 145.320 413.880 145.640 ; 
                RECT 2.880 146.680 22.560 147.000 ; 
                RECT 43.320 146.680 55.200 147.000 ; 
                RECT 63.040 146.680 72.880 147.000 ; 
                RECT 409.160 146.680 413.880 147.000 ; 
                RECT 2.880 148.040 36.840 148.360 ; 
                RECT 41.960 148.040 55.200 148.360 ; 
                RECT 63.040 148.040 72.880 148.360 ; 
                RECT 409.160 148.040 413.880 148.360 ; 
                RECT 2.880 149.400 22.560 149.720 ; 
                RECT 33.120 149.400 55.200 149.720 ; 
                RECT 63.040 149.400 72.880 149.720 ; 
                RECT 409.160 149.400 413.880 149.720 ; 
                RECT 2.880 150.760 22.560 151.080 ; 
                RECT 33.120 150.760 55.200 151.080 ; 
                RECT 63.040 150.760 72.880 151.080 ; 
                RECT 409.160 150.760 413.880 151.080 ; 
                RECT 2.880 152.120 22.560 152.440 ; 
                RECT 33.120 152.120 55.200 152.440 ; 
                RECT 59.640 152.120 72.880 152.440 ; 
                RECT 409.160 152.120 413.880 152.440 ; 
                RECT 2.880 153.480 72.880 153.800 ; 
                RECT 409.160 153.480 413.880 153.800 ; 
                RECT 2.880 154.840 55.200 155.160 ; 
                RECT 63.040 154.840 72.880 155.160 ; 
                RECT 409.160 154.840 413.880 155.160 ; 
                RECT 2.880 156.200 55.200 156.520 ; 
                RECT 63.040 156.200 72.880 156.520 ; 
                RECT 409.160 156.200 413.880 156.520 ; 
                RECT 2.880 157.560 15.760 157.880 ; 
                RECT 18.160 157.560 31.400 157.880 ; 
                RECT 34.480 157.560 60.640 157.880 ; 
                RECT 63.040 157.560 72.880 157.880 ; 
                RECT 409.160 157.560 413.880 157.880 ; 
                RECT 2.880 158.920 15.080 159.240 ; 
                RECT 18.160 158.920 55.200 159.240 ; 
                RECT 63.040 158.920 72.880 159.240 ; 
                RECT 409.160 158.920 413.880 159.240 ; 
                RECT 2.880 160.280 14.400 160.600 ; 
                RECT 18.160 160.280 55.200 160.600 ; 
                RECT 60.320 160.280 72.880 160.600 ; 
                RECT 409.160 160.280 413.880 160.600 ; 
                RECT 2.880 161.640 13.720 161.960 ; 
                RECT 18.160 161.640 57.240 161.960 ; 
                RECT 63.040 161.640 72.880 161.960 ; 
                RECT 409.160 161.640 413.880 161.960 ; 
                RECT 2.880 163.000 55.200 163.320 ; 
                RECT 56.920 163.000 72.880 163.320 ; 
                RECT 409.160 163.000 413.880 163.320 ; 
                RECT 2.880 164.360 13.040 164.680 ; 
                RECT 18.160 164.360 55.200 164.680 ; 
                RECT 61.000 164.360 72.880 164.680 ; 
                RECT 409.160 164.360 413.880 164.680 ; 
                RECT 2.880 165.720 55.200 166.040 ; 
                RECT 63.040 165.720 72.880 166.040 ; 
                RECT 409.160 165.720 413.880 166.040 ; 
                RECT 2.880 167.080 12.360 167.400 ; 
                RECT 18.160 167.080 31.400 167.400 ; 
                RECT 37.880 167.080 55.200 167.400 ; 
                RECT 63.040 167.080 72.880 167.400 ; 
                RECT 409.160 167.080 413.880 167.400 ; 
                RECT 2.880 168.440 11.680 168.760 ; 
                RECT 18.160 168.440 31.400 168.760 ; 
                RECT 36.520 168.440 55.200 168.760 ; 
                RECT 61.680 168.440 72.880 168.760 ; 
                RECT 409.160 168.440 413.880 168.760 ; 
                RECT 2.880 169.800 11.000 170.120 ; 
                RECT 18.160 169.800 31.400 170.120 ; 
                RECT 35.840 169.800 59.280 170.120 ; 
                RECT 63.040 169.800 72.880 170.120 ; 
                RECT 409.160 169.800 413.880 170.120 ; 
                RECT 2.880 171.160 55.200 171.480 ; 
                RECT 63.040 171.160 72.880 171.480 ; 
                RECT 409.160 171.160 413.880 171.480 ; 
                RECT 2.880 172.520 10.320 172.840 ; 
                RECT 18.160 172.520 31.400 172.840 ; 
                RECT 35.160 172.520 55.200 172.840 ; 
                RECT 62.360 172.520 72.880 172.840 ; 
                RECT 409.160 172.520 413.880 172.840 ; 
                RECT 2.880 173.880 9.640 174.200 ; 
                RECT 18.160 173.880 31.400 174.200 ; 
                RECT 34.480 173.880 55.200 174.200 ; 
                RECT 56.920 173.880 72.880 174.200 ; 
                RECT 409.160 173.880 413.880 174.200 ; 
                RECT 2.880 175.240 55.200 175.560 ; 
                RECT 63.040 175.240 72.880 175.560 ; 
                RECT 409.160 175.240 413.880 175.560 ; 
                RECT 2.880 176.600 72.880 176.920 ; 
                RECT 409.160 176.600 413.880 176.920 ; 
                RECT 2.880 177.960 57.240 178.280 ; 
                RECT 63.040 177.960 72.880 178.280 ; 
                RECT 409.160 177.960 413.880 178.280 ; 
                RECT 2.880 179.320 57.920 179.640 ; 
                RECT 63.040 179.320 72.880 179.640 ; 
                RECT 409.160 179.320 413.880 179.640 ; 
                RECT 2.880 180.680 58.600 181.000 ; 
                RECT 63.040 180.680 72.880 181.000 ; 
                RECT 409.160 180.680 413.880 181.000 ; 
                RECT 2.880 182.040 59.280 182.360 ; 
                RECT 63.040 182.040 72.880 182.360 ; 
                RECT 409.160 182.040 413.880 182.360 ; 
                RECT 2.880 183.400 72.880 183.720 ; 
                RECT 409.160 183.400 413.880 183.720 ; 
                RECT 2.880 184.760 34.800 185.080 ; 
                RECT 43.320 184.760 72.880 185.080 ; 
                RECT 409.160 184.760 413.880 185.080 ; 
                RECT 2.880 186.120 33.440 186.440 ; 
                RECT 42.640 186.120 55.200 186.440 ; 
                RECT 63.040 186.120 72.880 186.440 ; 
                RECT 409.160 186.120 413.880 186.440 ; 
                RECT 2.880 187.480 55.200 187.800 ; 
                RECT 63.040 187.480 72.880 187.800 ; 
                RECT 409.160 187.480 413.880 187.800 ; 
                RECT 2.880 188.840 55.200 189.160 ; 
                RECT 63.040 188.840 72.880 189.160 ; 
                RECT 409.160 188.840 413.880 189.160 ; 
                RECT 2.880 190.200 55.200 190.520 ; 
                RECT 63.040 190.200 72.880 190.520 ; 
                RECT 409.160 190.200 413.880 190.520 ; 
                RECT 2.880 191.560 55.200 191.880 ; 
                RECT 58.960 191.560 72.880 191.880 ; 
                RECT 409.160 191.560 413.880 191.880 ; 
                RECT 2.880 192.920 72.880 193.240 ; 
                RECT 409.160 192.920 413.880 193.240 ; 
                RECT 2.880 194.280 57.240 194.600 ; 
                RECT 63.040 194.280 72.880 194.600 ; 
                RECT 409.160 194.280 413.880 194.600 ; 
                RECT 2.880 195.640 57.920 195.960 ; 
                RECT 63.040 195.640 72.880 195.960 ; 
                RECT 409.160 195.640 413.880 195.960 ; 
                RECT 2.880 197.000 58.600 197.320 ; 
                RECT 63.040 197.000 72.880 197.320 ; 
                RECT 409.160 197.000 413.880 197.320 ; 
                RECT 2.880 198.360 59.280 198.680 ; 
                RECT 63.040 198.360 72.880 198.680 ; 
                RECT 409.160 198.360 413.880 198.680 ; 
                RECT 2.880 199.720 72.880 200.040 ; 
                RECT 409.160 199.720 413.880 200.040 ; 
                RECT 2.880 201.080 59.280 201.400 ; 
                RECT 63.040 201.080 72.880 201.400 ; 
                RECT 409.160 201.080 413.880 201.400 ; 
                RECT 2.880 202.440 72.880 202.760 ; 
                RECT 409.160 202.440 413.880 202.760 ; 
                RECT 2.880 203.800 59.960 204.120 ; 
                RECT 63.040 203.800 72.880 204.120 ; 
                RECT 409.160 203.800 413.880 204.120 ; 
                RECT 2.880 205.160 60.640 205.480 ; 
                RECT 63.040 205.160 72.880 205.480 ; 
                RECT 409.160 205.160 413.880 205.480 ; 
                RECT 2.880 206.520 60.640 206.840 ; 
                RECT 63.040 206.520 72.880 206.840 ; 
                RECT 409.160 206.520 413.880 206.840 ; 
                RECT 2.880 207.880 72.880 208.200 ; 
                RECT 409.160 207.880 413.880 208.200 ; 
                RECT 2.880 209.240 72.880 209.560 ; 
                RECT 409.160 209.240 413.880 209.560 ; 
                RECT 2.880 210.600 194.600 210.920 ; 
                RECT 409.160 210.600 413.880 210.920 ; 
                RECT 2.880 211.960 194.600 212.280 ; 
                RECT 409.160 211.960 413.880 212.280 ; 
                RECT 2.880 213.320 413.880 213.640 ; 
                RECT 2.880 214.680 413.880 215.000 ; 
                RECT 2.880 216.040 413.880 216.360 ; 
                RECT 2.880 217.400 413.880 217.720 ; 
                RECT 2.880 218.760 413.880 219.080 ; 
                RECT 2.880 2.880 413.880 4.240 ; 
                RECT 2.880 220.080 413.880 221.440 ; 
                RECT 198.740 38.075 204.540 39.195 ; 
                RECT 399.440 38.075 405.240 39.195 ; 
                RECT 198.740 43.875 204.540 44.525 ; 
                RECT 399.440 43.875 405.240 44.525 ; 
                RECT 198.740 49.085 204.540 49.775 ; 
                RECT 399.440 49.085 405.240 49.775 ; 
                RECT 198.740 54.555 204.540 55.245 ; 
                RECT 399.440 54.555 405.240 55.245 ; 
                RECT 198.740 77.820 405.240 78.620 ; 
                RECT 198.740 107.565 405.240 107.855 ; 
                RECT 198.740 85.720 405.240 86.520 ; 
                RECT 198.740 88.845 405.240 89.915 ; 
                RECT 198.740 121.790 405.240 122.160 ; 
                RECT 198.740 82.510 405.240 83.310 ; 
                RECT 198.740 68.770 405.240 70.570 ; 
                RECT 198.740 80.830 405.240 81.630 ; 
                RECT 198.740 28.705 405.240 30.505 ; 
                RECT 73.765 144.355 75.085 209.135 ; 
                RECT 84.310 144.355 86.230 209.135 ; 
                RECT 102.050 144.355 103.970 209.135 ; 
                RECT 105.890 144.355 107.810 209.135 ; 
                RECT 135.070 144.355 136.990 209.135 ; 
                RECT 138.910 144.355 140.830 209.135 ; 
                RECT 142.750 144.355 144.670 209.135 ; 
                RECT 146.590 144.355 148.510 209.135 ; 
                RECT 153.415 65.060 154.525 91.860 ; 
                RECT 160.930 65.060 161.820 91.860 ; 
                RECT 168.250 65.060 170.170 91.860 ; 
                RECT 158.125 119.500 159.235 137.720 ; 
                RECT 166.500 119.500 167.390 137.720 ; 
                RECT 173.045 119.500 174.365 137.720 ; 
                RECT 157.695 97.860 158.805 113.500 ; 
                RECT 166.070 97.860 166.960 113.500 ; 
                RECT 172.615 97.860 173.935 113.500 ; 
                RECT 174.245 55.480 175.355 59.060 ; 
                RECT 23.460 145.420 32.620 145.790 ; 
                RECT 23.460 148.755 32.620 149.645 ; 
                RECT 79.880 131.580 94.720 132.250 ; 
                RECT 79.880 132.930 94.720 133.940 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 416.760 224.320 ; 
        LAYER met2 ;
            RECT 0.000 0.000 416.760 224.320 ; 
    END 
END sram22_128x32m4w8 
END LIBRARY 

