VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sramgen_sram_512x32m4w8_replica_v1
  CLASS BLOCK ;
  ORIGIN 79.615 342.35 ;
  FOREIGN sramgen_sram_512x32m4w8_replica_v1 -79.615 -342.35 ;
  SIZE 422.075 BY 354.065 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT -73.8 -341.95 -73.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.2 -341.95 -71.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.6 -341.95 -70.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -69 -341.95 -68.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.4 -341.95 -67 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -65.8 -341.95 -65.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.2 -313.02 -63.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.6 -328.92 -62.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -61 -341.95 -60.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.4 -323.62 -59 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.4 -341.95 -59 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.8 -328.92 -57.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.2 -328.92 -55.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.2 -341.95 -55.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.6 -341.95 -54.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -53 -322.56 -52.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -53 -341.95 -52.6 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.4 -328.92 -51 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.8 -328.92 -49.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.8 -341.95 -49.4 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.2 -341.95 -47.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.6 -322.56 -46.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.6 -341.95 -46.2 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -328.92 -44.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -45 -341.95 -44.6 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.4 -341.95 -43 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -320.44 -41.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.8 -341.95 -41.4 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.2 -328.92 -39.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -328.92 -38.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.6 -341.95 -38.2 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -37 -341.95 -36.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -319.38 -35 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.4 -341.95 -35 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.8 -328.92 -33.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.2 -341.95 -31.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -319.38 -30.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.6 -341.95 -30.2 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -319.38 -28.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -29 -341.95 -28.6 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -328.92 -27 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.4 -341.95 -27 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.8 -341.95 -25.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -318.32 -23.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.2 -341.95 -23.8 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.6 -328.92 -22.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -328.92 -20.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -21 -341.95 -20.6 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.4 -341.95 -19 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -317.26 -17.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.8 -341.95 -17.4 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.2 -328.92 -15.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.6 -341.95 -14.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -316.2 -12.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -13 -341.95 -12.6 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -316.2 -11 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.4 -341.95 -11 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -212.32 -9.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -328.92 -9.4 -295.42 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.8 -341.95 -9.4 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.2 -341.95 -7.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -311.96 -6.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.6 -341.95 -6.2 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -5 -341.95 -4.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.4 -341.95 -3 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 2.86 -1.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.8 -341.95 -1.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 2.86 0.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.2 -341.95 0.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 2.86 1.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.4 -341.95 1.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 2.86 3.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 3 -341.95 3.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 2.86 5 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.6 -341.95 5 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 2.86 6.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 -254.72 6.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.2 -341.95 6.6 -293.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 2.86 8.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 -221.86 8.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.8 -290.76 8.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 2.86 9.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 -230.34 9.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.4 -341.95 9.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 2.86 11.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 11 -341.95 11.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 2.86 13 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.6 -296.06 13 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 2.86 14.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.2 -313.02 14.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 2.86 16.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.8 -341.95 16.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 2.86 17.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.4 -341.95 17.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 2.86 19.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 -230.34 19.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 19 -341.95 19.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 2.86 21 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 -221.86 21 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.6 -341.95 21 -314.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 2.86 22.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.2 -341.95 22.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 2.86 24.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.8 -341.95 24.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 2.86 25.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.4 -341.95 25.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 2.86 27.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 27 -341.95 27.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 2.86 29 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 -221.86 29 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.6 -290.76 29 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 2.86 30.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 -221.86 30.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.2 -341.95 30.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 2.86 32.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.8 -297.12 32.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 2.86 33.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -296.06 33.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.4 -341.95 33.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 2.86 35.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 35 -341.95 35.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 2.86 37 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.6 -341.95 37 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 2.86 38.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 -221.86 38.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.2 -290.76 38.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 2.86 40.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 -221.86 40.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.8 -341.95 40.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 2.86 41.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.4 -341.95 41.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 2.86 43.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 43 -341.95 43.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 2.86 45 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.6 -341.95 45 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 2.86 46.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.2 -341.95 46.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 2.86 48.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 -221.86 48.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.8 -290.76 48.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 2.86 49.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 -230.34 49.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.4 -341.95 49.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 2.86 51.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 51 -341.95 51.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 2.86 53 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.6 -296.06 53 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 2.86 54.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.2 -341.95 54.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 2.86 56.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.8 -341.95 56.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 2.86 57.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.4 -341.95 57.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 2.86 59.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 -230.34 59.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 59 -341.95 59.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 2.86 61 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 -221.86 61 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.6 -341.95 61 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 2.86 62.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.2 -341.95 62.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 2.86 64.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.8 -341.95 64.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 2.86 65.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.4 -341.95 65.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 2.86 67.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 67 -341.95 67.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 2.86 69 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 -221.86 69 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.6 -290.76 69 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 2.86 70.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 -221.86 70.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.2 -341.95 70.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 2.86 72.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.8 -297.12 72.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 2.86 73.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -296.06 73.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.4 -341.95 73.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 2.86 75.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 75 -341.95 75.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 2.86 77 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.6 -341.95 77 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 2.86 78.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 -221.86 78.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.2 -290.76 78.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 2.86 80.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 -221.86 80.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.8 -341.95 80.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 2.86 81.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.4 -341.95 81.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 2.86 83.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 83 -341.95 83.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 2.86 85 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.6 -341.95 85 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 2.86 86.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.2 -341.95 86.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 2.86 88.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 -221.86 88.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.8 -290.76 88.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 2.86 89.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 -230.34 89.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.4 -341.95 89.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 2.86 91.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 91 -341.95 91.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 2.86 93 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.6 -296.06 93 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 2.86 94.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.2 -313.02 94.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 2.86 96.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.8 -341.95 96.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 2.86 97.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.4 -341.95 97.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 2.86 99.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 -230.34 99.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 99 -341.95 99.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 2.86 101 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 -221.86 101 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.6 -341.95 101 -314.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 2.86 102.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.2 -341.95 102.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 2.86 104.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.8 -341.95 104.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 2.86 105.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.4 -341.95 105.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 2.86 107.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 107 -341.95 107.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 2.86 109 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 -221.86 109 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.6 -290.76 109 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 2.86 110.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 -221.86 110.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.2 -341.95 110.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 2.86 112.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.8 -297.12 112.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 2.86 113.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -296.06 113.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.4 -341.95 113.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 2.86 115.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 115 -341.95 115.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 2.86 117 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.6 -341.95 117 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 2.86 118.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 -221.86 118.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.2 -290.76 118.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 2.86 120.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 -221.86 120.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.8 -341.95 120.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 2.86 121.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.4 -341.95 121.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 2.86 123.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 123 -341.95 123.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 2.86 125 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.6 -341.95 125 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 2.86 126.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.2 -341.95 126.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 2.86 128.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 -221.86 128.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.8 -290.76 128.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 2.86 129.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 -230.34 129.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.4 -341.95 129.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 2.86 131.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 131 -341.95 131.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 2.86 133 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.6 -296.06 133 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 2.86 134.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.2 -341.95 134.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 2.86 136.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.8 -341.95 136.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 2.86 137.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.4 -341.95 137.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 2.86 139.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 -230.34 139.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 139 -341.95 139.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 2.86 141 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 -221.86 141 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.6 -341.95 141 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 2.86 142.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.2 -341.95 142.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 2.86 144.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.8 -341.95 144.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 2.86 145.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.4 -341.95 145.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 2.86 147.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 147 -341.95 147.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 2.86 149 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 -221.86 149 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.6 -290.76 149 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 2.86 150.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 -221.86 150.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.2 -341.95 150.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 2.86 152.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.8 -297.12 152.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 2.86 153.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -296.06 153.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.4 -341.95 153.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 2.86 155.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 155 -341.95 155.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 2.86 157 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.6 -341.95 157 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 2.86 158.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 -221.86 158.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.2 -290.76 158.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 2.86 160.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 -221.86 160.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.8 -341.95 160.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 2.86 161.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.4 -341.95 161.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 2.86 163.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 163 -341.95 163.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 2.86 165 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.6 -341.95 165 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 2.86 166.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.2 -341.95 166.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 2.86 168.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 -221.86 168.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.8 -290.76 168.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 2.86 169.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 -230.34 169.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.4 -341.95 169.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 171 2.86 171.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 171 -341.95 171.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 2.86 173 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.6 -296.06 173 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 2.86 174.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.2 -313.02 174.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.8 2.86 176.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.8 -341.95 176.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.4 2.86 177.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.4 -341.95 177.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 179 2.86 179.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 179 -230.34 179.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 179 -341.95 179.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.6 2.86 181 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.6 -221.86 181 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.6 -341.95 181 -314.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.2 2.86 182.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.2 -341.95 182.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.8 2.86 184.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.8 -341.95 184.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.4 2.86 185.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.4 -341.95 185.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 187 2.86 187.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 187 -341.95 187.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.6 2.86 189 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.6 -221.86 189 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.6 -290.76 189 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.2 2.86 190.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.2 -221.86 190.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.2 -341.95 190.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.8 2.86 192.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.8 -297.12 192.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 2.86 193.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 -296.06 193.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.4 -341.95 193.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 2.86 195.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 195 -341.95 195.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 2.86 197 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.6 -341.95 197 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.2 2.86 198.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.2 -221.86 198.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.2 -290.76 198.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.8 2.86 200.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.8 -221.86 200.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.8 -341.95 200.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.4 2.86 201.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.4 -341.95 201.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 203 2.86 203.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 203 -341.95 203.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.6 2.86 205 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.6 -341.95 205 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.2 2.86 206.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.2 -341.95 206.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.8 2.86 208.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.8 -221.86 208.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.8 -290.76 208.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.4 2.86 209.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.4 -230.34 209.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.4 -341.95 209.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 211 2.86 211.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 211 -341.95 211.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 2.86 213 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.6 -296.06 213 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 2.86 214.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.2 -341.95 214.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.8 2.86 216.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.8 -341.95 216.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.4 2.86 217.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.4 -341.95 217.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 219 2.86 219.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 219 -230.34 219.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 219 -341.95 219.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.6 2.86 221 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.6 -221.86 221 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.6 -341.95 221 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.2 2.86 222.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.2 -341.95 222.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 2.86 224.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.8 -341.95 224.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.4 2.86 225.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.4 -341.95 225.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 227 2.86 227.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 227 -341.95 227.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.6 2.86 229 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.6 -221.86 229 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.6 -290.76 229 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.2 2.86 230.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.2 -221.86 230.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.2 -341.95 230.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.8 2.86 232.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.8 -297.12 232.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 2.86 233.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 -296.06 233.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.4 -341.95 233.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 2.86 235.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 235 -341.95 235.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.6 2.86 237 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.6 -341.95 237 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.2 2.86 238.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.2 -221.86 238.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.2 -290.76 238.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.8 2.86 240.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.8 -221.86 240.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.8 -341.95 240.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.4 2.86 241.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.4 -341.95 241.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 243 2.86 243.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 243 -341.95 243.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.6 2.86 245 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.6 -341.95 245 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.2 2.86 246.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.2 -341.95 246.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.8 2.86 248.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.8 -221.86 248.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.8 -290.76 248.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 2.86 249.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 -230.34 249.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.4 -341.95 249.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 251 2.86 251.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 251 -341.95 251.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 2.86 253 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.6 -296.06 253 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 2.86 254.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.2 -313.02 254.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.8 2.86 256.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.8 -341.95 256.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.4 2.86 257.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.4 -341.95 257.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 259 2.86 259.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 259 -230.34 259.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 259 -341.95 259.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.6 2.86 261 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.6 -221.86 261 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.6 -341.95 261 -314.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.2 2.86 262.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.2 -341.95 262.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 2.86 264.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.8 -341.95 264.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.4 2.86 265.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.4 -341.95 265.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 267 2.86 267.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 267 -341.95 267.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.6 2.86 269 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.6 -221.86 269 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.6 -290.76 269 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.2 2.86 270.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.2 -221.86 270.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.2 -341.95 270.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.8 2.86 272.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.8 -297.12 272.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 2.86 273.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 -296.06 273.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.4 -341.95 273.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 2.86 275.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 275 -341.95 275.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.6 2.86 277 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.6 -341.95 277 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.2 2.86 278.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.2 -221.86 278.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.2 -290.76 278.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.8 2.86 280.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.8 -221.86 280.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.8 -341.95 280.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.4 2.86 281.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.4 -341.95 281.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 283 2.86 283.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 283 -341.95 283.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.6 2.86 285 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.6 -341.95 285 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.2 2.86 286.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.2 -341.95 286.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.8 2.86 288.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.8 -221.86 288.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.8 -290.76 288.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.4 2.86 289.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.4 -230.34 289.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.4 -341.95 289.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 291 2.86 291.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 291 -341.95 291.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 2.86 293 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.6 -296.06 293 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 2.86 294.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.2 -341.95 294.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.8 2.86 296.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.8 -341.95 296.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.4 2.86 297.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.4 -341.95 297.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 299 2.86 299.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 299 -230.34 299.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 299 -341.95 299.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.6 2.86 301 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.6 -221.86 301 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.6 -341.95 301 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.2 2.86 302.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.2 -341.95 302.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 2.86 304.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.8 -341.95 304.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.4 2.86 305.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.4 -341.95 305.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 307 2.86 307.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 307 -341.95 307.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.6 2.86 309 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.6 -221.86 309 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.6 -290.76 309 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.2 2.86 310.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.2 -221.86 310.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.2 -341.95 310.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.8 2.86 312.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.8 -297.12 312.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 2.86 313.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 -296.06 313.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.4 -341.95 313.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 2.86 315.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 315 -341.95 315.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.6 2.86 317 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.6 -341.95 317 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.2 2.86 318.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.2 -221.86 318.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.2 -290.76 318.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.8 2.86 320.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.8 -221.86 320.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.8 -341.95 320.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.4 2.86 321.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.4 -341.95 321.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 323 2.86 323.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 323 -341.95 323.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.6 2.86 325 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.6 -341.95 325 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.2 2.86 326.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.2 -341.95 326.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.8 2.86 328.2 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.8 -341.95 328.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.4 2.86 329.8 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.4 -341.95 329.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 331 -341.95 331.4 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.6 -341.95 333 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.2 -341.95 334.6 11.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.8 -341.95 336.2 11.315 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT -74.6 -340.41 -74.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -73 -340.41 -72.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.4 -340.41 -71 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -69.8 -340.41 -69.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.2 -340.41 -67.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.6 -340.41 -66.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -65 -340.41 -64.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -63.4 -313.02 -63 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.8 -328.92 -61.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.8 -340.41 -61.4 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.2 -340.41 -59.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.6 -323.62 -58.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.6 -340.41 -58.2 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -57 -328.92 -56.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.4 -340.41 -55 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.8 -322.56 -53.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.8 -340.41 -53.4 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.2 -323.62 -51.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.6 -328.92 -50.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.6 -340.41 -50.2 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -49 -340.41 -48.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.4 -321.5 -47 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.4 -340.41 -47 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.8 -328.92 -45.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -328.92 -43.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.2 -340.41 -43.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.6 -340.41 -42.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -320.44 -40.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -41 -340.41 -40.6 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.4 -328.92 -39 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.8 -340.41 -37.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -319.38 -35.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.2 -340.41 -35.8 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.6 -320.44 -34.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -328.92 -32.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -33 -340.41 -32.6 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.4 -340.41 -31 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -319.38 -29.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.8 -340.41 -29.4 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.2 -328.92 -27.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -328.92 -26.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.6 -340.41 -26.2 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -25 -340.41 -24.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -318.32 -23 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.4 -340.41 -23 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.8 -328.92 -21.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.2 -340.41 -19.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -317.26 -18.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.6 -340.41 -18.2 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -17 -317.26 -16.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -328.92 -15 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.4 -340.41 -15 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.8 -340.41 -13.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -316.2 -11.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.2 -340.41 -11.8 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -212.32 -10.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.6 -328.92 -10.2 -295.42 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -328.92 -8.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -9 -340.41 -8.6 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.4 -340.41 -7 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -311.96 -5.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.8 -340.41 -5.4 -331.46 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.2 -340.41 -3.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.6 -340.41 -2.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 2.86 -0.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT -1 -340.41 -0.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 2.86 1 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.6 -340.41 1 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 2.86 2.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.2 -340.41 2.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 2.86 4.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.8 -340.41 4.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 2.86 5.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 -254.72 5.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.4 -340.41 5.8 -293.3 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 2.86 7.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 7 -340.41 7.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 2.86 9 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 -221.86 9 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.6 -290.76 9 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 2.86 10.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 -221.86 10.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.2 -340.41 10.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 2.86 12.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.8 -297.12 12.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 2.86 13.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -296.06 13.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.4 -340.41 13.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 2.86 15.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 15 -340.41 15.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 2.86 17 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.6 -340.41 17 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 2.86 18.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 -221.86 18.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.2 -290.76 18.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 2.86 20.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 -221.86 20.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.8 -340.41 20.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 2.86 21.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 -235.64 21.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.4 -340.41 21.8 -314.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 2.86 23.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 23 -340.41 23.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 2.86 25 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.6 -340.41 25 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 2.86 26.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.2 -340.41 26.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 2.86 28.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 -221.86 28.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.8 -290.76 28.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 2.86 29.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 -230.34 29.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.4 -340.41 29.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 2.86 31.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 31 -340.41 31.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 2.86 33 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.6 -296.06 33 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 2.86 34.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.2 -340.41 34.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 2.86 36.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.8 -340.41 36.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 2.86 37.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.4 -340.41 37.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 2.86 39.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 -230.34 39.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 39 -340.41 39.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 2.86 41 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 -221.86 41 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.6 -340.41 41 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 2.86 42.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.2 -340.41 42.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 2.86 44.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.8 -340.41 44.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 2.86 45.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.4 -340.41 45.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 2.86 47.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 47 -340.41 47.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 2.86 49 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 -221.86 49 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.6 -290.76 49 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 2.86 50.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 -221.86 50.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.2 -340.41 50.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 2.86 52.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.8 -297.12 52.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 2.86 53.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -296.06 53.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.4 -340.41 53.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 2.86 55.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 55 -340.41 55.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 2.86 57 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.6 -340.41 57 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 2.86 58.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 -221.86 58.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.2 -290.76 58.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 2.86 60.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 -221.86 60.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.8 -340.41 60.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 2.86 61.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.4 -340.41 61.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 2.86 63.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 63 -340.41 63.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 2.86 65 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.6 -340.41 65 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 2.86 66.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.2 -340.41 66.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 2.86 68.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 -221.86 68.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.8 -290.76 68.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 2.86 69.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 -230.34 69.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.4 -340.41 69.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 2.86 71.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 71 -340.41 71.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 2.86 73 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.6 -296.06 73 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 2.86 74.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.2 -340.41 74.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 2.86 76.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.8 -340.41 76.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 2.86 77.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.4 -340.41 77.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 2.86 79.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 -230.34 79.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 79 -340.41 79.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 2.86 81 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 -221.86 81 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.6 -340.41 81 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 2.86 82.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.2 -340.41 82.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 2.86 84.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.8 -340.41 84.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 2.86 85.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.4 -340.41 85.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 2.86 87.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 87 -340.41 87.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 2.86 89 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 -221.86 89 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.6 -290.76 89 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 2.86 90.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 -221.86 90.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.2 -340.41 90.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 2.86 92.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.8 -297.12 92.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 2.86 93.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -296.06 93.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.4 -340.41 93.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 2.86 95.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 95 -340.41 95.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 2.86 97 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.6 -340.41 97 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 2.86 98.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 -221.86 98.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.2 -290.76 98.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 2.86 100.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 -221.86 100.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.8 -340.41 100.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 2.86 101.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 -235.64 101.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.4 -340.41 101.8 -314.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 2.86 103.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 103 -340.41 103.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 2.86 105 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.6 -340.41 105 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 2.86 106.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.2 -340.41 106.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 2.86 108.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 -221.86 108.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.8 -290.76 108.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 2.86 109.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 -230.34 109.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.4 -340.41 109.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 2.86 111.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 111 -340.41 111.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 2.86 113 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.6 -296.06 113 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 2.86 114.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.2 -340.41 114.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 2.86 116.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.8 -340.41 116.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 2.86 117.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.4 -340.41 117.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 2.86 119.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 -230.34 119.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 119 -340.41 119.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 2.86 121 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 -221.86 121 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.6 -340.41 121 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 2.86 122.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.2 -340.41 122.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 2.86 124.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.8 -340.41 124.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 2.86 125.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.4 -340.41 125.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 2.86 127.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 127 -340.41 127.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 2.86 129 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 -221.86 129 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.6 -290.76 129 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 2.86 130.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 -221.86 130.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.2 -340.41 130.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 2.86 132.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.8 -297.12 132.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 2.86 133.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -296.06 133.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.4 -340.41 133.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 2.86 135.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 135 -340.41 135.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 2.86 137 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.6 -340.41 137 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 2.86 138.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 -221.86 138.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.2 -290.76 138.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 2.86 140.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 -221.86 140.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.8 -340.41 140.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 2.86 141.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.4 -340.41 141.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 2.86 143.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 143 -340.41 143.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 2.86 145 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.6 -340.41 145 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 2.86 146.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.2 -340.41 146.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 2.86 148.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 -221.86 148.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.8 -290.76 148.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 2.86 149.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 -230.34 149.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.4 -340.41 149.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 2.86 151.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 151 -340.41 151.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 2.86 153 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.6 -296.06 153 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 2.86 154.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.2 -340.41 154.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 2.86 156.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.8 -340.41 156.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 2.86 157.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.4 -340.41 157.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 2.86 159.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 -230.34 159.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 159 -340.41 159.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 2.86 161 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 -221.86 161 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.6 -340.41 161 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 2.86 162.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.2 -340.41 162.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 2.86 164.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.8 -340.41 164.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 2.86 165.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.4 -340.41 165.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 2.86 167.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 167 -340.41 167.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 2.86 169 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 -221.86 169 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.6 -290.76 169 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 2.86 170.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 -221.86 170.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.2 -340.41 170.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.8 2.86 172.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.8 -297.12 172.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 2.86 173.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 -296.06 173.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.4 -340.41 173.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 2.86 175.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 175 -340.41 175.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.6 2.86 177 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.6 -340.41 177 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.2 2.86 178.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.2 -221.86 178.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.2 -290.76 178.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.8 2.86 180.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.8 -221.86 180.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.8 -340.41 180.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.4 2.86 181.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.4 -235.64 181.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.4 -340.41 181.8 -314.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 183 2.86 183.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 183 -340.41 183.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.6 2.86 185 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.6 -340.41 185 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.2 2.86 186.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.2 -340.41 186.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.8 2.86 188.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.8 -221.86 188.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.8 -290.76 188.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.4 2.86 189.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.4 -230.34 189.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.4 -340.41 189.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 191 2.86 191.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 191 -340.41 191.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 2.86 193 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.6 -296.06 193 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 2.86 194.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.2 -340.41 194.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 2.86 196.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.8 -340.41 196.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.4 2.86 197.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.4 -340.41 197.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 199 2.86 199.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 199 -230.34 199.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 199 -340.41 199.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.6 2.86 201 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.6 -221.86 201 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.6 -340.41 201 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.2 2.86 202.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.2 -340.41 202.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.8 2.86 204.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.8 -340.41 204.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.4 2.86 205.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.4 -340.41 205.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 207 2.86 207.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 207 -340.41 207.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.6 2.86 209 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.6 -221.86 209 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.6 -290.76 209 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.2 2.86 210.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.2 -221.86 210.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.2 -340.41 210.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.8 2.86 212.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.8 -297.12 212.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 2.86 213.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 -296.06 213.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.4 -340.41 213.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 2.86 215.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 215 -340.41 215.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.6 2.86 217 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.6 -340.41 217 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.2 2.86 218.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.2 -221.86 218.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.2 -290.76 218.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.8 2.86 220.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.8 -221.86 220.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.8 -340.41 220.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.4 2.86 221.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.4 -340.41 221.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 223 2.86 223.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 223 -340.41 223.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.6 2.86 225 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.6 -340.41 225 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.2 2.86 226.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.2 -340.41 226.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.8 2.86 228.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.8 -221.86 228.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.8 -290.76 228.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.4 2.86 229.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.4 -230.34 229.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.4 -340.41 229.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 231 2.86 231.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 231 -340.41 231.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 2.86 233 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.6 -296.06 233 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 2.86 234.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.2 -340.41 234.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.8 2.86 236.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.8 -340.41 236.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.4 2.86 237.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.4 -340.41 237.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 239 2.86 239.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 239 -230.34 239.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 239 -340.41 239.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.6 2.86 241 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.6 -221.86 241 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.6 -340.41 241 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.2 2.86 242.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.2 -340.41 242.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.8 2.86 244.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.8 -340.41 244.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.4 2.86 245.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.4 -340.41 245.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 247 2.86 247.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 247 -340.41 247.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.6 2.86 249 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.6 -221.86 249 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.6 -290.76 249 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.2 2.86 250.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.2 -221.86 250.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.2 -340.41 250.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.8 2.86 252.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.8 -297.12 252.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 2.86 253.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 -296.06 253.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.4 -340.41 253.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 2.86 255.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 255 -340.41 255.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.6 2.86 257 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.6 -340.41 257 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.2 2.86 258.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.2 -221.86 258.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.2 -290.76 258.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.8 2.86 260.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.8 -221.86 260.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.8 -340.41 260.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.4 2.86 261.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.4 -235.64 261.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.4 -340.41 261.8 -314.5 ;
    END
    PORT
      LAYER met3 ;
        RECT 263 2.86 263.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 263 -340.41 263.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.6 2.86 265 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.6 -340.41 265 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.2 2.86 266.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.2 -340.41 266.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.8 2.86 268.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.8 -221.86 268.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.8 -290.76 268.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.4 2.86 269.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.4 -230.34 269.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.4 -340.41 269.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 271 2.86 271.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 271 -340.41 271.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 2.86 273 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.6 -296.06 273 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 2.86 274.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.2 -340.41 274.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.8 2.86 276.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.8 -340.41 276.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.4 2.86 277.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.4 -340.41 277.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 279 2.86 279.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 279 -230.34 279.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 279 -340.41 279.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.6 2.86 281 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.6 -221.86 281 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.6 -340.41 281 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.2 2.86 282.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.2 -340.41 282.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.8 2.86 284.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.8 -340.41 284.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.4 2.86 285.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.4 -340.41 285.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 287 2.86 287.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 287 -340.41 287.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.6 2.86 289 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.6 -221.86 289 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.6 -290.76 289 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 2.86 290.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 -221.86 290.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.2 -340.41 290.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.8 2.86 292.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.8 -297.12 292.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 2.86 293.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 -296.06 293.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.4 -340.41 293.8 -334.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 2.86 295.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 295 -340.41 295.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.6 2.86 297 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.6 -340.41 297 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.2 2.86 298.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.2 -221.86 298.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.2 -290.76 298.6 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.8 2.86 300.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.8 -221.86 300.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.8 -340.41 300.2 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.4 2.86 301.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.4 -340.41 301.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 303 2.86 303.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 303 -340.41 303.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.6 2.86 305 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.6 -340.41 305 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.2 2.86 306.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.2 -340.41 306.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.8 2.86 308.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.8 -221.86 308.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.8 -290.76 308.2 -281.64 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.4 2.86 309.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.4 -230.34 309.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.4 -340.41 309.8 -297.54 ;
    END
    PORT
      LAYER met3 ;
        RECT 311 2.86 311.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 311 -340.41 311.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 2.86 313 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.6 -296.06 313 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 2.86 314.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.2 -340.41 314.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.8 2.86 316.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.8 -340.41 316.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.4 2.86 317.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.4 -340.41 317.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 319 2.86 319.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 319 -230.34 319.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 319 -340.41 319.4 -304.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.6 2.86 321 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.6 -221.86 321 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.6 -340.41 321 -281.64 ;
        RECT 320.58 -287.06 321 -286.73 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.2 2.86 322.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.2 -340.41 322.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.8 2.86 324.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.8 -340.41 324.2 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.4 2.86 325.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.4 -340.41 325.8 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 327 2.86 327.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 327 -340.41 327.4 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.6 2.86 329 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.6 -340.41 329 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.2 2.86 330.6 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.2 -340.41 330.6 -211.68 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.8 -340.41 332.2 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.4 -340.41 333.8 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 335 -340.41 335.4 9.775 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.6 -340.41 337 9.775 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -16.46 -342.35 -16.16 -342.05 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -22.3 -342.35 -22 -342.05 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -28.14 -342.35 -27.84 -342.05 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -33.98 -342.35 -33.68 -342.05 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -39.82 -342.35 -39.52 -342.05 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -45.66 -342.35 -45.36 -342.05 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -51.5 -342.35 -51.2 -342.05 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -57.34 -342.35 -57.04 -342.05 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -63.18 -342.35 -62.88 -342.05 ;
    END
  END addr[8]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -64.2 -342.35 -63.78 -341.93 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 12.015 -342.35 12.315 -342.05 ;
    END
  END din[0]
  PIN din[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 112.015 -342.35 112.315 -342.05 ;
    END
  END din[10]
  PIN din[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 112.63 -342.35 112.93 -342.05 ;
    END
  END din[11]
  PIN din[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 132.015 -342.35 132.315 -342.05 ;
    END
  END din[12]
  PIN din[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 132.63 -342.35 132.93 -342.05 ;
    END
  END din[13]
  PIN din[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 152.015 -342.35 152.315 -342.05 ;
    END
  END din[14]
  PIN din[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 152.63 -342.35 152.93 -342.05 ;
    END
  END din[15]
  PIN din[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 172.015 -342.35 172.315 -342.05 ;
    END
  END din[16]
  PIN din[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 172.63 -342.35 172.93 -342.05 ;
    END
  END din[17]
  PIN din[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 192.015 -342.35 192.315 -342.05 ;
    END
  END din[18]
  PIN din[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 192.63 -342.35 192.93 -342.05 ;
    END
  END din[19]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 12.63 -342.35 12.93 -342.05 ;
    END
  END din[1]
  PIN din[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.015 -342.35 212.315 -342.05 ;
    END
  END din[20]
  PIN din[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.63 -342.35 212.93 -342.05 ;
    END
  END din[21]
  PIN din[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 232.015 -342.35 232.315 -342.05 ;
    END
  END din[22]
  PIN din[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 232.63 -342.35 232.93 -342.05 ;
    END
  END din[23]
  PIN din[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 252.015 -342.35 252.315 -342.05 ;
    END
  END din[24]
  PIN din[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 252.63 -342.35 252.93 -342.05 ;
    END
  END din[25]
  PIN din[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 272.015 -342.35 272.315 -342.05 ;
    END
  END din[26]
  PIN din[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 272.63 -342.35 272.93 -342.05 ;
    END
  END din[27]
  PIN din[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 292.015 -342.35 292.315 -342.05 ;
    END
  END din[28]
  PIN din[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 292.63 -342.35 292.93 -342.05 ;
    END
  END din[29]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 32.015 -342.35 32.315 -342.05 ;
    END
  END din[2]
  PIN din[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 312.015 -342.35 312.315 -342.05 ;
    END
  END din[30]
  PIN din[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 312.63 -342.35 312.93 -342.05 ;
    END
  END din[31]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 32.63 -342.35 32.93 -342.05 ;
    END
  END din[3]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 52.015 -342.35 52.315 -342.05 ;
    END
  END din[4]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 52.63 -342.35 52.93 -342.05 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.015 -342.35 72.315 -342.05 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 72.63 -342.35 72.93 -342.05 ;
    END
  END din[7]
  PIN din[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 92.015 -342.35 92.315 -342.05 ;
    END
  END din[8]
  PIN din[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 92.63 -342.35 92.93 -342.05 ;
    END
  END din[9]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 8.285 -342.35 8.585 -342.05 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 108.285 -342.35 108.585 -342.05 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 118.285 -342.35 118.585 -342.05 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.285 -342.35 128.585 -342.05 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 138.285 -342.35 138.585 -342.05 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 148.285 -342.35 148.585 -342.05 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.285 -342.35 158.585 -342.05 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 168.285 -342.35 168.585 -342.05 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.285 -342.35 178.585 -342.05 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 188.285 -342.35 188.585 -342.05 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 198.285 -342.35 198.585 -342.05 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 18.285 -342.35 18.585 -342.05 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 208.285 -342.35 208.585 -342.05 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 218.285 -342.35 218.585 -342.05 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 228.285 -342.35 228.585 -342.05 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 238.285 -342.35 238.585 -342.05 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 248.285 -342.35 248.585 -342.05 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 258.285 -342.35 258.585 -342.05 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 268.285 -342.35 268.585 -342.05 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 278.285 -342.35 278.585 -342.05 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 288.285 -342.35 288.585 -342.05 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 298.285 -342.35 298.585 -342.05 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 28.285 -342.35 28.585 -342.05 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 308.285 -342.35 308.585 -342.05 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 318.285 -342.35 318.585 -342.05 ;
    END
  END dout[31]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 38.285 -342.35 38.585 -342.05 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 48.285 -342.35 48.585 -342.05 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.285 -342.35 58.585 -342.05 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 68.285 -342.35 68.585 -342.05 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 78.285 -342.35 78.585 -342.05 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 88.285 -342.35 88.585 -342.05 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 98.285 -342.35 98.585 -342.05 ;
    END
  END dout[9]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -10.62 -342.35 -10.32 -342.05 ;
    END
  END we
  PIN wmask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 14.125 -342.35 14.425 -342.05 ;
    END
  END wmask[0]
  PIN wmask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 94.125 -342.35 94.425 -342.05 ;
    END
  END wmask[1]
  PIN wmask[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 174.125 -342.35 174.425 -342.05 ;
    END
  END wmask[2]
  PIN wmask[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.125 -342.35 254.425 -342.05 ;
    END
  END wmask[3]
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -79.615 -342.35 342.46 11.715 ;
    LAYER met2 SPACING 0.14 ;
      RECT -79.615 -342.35 342.46 11.715 ;
    LAYER met3 SPACING 0.3 ;
      RECT 320.115 -265.25 320.445 -264.92 ;
      RECT 320.13 -280.68 320.43 -264.92 ;
      RECT 320.115 -280.68 320.445 -280.35 ;
      RECT 320.13 -261.465 320.43 -222.48 ;
      RECT 320.115 -224.455 320.445 -224.125 ;
      RECT 320.115 -261.055 320.445 -260.725 ;
      RECT 319.515 -304.57 319.815 -231.5 ;
      RECT 319.5 -231.875 319.83 -231.545 ;
      RECT 319.5 -248.835 319.83 -248.505 ;
      RECT 319.5 -304.57 319.83 -304.24 ;
      RECT 318.9 -244.175 319.2 -232.13 ;
      RECT 318.885 -232.505 319.215 -232.175 ;
      RECT 318.885 -244.175 319.215 -243.845 ;
      RECT 318.27 -291.655 318.6 -291.325 ;
      RECT 318.285 -341.56 318.585 -291.325 ;
      RECT 318.27 -265.71 318.6 -265.38 ;
      RECT 318.285 -280.68 318.585 -265.38 ;
      RECT 318.27 -280.68 318.6 -280.35 ;
      RECT 318.285 -261.485 318.585 -222.48 ;
      RECT 318.27 -222.855 318.6 -222.525 ;
      RECT 318.27 -261.485 318.6 -261.155 ;
      RECT 313.245 -297.045 313.575 -296.715 ;
      RECT 313.26 -334.29 313.56 -296.715 ;
      RECT 313.245 -304.285 313.575 -303.955 ;
      RECT 313.245 -334.245 313.575 -333.915 ;
      RECT 312.615 -303.485 312.945 -303.155 ;
      RECT 312.63 -341.56 312.93 -303.155 ;
      RECT 312 -297.845 312.33 -297.515 ;
      RECT 312.015 -341.56 312.315 -297.515 ;
      RECT 310.115 -265.25 310.445 -264.92 ;
      RECT 310.13 -280.68 310.43 -264.92 ;
      RECT 310.115 -280.68 310.445 -280.35 ;
      RECT 310.13 -261.465 310.43 -222.48 ;
      RECT 310.115 -224.455 310.445 -224.125 ;
      RECT 310.115 -261.055 310.445 -260.725 ;
      RECT 309.515 -296.56 309.815 -231.5 ;
      RECT 309.5 -231.875 309.83 -231.545 ;
      RECT 309.5 -248.835 309.83 -248.505 ;
      RECT 309.5 -296.56 309.83 -296.23 ;
      RECT 308.9 -244.175 309.2 -232.13 ;
      RECT 308.885 -232.505 309.215 -232.175 ;
      RECT 308.885 -244.175 309.215 -243.845 ;
      RECT 308.27 -291.655 308.6 -291.325 ;
      RECT 308.285 -341.56 308.585 -291.325 ;
      RECT 308.27 -265.71 308.6 -265.38 ;
      RECT 308.285 -280.68 308.585 -265.38 ;
      RECT 308.27 -280.68 308.6 -280.35 ;
      RECT 308.285 -261.485 308.585 -222.48 ;
      RECT 308.27 -222.855 308.6 -222.525 ;
      RECT 308.27 -261.485 308.6 -261.155 ;
      RECT 300.115 -265.25 300.445 -264.92 ;
      RECT 300.13 -280.68 300.43 -264.92 ;
      RECT 300.115 -280.68 300.445 -280.35 ;
      RECT 300.13 -261.465 300.43 -222.48 ;
      RECT 300.115 -224.455 300.445 -224.125 ;
      RECT 300.115 -261.055 300.445 -260.725 ;
      RECT 299.515 -304.57 299.815 -231.5 ;
      RECT 299.5 -231.875 299.83 -231.545 ;
      RECT 299.5 -248.835 299.83 -248.505 ;
      RECT 299.5 -304.57 299.83 -304.24 ;
      RECT 298.9 -244.175 299.2 -232.13 ;
      RECT 298.885 -232.505 299.215 -232.175 ;
      RECT 298.885 -244.175 299.215 -243.845 ;
      RECT 298.27 -291.655 298.6 -291.325 ;
      RECT 298.285 -341.56 298.585 -291.325 ;
      RECT 298.27 -265.71 298.6 -265.38 ;
      RECT 298.285 -280.68 298.585 -265.38 ;
      RECT 298.27 -280.68 298.6 -280.35 ;
      RECT 298.285 -261.485 298.585 -222.48 ;
      RECT 298.27 -222.855 298.6 -222.525 ;
      RECT 298.27 -261.485 298.6 -261.155 ;
      RECT 293.245 -297.045 293.575 -296.715 ;
      RECT 293.26 -334.29 293.56 -296.715 ;
      RECT 293.245 -304.285 293.575 -303.955 ;
      RECT 293.245 -334.245 293.575 -333.915 ;
      RECT 292.615 -303.485 292.945 -303.155 ;
      RECT 292.63 -341.56 292.93 -303.155 ;
      RECT 292 -297.845 292.33 -297.515 ;
      RECT 292.015 -341.56 292.315 -297.515 ;
      RECT 290.115 -265.25 290.445 -264.92 ;
      RECT 290.13 -280.68 290.43 -264.92 ;
      RECT 290.115 -280.68 290.445 -280.35 ;
      RECT 290.13 -261.465 290.43 -222.48 ;
      RECT 290.115 -224.455 290.445 -224.125 ;
      RECT 290.115 -261.055 290.445 -260.725 ;
      RECT 289.515 -296.56 289.815 -231.5 ;
      RECT 289.5 -231.875 289.83 -231.545 ;
      RECT 289.5 -248.835 289.83 -248.505 ;
      RECT 289.5 -296.56 289.83 -296.23 ;
      RECT 288.9 -244.175 289.2 -232.13 ;
      RECT 288.885 -232.505 289.215 -232.175 ;
      RECT 288.885 -244.175 289.215 -243.845 ;
      RECT 288.27 -291.655 288.6 -291.325 ;
      RECT 288.285 -341.56 288.585 -291.325 ;
      RECT 288.27 -265.71 288.6 -265.38 ;
      RECT 288.285 -280.68 288.585 -265.38 ;
      RECT 288.27 -280.68 288.6 -280.35 ;
      RECT 288.285 -261.485 288.585 -222.48 ;
      RECT 288.27 -222.855 288.6 -222.525 ;
      RECT 288.27 -261.485 288.6 -261.155 ;
      RECT 280.115 -265.25 280.445 -264.92 ;
      RECT 280.13 -280.68 280.43 -264.92 ;
      RECT 280.115 -280.68 280.445 -280.35 ;
      RECT 280.13 -261.465 280.43 -222.48 ;
      RECT 280.115 -224.455 280.445 -224.125 ;
      RECT 280.115 -261.055 280.445 -260.725 ;
      RECT 279.515 -304.57 279.815 -231.5 ;
      RECT 279.5 -231.875 279.83 -231.545 ;
      RECT 279.5 -248.835 279.83 -248.505 ;
      RECT 279.5 -304.57 279.83 -304.24 ;
      RECT 278.9 -244.175 279.2 -232.13 ;
      RECT 278.885 -232.505 279.215 -232.175 ;
      RECT 278.885 -244.175 279.215 -243.845 ;
      RECT 278.27 -291.655 278.6 -291.325 ;
      RECT 278.285 -341.56 278.585 -291.325 ;
      RECT 278.27 -265.71 278.6 -265.38 ;
      RECT 278.285 -280.68 278.585 -265.38 ;
      RECT 278.27 -280.68 278.6 -280.35 ;
      RECT 278.285 -261.485 278.585 -222.48 ;
      RECT 278.27 -222.855 278.6 -222.525 ;
      RECT 278.27 -261.485 278.6 -261.155 ;
      RECT 273.245 -297.045 273.575 -296.715 ;
      RECT 273.26 -334.29 273.56 -296.715 ;
      RECT 273.245 -304.285 273.575 -303.955 ;
      RECT 273.245 -334.245 273.575 -333.915 ;
      RECT 272.615 -303.485 272.945 -303.155 ;
      RECT 272.63 -341.56 272.93 -303.155 ;
      RECT 272 -297.845 272.33 -297.515 ;
      RECT 272.015 -341.56 272.315 -297.515 ;
      RECT 270.115 -265.25 270.445 -264.92 ;
      RECT 270.13 -280.68 270.43 -264.92 ;
      RECT 270.115 -280.68 270.445 -280.35 ;
      RECT 270.13 -261.465 270.43 -222.48 ;
      RECT 270.115 -224.455 270.445 -224.125 ;
      RECT 270.115 -261.055 270.445 -260.725 ;
      RECT 269.515 -296.56 269.815 -231.5 ;
      RECT 269.5 -231.875 269.83 -231.545 ;
      RECT 269.5 -248.835 269.83 -248.505 ;
      RECT 269.5 -296.56 269.83 -296.23 ;
      RECT 268.9 -244.175 269.2 -232.13 ;
      RECT 268.885 -232.505 269.215 -232.175 ;
      RECT 268.885 -244.175 269.215 -243.845 ;
      RECT 268.27 -291.655 268.6 -291.325 ;
      RECT 268.285 -341.56 268.585 -291.325 ;
      RECT 268.27 -265.71 268.6 -265.38 ;
      RECT 268.285 -280.68 268.585 -265.38 ;
      RECT 268.27 -280.68 268.6 -280.35 ;
      RECT 268.285 -261.485 268.585 -222.48 ;
      RECT 268.27 -222.855 268.6 -222.525 ;
      RECT 268.27 -261.485 268.6 -261.155 ;
      RECT 261.3 -313.41 261.6 -236.225 ;
      RECT 261.285 -236.6 261.615 -236.27 ;
      RECT 261.285 -313.41 261.615 -313.08 ;
      RECT 260.115 -265.25 260.445 -264.92 ;
      RECT 260.13 -280.68 260.43 -264.92 ;
      RECT 260.115 -280.68 260.445 -280.35 ;
      RECT 260.13 -261.465 260.43 -222.48 ;
      RECT 260.115 -224.455 260.445 -224.125 ;
      RECT 260.115 -261.055 260.445 -260.725 ;
      RECT 259.515 -304.57 259.815 -231.5 ;
      RECT 259.5 -231.875 259.83 -231.545 ;
      RECT 259.5 -248.835 259.83 -248.505 ;
      RECT 259.5 -304.57 259.83 -304.24 ;
      RECT 258.9 -244.175 259.2 -232.13 ;
      RECT 258.885 -232.505 259.215 -232.175 ;
      RECT 258.885 -244.175 259.215 -243.845 ;
      RECT 258.27 -291.655 258.6 -291.325 ;
      RECT 258.285 -341.56 258.585 -291.325 ;
      RECT 258.27 -265.71 258.6 -265.38 ;
      RECT 258.285 -280.68 258.585 -265.38 ;
      RECT 258.27 -280.68 258.6 -280.35 ;
      RECT 258.285 -261.485 258.585 -222.48 ;
      RECT 258.27 -222.855 258.6 -222.525 ;
      RECT 258.27 -261.485 258.6 -261.155 ;
      RECT 254.11 -313.785 254.44 -313.455 ;
      RECT 254.125 -341.56 254.425 -313.455 ;
      RECT 253.245 -297.045 253.575 -296.715 ;
      RECT 253.26 -334.29 253.56 -296.715 ;
      RECT 253.245 -304.285 253.575 -303.955 ;
      RECT 253.245 -312.985 253.575 -312.655 ;
      RECT 253.245 -334.245 253.575 -333.915 ;
      RECT 252.615 -303.485 252.945 -303.155 ;
      RECT 252.63 -341.56 252.93 -303.155 ;
      RECT 252 -297.845 252.33 -297.515 ;
      RECT 252.015 -341.56 252.315 -297.515 ;
      RECT 250.115 -265.25 250.445 -264.92 ;
      RECT 250.13 -280.68 250.43 -264.92 ;
      RECT 250.115 -280.68 250.445 -280.35 ;
      RECT 250.13 -261.465 250.43 -222.48 ;
      RECT 250.115 -224.455 250.445 -224.125 ;
      RECT 250.115 -261.055 250.445 -260.725 ;
      RECT 249.515 -296.56 249.815 -231.5 ;
      RECT 249.5 -231.875 249.83 -231.545 ;
      RECT 249.5 -248.835 249.83 -248.505 ;
      RECT 249.5 -296.56 249.83 -296.23 ;
      RECT 248.9 -244.175 249.2 -232.13 ;
      RECT 248.885 -232.505 249.215 -232.175 ;
      RECT 248.885 -244.175 249.215 -243.845 ;
      RECT 248.27 -291.655 248.6 -291.325 ;
      RECT 248.285 -341.56 248.585 -291.325 ;
      RECT 248.27 -265.71 248.6 -265.38 ;
      RECT 248.285 -280.68 248.585 -265.38 ;
      RECT 248.27 -280.68 248.6 -280.35 ;
      RECT 248.285 -261.485 248.585 -222.48 ;
      RECT 248.27 -222.855 248.6 -222.525 ;
      RECT 248.27 -261.485 248.6 -261.155 ;
      RECT 240.115 -265.25 240.445 -264.92 ;
      RECT 240.13 -280.68 240.43 -264.92 ;
      RECT 240.115 -280.68 240.445 -280.35 ;
      RECT 240.13 -261.465 240.43 -222.48 ;
      RECT 240.115 -224.455 240.445 -224.125 ;
      RECT 240.115 -261.055 240.445 -260.725 ;
      RECT 239.515 -304.57 239.815 -231.5 ;
      RECT 239.5 -231.875 239.83 -231.545 ;
      RECT 239.5 -248.835 239.83 -248.505 ;
      RECT 239.5 -304.57 239.83 -304.24 ;
      RECT 238.9 -244.175 239.2 -232.13 ;
      RECT 238.885 -232.505 239.215 -232.175 ;
      RECT 238.885 -244.175 239.215 -243.845 ;
      RECT 238.27 -291.655 238.6 -291.325 ;
      RECT 238.285 -341.56 238.585 -291.325 ;
      RECT 238.27 -265.71 238.6 -265.38 ;
      RECT 238.285 -280.68 238.585 -265.38 ;
      RECT 238.27 -280.68 238.6 -280.35 ;
      RECT 238.285 -261.485 238.585 -222.48 ;
      RECT 238.27 -222.855 238.6 -222.525 ;
      RECT 238.27 -261.485 238.6 -261.155 ;
      RECT 233.245 -297.045 233.575 -296.715 ;
      RECT 233.26 -334.29 233.56 -296.715 ;
      RECT 233.245 -304.285 233.575 -303.955 ;
      RECT 233.245 -334.245 233.575 -333.915 ;
      RECT 232.615 -303.485 232.945 -303.155 ;
      RECT 232.63 -341.56 232.93 -303.155 ;
      RECT 232 -297.845 232.33 -297.515 ;
      RECT 232.015 -341.56 232.315 -297.515 ;
      RECT 230.115 -265.25 230.445 -264.92 ;
      RECT 230.13 -280.68 230.43 -264.92 ;
      RECT 230.115 -280.68 230.445 -280.35 ;
      RECT 230.13 -261.465 230.43 -222.48 ;
      RECT 230.115 -224.455 230.445 -224.125 ;
      RECT 230.115 -261.055 230.445 -260.725 ;
      RECT 229.515 -296.56 229.815 -231.5 ;
      RECT 229.5 -231.875 229.83 -231.545 ;
      RECT 229.5 -248.835 229.83 -248.505 ;
      RECT 229.5 -296.56 229.83 -296.23 ;
      RECT 228.9 -244.175 229.2 -232.13 ;
      RECT 228.885 -232.505 229.215 -232.175 ;
      RECT 228.885 -244.175 229.215 -243.845 ;
      RECT 228.27 -291.655 228.6 -291.325 ;
      RECT 228.285 -341.56 228.585 -291.325 ;
      RECT 228.27 -265.71 228.6 -265.38 ;
      RECT 228.285 -280.68 228.585 -265.38 ;
      RECT 228.27 -280.68 228.6 -280.35 ;
      RECT 228.285 -261.485 228.585 -222.48 ;
      RECT 228.27 -222.855 228.6 -222.525 ;
      RECT 228.27 -261.485 228.6 -261.155 ;
      RECT 220.115 -265.25 220.445 -264.92 ;
      RECT 220.13 -280.68 220.43 -264.92 ;
      RECT 220.115 -280.68 220.445 -280.35 ;
      RECT 220.13 -261.465 220.43 -222.48 ;
      RECT 220.115 -224.455 220.445 -224.125 ;
      RECT 220.115 -261.055 220.445 -260.725 ;
      RECT 219.515 -304.57 219.815 -231.5 ;
      RECT 219.5 -231.875 219.83 -231.545 ;
      RECT 219.5 -248.835 219.83 -248.505 ;
      RECT 219.5 -304.57 219.83 -304.24 ;
      RECT 218.9 -244.175 219.2 -232.13 ;
      RECT 218.885 -232.505 219.215 -232.175 ;
      RECT 218.885 -244.175 219.215 -243.845 ;
      RECT 218.27 -291.655 218.6 -291.325 ;
      RECT 218.285 -341.56 218.585 -291.325 ;
      RECT 218.27 -265.71 218.6 -265.38 ;
      RECT 218.285 -280.68 218.585 -265.38 ;
      RECT 218.27 -280.68 218.6 -280.35 ;
      RECT 218.285 -261.485 218.585 -222.48 ;
      RECT 218.27 -222.855 218.6 -222.525 ;
      RECT 218.27 -261.485 218.6 -261.155 ;
      RECT 213.245 -297.045 213.575 -296.715 ;
      RECT 213.26 -334.29 213.56 -296.715 ;
      RECT 213.245 -304.285 213.575 -303.955 ;
      RECT 213.245 -334.245 213.575 -333.915 ;
      RECT 212.615 -303.485 212.945 -303.155 ;
      RECT 212.63 -341.56 212.93 -303.155 ;
      RECT 212 -297.845 212.33 -297.515 ;
      RECT 212.015 -341.56 212.315 -297.515 ;
      RECT 210.115 -265.25 210.445 -264.92 ;
      RECT 210.13 -280.68 210.43 -264.92 ;
      RECT 210.115 -280.68 210.445 -280.35 ;
      RECT 210.13 -261.465 210.43 -222.48 ;
      RECT 210.115 -224.455 210.445 -224.125 ;
      RECT 210.115 -261.055 210.445 -260.725 ;
      RECT 209.515 -296.56 209.815 -231.5 ;
      RECT 209.5 -231.875 209.83 -231.545 ;
      RECT 209.5 -248.835 209.83 -248.505 ;
      RECT 209.5 -296.56 209.83 -296.23 ;
      RECT 208.9 -244.175 209.2 -232.13 ;
      RECT 208.885 -232.505 209.215 -232.175 ;
      RECT 208.885 -244.175 209.215 -243.845 ;
      RECT 208.27 -291.655 208.6 -291.325 ;
      RECT 208.285 -341.56 208.585 -291.325 ;
      RECT 208.27 -265.71 208.6 -265.38 ;
      RECT 208.285 -280.68 208.585 -265.38 ;
      RECT 208.27 -280.68 208.6 -280.35 ;
      RECT 208.285 -261.485 208.585 -222.48 ;
      RECT 208.27 -222.855 208.6 -222.525 ;
      RECT 208.27 -261.485 208.6 -261.155 ;
      RECT 200.115 -265.25 200.445 -264.92 ;
      RECT 200.13 -280.68 200.43 -264.92 ;
      RECT 200.115 -280.68 200.445 -280.35 ;
      RECT 200.13 -261.465 200.43 -222.48 ;
      RECT 200.115 -224.455 200.445 -224.125 ;
      RECT 200.115 -261.055 200.445 -260.725 ;
      RECT 199.515 -304.57 199.815 -231.5 ;
      RECT 199.5 -231.875 199.83 -231.545 ;
      RECT 199.5 -248.835 199.83 -248.505 ;
      RECT 199.5 -304.57 199.83 -304.24 ;
      RECT 198.9 -244.175 199.2 -232.13 ;
      RECT 198.885 -232.505 199.215 -232.175 ;
      RECT 198.885 -244.175 199.215 -243.845 ;
      RECT 198.27 -291.655 198.6 -291.325 ;
      RECT 198.285 -341.56 198.585 -291.325 ;
      RECT 198.27 -265.71 198.6 -265.38 ;
      RECT 198.285 -280.68 198.585 -265.38 ;
      RECT 198.27 -280.68 198.6 -280.35 ;
      RECT 198.285 -261.485 198.585 -222.48 ;
      RECT 198.27 -222.855 198.6 -222.525 ;
      RECT 198.27 -261.485 198.6 -261.155 ;
      RECT 193.245 -297.045 193.575 -296.715 ;
      RECT 193.26 -334.29 193.56 -296.715 ;
      RECT 193.245 -304.285 193.575 -303.955 ;
      RECT 193.245 -334.245 193.575 -333.915 ;
      RECT 192.615 -303.485 192.945 -303.155 ;
      RECT 192.63 -341.56 192.93 -303.155 ;
      RECT 192 -297.845 192.33 -297.515 ;
      RECT 192.015 -341.56 192.315 -297.515 ;
      RECT 190.115 -265.25 190.445 -264.92 ;
      RECT 190.13 -280.68 190.43 -264.92 ;
      RECT 190.115 -280.68 190.445 -280.35 ;
      RECT 190.13 -261.465 190.43 -222.48 ;
      RECT 190.115 -224.455 190.445 -224.125 ;
      RECT 190.115 -261.055 190.445 -260.725 ;
      RECT 189.515 -296.56 189.815 -231.5 ;
      RECT 189.5 -231.875 189.83 -231.545 ;
      RECT 189.5 -248.835 189.83 -248.505 ;
      RECT 189.5 -296.56 189.83 -296.23 ;
      RECT 188.9 -244.175 189.2 -232.13 ;
      RECT 188.885 -232.505 189.215 -232.175 ;
      RECT 188.885 -244.175 189.215 -243.845 ;
      RECT 188.27 -291.655 188.6 -291.325 ;
      RECT 188.285 -341.56 188.585 -291.325 ;
      RECT 188.27 -265.71 188.6 -265.38 ;
      RECT 188.285 -280.68 188.585 -265.38 ;
      RECT 188.27 -280.68 188.6 -280.35 ;
      RECT 188.285 -261.485 188.585 -222.48 ;
      RECT 188.27 -222.855 188.6 -222.525 ;
      RECT 188.27 -261.485 188.6 -261.155 ;
      RECT 181.3 -313.41 181.6 -236.225 ;
      RECT 181.285 -236.6 181.615 -236.27 ;
      RECT 181.285 -313.41 181.615 -313.08 ;
      RECT 180.115 -265.25 180.445 -264.92 ;
      RECT 180.13 -280.68 180.43 -264.92 ;
      RECT 180.115 -280.68 180.445 -280.35 ;
      RECT 180.13 -261.465 180.43 -222.48 ;
      RECT 180.115 -224.455 180.445 -224.125 ;
      RECT 180.115 -261.055 180.445 -260.725 ;
      RECT 179.515 -304.57 179.815 -231.5 ;
      RECT 179.5 -231.875 179.83 -231.545 ;
      RECT 179.5 -248.835 179.83 -248.505 ;
      RECT 179.5 -304.57 179.83 -304.24 ;
      RECT 178.9 -244.175 179.2 -232.13 ;
      RECT 178.885 -232.505 179.215 -232.175 ;
      RECT 178.885 -244.175 179.215 -243.845 ;
      RECT 178.27 -291.655 178.6 -291.325 ;
      RECT 178.285 -341.56 178.585 -291.325 ;
      RECT 178.27 -265.71 178.6 -265.38 ;
      RECT 178.285 -280.68 178.585 -265.38 ;
      RECT 178.27 -280.68 178.6 -280.35 ;
      RECT 178.285 -261.485 178.585 -222.48 ;
      RECT 178.27 -222.855 178.6 -222.525 ;
      RECT 178.27 -261.485 178.6 -261.155 ;
      RECT 174.11 -313.785 174.44 -313.455 ;
      RECT 174.125 -341.56 174.425 -313.455 ;
      RECT 173.245 -297.045 173.575 -296.715 ;
      RECT 173.26 -334.29 173.56 -296.715 ;
      RECT 173.245 -304.285 173.575 -303.955 ;
      RECT 173.245 -312.985 173.575 -312.655 ;
      RECT 173.245 -334.245 173.575 -333.915 ;
      RECT 172.615 -303.485 172.945 -303.155 ;
      RECT 172.63 -341.56 172.93 -303.155 ;
      RECT 172 -297.845 172.33 -297.515 ;
      RECT 172.015 -341.56 172.315 -297.515 ;
      RECT 170.115 -265.25 170.445 -264.92 ;
      RECT 170.13 -280.68 170.43 -264.92 ;
      RECT 170.115 -280.68 170.445 -280.35 ;
      RECT 170.13 -261.465 170.43 -222.48 ;
      RECT 170.115 -224.455 170.445 -224.125 ;
      RECT 170.115 -261.055 170.445 -260.725 ;
      RECT 169.515 -296.56 169.815 -231.5 ;
      RECT 169.5 -231.875 169.83 -231.545 ;
      RECT 169.5 -248.835 169.83 -248.505 ;
      RECT 169.5 -296.56 169.83 -296.23 ;
      RECT 168.9 -244.175 169.2 -232.13 ;
      RECT 168.885 -232.505 169.215 -232.175 ;
      RECT 168.885 -244.175 169.215 -243.845 ;
      RECT 168.27 -291.655 168.6 -291.325 ;
      RECT 168.285 -341.56 168.585 -291.325 ;
      RECT 168.27 -265.71 168.6 -265.38 ;
      RECT 168.285 -280.68 168.585 -265.38 ;
      RECT 168.27 -280.68 168.6 -280.35 ;
      RECT 168.285 -261.485 168.585 -222.48 ;
      RECT 168.27 -222.855 168.6 -222.525 ;
      RECT 168.27 -261.485 168.6 -261.155 ;
      RECT 160.115 -265.25 160.445 -264.92 ;
      RECT 160.13 -280.68 160.43 -264.92 ;
      RECT 160.115 -280.68 160.445 -280.35 ;
      RECT 160.13 -261.465 160.43 -222.48 ;
      RECT 160.115 -224.455 160.445 -224.125 ;
      RECT 160.115 -261.055 160.445 -260.725 ;
      RECT 159.515 -304.57 159.815 -231.5 ;
      RECT 159.5 -231.875 159.83 -231.545 ;
      RECT 159.5 -248.835 159.83 -248.505 ;
      RECT 159.5 -304.57 159.83 -304.24 ;
      RECT 158.9 -244.175 159.2 -232.13 ;
      RECT 158.885 -232.505 159.215 -232.175 ;
      RECT 158.885 -244.175 159.215 -243.845 ;
      RECT 158.27 -291.655 158.6 -291.325 ;
      RECT 158.285 -341.56 158.585 -291.325 ;
      RECT 158.27 -265.71 158.6 -265.38 ;
      RECT 158.285 -280.68 158.585 -265.38 ;
      RECT 158.27 -280.68 158.6 -280.35 ;
      RECT 158.285 -261.485 158.585 -222.48 ;
      RECT 158.27 -222.855 158.6 -222.525 ;
      RECT 158.27 -261.485 158.6 -261.155 ;
      RECT 153.245 -297.045 153.575 -296.715 ;
      RECT 153.26 -334.29 153.56 -296.715 ;
      RECT 153.245 -304.285 153.575 -303.955 ;
      RECT 153.245 -334.245 153.575 -333.915 ;
      RECT 152.615 -303.485 152.945 -303.155 ;
      RECT 152.63 -341.56 152.93 -303.155 ;
      RECT 152 -297.845 152.33 -297.515 ;
      RECT 152.015 -341.56 152.315 -297.515 ;
      RECT 150.115 -265.25 150.445 -264.92 ;
      RECT 150.13 -280.68 150.43 -264.92 ;
      RECT 150.115 -280.68 150.445 -280.35 ;
      RECT 150.13 -261.465 150.43 -222.48 ;
      RECT 150.115 -224.455 150.445 -224.125 ;
      RECT 150.115 -261.055 150.445 -260.725 ;
      RECT 149.515 -296.56 149.815 -231.5 ;
      RECT 149.5 -231.875 149.83 -231.545 ;
      RECT 149.5 -248.835 149.83 -248.505 ;
      RECT 149.5 -296.56 149.83 -296.23 ;
      RECT 148.9 -244.175 149.2 -232.13 ;
      RECT 148.885 -232.505 149.215 -232.175 ;
      RECT 148.885 -244.175 149.215 -243.845 ;
      RECT 148.27 -291.655 148.6 -291.325 ;
      RECT 148.285 -341.56 148.585 -291.325 ;
      RECT 148.27 -265.71 148.6 -265.38 ;
      RECT 148.285 -280.68 148.585 -265.38 ;
      RECT 148.27 -280.68 148.6 -280.35 ;
      RECT 148.285 -261.485 148.585 -222.48 ;
      RECT 148.27 -222.855 148.6 -222.525 ;
      RECT 148.27 -261.485 148.6 -261.155 ;
      RECT 140.115 -265.25 140.445 -264.92 ;
      RECT 140.13 -280.68 140.43 -264.92 ;
      RECT 140.115 -280.68 140.445 -280.35 ;
      RECT 140.13 -261.465 140.43 -222.48 ;
      RECT 140.115 -224.455 140.445 -224.125 ;
      RECT 140.115 -261.055 140.445 -260.725 ;
      RECT 139.515 -304.57 139.815 -231.5 ;
      RECT 139.5 -231.875 139.83 -231.545 ;
      RECT 139.5 -248.835 139.83 -248.505 ;
      RECT 139.5 -304.57 139.83 -304.24 ;
      RECT 138.9 -244.175 139.2 -232.13 ;
      RECT 138.885 -232.505 139.215 -232.175 ;
      RECT 138.885 -244.175 139.215 -243.845 ;
      RECT 138.27 -291.655 138.6 -291.325 ;
      RECT 138.285 -341.56 138.585 -291.325 ;
      RECT 138.27 -265.71 138.6 -265.38 ;
      RECT 138.285 -280.68 138.585 -265.38 ;
      RECT 138.27 -280.68 138.6 -280.35 ;
      RECT 138.285 -261.485 138.585 -222.48 ;
      RECT 138.27 -222.855 138.6 -222.525 ;
      RECT 138.27 -261.485 138.6 -261.155 ;
      RECT 133.245 -297.045 133.575 -296.715 ;
      RECT 133.26 -334.29 133.56 -296.715 ;
      RECT 133.245 -304.285 133.575 -303.955 ;
      RECT 133.245 -334.245 133.575 -333.915 ;
      RECT 132.615 -303.485 132.945 -303.155 ;
      RECT 132.63 -341.56 132.93 -303.155 ;
      RECT 132 -297.845 132.33 -297.515 ;
      RECT 132.015 -341.56 132.315 -297.515 ;
      RECT 130.115 -265.25 130.445 -264.92 ;
      RECT 130.13 -280.68 130.43 -264.92 ;
      RECT 130.115 -280.68 130.445 -280.35 ;
      RECT 130.13 -261.465 130.43 -222.48 ;
      RECT 130.115 -224.455 130.445 -224.125 ;
      RECT 130.115 -261.055 130.445 -260.725 ;
      RECT 129.515 -296.56 129.815 -231.5 ;
      RECT 129.5 -231.875 129.83 -231.545 ;
      RECT 129.5 -248.835 129.83 -248.505 ;
      RECT 129.5 -296.56 129.83 -296.23 ;
      RECT 128.9 -244.175 129.2 -232.13 ;
      RECT 128.885 -232.505 129.215 -232.175 ;
      RECT 128.885 -244.175 129.215 -243.845 ;
      RECT 128.27 -291.655 128.6 -291.325 ;
      RECT 128.285 -341.56 128.585 -291.325 ;
      RECT 128.27 -265.71 128.6 -265.38 ;
      RECT 128.285 -280.68 128.585 -265.38 ;
      RECT 128.27 -280.68 128.6 -280.35 ;
      RECT 128.285 -261.485 128.585 -222.48 ;
      RECT 128.27 -222.855 128.6 -222.525 ;
      RECT 128.27 -261.485 128.6 -261.155 ;
      RECT 120.115 -265.25 120.445 -264.92 ;
      RECT 120.13 -280.68 120.43 -264.92 ;
      RECT 120.115 -280.68 120.445 -280.35 ;
      RECT 120.13 -261.465 120.43 -222.48 ;
      RECT 120.115 -224.455 120.445 -224.125 ;
      RECT 120.115 -261.055 120.445 -260.725 ;
      RECT 119.515 -304.57 119.815 -231.5 ;
      RECT 119.5 -231.875 119.83 -231.545 ;
      RECT 119.5 -248.835 119.83 -248.505 ;
      RECT 119.5 -304.57 119.83 -304.24 ;
      RECT 118.9 -244.175 119.2 -232.13 ;
      RECT 118.885 -232.505 119.215 -232.175 ;
      RECT 118.885 -244.175 119.215 -243.845 ;
      RECT 118.27 -291.655 118.6 -291.325 ;
      RECT 118.285 -341.56 118.585 -291.325 ;
      RECT 118.27 -265.71 118.6 -265.38 ;
      RECT 118.285 -280.68 118.585 -265.38 ;
      RECT 118.27 -280.68 118.6 -280.35 ;
      RECT 118.285 -261.485 118.585 -222.48 ;
      RECT 118.27 -222.855 118.6 -222.525 ;
      RECT 118.27 -261.485 118.6 -261.155 ;
      RECT 113.245 -297.045 113.575 -296.715 ;
      RECT 113.26 -334.29 113.56 -296.715 ;
      RECT 113.245 -304.285 113.575 -303.955 ;
      RECT 113.245 -334.245 113.575 -333.915 ;
      RECT 112.615 -303.485 112.945 -303.155 ;
      RECT 112.63 -341.56 112.93 -303.155 ;
      RECT 112 -297.845 112.33 -297.515 ;
      RECT 112.015 -341.56 112.315 -297.515 ;
      RECT 110.115 -265.25 110.445 -264.92 ;
      RECT 110.13 -280.68 110.43 -264.92 ;
      RECT 110.115 -280.68 110.445 -280.35 ;
      RECT 110.13 -261.465 110.43 -222.48 ;
      RECT 110.115 -224.455 110.445 -224.125 ;
      RECT 110.115 -261.055 110.445 -260.725 ;
      RECT 109.515 -296.56 109.815 -231.5 ;
      RECT 109.5 -231.875 109.83 -231.545 ;
      RECT 109.5 -248.835 109.83 -248.505 ;
      RECT 109.5 -296.56 109.83 -296.23 ;
      RECT 108.9 -244.175 109.2 -232.13 ;
      RECT 108.885 -232.505 109.215 -232.175 ;
      RECT 108.885 -244.175 109.215 -243.845 ;
      RECT 108.27 -291.655 108.6 -291.325 ;
      RECT 108.285 -341.56 108.585 -291.325 ;
      RECT 108.27 -265.71 108.6 -265.38 ;
      RECT 108.285 -280.68 108.585 -265.38 ;
      RECT 108.27 -280.68 108.6 -280.35 ;
      RECT 108.285 -261.485 108.585 -222.48 ;
      RECT 108.27 -222.855 108.6 -222.525 ;
      RECT 108.27 -261.485 108.6 -261.155 ;
      RECT 101.3 -313.41 101.6 -236.225 ;
      RECT 101.285 -236.6 101.615 -236.27 ;
      RECT 101.285 -313.41 101.615 -313.08 ;
      RECT 100.115 -265.25 100.445 -264.92 ;
      RECT 100.13 -280.68 100.43 -264.92 ;
      RECT 100.115 -280.68 100.445 -280.35 ;
      RECT 100.13 -261.465 100.43 -222.48 ;
      RECT 100.115 -224.455 100.445 -224.125 ;
      RECT 100.115 -261.055 100.445 -260.725 ;
      RECT 99.515 -304.57 99.815 -231.5 ;
      RECT 99.5 -231.875 99.83 -231.545 ;
      RECT 99.5 -248.835 99.83 -248.505 ;
      RECT 99.5 -304.57 99.83 -304.24 ;
      RECT 98.9 -244.175 99.2 -232.13 ;
      RECT 98.885 -232.505 99.215 -232.175 ;
      RECT 98.885 -244.175 99.215 -243.845 ;
      RECT 98.27 -291.655 98.6 -291.325 ;
      RECT 98.285 -341.56 98.585 -291.325 ;
      RECT 98.27 -265.71 98.6 -265.38 ;
      RECT 98.285 -280.68 98.585 -265.38 ;
      RECT 98.27 -280.68 98.6 -280.35 ;
      RECT 98.285 -261.485 98.585 -222.48 ;
      RECT 98.27 -222.855 98.6 -222.525 ;
      RECT 98.27 -261.485 98.6 -261.155 ;
      RECT 94.11 -313.785 94.44 -313.455 ;
      RECT 94.125 -341.56 94.425 -313.455 ;
      RECT 93.245 -297.045 93.575 -296.715 ;
      RECT 93.26 -334.29 93.56 -296.715 ;
      RECT 93.245 -304.285 93.575 -303.955 ;
      RECT 93.245 -312.985 93.575 -312.655 ;
      RECT 93.245 -334.245 93.575 -333.915 ;
      RECT 92.615 -303.485 92.945 -303.155 ;
      RECT 92.63 -341.56 92.93 -303.155 ;
      RECT 92 -297.845 92.33 -297.515 ;
      RECT 92.015 -341.56 92.315 -297.515 ;
      RECT 90.115 -265.25 90.445 -264.92 ;
      RECT 90.13 -280.68 90.43 -264.92 ;
      RECT 90.115 -280.68 90.445 -280.35 ;
      RECT 90.13 -261.465 90.43 -222.48 ;
      RECT 90.115 -224.455 90.445 -224.125 ;
      RECT 90.115 -261.055 90.445 -260.725 ;
      RECT 89.515 -296.56 89.815 -231.5 ;
      RECT 89.5 -231.875 89.83 -231.545 ;
      RECT 89.5 -248.835 89.83 -248.505 ;
      RECT 89.5 -296.56 89.83 -296.23 ;
      RECT 88.9 -244.175 89.2 -232.13 ;
      RECT 88.885 -232.505 89.215 -232.175 ;
      RECT 88.885 -244.175 89.215 -243.845 ;
      RECT 88.27 -291.655 88.6 -291.325 ;
      RECT 88.285 -341.56 88.585 -291.325 ;
      RECT 88.27 -265.71 88.6 -265.38 ;
      RECT 88.285 -280.68 88.585 -265.38 ;
      RECT 88.27 -280.68 88.6 -280.35 ;
      RECT 88.285 -261.485 88.585 -222.48 ;
      RECT 88.27 -222.855 88.6 -222.525 ;
      RECT 88.27 -261.485 88.6 -261.155 ;
      RECT 80.115 -265.25 80.445 -264.92 ;
      RECT 80.13 -280.68 80.43 -264.92 ;
      RECT 80.115 -280.68 80.445 -280.35 ;
      RECT 80.13 -261.465 80.43 -222.48 ;
      RECT 80.115 -224.455 80.445 -224.125 ;
      RECT 80.115 -261.055 80.445 -260.725 ;
      RECT 79.515 -304.57 79.815 -231.5 ;
      RECT 79.5 -231.875 79.83 -231.545 ;
      RECT 79.5 -248.835 79.83 -248.505 ;
      RECT 79.5 -304.57 79.83 -304.24 ;
      RECT 78.9 -244.175 79.2 -232.13 ;
      RECT 78.885 -232.505 79.215 -232.175 ;
      RECT 78.885 -244.175 79.215 -243.845 ;
      RECT 78.27 -291.655 78.6 -291.325 ;
      RECT 78.285 -341.56 78.585 -291.325 ;
      RECT 78.27 -265.71 78.6 -265.38 ;
      RECT 78.285 -280.68 78.585 -265.38 ;
      RECT 78.27 -280.68 78.6 -280.35 ;
      RECT 78.285 -261.485 78.585 -222.48 ;
      RECT 78.27 -222.855 78.6 -222.525 ;
      RECT 78.27 -261.485 78.6 -261.155 ;
      RECT 73.245 -297.045 73.575 -296.715 ;
      RECT 73.26 -334.29 73.56 -296.715 ;
      RECT 73.245 -304.285 73.575 -303.955 ;
      RECT 73.245 -334.245 73.575 -333.915 ;
      RECT 72.615 -303.485 72.945 -303.155 ;
      RECT 72.63 -341.56 72.93 -303.155 ;
      RECT 72 -297.845 72.33 -297.515 ;
      RECT 72.015 -341.56 72.315 -297.515 ;
      RECT 70.115 -265.25 70.445 -264.92 ;
      RECT 70.13 -280.68 70.43 -264.92 ;
      RECT 70.115 -280.68 70.445 -280.35 ;
      RECT 70.13 -261.465 70.43 -222.48 ;
      RECT 70.115 -224.455 70.445 -224.125 ;
      RECT 70.115 -261.055 70.445 -260.725 ;
      RECT 69.515 -296.56 69.815 -231.5 ;
      RECT 69.5 -231.875 69.83 -231.545 ;
      RECT 69.5 -248.835 69.83 -248.505 ;
      RECT 69.5 -296.56 69.83 -296.23 ;
      RECT 68.9 -244.175 69.2 -232.13 ;
      RECT 68.885 -232.505 69.215 -232.175 ;
      RECT 68.885 -244.175 69.215 -243.845 ;
      RECT 68.27 -291.655 68.6 -291.325 ;
      RECT 68.285 -341.56 68.585 -291.325 ;
      RECT 68.27 -265.71 68.6 -265.38 ;
      RECT 68.285 -280.68 68.585 -265.38 ;
      RECT 68.27 -280.68 68.6 -280.35 ;
      RECT 68.285 -261.485 68.585 -222.48 ;
      RECT 68.27 -222.855 68.6 -222.525 ;
      RECT 68.27 -261.485 68.6 -261.155 ;
      RECT 60.115 -265.25 60.445 -264.92 ;
      RECT 60.13 -280.68 60.43 -264.92 ;
      RECT 60.115 -280.68 60.445 -280.35 ;
      RECT 60.13 -261.465 60.43 -222.48 ;
      RECT 60.115 -224.455 60.445 -224.125 ;
      RECT 60.115 -261.055 60.445 -260.725 ;
      RECT 59.515 -304.57 59.815 -231.5 ;
      RECT 59.5 -231.875 59.83 -231.545 ;
      RECT 59.5 -248.835 59.83 -248.505 ;
      RECT 59.5 -304.57 59.83 -304.24 ;
      RECT 58.9 -244.175 59.2 -232.13 ;
      RECT 58.885 -232.505 59.215 -232.175 ;
      RECT 58.885 -244.175 59.215 -243.845 ;
      RECT 58.27 -291.655 58.6 -291.325 ;
      RECT 58.285 -341.56 58.585 -291.325 ;
      RECT 58.27 -265.71 58.6 -265.38 ;
      RECT 58.285 -280.68 58.585 -265.38 ;
      RECT 58.27 -280.68 58.6 -280.35 ;
      RECT 58.285 -261.485 58.585 -222.48 ;
      RECT 58.27 -222.855 58.6 -222.525 ;
      RECT 58.27 -261.485 58.6 -261.155 ;
      RECT 53.245 -297.045 53.575 -296.715 ;
      RECT 53.26 -334.29 53.56 -296.715 ;
      RECT 53.245 -304.285 53.575 -303.955 ;
      RECT 53.245 -334.245 53.575 -333.915 ;
      RECT 52.615 -303.485 52.945 -303.155 ;
      RECT 52.63 -341.56 52.93 -303.155 ;
      RECT 52 -297.845 52.33 -297.515 ;
      RECT 52.015 -341.56 52.315 -297.515 ;
      RECT 50.115 -265.25 50.445 -264.92 ;
      RECT 50.13 -280.68 50.43 -264.92 ;
      RECT 50.115 -280.68 50.445 -280.35 ;
      RECT 50.13 -261.465 50.43 -222.48 ;
      RECT 50.115 -224.455 50.445 -224.125 ;
      RECT 50.115 -261.055 50.445 -260.725 ;
      RECT 49.515 -296.56 49.815 -231.5 ;
      RECT 49.5 -231.875 49.83 -231.545 ;
      RECT 49.5 -248.835 49.83 -248.505 ;
      RECT 49.5 -296.56 49.83 -296.23 ;
      RECT 48.9 -244.175 49.2 -232.13 ;
      RECT 48.885 -232.505 49.215 -232.175 ;
      RECT 48.885 -244.175 49.215 -243.845 ;
      RECT 48.27 -291.655 48.6 -291.325 ;
      RECT 48.285 -341.56 48.585 -291.325 ;
      RECT 48.27 -265.71 48.6 -265.38 ;
      RECT 48.285 -280.68 48.585 -265.38 ;
      RECT 48.27 -280.68 48.6 -280.35 ;
      RECT 48.285 -261.485 48.585 -222.48 ;
      RECT 48.27 -222.855 48.6 -222.525 ;
      RECT 48.27 -261.485 48.6 -261.155 ;
      RECT 40.115 -265.25 40.445 -264.92 ;
      RECT 40.13 -280.68 40.43 -264.92 ;
      RECT 40.115 -280.68 40.445 -280.35 ;
      RECT 40.13 -261.465 40.43 -222.48 ;
      RECT 40.115 -224.455 40.445 -224.125 ;
      RECT 40.115 -261.055 40.445 -260.725 ;
      RECT 39.515 -304.57 39.815 -231.5 ;
      RECT 39.5 -231.875 39.83 -231.545 ;
      RECT 39.5 -248.835 39.83 -248.505 ;
      RECT 39.5 -304.57 39.83 -304.24 ;
      RECT 38.9 -244.175 39.2 -232.13 ;
      RECT 38.885 -232.505 39.215 -232.175 ;
      RECT 38.885 -244.175 39.215 -243.845 ;
      RECT 38.27 -291.655 38.6 -291.325 ;
      RECT 38.285 -341.56 38.585 -291.325 ;
      RECT 38.27 -265.71 38.6 -265.38 ;
      RECT 38.285 -280.68 38.585 -265.38 ;
      RECT 38.27 -280.68 38.6 -280.35 ;
      RECT 38.285 -261.485 38.585 -222.48 ;
      RECT 38.27 -222.855 38.6 -222.525 ;
      RECT 38.27 -261.485 38.6 -261.155 ;
      RECT 33.245 -297.045 33.575 -296.715 ;
      RECT 33.26 -334.29 33.56 -296.715 ;
      RECT 33.245 -304.285 33.575 -303.955 ;
      RECT 33.245 -334.245 33.575 -333.915 ;
      RECT 32.615 -303.485 32.945 -303.155 ;
      RECT 32.63 -341.56 32.93 -303.155 ;
      RECT 32 -297.845 32.33 -297.515 ;
      RECT 32.015 -341.56 32.315 -297.515 ;
      RECT 30.115 -265.25 30.445 -264.92 ;
      RECT 30.13 -280.68 30.43 -264.92 ;
      RECT 30.115 -280.68 30.445 -280.35 ;
      RECT 30.13 -261.465 30.43 -222.48 ;
      RECT 30.115 -224.455 30.445 -224.125 ;
      RECT 30.115 -261.055 30.445 -260.725 ;
      RECT 29.515 -296.56 29.815 -231.5 ;
      RECT 29.5 -231.875 29.83 -231.545 ;
      RECT 29.5 -248.835 29.83 -248.505 ;
      RECT 29.5 -296.56 29.83 -296.23 ;
      RECT 28.9 -244.175 29.2 -232.13 ;
      RECT 28.885 -232.505 29.215 -232.175 ;
      RECT 28.885 -244.175 29.215 -243.845 ;
      RECT 28.27 -291.655 28.6 -291.325 ;
      RECT 28.285 -341.56 28.585 -291.325 ;
      RECT 28.27 -265.71 28.6 -265.38 ;
      RECT 28.285 -280.68 28.585 -265.38 ;
      RECT 28.27 -280.68 28.6 -280.35 ;
      RECT 28.285 -261.485 28.585 -222.48 ;
      RECT 28.27 -222.855 28.6 -222.525 ;
      RECT 28.27 -261.485 28.6 -261.155 ;
      RECT 21.3 -313.41 21.6 -236.225 ;
      RECT 21.285 -236.6 21.615 -236.27 ;
      RECT 21.285 -313.41 21.615 -313.08 ;
      RECT 20.115 -265.25 20.445 -264.92 ;
      RECT 20.13 -280.68 20.43 -264.92 ;
      RECT 20.115 -280.68 20.445 -280.35 ;
      RECT 20.13 -261.465 20.43 -222.48 ;
      RECT 20.115 -224.455 20.445 -224.125 ;
      RECT 20.115 -261.055 20.445 -260.725 ;
      RECT 19.515 -304.57 19.815 -231.5 ;
      RECT 19.5 -231.875 19.83 -231.545 ;
      RECT 19.5 -248.835 19.83 -248.505 ;
      RECT 19.5 -304.57 19.83 -304.24 ;
      RECT 18.9 -244.175 19.2 -232.13 ;
      RECT 18.885 -232.505 19.215 -232.175 ;
      RECT 18.885 -244.175 19.215 -243.845 ;
      RECT 18.27 -291.655 18.6 -291.325 ;
      RECT 18.285 -341.56 18.585 -291.325 ;
      RECT 18.27 -265.71 18.6 -265.38 ;
      RECT 18.285 -280.68 18.585 -265.38 ;
      RECT 18.27 -280.68 18.6 -280.35 ;
      RECT 18.285 -261.485 18.585 -222.48 ;
      RECT 18.27 -222.855 18.6 -222.525 ;
      RECT 18.27 -261.485 18.6 -261.155 ;
      RECT 14.11 -313.785 14.44 -313.455 ;
      RECT 14.125 -341.56 14.425 -313.455 ;
      RECT 13.245 -297.045 13.575 -296.715 ;
      RECT 13.26 -334.29 13.56 -296.715 ;
      RECT 13.245 -304.285 13.575 -303.955 ;
      RECT 13.245 -312.985 13.575 -312.655 ;
      RECT 13.245 -334.245 13.575 -333.915 ;
      RECT 12.615 -303.485 12.945 -303.155 ;
      RECT 12.63 -341.56 12.93 -303.155 ;
      RECT 12 -297.845 12.33 -297.515 ;
      RECT 12.015 -341.56 12.315 -297.515 ;
      RECT 10.115 -265.25 10.445 -264.92 ;
      RECT 10.13 -280.68 10.43 -264.92 ;
      RECT 10.115 -280.68 10.445 -280.35 ;
      RECT 10.13 -261.465 10.43 -222.48 ;
      RECT 10.115 -224.455 10.445 -224.125 ;
      RECT 10.115 -261.055 10.445 -260.725 ;
      RECT 9.515 -296.56 9.815 -231.5 ;
      RECT 9.5 -231.875 9.83 -231.545 ;
      RECT 9.5 -248.835 9.83 -248.505 ;
      RECT 9.5 -296.56 9.83 -296.23 ;
      RECT 8.9 -244.175 9.2 -232.13 ;
      RECT 8.885 -232.505 9.215 -232.175 ;
      RECT 8.885 -244.175 9.215 -243.845 ;
      RECT 8.27 -291.655 8.6 -291.325 ;
      RECT 8.285 -341.56 8.585 -291.325 ;
      RECT 8.27 -265.71 8.6 -265.38 ;
      RECT 8.285 -280.68 8.585 -265.38 ;
      RECT 8.27 -280.68 8.6 -280.35 ;
      RECT 8.285 -261.485 8.585 -222.48 ;
      RECT 8.27 -222.855 8.6 -222.525 ;
      RECT 8.27 -261.485 8.6 -261.155 ;
      RECT 6.005 -255.47 6.335 -255.14 ;
      RECT 6.02 -292.36 6.32 -255.14 ;
      RECT 6.005 -292.36 6.335 -292.03 ;
      RECT -5.91 -312.795 -5.58 -312.465 ;
      RECT -5.895 -330.23 -5.595 -312.465 ;
      RECT -5.91 -330.23 -5.58 -329.9 ;
      RECT -9.505 -329.785 -9.175 -329.455 ;
      RECT -9.49 -334.29 -9.19 -329.455 ;
      RECT -9.505 -334.245 -9.175 -333.915 ;
      RECT -10.34 -213.02 -10.01 -212.69 ;
      RECT -10.325 -294.15 -10.025 -212.69 ;
      RECT -10.34 -294.15 -10.01 -293.82 ;
      RECT -10.635 -330.585 -10.305 -330.255 ;
      RECT -10.62 -341.56 -10.32 -330.255 ;
      RECT -11.75 -317.56 -11.42 -317.23 ;
      RECT -11.735 -330.23 -11.435 -317.23 ;
      RECT -11.75 -330.23 -11.42 -329.9 ;
      RECT -12.385 -317.06 -12.055 -316.73 ;
      RECT -12.37 -330.985 -12.07 -316.73 ;
      RECT -12.385 -330.985 -12.055 -330.655 ;
      RECT -15.345 -329.785 -15.015 -329.455 ;
      RECT -15.33 -334.29 -15.03 -329.455 ;
      RECT -15.345 -334.245 -15.015 -333.915 ;
      RECT -16.475 -330.585 -16.145 -330.255 ;
      RECT -16.46 -341.56 -16.16 -330.255 ;
      RECT -17.59 -318.56 -17.26 -318.23 ;
      RECT -17.575 -330.23 -17.275 -318.23 ;
      RECT -17.59 -330.23 -17.26 -329.9 ;
      RECT -18.225 -318.06 -17.895 -317.73 ;
      RECT -18.21 -330.985 -17.91 -317.73 ;
      RECT -18.225 -330.985 -17.895 -330.655 ;
      RECT -21.185 -329.785 -20.855 -329.455 ;
      RECT -21.17 -334.29 -20.87 -329.455 ;
      RECT -21.185 -334.245 -20.855 -333.915 ;
      RECT -22.315 -330.585 -21.985 -330.255 ;
      RECT -22.3 -341.56 -22 -330.255 ;
      RECT -23.43 -319.56 -23.1 -319.23 ;
      RECT -23.415 -330.23 -23.115 -319.23 ;
      RECT -23.43 -330.23 -23.1 -329.9 ;
      RECT -24.065 -319.06 -23.735 -318.73 ;
      RECT -24.05 -330.985 -23.75 -318.73 ;
      RECT -24.065 -330.985 -23.735 -330.655 ;
      RECT -27.025 -329.785 -26.695 -329.455 ;
      RECT -27.01 -334.29 -26.71 -329.455 ;
      RECT -27.025 -334.245 -26.695 -333.915 ;
      RECT -28.155 -330.585 -27.825 -330.255 ;
      RECT -28.14 -341.56 -27.84 -330.255 ;
      RECT -29.27 -320.56 -28.94 -320.23 ;
      RECT -29.255 -330.23 -28.955 -320.23 ;
      RECT -29.27 -330.23 -28.94 -329.9 ;
      RECT -29.905 -320.06 -29.575 -319.73 ;
      RECT -29.89 -330.985 -29.59 -319.73 ;
      RECT -29.905 -330.985 -29.575 -330.655 ;
      RECT -32.865 -329.785 -32.535 -329.455 ;
      RECT -32.85 -334.29 -32.55 -329.455 ;
      RECT -32.865 -334.245 -32.535 -333.915 ;
      RECT -33.995 -330.585 -33.665 -330.255 ;
      RECT -33.98 -341.56 -33.68 -330.255 ;
      RECT -35.11 -321.56 -34.78 -321.23 ;
      RECT -35.095 -330.23 -34.795 -321.23 ;
      RECT -35.11 -330.23 -34.78 -329.9 ;
      RECT -35.745 -321.06 -35.415 -320.73 ;
      RECT -35.73 -330.985 -35.43 -320.73 ;
      RECT -35.745 -330.985 -35.415 -330.655 ;
      RECT -38.705 -329.785 -38.375 -329.455 ;
      RECT -38.69 -334.29 -38.39 -329.455 ;
      RECT -38.705 -334.245 -38.375 -333.915 ;
      RECT -39.835 -330.585 -39.505 -330.255 ;
      RECT -39.82 -341.56 -39.52 -330.255 ;
      RECT -40.95 -322.56 -40.62 -322.23 ;
      RECT -40.935 -330.23 -40.635 -322.23 ;
      RECT -40.95 -330.23 -40.62 -329.9 ;
      RECT -41.585 -322.06 -41.255 -321.73 ;
      RECT -41.57 -330.985 -41.27 -321.73 ;
      RECT -41.585 -330.985 -41.255 -330.655 ;
      RECT -44.545 -329.785 -44.215 -329.455 ;
      RECT -44.53 -334.29 -44.23 -329.455 ;
      RECT -44.545 -334.245 -44.215 -333.915 ;
      RECT -45.675 -330.585 -45.345 -330.255 ;
      RECT -45.66 -341.56 -45.36 -330.255 ;
      RECT -46.79 -323.56 -46.46 -323.23 ;
      RECT -46.775 -330.23 -46.475 -323.23 ;
      RECT -46.79 -330.23 -46.46 -329.9 ;
      RECT -47.425 -323.06 -47.095 -322.73 ;
      RECT -47.41 -330.985 -47.11 -322.73 ;
      RECT -47.425 -330.985 -47.095 -330.655 ;
      RECT -50.385 -329.785 -50.055 -329.455 ;
      RECT -50.37 -334.29 -50.07 -329.455 ;
      RECT -50.385 -334.245 -50.055 -333.915 ;
      RECT -51.515 -330.585 -51.185 -330.255 ;
      RECT -51.5 -341.56 -51.2 -330.255 ;
      RECT -52.63 -324.56 -52.3 -324.23 ;
      RECT -52.615 -330.23 -52.315 -324.23 ;
      RECT -52.63 -330.23 -52.3 -329.9 ;
      RECT -53.265 -324.06 -52.935 -323.73 ;
      RECT -53.25 -330.985 -52.95 -323.73 ;
      RECT -53.265 -330.985 -52.935 -330.655 ;
      RECT -56.225 -329.785 -55.895 -329.455 ;
      RECT -56.21 -334.29 -55.91 -329.455 ;
      RECT -56.225 -334.245 -55.895 -333.915 ;
      RECT -57.355 -330.585 -57.025 -330.255 ;
      RECT -57.34 -341.56 -57.04 -330.255 ;
      RECT -58.47 -325.56 -58.14 -325.23 ;
      RECT -58.455 -330.23 -58.155 -325.23 ;
      RECT -58.47 -330.23 -58.14 -329.9 ;
      RECT -59.105 -325.06 -58.775 -324.73 ;
      RECT -59.09 -330.985 -58.79 -324.73 ;
      RECT -59.105 -330.985 -58.775 -330.655 ;
      RECT -62.065 -329.785 -61.735 -329.455 ;
      RECT -62.05 -334.29 -61.75 -329.455 ;
      RECT -62.065 -334.245 -61.735 -333.915 ;
      RECT -63.195 -330.585 -62.865 -330.255 ;
      RECT -63.18 -341.56 -62.88 -330.255 ;
      RECT -64.06 -334.29 -63.66 -314.105 ;
      RECT -64.2 -341.44 -63.78 -333.87 ;
  END
END sramgen_sram_512x32m4w8_replica_v1

END LIBRARY
