VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_512x32m4w8
    CLASS BLOCK  ;
    FOREIGN sram22_512x32m4w8   ;
    SIZE 443.280 BY 448.720 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 235.030 0.000 235.170 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 241.130 0.000 241.270 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 247.230 0.000 247.370 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 253.330 0.000 253.470 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 259.430 0.000 259.570 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 265.530 0.000 265.670 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 271.630 0.000 271.770 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 277.730 0.000 277.870 0.140 ; 
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 283.830 0.000 283.970 0.140 ; 
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 289.930 0.000 290.070 0.140 ; 
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 296.030 0.000 296.170 0.140 ; 
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 302.130 0.000 302.270 0.140 ; 
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 308.230 0.000 308.370 0.140 ; 
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 314.330 0.000 314.470 0.140 ; 
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 320.430 0.000 320.570 0.140 ; 
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 326.530 0.000 326.670 0.140 ; 
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 332.630 0.000 332.770 0.140 ; 
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 338.730 0.000 338.870 0.140 ; 
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 344.830 0.000 344.970 0.140 ; 
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 350.930 0.000 351.070 0.140 ; 
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 357.030 0.000 357.170 0.140 ; 
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 363.130 0.000 363.270 0.140 ; 
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 369.230 0.000 369.370 0.140 ; 
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 375.330 0.000 375.470 0.140 ; 
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 381.430 0.000 381.570 0.140 ; 
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 387.530 0.000 387.670 0.140 ; 
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 393.630 0.000 393.770 0.140 ; 
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 399.730 0.000 399.870 0.140 ; 
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 405.830 0.000 405.970 0.140 ; 
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 411.930 0.000 412.070 0.140 ; 
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 418.030 0.000 418.170 0.140 ; 
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 424.130 0.000 424.270 0.140 ; 
        END 
    END dout[31] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 234.610 0.000 234.750 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 240.710 0.000 240.850 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 246.810 0.000 246.950 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 252.910 0.000 253.050 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 259.010 0.000 259.150 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 265.110 0.000 265.250 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 271.210 0.000 271.350 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 277.310 0.000 277.450 0.140 ; 
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 283.410 0.000 283.550 0.140 ; 
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 289.510 0.000 289.650 0.140 ; 
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 295.610 0.000 295.750 0.140 ; 
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 301.710 0.000 301.850 0.140 ; 
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 307.810 0.000 307.950 0.140 ; 
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 313.910 0.000 314.050 0.140 ; 
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 320.010 0.000 320.150 0.140 ; 
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 326.110 0.000 326.250 0.140 ; 
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 332.210 0.000 332.350 0.140 ; 
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 338.310 0.000 338.450 0.140 ; 
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 344.410 0.000 344.550 0.140 ; 
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 350.510 0.000 350.650 0.140 ; 
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 356.610 0.000 356.750 0.140 ; 
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 362.710 0.000 362.850 0.140 ; 
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 368.810 0.000 368.950 0.140 ; 
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 374.910 0.000 375.050 0.140 ; 
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 381.010 0.000 381.150 0.140 ; 
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 387.110 0.000 387.250 0.140 ; 
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 393.210 0.000 393.350 0.140 ; 
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 399.310 0.000 399.450 0.140 ; 
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 405.410 0.000 405.550 0.140 ; 
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 411.510 0.000 411.650 0.140 ; 
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 417.610 0.000 417.750 0.140 ; 
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.851800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 423.710 0.000 423.850 0.140 ; 
        END 
    END din[31] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.662200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 234.260 0.000 234.400 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.662200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 283.060 0.000 283.200 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.662200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 331.860 0.000 332.000 0.140 ; 
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.662200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 380.660 0.000 380.800 0.140 ; 
        END 
    END wmask[3] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.616700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 192.920 0.000 193.240 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.616700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 186.800 0.000 187.120 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.616700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 180.680 0.000 181.000 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.616700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 174.560 0.000 174.880 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.616700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 168.440 0.000 168.760 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.616700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 162.320 0.000 162.640 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.616700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 156.200 0.000 156.520 0.320 ; 
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.616700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 150.080 0.000 150.400 0.320 ; 
        END 
    END addr[7] 
    PIN addr[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.616700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 143.960 0.000 144.280 0.320 ; 
        END 
    END addr[8] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.616700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 205.160 0.000 205.480 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.616700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 199.040 0.000 199.360 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 22.599000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 207.880 0.000 208.200 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 26.505000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 208.560 0.000 208.880 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 234.040 6.240 ; 
                RECT 424.800 5.920 443.120 6.240 ; 
                RECT 0.160 7.280 443.120 7.600 ; 
                RECT 0.160 8.640 443.120 8.960 ; 
                RECT 0.160 10.000 207.520 10.320 ; 
                RECT 381.280 10.000 443.120 10.320 ; 
                RECT 0.160 11.360 223.840 11.680 ; 
                RECT 433.640 11.360 443.120 11.680 ; 
                RECT 0.160 12.720 223.840 13.040 ; 
                RECT 433.640 12.720 443.120 13.040 ; 
                RECT 0.160 14.080 223.840 14.400 ; 
                RECT 433.640 14.080 443.120 14.400 ; 
                RECT 0.160 15.440 223.840 15.760 ; 
                RECT 433.640 15.440 443.120 15.760 ; 
                RECT 0.160 16.800 223.840 17.120 ; 
                RECT 433.640 16.800 443.120 17.120 ; 
                RECT 0.160 18.160 223.840 18.480 ; 
                RECT 433.640 18.160 443.120 18.480 ; 
                RECT 0.160 19.520 223.840 19.840 ; 
                RECT 433.640 19.520 443.120 19.840 ; 
                RECT 0.160 20.880 223.840 21.200 ; 
                RECT 433.640 20.880 443.120 21.200 ; 
                RECT 0.160 22.240 140.200 22.560 ; 
                RECT 209.240 22.240 223.840 22.560 ; 
                RECT 433.640 22.240 443.120 22.560 ; 
                RECT 0.160 23.600 223.840 23.920 ; 
                RECT 433.640 23.600 443.120 23.920 ; 
                RECT 0.160 24.960 223.840 25.280 ; 
                RECT 433.640 24.960 443.120 25.280 ; 
                RECT 0.160 26.320 140.200 26.640 ; 
                RECT 208.560 26.320 223.840 26.640 ; 
                RECT 433.640 26.320 443.120 26.640 ; 
                RECT 0.160 27.680 223.160 28.000 ; 
                RECT 433.640 27.680 443.120 28.000 ; 
                RECT 0.160 29.040 223.840 29.360 ; 
                RECT 433.640 29.040 443.120 29.360 ; 
                RECT 0.160 30.400 223.840 30.720 ; 
                RECT 433.640 30.400 443.120 30.720 ; 
                RECT 0.160 31.760 223.840 32.080 ; 
                RECT 433.640 31.760 443.120 32.080 ; 
                RECT 0.160 33.120 223.840 33.440 ; 
                RECT 433.640 33.120 443.120 33.440 ; 
                RECT 0.160 34.480 223.840 34.800 ; 
                RECT 433.640 34.480 443.120 34.800 ; 
                RECT 0.160 35.840 223.840 36.160 ; 
                RECT 433.640 35.840 443.120 36.160 ; 
                RECT 0.160 37.200 223.840 37.520 ; 
                RECT 433.640 37.200 443.120 37.520 ; 
                RECT 0.160 38.560 223.840 38.880 ; 
                RECT 433.640 38.560 443.120 38.880 ; 
                RECT 0.160 39.920 223.840 40.240 ; 
                RECT 433.640 39.920 443.120 40.240 ; 
                RECT 0.160 41.280 223.840 41.600 ; 
                RECT 433.640 41.280 443.120 41.600 ; 
                RECT 0.160 42.640 223.840 42.960 ; 
                RECT 433.640 42.640 443.120 42.960 ; 
                RECT 0.160 44.000 138.840 44.320 ; 
                RECT 187.480 44.000 223.840 44.320 ; 
                RECT 433.640 44.000 443.120 44.320 ; 
                RECT 0.160 45.360 137.480 45.680 ; 
                RECT 193.600 45.360 223.840 45.680 ; 
                RECT 433.640 45.360 443.120 45.680 ; 
                RECT 0.160 46.720 115.040 47.040 ; 
                RECT 208.560 46.720 223.840 47.040 ; 
                RECT 433.640 46.720 443.120 47.040 ; 
                RECT 0.160 48.080 115.720 48.400 ; 
                RECT 199.040 48.080 223.840 48.400 ; 
                RECT 433.640 48.080 443.120 48.400 ; 
                RECT 0.160 49.440 223.840 49.760 ; 
                RECT 433.640 49.440 443.120 49.760 ; 
                RECT 0.160 50.800 223.840 51.120 ; 
                RECT 433.640 50.800 443.120 51.120 ; 
                RECT 0.160 52.160 200.040 52.480 ; 
                RECT 206.520 52.160 223.840 52.480 ; 
                RECT 433.640 52.160 443.120 52.480 ; 
                RECT 0.160 53.520 200.040 53.840 ; 
                RECT 433.640 53.520 443.120 53.840 ; 
                RECT 0.160 54.880 135.440 55.200 ; 
                RECT 197.000 54.880 200.040 55.200 ; 
                RECT 206.520 54.880 223.840 55.200 ; 
                RECT 433.640 54.880 443.120 55.200 ; 
                RECT 0.160 56.240 223.840 56.560 ; 
                RECT 433.640 56.240 443.120 56.560 ; 
                RECT 0.160 57.600 223.840 57.920 ; 
                RECT 433.640 57.600 443.120 57.920 ; 
                RECT 0.160 58.960 223.840 59.280 ; 
                RECT 433.640 58.960 443.120 59.280 ; 
                RECT 0.160 60.320 223.840 60.640 ; 
                RECT 433.640 60.320 443.120 60.640 ; 
                RECT 0.160 61.680 136.800 62.000 ; 
                RECT 143.280 61.680 148.360 62.000 ; 
                RECT 205.840 61.680 223.840 62.000 ; 
                RECT 433.640 61.680 443.120 62.000 ; 
                RECT 0.160 63.040 138.160 63.360 ; 
                RECT 141.920 63.040 148.360 63.360 ; 
                RECT 216.040 63.040 223.840 63.360 ; 
                RECT 433.640 63.040 443.120 63.360 ; 
                RECT 0.160 64.400 148.360 64.720 ; 
                RECT 214.680 64.400 223.840 64.720 ; 
                RECT 433.640 64.400 443.120 64.720 ; 
                RECT 0.160 65.760 148.360 66.080 ; 
                RECT 216.040 65.760 223.840 66.080 ; 
                RECT 433.640 65.760 443.120 66.080 ; 
                RECT 0.160 67.120 148.360 67.440 ; 
                RECT 216.040 67.120 223.840 67.440 ; 
                RECT 433.640 67.120 443.120 67.440 ; 
                RECT 0.160 68.480 148.360 68.800 ; 
                RECT 216.040 68.480 223.840 68.800 ; 
                RECT 433.640 68.480 443.120 68.800 ; 
                RECT 0.160 69.840 148.360 70.160 ; 
                RECT 214.680 69.840 223.840 70.160 ; 
                RECT 433.640 69.840 443.120 70.160 ; 
                RECT 0.160 71.200 148.360 71.520 ; 
                RECT 205.840 71.200 223.840 71.520 ; 
                RECT 433.640 71.200 443.120 71.520 ; 
                RECT 0.160 72.560 113.000 72.880 ; 
                RECT 123.560 72.560 148.360 72.880 ; 
                RECT 214.680 72.560 223.840 72.880 ; 
                RECT 433.640 72.560 443.120 72.880 ; 
                RECT 0.160 73.920 114.360 74.240 ; 
                RECT 120.160 73.920 127.960 74.240 ; 
                RECT 130.360 73.920 148.360 74.240 ; 
                RECT 216.040 73.920 223.840 74.240 ; 
                RECT 433.640 73.920 443.120 74.240 ; 
                RECT 0.160 75.280 115.720 75.600 ; 
                RECT 119.480 75.280 148.360 75.600 ; 
                RECT 218.760 75.280 223.840 75.600 ; 
                RECT 433.640 75.280 443.120 75.600 ; 
                RECT 0.160 76.640 122.520 76.960 ; 
                RECT 129.680 76.640 148.360 76.960 ; 
                RECT 217.400 76.640 223.840 76.960 ; 
                RECT 433.640 76.640 443.120 76.960 ; 
                RECT 0.160 78.000 117.760 78.320 ; 
                RECT 131.040 78.000 148.360 78.320 ; 
                RECT 218.760 78.000 223.840 78.320 ; 
                RECT 433.640 78.000 443.120 78.320 ; 
                RECT 0.160 79.360 115.040 79.680 ; 
                RECT 123.560 79.360 148.360 79.680 ; 
                RECT 205.840 79.360 223.840 79.680 ; 
                RECT 433.640 79.360 443.120 79.680 ; 
                RECT 0.160 80.720 148.360 81.040 ; 
                RECT 218.760 80.720 223.840 81.040 ; 
                RECT 433.640 80.720 443.120 81.040 ; 
                RECT 0.160 82.080 114.360 82.400 ; 
                RECT 116.760 82.080 148.360 82.400 ; 
                RECT 218.760 82.080 223.840 82.400 ; 
                RECT 433.640 82.080 443.120 82.400 ; 
                RECT 0.160 83.440 112.320 83.760 ; 
                RECT 129.680 83.440 148.360 83.760 ; 
                RECT 217.400 83.440 223.840 83.760 ; 
                RECT 433.640 83.440 443.120 83.760 ; 
                RECT 0.160 84.800 121.160 85.120 ; 
                RECT 123.560 84.800 148.360 85.120 ; 
                RECT 218.760 84.800 223.840 85.120 ; 
                RECT 433.640 84.800 443.120 85.120 ; 
                RECT 0.160 86.160 148.360 86.480 ; 
                RECT 218.760 86.160 223.840 86.480 ; 
                RECT 433.640 86.160 443.120 86.480 ; 
                RECT 0.160 87.520 122.520 87.840 ; 
                RECT 130.360 87.520 148.360 87.840 ; 
                RECT 205.840 87.520 223.840 87.840 ; 
                RECT 433.640 87.520 443.120 87.840 ; 
                RECT 0.160 88.880 119.120 89.200 ; 
                RECT 123.560 88.880 148.360 89.200 ; 
                RECT 221.480 88.880 223.840 89.200 ; 
                RECT 433.640 88.880 443.120 89.200 ; 
                RECT 0.160 90.240 121.160 90.560 ; 
                RECT 123.560 90.240 148.360 90.560 ; 
                RECT 220.120 90.240 223.840 90.560 ; 
                RECT 433.640 90.240 443.120 90.560 ; 
                RECT 0.160 91.600 148.360 91.920 ; 
                RECT 221.480 91.600 223.840 91.920 ; 
                RECT 433.640 91.600 443.120 91.920 ; 
                RECT 0.160 92.960 112.320 93.280 ; 
                RECT 135.120 92.960 148.360 93.280 ; 
                RECT 221.480 92.960 223.840 93.280 ; 
                RECT 433.640 92.960 443.120 93.280 ; 
                RECT 0.160 94.320 130.680 94.640 ; 
                RECT 136.480 94.320 148.360 94.640 ; 
                RECT 221.480 94.320 223.840 94.640 ; 
                RECT 433.640 94.320 443.120 94.640 ; 
                RECT 0.160 95.680 121.160 96.000 ; 
                RECT 123.560 95.680 133.400 96.000 ; 
                RECT 137.160 95.680 148.360 96.000 ; 
                RECT 220.120 95.680 223.840 96.000 ; 
                RECT 433.640 95.680 443.120 96.000 ; 
                RECT 0.160 97.040 113.000 97.360 ; 
                RECT 126.960 97.040 148.360 97.360 ; 
                RECT 205.840 97.040 223.840 97.360 ; 
                RECT 433.640 97.040 443.120 97.360 ; 
                RECT 0.160 98.400 121.840 98.720 ; 
                RECT 130.360 98.400 148.360 98.720 ; 
                RECT 220.120 98.400 223.840 98.720 ; 
                RECT 433.640 98.400 443.120 98.720 ; 
                RECT 0.160 99.760 119.120 100.080 ; 
                RECT 123.560 99.760 148.360 100.080 ; 
                RECT 221.480 99.760 223.840 100.080 ; 
                RECT 433.640 99.760 443.120 100.080 ; 
                RECT 0.160 101.120 122.520 101.440 ; 
                RECT 131.040 101.120 148.360 101.440 ; 
                RECT 433.640 101.120 443.120 101.440 ; 
                RECT 0.160 102.480 148.360 102.800 ; 
                RECT 433.640 102.480 443.120 102.800 ; 
                RECT 0.160 103.840 115.040 104.160 ; 
                RECT 118.120 103.840 148.360 104.160 ; 
                RECT 433.640 103.840 443.120 104.160 ; 
                RECT 0.160 105.200 115.040 105.520 ; 
                RECT 123.560 105.200 148.360 105.520 ; 
                RECT 205.840 105.200 223.840 105.520 ; 
                RECT 433.640 105.200 443.120 105.520 ; 
                RECT 0.160 106.560 148.360 106.880 ; 
                RECT 433.640 106.560 443.120 106.880 ; 
                RECT 0.160 107.920 121.160 108.240 ; 
                RECT 123.560 107.920 148.360 108.240 ; 
                RECT 433.640 107.920 443.120 108.240 ; 
                RECT 0.160 109.280 114.360 109.600 ; 
                RECT 120.160 109.280 122.520 109.600 ; 
                RECT 124.240 109.280 148.360 109.600 ; 
                RECT 433.640 109.280 443.120 109.600 ; 
                RECT 0.160 110.640 118.440 110.960 ; 
                RECT 129.680 110.640 148.360 110.960 ; 
                RECT 433.640 110.640 443.120 110.960 ; 
                RECT 0.160 112.000 121.160 112.320 ; 
                RECT 123.560 112.000 148.360 112.320 ; 
                RECT 433.640 112.000 443.120 112.320 ; 
                RECT 0.160 113.360 116.400 113.680 ; 
                RECT 123.560 113.360 148.360 113.680 ; 
                RECT 205.840 113.360 223.840 113.680 ; 
                RECT 433.640 113.360 443.120 113.680 ; 
                RECT 0.160 114.720 121.840 115.040 ; 
                RECT 124.240 114.720 223.840 115.040 ; 
                RECT 433.640 114.720 443.120 115.040 ; 
                RECT 0.160 116.080 113.000 116.400 ; 
                RECT 120.160 116.080 223.840 116.400 ; 
                RECT 433.640 116.080 443.120 116.400 ; 
                RECT 0.160 117.440 112.320 117.760 ; 
                RECT 130.360 117.440 210.240 117.760 ; 
                RECT 433.640 117.440 443.120 117.760 ; 
                RECT 0.160 118.800 109.600 119.120 ; 
                RECT 130.360 118.800 221.120 119.120 ; 
                RECT 433.640 118.800 443.120 119.120 ; 
                RECT 0.160 120.160 113.000 120.480 ; 
                RECT 126.960 120.160 218.400 120.480 ; 
                RECT 433.640 120.160 443.120 120.480 ; 
                RECT 0.160 121.520 91.240 121.840 ; 
                RECT 109.960 121.520 215.680 121.840 ; 
                RECT 433.640 121.520 443.120 121.840 ; 
                RECT 0.160 122.880 91.240 123.200 ; 
                RECT 109.960 122.880 212.960 123.200 ; 
                RECT 433.640 122.880 443.120 123.200 ; 
                RECT 0.160 124.240 91.240 124.560 ; 
                RECT 109.960 124.240 125.240 124.560 ; 
                RECT 132.400 124.240 223.840 124.560 ; 
                RECT 433.640 124.240 443.120 124.560 ; 
                RECT 0.160 125.600 91.240 125.920 ; 
                RECT 109.960 125.600 223.840 125.920 ; 
                RECT 433.640 125.600 443.120 125.920 ; 
                RECT 0.160 126.960 91.240 127.280 ; 
                RECT 109.960 126.960 136.120 127.280 ; 
                RECT 165.720 126.960 168.760 127.280 ; 
                RECT 205.160 126.960 223.840 127.280 ; 
                RECT 433.640 126.960 443.120 127.280 ; 
                RECT 0.160 128.320 91.240 128.640 ; 
                RECT 109.960 128.320 168.760 128.640 ; 
                RECT 205.160 128.320 223.840 128.640 ; 
                RECT 433.640 128.320 443.120 128.640 ; 
                RECT 0.160 129.680 91.240 130.000 ; 
                RECT 109.960 129.680 112.320 130.000 ; 
                RECT 118.120 129.680 168.760 130.000 ; 
                RECT 205.160 129.680 223.840 130.000 ; 
                RECT 433.640 129.680 443.120 130.000 ; 
                RECT 0.160 131.040 91.240 131.360 ; 
                RECT 109.960 131.040 117.760 131.360 ; 
                RECT 130.360 131.040 168.760 131.360 ; 
                RECT 205.160 131.040 223.840 131.360 ; 
                RECT 433.640 131.040 443.120 131.360 ; 
                RECT 0.160 132.400 91.240 132.720 ; 
                RECT 109.960 132.400 168.760 132.720 ; 
                RECT 205.160 132.400 223.840 132.720 ; 
                RECT 433.640 132.400 443.120 132.720 ; 
                RECT 0.160 133.760 91.240 134.080 ; 
                RECT 109.960 133.760 168.760 134.080 ; 
                RECT 205.160 133.760 223.840 134.080 ; 
                RECT 433.640 133.760 443.120 134.080 ; 
                RECT 0.160 135.120 91.240 135.440 ; 
                RECT 109.960 135.120 223.840 135.440 ; 
                RECT 433.640 135.120 443.120 135.440 ; 
                RECT 0.160 136.480 91.240 136.800 ; 
                RECT 109.960 136.480 223.840 136.800 ; 
                RECT 433.640 136.480 443.120 136.800 ; 
                RECT 0.160 137.840 91.240 138.160 ; 
                RECT 109.960 137.840 223.840 138.160 ; 
                RECT 433.640 137.840 443.120 138.160 ; 
                RECT 0.160 139.200 91.240 139.520 ; 
                RECT 109.960 139.200 115.040 139.520 ; 
                RECT 119.480 139.200 127.960 139.520 ; 
                RECT 131.040 139.200 161.280 139.520 ; 
                RECT 207.200 139.200 223.840 139.520 ; 
                RECT 433.640 139.200 443.120 139.520 ; 
                RECT 0.160 140.560 91.240 140.880 ; 
                RECT 110.640 140.560 161.280 140.880 ; 
                RECT 207.200 140.560 223.840 140.880 ; 
                RECT 433.640 140.560 443.120 140.880 ; 
                RECT 0.160 141.920 91.240 142.240 ; 
                RECT 109.960 141.920 161.280 142.240 ; 
                RECT 207.200 141.920 223.840 142.240 ; 
                RECT 433.640 141.920 443.120 142.240 ; 
                RECT 0.160 143.280 91.240 143.600 ; 
                RECT 109.960 143.280 161.280 143.600 ; 
                RECT 207.200 143.280 223.840 143.600 ; 
                RECT 433.640 143.280 443.120 143.600 ; 
                RECT 0.160 144.640 91.240 144.960 ; 
                RECT 109.960 144.640 161.280 144.960 ; 
                RECT 207.200 144.640 223.840 144.960 ; 
                RECT 433.640 144.640 443.120 144.960 ; 
                RECT 0.160 146.000 91.240 146.320 ; 
                RECT 109.960 146.000 114.360 146.320 ; 
                RECT 117.440 146.000 161.280 146.320 ; 
                RECT 207.200 146.000 223.840 146.320 ; 
                RECT 433.640 146.000 443.120 146.320 ; 
                RECT 0.160 147.360 91.240 147.680 ; 
                RECT 109.960 147.360 121.160 147.680 ; 
                RECT 129.680 147.360 161.280 147.680 ; 
                RECT 207.200 147.360 223.840 147.680 ; 
                RECT 433.640 147.360 443.120 147.680 ; 
                RECT 0.160 148.720 91.240 149.040 ; 
                RECT 109.960 148.720 161.280 149.040 ; 
                RECT 207.200 148.720 214.320 149.040 ; 
                RECT 433.640 148.720 443.120 149.040 ; 
                RECT 0.160 150.080 91.240 150.400 ; 
                RECT 109.960 150.080 117.760 150.400 ; 
                RECT 120.160 150.080 161.280 150.400 ; 
                RECT 207.200 150.080 214.320 150.400 ; 
                RECT 433.640 150.080 443.120 150.400 ; 
                RECT 0.160 151.440 91.240 151.760 ; 
                RECT 109.960 151.440 161.280 151.760 ; 
                RECT 207.200 151.440 217.040 151.760 ; 
                RECT 433.640 151.440 443.120 151.760 ; 
                RECT 0.160 152.800 91.240 153.120 ; 
                RECT 109.960 152.800 161.280 153.120 ; 
                RECT 207.200 152.800 219.760 153.120 ; 
                RECT 433.640 152.800 443.120 153.120 ; 
                RECT 0.160 154.160 91.240 154.480 ; 
                RECT 109.960 154.160 161.280 154.480 ; 
                RECT 433.640 154.160 443.120 154.480 ; 
                RECT 0.160 155.520 91.240 155.840 ; 
                RECT 109.960 155.520 161.280 155.840 ; 
                RECT 433.640 155.520 443.120 155.840 ; 
                RECT 0.160 156.880 91.240 157.200 ; 
                RECT 109.960 156.880 161.280 157.200 ; 
                RECT 207.200 156.880 223.840 157.200 ; 
                RECT 433.640 156.880 443.120 157.200 ; 
                RECT 0.160 158.240 91.240 158.560 ; 
                RECT 109.960 158.240 161.280 158.560 ; 
                RECT 207.200 158.240 223.840 158.560 ; 
                RECT 433.640 158.240 443.120 158.560 ; 
                RECT 0.160 159.600 91.240 159.920 ; 
                RECT 109.960 159.600 161.280 159.920 ; 
                RECT 207.200 159.600 223.840 159.920 ; 
                RECT 433.640 159.600 443.120 159.920 ; 
                RECT 0.160 160.960 91.240 161.280 ; 
                RECT 109.960 160.960 116.400 161.280 ; 
                RECT 120.160 160.960 161.280 161.280 ; 
                RECT 207.200 160.960 223.840 161.280 ; 
                RECT 433.640 160.960 443.120 161.280 ; 
                RECT 0.160 162.320 161.280 162.640 ; 
                RECT 207.200 162.320 223.840 162.640 ; 
                RECT 433.640 162.320 443.120 162.640 ; 
                RECT 0.160 163.680 161.280 164.000 ; 
                RECT 207.200 163.680 223.840 164.000 ; 
                RECT 433.640 163.680 443.120 164.000 ; 
                RECT 0.160 165.040 72.880 165.360 ; 
                RECT 90.920 165.040 161.280 165.360 ; 
                RECT 207.200 165.040 223.840 165.360 ; 
                RECT 433.640 165.040 443.120 165.360 ; 
                RECT 0.160 166.400 72.880 166.720 ; 
                RECT 90.920 166.400 118.440 166.720 ; 
                RECT 124.240 166.400 161.280 166.720 ; 
                RECT 207.200 166.400 223.840 166.720 ; 
                RECT 433.640 166.400 443.120 166.720 ; 
                RECT 0.160 167.760 72.880 168.080 ; 
                RECT 90.920 167.760 97.360 168.080 ; 
                RECT 104.520 167.760 161.280 168.080 ; 
                RECT 207.200 167.760 223.840 168.080 ; 
                RECT 433.640 167.760 443.120 168.080 ; 
                RECT 0.160 169.120 72.880 169.440 ; 
                RECT 90.920 169.120 91.920 169.440 ; 
                RECT 109.280 169.120 161.280 169.440 ; 
                RECT 207.200 169.120 223.840 169.440 ; 
                RECT 433.640 169.120 443.120 169.440 ; 
                RECT 0.160 170.480 72.880 170.800 ; 
                RECT 90.920 170.480 161.280 170.800 ; 
                RECT 433.640 170.480 443.120 170.800 ; 
                RECT 0.160 171.840 69.480 172.160 ; 
                RECT 104.520 171.840 113.000 172.160 ; 
                RECT 122.880 171.840 161.280 172.160 ; 
                RECT 207.200 171.840 223.840 172.160 ; 
                RECT 433.640 171.840 443.120 172.160 ; 
                RECT 0.160 173.200 97.360 173.520 ; 
                RECT 117.440 173.200 443.120 173.520 ; 
                RECT 0.160 174.560 32.080 174.880 ; 
                RECT 116.760 174.560 443.120 174.880 ; 
                RECT 0.160 175.920 221.120 176.240 ; 
                RECT 435.680 175.920 443.120 176.240 ; 
                RECT 0.160 177.280 221.120 177.600 ; 
                RECT 435.680 177.280 443.120 177.600 ; 
                RECT 0.160 178.640 27.320 178.960 ; 
                RECT 33.800 178.640 99.400 178.960 ; 
                RECT 435.680 178.640 443.120 178.960 ; 
                RECT 0.160 180.000 25.280 180.320 ; 
                RECT 35.840 180.000 36.840 180.320 ; 
                RECT 48.760 180.000 99.400 180.320 ; 
                RECT 435.680 180.000 443.120 180.320 ; 
                RECT 0.160 181.360 25.280 181.680 ; 
                RECT 35.840 181.360 38.200 181.680 ; 
                RECT 47.400 181.360 59.280 181.680 ; 
                RECT 61.000 181.360 75.600 181.680 ; 
                RECT 89.560 181.360 99.400 181.680 ; 
                RECT 435.680 181.360 443.120 181.680 ; 
                RECT 0.160 182.720 59.280 183.040 ; 
                RECT 61.000 182.720 75.600 183.040 ; 
                RECT 89.560 182.720 99.400 183.040 ; 
                RECT 435.680 182.720 443.120 183.040 ; 
                RECT 0.160 184.080 25.280 184.400 ; 
                RECT 35.840 184.080 59.280 184.400 ; 
                RECT 63.720 184.080 75.600 184.400 ; 
                RECT 89.560 184.080 99.400 184.400 ; 
                RECT 435.680 184.080 443.120 184.400 ; 
                RECT 0.160 185.440 25.280 185.760 ; 
                RECT 35.840 185.440 59.280 185.760 ; 
                RECT 64.400 185.440 75.600 185.760 ; 
                RECT 89.560 185.440 99.400 185.760 ; 
                RECT 435.680 185.440 443.120 185.760 ; 
                RECT 0.160 186.800 25.280 187.120 ; 
                RECT 35.840 186.800 59.280 187.120 ; 
                RECT 65.080 186.800 75.600 187.120 ; 
                RECT 89.560 186.800 99.400 187.120 ; 
                RECT 435.680 186.800 443.120 187.120 ; 
                RECT 0.160 188.160 25.280 188.480 ; 
                RECT 35.840 188.160 99.400 188.480 ; 
                RECT 435.680 188.160 443.120 188.480 ; 
                RECT 0.160 189.520 75.600 189.840 ; 
                RECT 89.560 189.520 99.400 189.840 ; 
                RECT 435.680 189.520 443.120 189.840 ; 
                RECT 0.160 190.880 75.600 191.200 ; 
                RECT 89.560 190.880 99.400 191.200 ; 
                RECT 435.680 190.880 443.120 191.200 ; 
                RECT 0.160 192.240 18.480 192.560 ; 
                RECT 20.880 192.240 75.600 192.560 ; 
                RECT 89.560 192.240 99.400 192.560 ; 
                RECT 435.680 192.240 443.120 192.560 ; 
                RECT 0.160 193.600 17.800 193.920 ; 
                RECT 20.880 193.600 75.600 193.920 ; 
                RECT 89.560 193.600 99.400 193.920 ; 
                RECT 435.680 193.600 443.120 193.920 ; 
                RECT 0.160 194.960 38.880 195.280 ; 
                RECT 48.760 194.960 75.600 195.280 ; 
                RECT 83.440 194.960 99.400 195.280 ; 
                RECT 435.680 194.960 443.120 195.280 ; 
                RECT 0.160 196.320 17.120 196.640 ; 
                RECT 20.880 196.320 34.120 196.640 ; 
                RECT 48.080 196.320 83.760 196.640 ; 
                RECT 89.560 196.320 99.400 196.640 ; 
                RECT 435.680 196.320 443.120 196.640 ; 
                RECT 0.160 197.680 16.440 198.000 ; 
                RECT 20.880 197.680 34.120 198.000 ; 
                RECT 39.240 197.680 59.280 198.000 ; 
                RECT 61.680 197.680 75.600 198.000 ; 
                RECT 89.560 197.680 99.400 198.000 ; 
                RECT 435.680 197.680 443.120 198.000 ; 
                RECT 0.160 199.040 59.280 199.360 ; 
                RECT 62.360 199.040 75.600 199.360 ; 
                RECT 89.560 199.040 99.400 199.360 ; 
                RECT 435.680 199.040 443.120 199.360 ; 
                RECT 0.160 200.400 15.760 200.720 ; 
                RECT 20.880 200.400 34.120 200.720 ; 
                RECT 39.920 200.400 59.280 200.720 ; 
                RECT 62.360 200.400 75.600 200.720 ; 
                RECT 89.560 200.400 99.400 200.720 ; 
                RECT 435.680 200.400 443.120 200.720 ; 
                RECT 0.160 201.760 15.080 202.080 ; 
                RECT 20.880 201.760 34.120 202.080 ; 
                RECT 40.600 201.760 59.280 202.080 ; 
                RECT 61.000 201.760 75.600 202.080 ; 
                RECT 89.560 201.760 99.400 202.080 ; 
                RECT 435.680 201.760 443.120 202.080 ; 
                RECT 0.160 203.120 14.400 203.440 ; 
                RECT 20.880 203.120 34.120 203.440 ; 
                RECT 41.280 203.120 59.280 203.440 ; 
                RECT 63.040 203.120 75.600 203.440 ; 
                RECT 84.120 203.120 99.400 203.440 ; 
                RECT 435.680 203.120 443.120 203.440 ; 
                RECT 0.160 204.480 13.720 204.800 ; 
                RECT 20.880 204.480 75.600 204.800 ; 
                RECT 89.560 204.480 99.400 204.800 ; 
                RECT 435.680 204.480 443.120 204.800 ; 
                RECT 0.160 205.840 75.600 206.160 ; 
                RECT 89.560 205.840 99.400 206.160 ; 
                RECT 435.680 205.840 443.120 206.160 ; 
                RECT 0.160 207.200 13.040 207.520 ; 
                RECT 20.880 207.200 75.600 207.520 ; 
                RECT 89.560 207.200 99.400 207.520 ; 
                RECT 435.680 207.200 443.120 207.520 ; 
                RECT 0.160 208.560 12.360 208.880 ; 
                RECT 20.880 208.560 75.600 208.880 ; 
                RECT 89.560 208.560 99.400 208.880 ; 
                RECT 435.680 208.560 443.120 208.880 ; 
                RECT 0.160 209.920 11.680 210.240 ; 
                RECT 20.880 209.920 75.600 210.240 ; 
                RECT 89.560 209.920 99.400 210.240 ; 
                RECT 435.680 209.920 443.120 210.240 ; 
                RECT 0.160 211.280 99.400 211.600 ; 
                RECT 435.680 211.280 443.120 211.600 ; 
                RECT 0.160 212.640 11.000 212.960 ; 
                RECT 20.880 212.640 34.120 212.960 ; 
                RECT 38.560 212.640 75.600 212.960 ; 
                RECT 89.560 212.640 99.400 212.960 ; 
                RECT 435.680 212.640 443.120 212.960 ; 
                RECT 0.160 214.000 10.320 214.320 ; 
                RECT 20.880 214.000 75.600 214.320 ; 
                RECT 89.560 214.000 99.400 214.320 ; 
                RECT 435.680 214.000 443.120 214.320 ; 
                RECT 0.160 215.360 75.600 215.680 ; 
                RECT 89.560 215.360 99.400 215.680 ; 
                RECT 435.680 215.360 443.120 215.680 ; 
                RECT 0.160 216.720 9.640 217.040 ; 
                RECT 20.880 216.720 34.120 217.040 ; 
                RECT 37.200 216.720 75.600 217.040 ; 
                RECT 89.560 216.720 99.400 217.040 ; 
                RECT 435.680 216.720 443.120 217.040 ; 
                RECT 0.160 218.080 75.600 218.400 ; 
                RECT 89.560 218.080 99.400 218.400 ; 
                RECT 435.680 218.080 443.120 218.400 ; 
                RECT 0.160 219.440 99.400 219.760 ; 
                RECT 435.680 219.440 443.120 219.760 ; 
                RECT 0.160 220.800 75.600 221.120 ; 
                RECT 89.560 220.800 99.400 221.120 ; 
                RECT 435.680 220.800 443.120 221.120 ; 
                RECT 0.160 222.160 75.600 222.480 ; 
                RECT 89.560 222.160 99.400 222.480 ; 
                RECT 435.680 222.160 443.120 222.480 ; 
                RECT 0.160 223.520 75.600 223.840 ; 
                RECT 89.560 223.520 99.400 223.840 ; 
                RECT 435.680 223.520 443.120 223.840 ; 
                RECT 0.160 224.880 75.600 225.200 ; 
                RECT 89.560 224.880 99.400 225.200 ; 
                RECT 435.680 224.880 443.120 225.200 ; 
                RECT 0.160 226.240 75.600 226.560 ; 
                RECT 89.560 226.240 99.400 226.560 ; 
                RECT 435.680 226.240 443.120 226.560 ; 
                RECT 0.160 227.600 99.400 227.920 ; 
                RECT 435.680 227.600 443.120 227.920 ; 
                RECT 0.160 228.960 75.600 229.280 ; 
                RECT 89.560 228.960 99.400 229.280 ; 
                RECT 435.680 228.960 443.120 229.280 ; 
                RECT 0.160 230.320 75.600 230.640 ; 
                RECT 89.560 230.320 99.400 230.640 ; 
                RECT 435.680 230.320 443.120 230.640 ; 
                RECT 0.160 231.680 75.600 232.000 ; 
                RECT 89.560 231.680 99.400 232.000 ; 
                RECT 435.680 231.680 443.120 232.000 ; 
                RECT 0.160 233.040 75.600 233.360 ; 
                RECT 89.560 233.040 99.400 233.360 ; 
                RECT 435.680 233.040 443.120 233.360 ; 
                RECT 0.160 234.400 75.600 234.720 ; 
                RECT 88.200 234.400 99.400 234.720 ; 
                RECT 435.680 234.400 443.120 234.720 ; 
                RECT 0.160 235.760 85.800 236.080 ; 
                RECT 89.560 235.760 99.400 236.080 ; 
                RECT 435.680 235.760 443.120 236.080 ; 
                RECT 0.160 237.120 75.600 237.440 ; 
                RECT 89.560 237.120 99.400 237.440 ; 
                RECT 435.680 237.120 443.120 237.440 ; 
                RECT 0.160 238.480 75.600 238.800 ; 
                RECT 89.560 238.480 99.400 238.800 ; 
                RECT 435.680 238.480 443.120 238.800 ; 
                RECT 0.160 239.840 75.600 240.160 ; 
                RECT 89.560 239.840 99.400 240.160 ; 
                RECT 435.680 239.840 443.120 240.160 ; 
                RECT 0.160 241.200 75.600 241.520 ; 
                RECT 89.560 241.200 99.400 241.520 ; 
                RECT 435.680 241.200 443.120 241.520 ; 
                RECT 0.160 242.560 75.600 242.880 ; 
                RECT 88.880 242.560 99.400 242.880 ; 
                RECT 435.680 242.560 443.120 242.880 ; 
                RECT 0.160 243.920 80.360 244.240 ; 
                RECT 89.560 243.920 99.400 244.240 ; 
                RECT 435.680 243.920 443.120 244.240 ; 
                RECT 0.160 245.280 77.640 245.600 ; 
                RECT 89.560 245.280 99.400 245.600 ; 
                RECT 435.680 245.280 443.120 245.600 ; 
                RECT 0.160 246.640 77.640 246.960 ; 
                RECT 89.560 246.640 99.400 246.960 ; 
                RECT 435.680 246.640 443.120 246.960 ; 
                RECT 0.160 248.000 77.640 248.320 ; 
                RECT 89.560 248.000 99.400 248.320 ; 
                RECT 435.680 248.000 443.120 248.320 ; 
                RECT 0.160 249.360 77.640 249.680 ; 
                RECT 89.560 249.360 99.400 249.680 ; 
                RECT 435.680 249.360 443.120 249.680 ; 
                RECT 0.160 250.720 39.560 251.040 ; 
                RECT 65.080 250.720 99.400 251.040 ; 
                RECT 435.680 250.720 443.120 251.040 ; 
                RECT 0.160 252.080 38.200 252.400 ; 
                RECT 64.400 252.080 77.640 252.400 ; 
                RECT 89.560 252.080 99.400 252.400 ; 
                RECT 435.680 252.080 443.120 252.400 ; 
                RECT 0.160 253.440 36.840 253.760 ; 
                RECT 63.040 253.440 75.600 253.760 ; 
                RECT 89.560 253.440 99.400 253.760 ; 
                RECT 435.680 253.440 443.120 253.760 ; 
                RECT 0.160 254.800 75.600 255.120 ; 
                RECT 89.560 254.800 99.400 255.120 ; 
                RECT 435.680 254.800 443.120 255.120 ; 
                RECT 0.160 256.160 75.600 256.480 ; 
                RECT 89.560 256.160 99.400 256.480 ; 
                RECT 435.680 256.160 443.120 256.480 ; 
                RECT 0.160 257.520 75.600 257.840 ; 
                RECT 89.560 257.520 99.400 257.840 ; 
                RECT 435.680 257.520 443.120 257.840 ; 
                RECT 0.160 258.880 99.400 259.200 ; 
                RECT 435.680 258.880 443.120 259.200 ; 
                RECT 0.160 260.240 77.640 260.560 ; 
                RECT 89.560 260.240 99.400 260.560 ; 
                RECT 435.680 260.240 443.120 260.560 ; 
                RECT 0.160 261.600 75.600 261.920 ; 
                RECT 89.560 261.600 99.400 261.920 ; 
                RECT 435.680 261.600 443.120 261.920 ; 
                RECT 0.160 262.960 75.600 263.280 ; 
                RECT 89.560 262.960 99.400 263.280 ; 
                RECT 435.680 262.960 443.120 263.280 ; 
                RECT 0.160 264.320 75.600 264.640 ; 
                RECT 89.560 264.320 99.400 264.640 ; 
                RECT 435.680 264.320 443.120 264.640 ; 
                RECT 0.160 265.680 75.600 266.000 ; 
                RECT 89.560 265.680 99.400 266.000 ; 
                RECT 435.680 265.680 443.120 266.000 ; 
                RECT 0.160 267.040 99.400 267.360 ; 
                RECT 435.680 267.040 443.120 267.360 ; 
                RECT 0.160 268.400 75.600 268.720 ; 
                RECT 89.560 268.400 99.400 268.720 ; 
                RECT 435.680 268.400 443.120 268.720 ; 
                RECT 0.160 269.760 75.600 270.080 ; 
                RECT 89.560 269.760 99.400 270.080 ; 
                RECT 435.680 269.760 443.120 270.080 ; 
                RECT 0.160 271.120 75.600 271.440 ; 
                RECT 89.560 271.120 99.400 271.440 ; 
                RECT 435.680 271.120 443.120 271.440 ; 
                RECT 0.160 272.480 75.600 272.800 ; 
                RECT 89.560 272.480 99.400 272.800 ; 
                RECT 435.680 272.480 443.120 272.800 ; 
                RECT 0.160 273.840 75.600 274.160 ; 
                RECT 78.680 273.840 99.400 274.160 ; 
                RECT 435.680 273.840 443.120 274.160 ; 
                RECT 0.160 275.200 80.360 275.520 ; 
                RECT 89.560 275.200 99.400 275.520 ; 
                RECT 435.680 275.200 443.120 275.520 ; 
                RECT 0.160 276.560 75.600 276.880 ; 
                RECT 89.560 276.560 99.400 276.880 ; 
                RECT 435.680 276.560 443.120 276.880 ; 
                RECT 0.160 277.920 75.600 278.240 ; 
                RECT 89.560 277.920 99.400 278.240 ; 
                RECT 435.680 277.920 443.120 278.240 ; 
                RECT 0.160 279.280 77.640 279.600 ; 
                RECT 89.560 279.280 99.400 279.600 ; 
                RECT 435.680 279.280 443.120 279.600 ; 
                RECT 0.160 280.640 75.600 280.960 ; 
                RECT 89.560 280.640 99.400 280.960 ; 
                RECT 435.680 280.640 443.120 280.960 ; 
                RECT 0.160 282.000 75.600 282.320 ; 
                RECT 79.360 282.000 99.400 282.320 ; 
                RECT 435.680 282.000 443.120 282.320 ; 
                RECT 0.160 283.360 82.400 283.680 ; 
                RECT 89.560 283.360 99.400 283.680 ; 
                RECT 435.680 283.360 443.120 283.680 ; 
                RECT 0.160 284.720 75.600 285.040 ; 
                RECT 89.560 284.720 99.400 285.040 ; 
                RECT 435.680 284.720 443.120 285.040 ; 
                RECT 0.160 286.080 75.600 286.400 ; 
                RECT 89.560 286.080 99.400 286.400 ; 
                RECT 435.680 286.080 443.120 286.400 ; 
                RECT 0.160 287.440 75.600 287.760 ; 
                RECT 89.560 287.440 99.400 287.760 ; 
                RECT 435.680 287.440 443.120 287.760 ; 
                RECT 0.160 288.800 75.600 289.120 ; 
                RECT 89.560 288.800 99.400 289.120 ; 
                RECT 435.680 288.800 443.120 289.120 ; 
                RECT 0.160 290.160 99.400 290.480 ; 
                RECT 435.680 290.160 443.120 290.480 ; 
                RECT 0.160 291.520 77.640 291.840 ; 
                RECT 89.560 291.520 99.400 291.840 ; 
                RECT 435.680 291.520 443.120 291.840 ; 
                RECT 0.160 292.880 75.600 293.200 ; 
                RECT 89.560 292.880 99.400 293.200 ; 
                RECT 435.680 292.880 443.120 293.200 ; 
                RECT 0.160 294.240 75.600 294.560 ; 
                RECT 89.560 294.240 99.400 294.560 ; 
                RECT 435.680 294.240 443.120 294.560 ; 
                RECT 0.160 295.600 75.600 295.920 ; 
                RECT 89.560 295.600 99.400 295.920 ; 
                RECT 435.680 295.600 443.120 295.920 ; 
                RECT 0.160 296.960 75.600 297.280 ; 
                RECT 89.560 296.960 99.400 297.280 ; 
                RECT 435.680 296.960 443.120 297.280 ; 
                RECT 0.160 298.320 99.400 298.640 ; 
                RECT 435.680 298.320 443.120 298.640 ; 
                RECT 0.160 299.680 77.640 300.000 ; 
                RECT 89.560 299.680 99.400 300.000 ; 
                RECT 435.680 299.680 443.120 300.000 ; 
                RECT 0.160 301.040 75.600 301.360 ; 
                RECT 89.560 301.040 99.400 301.360 ; 
                RECT 435.680 301.040 443.120 301.360 ; 
                RECT 0.160 302.400 75.600 302.720 ; 
                RECT 89.560 302.400 99.400 302.720 ; 
                RECT 435.680 302.400 443.120 302.720 ; 
                RECT 0.160 303.760 75.600 304.080 ; 
                RECT 89.560 303.760 99.400 304.080 ; 
                RECT 435.680 303.760 443.120 304.080 ; 
                RECT 0.160 305.120 75.600 305.440 ; 
                RECT 89.560 305.120 99.400 305.440 ; 
                RECT 435.680 305.120 443.120 305.440 ; 
                RECT 0.160 306.480 99.400 306.800 ; 
                RECT 435.680 306.480 443.120 306.800 ; 
                RECT 0.160 307.840 75.600 308.160 ; 
                RECT 89.560 307.840 99.400 308.160 ; 
                RECT 435.680 307.840 443.120 308.160 ; 
                RECT 0.160 309.200 75.600 309.520 ; 
                RECT 89.560 309.200 99.400 309.520 ; 
                RECT 435.680 309.200 443.120 309.520 ; 
                RECT 0.160 310.560 75.600 310.880 ; 
                RECT 89.560 310.560 99.400 310.880 ; 
                RECT 435.680 310.560 443.120 310.880 ; 
                RECT 0.160 311.920 75.600 312.240 ; 
                RECT 89.560 311.920 99.400 312.240 ; 
                RECT 435.680 311.920 443.120 312.240 ; 
                RECT 0.160 313.280 75.600 313.600 ; 
                RECT 81.400 313.280 99.400 313.600 ; 
                RECT 435.680 313.280 443.120 313.600 ; 
                RECT 0.160 314.640 99.400 314.960 ; 
                RECT 435.680 314.640 443.120 314.960 ; 
                RECT 0.160 316.000 78.320 316.320 ; 
                RECT 89.560 316.000 99.400 316.320 ; 
                RECT 435.680 316.000 443.120 316.320 ; 
                RECT 0.160 317.360 78.320 317.680 ; 
                RECT 89.560 317.360 99.400 317.680 ; 
                RECT 435.680 317.360 443.120 317.680 ; 
                RECT 0.160 318.720 78.320 319.040 ; 
                RECT 89.560 318.720 99.400 319.040 ; 
                RECT 435.680 318.720 443.120 319.040 ; 
                RECT 0.160 320.080 78.320 320.400 ; 
                RECT 89.560 320.080 99.400 320.400 ; 
                RECT 435.680 320.080 443.120 320.400 ; 
                RECT 0.160 321.440 99.400 321.760 ; 
                RECT 435.680 321.440 443.120 321.760 ; 
                RECT 0.160 322.800 83.760 323.120 ; 
                RECT 89.560 322.800 99.400 323.120 ; 
                RECT 435.680 322.800 443.120 323.120 ; 
                RECT 0.160 324.160 78.320 324.480 ; 
                RECT 89.560 324.160 99.400 324.480 ; 
                RECT 435.680 324.160 443.120 324.480 ; 
                RECT 0.160 325.520 78.320 325.840 ; 
                RECT 89.560 325.520 99.400 325.840 ; 
                RECT 435.680 325.520 443.120 325.840 ; 
                RECT 0.160 326.880 78.320 327.200 ; 
                RECT 89.560 326.880 99.400 327.200 ; 
                RECT 435.680 326.880 443.120 327.200 ; 
                RECT 0.160 328.240 78.320 328.560 ; 
                RECT 89.560 328.240 99.400 328.560 ; 
                RECT 435.680 328.240 443.120 328.560 ; 
                RECT 0.160 329.600 99.400 329.920 ; 
                RECT 435.680 329.600 443.120 329.920 ; 
                RECT 0.160 330.960 78.320 331.280 ; 
                RECT 89.560 330.960 99.400 331.280 ; 
                RECT 435.680 330.960 443.120 331.280 ; 
                RECT 0.160 332.320 86.480 332.640 ; 
                RECT 89.560 332.320 99.400 332.640 ; 
                RECT 435.680 332.320 443.120 332.640 ; 
                RECT 0.160 333.680 78.320 334.000 ; 
                RECT 89.560 333.680 99.400 334.000 ; 
                RECT 435.680 333.680 443.120 334.000 ; 
                RECT 0.160 335.040 78.320 335.360 ; 
                RECT 89.560 335.040 99.400 335.360 ; 
                RECT 435.680 335.040 443.120 335.360 ; 
                RECT 0.160 336.400 78.320 336.720 ; 
                RECT 89.560 336.400 99.400 336.720 ; 
                RECT 435.680 336.400 443.120 336.720 ; 
                RECT 0.160 337.760 99.400 338.080 ; 
                RECT 435.680 337.760 443.120 338.080 ; 
                RECT 0.160 339.120 79.000 339.440 ; 
                RECT 89.560 339.120 99.400 339.440 ; 
                RECT 435.680 339.120 443.120 339.440 ; 
                RECT 0.160 340.480 79.000 340.800 ; 
                RECT 89.560 340.480 99.400 340.800 ; 
                RECT 435.680 340.480 443.120 340.800 ; 
                RECT 0.160 341.840 81.040 342.160 ; 
                RECT 89.560 341.840 99.400 342.160 ; 
                RECT 435.680 341.840 443.120 342.160 ; 
                RECT 0.160 343.200 79.000 343.520 ; 
                RECT 89.560 343.200 99.400 343.520 ; 
                RECT 435.680 343.200 443.120 343.520 ; 
                RECT 0.160 344.560 79.000 344.880 ; 
                RECT 89.560 344.560 99.400 344.880 ; 
                RECT 435.680 344.560 443.120 344.880 ; 
                RECT 0.160 345.920 99.400 346.240 ; 
                RECT 435.680 345.920 443.120 346.240 ; 
                RECT 0.160 347.280 79.000 347.600 ; 
                RECT 89.560 347.280 99.400 347.600 ; 
                RECT 435.680 347.280 443.120 347.600 ; 
                RECT 0.160 348.640 79.000 348.960 ; 
                RECT 89.560 348.640 99.400 348.960 ; 
                RECT 435.680 348.640 443.120 348.960 ; 
                RECT 0.160 350.000 79.000 350.320 ; 
                RECT 89.560 350.000 99.400 350.320 ; 
                RECT 435.680 350.000 443.120 350.320 ; 
                RECT 0.160 351.360 83.760 351.680 ; 
                RECT 89.560 351.360 99.400 351.680 ; 
                RECT 435.680 351.360 443.120 351.680 ; 
                RECT 0.160 352.720 79.000 353.040 ; 
                RECT 89.560 352.720 99.400 353.040 ; 
                RECT 435.680 352.720 443.120 353.040 ; 
                RECT 0.160 354.080 99.400 354.400 ; 
                RECT 435.680 354.080 443.120 354.400 ; 
                RECT 0.160 355.440 79.000 355.760 ; 
                RECT 89.560 355.440 99.400 355.760 ; 
                RECT 435.680 355.440 443.120 355.760 ; 
                RECT 0.160 356.800 79.000 357.120 ; 
                RECT 89.560 356.800 99.400 357.120 ; 
                RECT 435.680 356.800 443.120 357.120 ; 
                RECT 0.160 358.160 79.000 358.480 ; 
                RECT 89.560 358.160 99.400 358.480 ; 
                RECT 435.680 358.160 443.120 358.480 ; 
                RECT 0.160 359.520 79.000 359.840 ; 
                RECT 89.560 359.520 99.400 359.840 ; 
                RECT 435.680 359.520 443.120 359.840 ; 
                RECT 0.160 360.880 99.400 361.200 ; 
                RECT 435.680 360.880 443.120 361.200 ; 
                RECT 0.160 362.240 85.800 362.560 ; 
                RECT 89.560 362.240 99.400 362.560 ; 
                RECT 435.680 362.240 443.120 362.560 ; 
                RECT 0.160 363.600 79.000 363.920 ; 
                RECT 89.560 363.600 99.400 363.920 ; 
                RECT 435.680 363.600 443.120 363.920 ; 
                RECT 0.160 364.960 79.000 365.280 ; 
                RECT 89.560 364.960 99.400 365.280 ; 
                RECT 435.680 364.960 443.120 365.280 ; 
                RECT 0.160 366.320 79.000 366.640 ; 
                RECT 89.560 366.320 99.400 366.640 ; 
                RECT 435.680 366.320 443.120 366.640 ; 
                RECT 0.160 367.680 79.000 368.000 ; 
                RECT 89.560 367.680 99.400 368.000 ; 
                RECT 435.680 367.680 443.120 368.000 ; 
                RECT 0.160 369.040 99.400 369.360 ; 
                RECT 435.680 369.040 443.120 369.360 ; 
                RECT 0.160 370.400 80.360 370.720 ; 
                RECT 89.560 370.400 99.400 370.720 ; 
                RECT 435.680 370.400 443.120 370.720 ; 
                RECT 0.160 371.760 80.360 372.080 ; 
                RECT 89.560 371.760 99.400 372.080 ; 
                RECT 435.680 371.760 443.120 372.080 ; 
                RECT 0.160 373.120 79.000 373.440 ; 
                RECT 89.560 373.120 99.400 373.440 ; 
                RECT 435.680 373.120 443.120 373.440 ; 
                RECT 0.160 374.480 79.000 374.800 ; 
                RECT 89.560 374.480 99.400 374.800 ; 
                RECT 435.680 374.480 443.120 374.800 ; 
                RECT 0.160 375.840 79.000 376.160 ; 
                RECT 89.560 375.840 99.400 376.160 ; 
                RECT 435.680 375.840 443.120 376.160 ; 
                RECT 0.160 377.200 99.400 377.520 ; 
                RECT 435.680 377.200 443.120 377.520 ; 
                RECT 0.160 378.560 79.000 378.880 ; 
                RECT 89.560 378.560 99.400 378.880 ; 
                RECT 435.680 378.560 443.120 378.880 ; 
                RECT 0.160 379.920 79.000 380.240 ; 
                RECT 89.560 379.920 99.400 380.240 ; 
                RECT 435.680 379.920 443.120 380.240 ; 
                RECT 0.160 381.280 83.080 381.600 ; 
                RECT 89.560 381.280 99.400 381.600 ; 
                RECT 435.680 381.280 443.120 381.600 ; 
                RECT 0.160 382.640 79.000 382.960 ; 
                RECT 89.560 382.640 99.400 382.960 ; 
                RECT 435.680 382.640 443.120 382.960 ; 
                RECT 0.160 384.000 79.000 384.320 ; 
                RECT 89.560 384.000 99.400 384.320 ; 
                RECT 435.680 384.000 443.120 384.320 ; 
                RECT 0.160 385.360 99.400 385.680 ; 
                RECT 435.680 385.360 443.120 385.680 ; 
                RECT 0.160 386.720 79.000 387.040 ; 
                RECT 89.560 386.720 99.400 387.040 ; 
                RECT 435.680 386.720 443.120 387.040 ; 
                RECT 0.160 388.080 79.000 388.400 ; 
                RECT 89.560 388.080 99.400 388.400 ; 
                RECT 435.680 388.080 443.120 388.400 ; 
                RECT 0.160 389.440 79.000 389.760 ; 
                RECT 89.560 389.440 99.400 389.760 ; 
                RECT 435.680 389.440 443.120 389.760 ; 
                RECT 0.160 390.800 85.800 391.120 ; 
                RECT 89.560 390.800 99.400 391.120 ; 
                RECT 435.680 390.800 443.120 391.120 ; 
                RECT 0.160 392.160 79.000 392.480 ; 
                RECT 89.560 392.160 99.400 392.480 ; 
                RECT 435.680 392.160 443.120 392.480 ; 
                RECT 0.160 393.520 99.400 393.840 ; 
                RECT 435.680 393.520 443.120 393.840 ; 
                RECT 0.160 394.880 79.000 395.200 ; 
                RECT 89.560 394.880 99.400 395.200 ; 
                RECT 435.680 394.880 443.120 395.200 ; 
                RECT 0.160 396.240 79.000 396.560 ; 
                RECT 89.560 396.240 99.400 396.560 ; 
                RECT 435.680 396.240 443.120 396.560 ; 
                RECT 0.160 397.600 79.000 397.920 ; 
                RECT 89.560 397.600 99.400 397.920 ; 
                RECT 435.680 397.600 443.120 397.920 ; 
                RECT 0.160 398.960 79.000 399.280 ; 
                RECT 89.560 398.960 99.400 399.280 ; 
                RECT 435.680 398.960 443.120 399.280 ; 
                RECT 0.160 400.320 99.400 400.640 ; 
                RECT 435.680 400.320 443.120 400.640 ; 
                RECT 0.160 401.680 80.360 402.000 ; 
                RECT 89.560 401.680 99.400 402.000 ; 
                RECT 435.680 401.680 443.120 402.000 ; 
                RECT 0.160 403.040 79.680 403.360 ; 
                RECT 89.560 403.040 99.400 403.360 ; 
                RECT 435.680 403.040 443.120 403.360 ; 
                RECT 0.160 404.400 79.680 404.720 ; 
                RECT 89.560 404.400 99.400 404.720 ; 
                RECT 435.680 404.400 443.120 404.720 ; 
                RECT 0.160 405.760 79.680 406.080 ; 
                RECT 89.560 405.760 99.400 406.080 ; 
                RECT 435.680 405.760 443.120 406.080 ; 
                RECT 0.160 407.120 79.680 407.440 ; 
                RECT 89.560 407.120 99.400 407.440 ; 
                RECT 435.680 407.120 443.120 407.440 ; 
                RECT 0.160 408.480 99.400 408.800 ; 
                RECT 435.680 408.480 443.120 408.800 ; 
                RECT 0.160 409.840 82.400 410.160 ; 
                RECT 89.560 409.840 99.400 410.160 ; 
                RECT 435.680 409.840 443.120 410.160 ; 
                RECT 0.160 411.200 79.680 411.520 ; 
                RECT 89.560 411.200 99.400 411.520 ; 
                RECT 435.680 411.200 443.120 411.520 ; 
                RECT 0.160 412.560 79.680 412.880 ; 
                RECT 89.560 412.560 99.400 412.880 ; 
                RECT 435.680 412.560 443.120 412.880 ; 
                RECT 0.160 413.920 79.680 414.240 ; 
                RECT 89.560 413.920 99.400 414.240 ; 
                RECT 435.680 413.920 443.120 414.240 ; 
                RECT 0.160 415.280 79.680 415.600 ; 
                RECT 89.560 415.280 99.400 415.600 ; 
                RECT 435.680 415.280 443.120 415.600 ; 
                RECT 0.160 416.640 99.400 416.960 ; 
                RECT 435.680 416.640 443.120 416.960 ; 
                RECT 0.160 418.000 79.680 418.320 ; 
                RECT 89.560 418.000 99.400 418.320 ; 
                RECT 435.680 418.000 443.120 418.320 ; 
                RECT 0.160 419.360 84.440 419.680 ; 
                RECT 89.560 419.360 99.400 419.680 ; 
                RECT 435.680 419.360 443.120 419.680 ; 
                RECT 0.160 420.720 85.120 421.040 ; 
                RECT 89.560 420.720 99.400 421.040 ; 
                RECT 435.680 420.720 443.120 421.040 ; 
                RECT 0.160 422.080 79.680 422.400 ; 
                RECT 89.560 422.080 99.400 422.400 ; 
                RECT 435.680 422.080 443.120 422.400 ; 
                RECT 0.160 423.440 79.680 423.760 ; 
                RECT 89.560 423.440 99.400 423.760 ; 
                RECT 435.680 423.440 443.120 423.760 ; 
                RECT 0.160 424.800 99.400 425.120 ; 
                RECT 435.680 424.800 443.120 425.120 ; 
                RECT 0.160 426.160 79.680 426.480 ; 
                RECT 89.560 426.160 99.400 426.480 ; 
                RECT 435.680 426.160 443.120 426.480 ; 
                RECT 0.160 427.520 79.680 427.840 ; 
                RECT 89.560 427.520 99.400 427.840 ; 
                RECT 435.680 427.520 443.120 427.840 ; 
                RECT 0.160 428.880 87.160 429.200 ; 
                RECT 89.560 428.880 99.400 429.200 ; 
                RECT 435.680 428.880 443.120 429.200 ; 
                RECT 0.160 430.240 87.160 430.560 ; 
                RECT 89.560 430.240 99.400 430.560 ; 
                RECT 435.680 430.240 443.120 430.560 ; 
                RECT 0.160 431.600 79.680 431.920 ; 
                RECT 89.560 431.600 99.400 431.920 ; 
                RECT 435.680 431.600 443.120 431.920 ; 
                RECT 0.160 432.960 99.400 433.280 ; 
                RECT 435.680 432.960 443.120 433.280 ; 
                RECT 0.160 434.320 221.120 434.640 ; 
                RECT 435.680 434.320 443.120 434.640 ; 
                RECT 0.160 435.680 221.120 436.000 ; 
                RECT 435.680 435.680 443.120 436.000 ; 
                RECT 0.160 437.040 221.120 437.360 ; 
                RECT 435.680 437.040 443.120 437.360 ; 
                RECT 0.160 438.400 443.120 438.720 ; 
                RECT 0.160 439.760 443.120 440.080 ; 
                RECT 0.160 441.120 443.120 441.440 ; 
                RECT 0.160 442.480 443.120 442.800 ; 
                RECT 0.160 0.160 443.120 1.520 ; 
                RECT 0.160 447.200 443.120 448.560 ; 
                RECT 225.260 32.370 231.060 33.740 ; 
                RECT 425.960 32.370 431.760 33.740 ; 
                RECT 225.260 37.405 231.060 38.765 ; 
                RECT 425.960 37.405 431.760 38.765 ; 
                RECT 225.260 42.470 231.060 43.870 ; 
                RECT 425.960 42.470 431.760 43.870 ; 
                RECT 225.260 47.645 231.060 49.085 ; 
                RECT 425.960 47.645 431.760 49.085 ; 
                RECT 225.260 52.740 231.060 54.070 ; 
                RECT 425.960 52.740 431.760 54.070 ; 
                RECT 225.260 57.670 231.060 59.000 ; 
                RECT 425.960 57.670 431.760 59.000 ; 
                RECT 225.260 95.705 431.760 99.305 ; 
                RECT 225.260 80.290 431.760 81.090 ; 
                RECT 225.260 130.125 431.760 131.925 ; 
                RECT 225.260 65.810 431.760 67.610 ; 
                RECT 225.260 77.280 431.760 78.080 ; 
                RECT 225.260 162.465 431.760 166.065 ; 
                RECT 225.260 85.180 431.760 85.980 ; 
                RECT 225.260 103.085 431.760 103.375 ; 
                RECT 225.260 16.615 431.760 18.415 ; 
                RECT 104.630 179.035 106.550 433.415 ; 
                RECT 115.505 179.035 117.425 433.415 ; 
                RECT 119.345 179.035 121.265 433.415 ; 
                RECT 123.185 179.035 125.105 433.415 ; 
                RECT 138.850 179.035 140.770 433.415 ; 
                RECT 142.690 179.035 144.610 433.415 ; 
                RECT 146.530 179.035 148.450 433.415 ; 
                RECT 150.370 179.035 152.290 433.415 ; 
                RECT 154.210 179.035 156.130 433.415 ; 
                RECT 178.810 179.035 180.730 433.415 ; 
                RECT 182.650 179.035 184.570 433.415 ; 
                RECT 186.490 179.035 188.410 433.415 ; 
                RECT 190.330 179.035 192.250 433.415 ; 
                RECT 194.170 179.035 196.090 433.415 ; 
                RECT 198.010 179.035 199.930 433.415 ; 
                RECT 201.850 179.035 203.770 433.415 ; 
                RECT 205.690 179.035 207.610 433.415 ; 
                RECT 209.530 179.035 211.450 433.415 ; 
                RECT 213.370 179.035 215.290 433.415 ; 
                RECT 217.210 179.035 219.130 433.415 ; 
                RECT 151.735 61.485 153.655 114.085 ; 
                RECT 158.255 61.485 159.795 114.085 ; 
                RECT 164.395 61.485 166.315 114.085 ; 
                RECT 173.105 61.485 175.025 114.085 ; 
                RECT 176.945 61.485 178.865 114.085 ; 
                RECT 191.505 61.485 193.425 114.085 ; 
                RECT 195.345 61.485 197.265 114.085 ; 
                RECT 199.185 61.485 201.105 114.085 ; 
                RECT 203.025 61.485 204.945 114.085 ; 
                RECT 164.830 139.540 166.750 172.400 ; 
                RECT 171.805 139.540 173.725 172.400 ; 
                RECT 178.435 139.540 180.185 172.400 ; 
                RECT 185.755 139.540 187.675 172.400 ; 
                RECT 196.630 139.540 198.550 172.400 ; 
                RECT 200.470 139.540 202.390 172.400 ; 
                RECT 204.310 139.540 206.230 172.400 ; 
                RECT 172.760 126.800 174.680 133.540 ; 
                RECT 181.240 126.800 183.160 133.540 ; 
                RECT 195.125 126.800 197.045 133.540 ; 
                RECT 198.965 126.800 200.885 133.540 ; 
                RECT 202.805 126.800 204.725 133.540 ; 
                RECT 204.145 51.905 206.065 55.485 ; 
                RECT 26.170 181.305 35.330 182.055 ; 
                RECT 26.170 186.060 35.330 187.980 ; 
                RECT 92.480 169.015 108.520 169.865 ; 
                RECT 73.280 169.355 90.520 171.385 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 234.040 5.560 ; 
                RECT 424.800 5.240 440.400 5.560 ; 
                RECT 2.880 6.600 440.400 6.920 ; 
                RECT 2.880 7.960 440.400 8.280 ; 
                RECT 2.880 9.320 208.200 9.640 ; 
                RECT 229.640 9.320 440.400 9.640 ; 
                RECT 2.880 10.680 223.840 11.000 ; 
                RECT 433.640 10.680 440.400 11.000 ; 
                RECT 2.880 12.040 223.840 12.360 ; 
                RECT 433.640 12.040 440.400 12.360 ; 
                RECT 2.880 13.400 223.840 13.720 ; 
                RECT 433.640 13.400 440.400 13.720 ; 
                RECT 2.880 14.760 223.840 15.080 ; 
                RECT 433.640 14.760 440.400 15.080 ; 
                RECT 2.880 16.120 223.840 16.440 ; 
                RECT 433.640 16.120 440.400 16.440 ; 
                RECT 2.880 17.480 223.840 17.800 ; 
                RECT 433.640 17.480 440.400 17.800 ; 
                RECT 2.880 18.840 223.840 19.160 ; 
                RECT 433.640 18.840 440.400 19.160 ; 
                RECT 2.880 20.200 223.840 20.520 ; 
                RECT 433.640 20.200 440.400 20.520 ; 
                RECT 2.880 21.560 140.200 21.880 ; 
                RECT 209.240 21.560 223.840 21.880 ; 
                RECT 433.640 21.560 440.400 21.880 ; 
                RECT 2.880 22.920 223.840 23.240 ; 
                RECT 433.640 22.920 440.400 23.240 ; 
                RECT 2.880 24.280 223.840 24.600 ; 
                RECT 433.640 24.280 440.400 24.600 ; 
                RECT 2.880 25.640 223.840 25.960 ; 
                RECT 433.640 25.640 440.400 25.960 ; 
                RECT 2.880 27.000 140.200 27.320 ; 
                RECT 208.560 27.000 223.840 27.320 ; 
                RECT 433.640 27.000 440.400 27.320 ; 
                RECT 2.880 28.360 223.160 28.680 ; 
                RECT 433.640 28.360 440.400 28.680 ; 
                RECT 2.880 29.720 223.840 30.040 ; 
                RECT 433.640 29.720 440.400 30.040 ; 
                RECT 2.880 31.080 223.840 31.400 ; 
                RECT 433.640 31.080 440.400 31.400 ; 
                RECT 2.880 32.440 223.840 32.760 ; 
                RECT 433.640 32.440 440.400 32.760 ; 
                RECT 2.880 33.800 223.840 34.120 ; 
                RECT 433.640 33.800 440.400 34.120 ; 
                RECT 2.880 35.160 223.840 35.480 ; 
                RECT 433.640 35.160 440.400 35.480 ; 
                RECT 2.880 36.520 223.840 36.840 ; 
                RECT 433.640 36.520 440.400 36.840 ; 
                RECT 2.880 37.880 223.840 38.200 ; 
                RECT 433.640 37.880 440.400 38.200 ; 
                RECT 2.880 39.240 223.840 39.560 ; 
                RECT 433.640 39.240 440.400 39.560 ; 
                RECT 2.880 40.600 223.840 40.920 ; 
                RECT 433.640 40.600 440.400 40.920 ; 
                RECT 2.880 41.960 223.840 42.280 ; 
                RECT 433.640 41.960 440.400 42.280 ; 
                RECT 2.880 43.320 223.840 43.640 ; 
                RECT 433.640 43.320 440.400 43.640 ; 
                RECT 2.880 44.680 138.160 45.000 ; 
                RECT 186.120 44.680 223.840 45.000 ; 
                RECT 433.640 44.680 440.400 45.000 ; 
                RECT 2.880 46.040 136.800 46.360 ; 
                RECT 192.240 46.040 223.840 46.360 ; 
                RECT 433.640 46.040 440.400 46.360 ; 
                RECT 2.880 47.400 117.760 47.720 ; 
                RECT 209.240 47.400 223.840 47.720 ; 
                RECT 433.640 47.400 440.400 47.720 ; 
                RECT 2.880 48.760 116.400 49.080 ; 
                RECT 205.160 48.760 223.840 49.080 ; 
                RECT 433.640 48.760 440.400 49.080 ; 
                RECT 2.880 50.120 223.840 50.440 ; 
                RECT 433.640 50.120 440.400 50.440 ; 
                RECT 2.880 51.480 200.040 51.800 ; 
                RECT 206.520 51.480 223.840 51.800 ; 
                RECT 433.640 51.480 440.400 51.800 ; 
                RECT 2.880 52.840 200.040 53.160 ; 
                RECT 206.520 52.840 223.840 53.160 ; 
                RECT 433.640 52.840 440.400 53.160 ; 
                RECT 2.880 54.200 200.040 54.520 ; 
                RECT 206.520 54.200 223.840 54.520 ; 
                RECT 433.640 54.200 440.400 54.520 ; 
                RECT 2.880 55.560 200.040 55.880 ; 
                RECT 206.520 55.560 223.840 55.880 ; 
                RECT 433.640 55.560 440.400 55.880 ; 
                RECT 2.880 56.920 223.840 57.240 ; 
                RECT 433.640 56.920 440.400 57.240 ; 
                RECT 2.880 58.280 223.840 58.600 ; 
                RECT 433.640 58.280 440.400 58.600 ; 
                RECT 2.880 59.640 223.840 59.960 ; 
                RECT 433.640 59.640 440.400 59.960 ; 
                RECT 2.880 61.000 148.360 61.320 ; 
                RECT 205.840 61.000 223.840 61.320 ; 
                RECT 433.640 61.000 440.400 61.320 ; 
                RECT 2.880 62.360 137.480 62.680 ; 
                RECT 142.600 62.360 148.360 62.680 ; 
                RECT 205.840 62.360 223.840 62.680 ; 
                RECT 433.640 62.360 440.400 62.680 ; 
                RECT 2.880 63.720 138.840 64.040 ; 
                RECT 141.240 63.720 148.360 64.040 ; 
                RECT 216.040 63.720 223.840 64.040 ; 
                RECT 433.640 63.720 440.400 64.040 ; 
                RECT 2.880 65.080 148.360 65.400 ; 
                RECT 216.040 65.080 223.840 65.400 ; 
                RECT 433.640 65.080 440.400 65.400 ; 
                RECT 2.880 66.440 148.360 66.760 ; 
                RECT 205.840 66.440 223.840 66.760 ; 
                RECT 433.640 66.440 440.400 66.760 ; 
                RECT 2.880 67.800 148.360 68.120 ; 
                RECT 214.680 67.800 223.840 68.120 ; 
                RECT 433.640 67.800 440.400 68.120 ; 
                RECT 2.880 69.160 148.360 69.480 ; 
                RECT 216.040 69.160 223.840 69.480 ; 
                RECT 433.640 69.160 440.400 69.480 ; 
                RECT 2.880 70.520 148.360 70.840 ; 
                RECT 205.840 70.520 223.840 70.840 ; 
                RECT 433.640 70.520 440.400 70.840 ; 
                RECT 2.880 71.880 113.000 72.200 ; 
                RECT 123.560 71.880 148.360 72.200 ; 
                RECT 216.040 71.880 223.840 72.200 ; 
                RECT 433.640 71.880 440.400 72.200 ; 
                RECT 2.880 73.240 114.360 73.560 ; 
                RECT 118.120 73.240 148.360 73.560 ; 
                RECT 216.040 73.240 223.840 73.560 ; 
                RECT 433.640 73.240 440.400 73.560 ; 
                RECT 2.880 74.600 115.720 74.920 ; 
                RECT 120.160 74.600 127.960 74.920 ; 
                RECT 130.360 74.600 148.360 74.920 ; 
                RECT 214.680 74.600 223.840 74.920 ; 
                RECT 433.640 74.600 440.400 74.920 ; 
                RECT 2.880 75.960 148.360 76.280 ; 
                RECT 218.760 75.960 223.840 76.280 ; 
                RECT 433.640 75.960 440.400 76.280 ; 
                RECT 2.880 77.320 122.520 77.640 ; 
                RECT 131.040 77.320 148.360 77.640 ; 
                RECT 218.760 77.320 223.840 77.640 ; 
                RECT 433.640 77.320 440.400 77.640 ; 
                RECT 2.880 78.680 115.040 79.000 ; 
                RECT 123.560 78.680 148.360 79.000 ; 
                RECT 217.400 78.680 223.840 79.000 ; 
                RECT 433.640 78.680 440.400 79.000 ; 
                RECT 2.880 80.040 118.440 80.360 ; 
                RECT 123.560 80.040 148.360 80.360 ; 
                RECT 218.760 80.040 223.840 80.360 ; 
                RECT 433.640 80.040 440.400 80.360 ; 
                RECT 2.880 81.400 148.360 81.720 ; 
                RECT 217.400 81.400 223.840 81.720 ; 
                RECT 433.640 81.400 440.400 81.720 ; 
                RECT 2.880 82.760 112.320 83.080 ; 
                RECT 123.560 82.760 148.360 83.080 ; 
                RECT 218.760 82.760 223.840 83.080 ; 
                RECT 433.640 82.760 440.400 83.080 ; 
                RECT 2.880 84.120 122.520 84.440 ; 
                RECT 129.680 84.120 148.360 84.440 ; 
                RECT 218.760 84.120 223.840 84.440 ; 
                RECT 433.640 84.120 440.400 84.440 ; 
                RECT 2.880 85.480 121.160 85.800 ; 
                RECT 123.560 85.480 148.360 85.800 ; 
                RECT 217.400 85.480 223.840 85.800 ; 
                RECT 433.640 85.480 440.400 85.800 ; 
                RECT 2.880 86.840 148.360 87.160 ; 
                RECT 218.760 86.840 223.840 87.160 ; 
                RECT 433.640 86.840 440.400 87.160 ; 
                RECT 2.880 88.200 122.520 88.520 ; 
                RECT 130.360 88.200 148.360 88.520 ; 
                RECT 205.840 88.200 223.840 88.520 ; 
                RECT 433.640 88.200 440.400 88.520 ; 
                RECT 2.880 89.560 119.120 89.880 ; 
                RECT 123.560 89.560 148.360 89.880 ; 
                RECT 221.480 89.560 223.840 89.880 ; 
                RECT 433.640 89.560 440.400 89.880 ; 
                RECT 2.880 90.920 121.160 91.240 ; 
                RECT 123.560 90.920 148.360 91.240 ; 
                RECT 221.480 90.920 223.840 91.240 ; 
                RECT 433.640 90.920 440.400 91.240 ; 
                RECT 2.880 92.280 125.240 92.600 ; 
                RECT 135.120 92.280 148.360 92.600 ; 
                RECT 221.480 92.280 223.840 92.600 ; 
                RECT 433.640 92.280 440.400 92.600 ; 
                RECT 2.880 93.640 112.320 93.960 ; 
                RECT 130.360 93.640 148.360 93.960 ; 
                RECT 220.120 93.640 223.840 93.960 ; 
                RECT 433.640 93.640 440.400 93.960 ; 
                RECT 2.880 95.000 121.160 95.320 ; 
                RECT 123.560 95.000 130.680 95.320 ; 
                RECT 136.480 95.000 148.360 95.320 ; 
                RECT 221.480 95.000 223.840 95.320 ; 
                RECT 433.640 95.000 440.400 95.320 ; 
                RECT 2.880 96.360 133.400 96.680 ; 
                RECT 137.160 96.360 148.360 96.680 ; 
                RECT 205.840 96.360 223.840 96.680 ; 
                RECT 433.640 96.360 440.400 96.680 ; 
                RECT 2.880 97.720 113.000 98.040 ; 
                RECT 126.960 97.720 148.360 98.040 ; 
                RECT 221.480 97.720 223.840 98.040 ; 
                RECT 433.640 97.720 440.400 98.040 ; 
                RECT 2.880 99.080 121.840 99.400 ; 
                RECT 130.360 99.080 148.360 99.400 ; 
                RECT 221.480 99.080 223.840 99.400 ; 
                RECT 433.640 99.080 440.400 99.400 ; 
                RECT 2.880 100.440 119.120 100.760 ; 
                RECT 131.040 100.440 148.360 100.760 ; 
                RECT 220.120 100.440 223.840 100.760 ; 
                RECT 433.640 100.440 440.400 100.760 ; 
                RECT 2.880 101.800 148.360 102.120 ; 
                RECT 433.640 101.800 440.400 102.120 ; 
                RECT 2.880 103.160 115.040 103.480 ; 
                RECT 118.120 103.160 148.360 103.480 ; 
                RECT 433.640 103.160 440.400 103.480 ; 
                RECT 2.880 104.520 115.040 104.840 ; 
                RECT 123.560 104.520 148.360 104.840 ; 
                RECT 433.640 104.520 440.400 104.840 ; 
                RECT 2.880 105.880 117.760 106.200 ; 
                RECT 120.840 105.880 148.360 106.200 ; 
                RECT 433.640 105.880 440.400 106.200 ; 
                RECT 2.880 107.240 148.360 107.560 ; 
                RECT 433.640 107.240 440.400 107.560 ; 
                RECT 2.880 108.600 121.160 108.920 ; 
                RECT 123.560 108.600 148.360 108.920 ; 
                RECT 433.640 108.600 440.400 108.920 ; 
                RECT 2.880 109.960 114.360 110.280 ; 
                RECT 129.680 109.960 148.360 110.280 ; 
                RECT 433.640 109.960 440.400 110.280 ; 
                RECT 2.880 111.320 121.160 111.640 ; 
                RECT 123.560 111.320 148.360 111.640 ; 
                RECT 205.840 111.320 223.840 111.640 ; 
                RECT 433.640 111.320 440.400 111.640 ; 
                RECT 2.880 112.680 148.360 113.000 ; 
                RECT 433.640 112.680 440.400 113.000 ; 
                RECT 2.880 114.040 116.400 114.360 ; 
                RECT 123.560 114.040 148.360 114.360 ; 
                RECT 205.840 114.040 223.840 114.360 ; 
                RECT 433.640 114.040 440.400 114.360 ; 
                RECT 2.880 115.400 113.000 115.720 ; 
                RECT 124.240 115.400 223.840 115.720 ; 
                RECT 433.640 115.400 440.400 115.720 ; 
                RECT 2.880 116.760 210.240 117.080 ; 
                RECT 433.640 116.760 440.400 117.080 ; 
                RECT 2.880 118.120 112.320 118.440 ; 
                RECT 130.360 118.120 221.120 118.440 ; 
                RECT 433.640 118.120 440.400 118.440 ; 
                RECT 2.880 119.480 109.600 119.800 ; 
                RECT 122.880 119.480 127.960 119.800 ; 
                RECT 130.360 119.480 218.400 119.800 ; 
                RECT 433.640 119.480 440.400 119.800 ; 
                RECT 2.880 120.840 113.000 121.160 ; 
                RECT 126.960 120.840 215.680 121.160 ; 
                RECT 433.640 120.840 440.400 121.160 ; 
                RECT 2.880 122.200 91.240 122.520 ; 
                RECT 109.960 122.200 212.960 122.520 ; 
                RECT 433.640 122.200 440.400 122.520 ; 
                RECT 2.880 123.560 91.240 123.880 ; 
                RECT 109.960 123.560 212.960 123.880 ; 
                RECT 433.640 123.560 440.400 123.880 ; 
                RECT 2.880 124.920 91.240 125.240 ; 
                RECT 109.960 124.920 125.240 125.240 ; 
                RECT 132.400 124.920 223.840 125.240 ; 
                RECT 433.640 124.920 440.400 125.240 ; 
                RECT 2.880 126.280 91.240 126.600 ; 
                RECT 109.960 126.280 168.760 126.600 ; 
                RECT 205.160 126.280 223.840 126.600 ; 
                RECT 433.640 126.280 440.400 126.600 ; 
                RECT 2.880 127.640 91.240 127.960 ; 
                RECT 109.960 127.640 168.760 127.960 ; 
                RECT 205.160 127.640 223.840 127.960 ; 
                RECT 433.640 127.640 440.400 127.960 ; 
                RECT 2.880 129.000 91.240 129.320 ; 
                RECT 109.960 129.000 115.040 129.320 ; 
                RECT 118.120 129.000 168.760 129.320 ; 
                RECT 205.160 129.000 223.840 129.320 ; 
                RECT 433.640 129.000 440.400 129.320 ; 
                RECT 2.880 130.360 91.240 130.680 ; 
                RECT 109.960 130.360 112.320 130.680 ; 
                RECT 130.360 130.360 168.760 130.680 ; 
                RECT 205.160 130.360 223.840 130.680 ; 
                RECT 433.640 130.360 440.400 130.680 ; 
                RECT 2.880 131.720 91.240 132.040 ; 
                RECT 109.960 131.720 168.760 132.040 ; 
                RECT 205.160 131.720 223.840 132.040 ; 
                RECT 433.640 131.720 440.400 132.040 ; 
                RECT 2.880 133.080 91.240 133.400 ; 
                RECT 109.960 133.080 168.760 133.400 ; 
                RECT 205.160 133.080 223.840 133.400 ; 
                RECT 433.640 133.080 440.400 133.400 ; 
                RECT 2.880 134.440 91.240 134.760 ; 
                RECT 109.960 134.440 223.840 134.760 ; 
                RECT 433.640 134.440 440.400 134.760 ; 
                RECT 2.880 135.800 91.240 136.120 ; 
                RECT 109.960 135.800 223.840 136.120 ; 
                RECT 433.640 135.800 440.400 136.120 ; 
                RECT 2.880 137.160 91.240 137.480 ; 
                RECT 109.960 137.160 223.840 137.480 ; 
                RECT 433.640 137.160 440.400 137.480 ; 
                RECT 2.880 138.520 91.240 138.840 ; 
                RECT 109.960 138.520 115.040 138.840 ; 
                RECT 119.480 138.520 127.960 138.840 ; 
                RECT 131.040 138.520 223.840 138.840 ; 
                RECT 433.640 138.520 440.400 138.840 ; 
                RECT 2.880 139.880 91.240 140.200 ; 
                RECT 110.640 139.880 161.280 140.200 ; 
                RECT 207.200 139.880 223.840 140.200 ; 
                RECT 433.640 139.880 440.400 140.200 ; 
                RECT 2.880 141.240 91.240 141.560 ; 
                RECT 109.960 141.240 161.280 141.560 ; 
                RECT 207.200 141.240 223.840 141.560 ; 
                RECT 433.640 141.240 440.400 141.560 ; 
                RECT 2.880 142.600 91.240 142.920 ; 
                RECT 109.960 142.600 161.280 142.920 ; 
                RECT 207.200 142.600 223.840 142.920 ; 
                RECT 433.640 142.600 440.400 142.920 ; 
                RECT 2.880 143.960 91.240 144.280 ; 
                RECT 109.960 143.960 161.280 144.280 ; 
                RECT 207.200 143.960 223.840 144.280 ; 
                RECT 433.640 143.960 440.400 144.280 ; 
                RECT 2.880 145.320 91.240 145.640 ; 
                RECT 109.960 145.320 114.360 145.640 ; 
                RECT 117.440 145.320 161.280 145.640 ; 
                RECT 207.200 145.320 223.840 145.640 ; 
                RECT 433.640 145.320 440.400 145.640 ; 
                RECT 2.880 146.680 91.240 147.000 ; 
                RECT 109.960 146.680 161.280 147.000 ; 
                RECT 207.200 146.680 223.840 147.000 ; 
                RECT 433.640 146.680 440.400 147.000 ; 
                RECT 2.880 148.040 91.240 148.360 ; 
                RECT 109.960 148.040 121.160 148.360 ; 
                RECT 129.680 148.040 161.280 148.360 ; 
                RECT 207.200 148.040 223.840 148.360 ; 
                RECT 433.640 148.040 440.400 148.360 ; 
                RECT 2.880 149.400 91.240 149.720 ; 
                RECT 109.960 149.400 161.280 149.720 ; 
                RECT 207.200 149.400 214.320 149.720 ; 
                RECT 433.640 149.400 440.400 149.720 ; 
                RECT 2.880 150.760 91.240 151.080 ; 
                RECT 109.960 150.760 117.760 151.080 ; 
                RECT 120.160 150.760 161.280 151.080 ; 
                RECT 207.200 150.760 217.040 151.080 ; 
                RECT 433.640 150.760 440.400 151.080 ; 
                RECT 2.880 152.120 91.240 152.440 ; 
                RECT 109.960 152.120 161.280 152.440 ; 
                RECT 207.200 152.120 219.760 152.440 ; 
                RECT 433.640 152.120 440.400 152.440 ; 
                RECT 2.880 153.480 91.240 153.800 ; 
                RECT 109.960 153.480 161.280 153.800 ; 
                RECT 207.200 153.480 222.480 153.800 ; 
                RECT 433.640 153.480 440.400 153.800 ; 
                RECT 2.880 154.840 91.240 155.160 ; 
                RECT 109.960 154.840 161.280 155.160 ; 
                RECT 433.640 154.840 440.400 155.160 ; 
                RECT 2.880 156.200 91.240 156.520 ; 
                RECT 109.960 156.200 161.280 156.520 ; 
                RECT 207.200 156.200 223.840 156.520 ; 
                RECT 433.640 156.200 440.400 156.520 ; 
                RECT 2.880 157.560 91.240 157.880 ; 
                RECT 109.960 157.560 161.280 157.880 ; 
                RECT 207.200 157.560 223.840 157.880 ; 
                RECT 433.640 157.560 440.400 157.880 ; 
                RECT 2.880 158.920 91.240 159.240 ; 
                RECT 109.960 158.920 161.280 159.240 ; 
                RECT 207.200 158.920 223.840 159.240 ; 
                RECT 433.640 158.920 440.400 159.240 ; 
                RECT 2.880 160.280 91.240 160.600 ; 
                RECT 109.960 160.280 161.280 160.600 ; 
                RECT 207.200 160.280 223.840 160.600 ; 
                RECT 433.640 160.280 440.400 160.600 ; 
                RECT 2.880 161.640 116.400 161.960 ; 
                RECT 120.160 161.640 161.280 161.960 ; 
                RECT 207.200 161.640 223.840 161.960 ; 
                RECT 433.640 161.640 440.400 161.960 ; 
                RECT 2.880 163.000 161.280 163.320 ; 
                RECT 207.200 163.000 223.840 163.320 ; 
                RECT 433.640 163.000 440.400 163.320 ; 
                RECT 2.880 164.360 161.280 164.680 ; 
                RECT 207.200 164.360 223.840 164.680 ; 
                RECT 433.640 164.360 440.400 164.680 ; 
                RECT 2.880 165.720 72.880 166.040 ; 
                RECT 90.920 165.720 118.440 166.040 ; 
                RECT 124.240 165.720 161.280 166.040 ; 
                RECT 207.200 165.720 223.840 166.040 ; 
                RECT 433.640 165.720 440.400 166.040 ; 
                RECT 2.880 167.080 72.880 167.400 ; 
                RECT 90.920 167.080 97.360 167.400 ; 
                RECT 104.520 167.080 161.280 167.400 ; 
                RECT 207.200 167.080 223.840 167.400 ; 
                RECT 433.640 167.080 440.400 167.400 ; 
                RECT 2.880 168.440 72.880 168.760 ; 
                RECT 90.920 168.440 91.920 168.760 ; 
                RECT 109.280 168.440 161.280 168.760 ; 
                RECT 207.200 168.440 223.840 168.760 ; 
                RECT 433.640 168.440 440.400 168.760 ; 
                RECT 2.880 169.800 72.880 170.120 ; 
                RECT 90.920 169.800 91.920 170.120 ; 
                RECT 109.280 169.800 161.280 170.120 ; 
                RECT 433.640 169.800 440.400 170.120 ; 
                RECT 2.880 171.160 72.880 171.480 ; 
                RECT 90.920 171.160 97.360 171.480 ; 
                RECT 104.520 171.160 113.000 171.480 ; 
                RECT 122.880 171.160 161.280 171.480 ; 
                RECT 433.640 171.160 440.400 171.480 ; 
                RECT 2.880 172.520 69.480 172.840 ; 
                RECT 103.840 172.520 161.280 172.840 ; 
                RECT 207.200 172.520 440.400 172.840 ; 
                RECT 2.880 173.880 103.480 174.200 ; 
                RECT 158.240 173.880 440.400 174.200 ; 
                RECT 2.880 175.240 221.120 175.560 ; 
                RECT 435.680 175.240 440.400 175.560 ; 
                RECT 2.880 176.600 221.120 176.920 ; 
                RECT 435.680 176.600 440.400 176.920 ; 
                RECT 2.880 177.960 221.120 178.280 ; 
                RECT 435.680 177.960 440.400 178.280 ; 
                RECT 2.880 179.320 27.320 179.640 ; 
                RECT 33.800 179.320 36.160 179.640 ; 
                RECT 48.760 179.320 99.400 179.640 ; 
                RECT 435.680 179.320 440.400 179.640 ; 
                RECT 2.880 180.680 25.280 181.000 ; 
                RECT 48.080 180.680 59.280 181.000 ; 
                RECT 61.000 180.680 75.600 181.000 ; 
                RECT 89.560 180.680 99.400 181.000 ; 
                RECT 435.680 180.680 440.400 181.000 ; 
                RECT 2.880 182.040 25.280 182.360 ; 
                RECT 35.840 182.040 59.280 182.360 ; 
                RECT 63.720 182.040 75.600 182.360 ; 
                RECT 89.560 182.040 99.400 182.360 ; 
                RECT 435.680 182.040 440.400 182.360 ; 
                RECT 2.880 183.400 25.280 183.720 ; 
                RECT 35.840 183.400 59.280 183.720 ; 
                RECT 63.720 183.400 75.600 183.720 ; 
                RECT 89.560 183.400 99.400 183.720 ; 
                RECT 435.680 183.400 440.400 183.720 ; 
                RECT 2.880 184.760 59.280 185.080 ; 
                RECT 64.400 184.760 75.600 185.080 ; 
                RECT 89.560 184.760 99.400 185.080 ; 
                RECT 435.680 184.760 440.400 185.080 ; 
                RECT 2.880 186.120 25.280 186.440 ; 
                RECT 35.840 186.120 59.280 186.440 ; 
                RECT 61.000 186.120 75.600 186.440 ; 
                RECT 89.560 186.120 99.400 186.440 ; 
                RECT 435.680 186.120 440.400 186.440 ; 
                RECT 2.880 187.480 25.280 187.800 ; 
                RECT 35.840 187.480 99.400 187.800 ; 
                RECT 435.680 187.480 440.400 187.800 ; 
                RECT 2.880 188.840 75.600 189.160 ; 
                RECT 89.560 188.840 99.400 189.160 ; 
                RECT 435.680 188.840 440.400 189.160 ; 
                RECT 2.880 190.200 75.600 190.520 ; 
                RECT 89.560 190.200 99.400 190.520 ; 
                RECT 435.680 190.200 440.400 190.520 ; 
                RECT 2.880 191.560 75.600 191.880 ; 
                RECT 89.560 191.560 99.400 191.880 ; 
                RECT 435.680 191.560 440.400 191.880 ; 
                RECT 2.880 192.920 18.480 193.240 ; 
                RECT 20.880 192.920 34.120 193.240 ; 
                RECT 37.200 192.920 75.600 193.240 ; 
                RECT 89.560 192.920 99.400 193.240 ; 
                RECT 435.680 192.920 440.400 193.240 ; 
                RECT 2.880 194.280 17.800 194.600 ; 
                RECT 20.880 194.280 34.120 194.600 ; 
                RECT 37.880 194.280 75.600 194.600 ; 
                RECT 89.560 194.280 99.400 194.600 ; 
                RECT 435.680 194.280 440.400 194.600 ; 
                RECT 2.880 195.640 17.120 195.960 ; 
                RECT 20.880 195.640 39.560 195.960 ; 
                RECT 48.760 195.640 99.400 195.960 ; 
                RECT 435.680 195.640 440.400 195.960 ; 
                RECT 2.880 197.000 16.440 197.320 ; 
                RECT 20.880 197.000 40.920 197.320 ; 
                RECT 47.400 197.000 59.280 197.320 ; 
                RECT 61.000 197.000 75.600 197.320 ; 
                RECT 89.560 197.000 99.400 197.320 ; 
                RECT 435.680 197.000 440.400 197.320 ; 
                RECT 2.880 198.360 59.280 198.680 ; 
                RECT 61.680 198.360 75.600 198.680 ; 
                RECT 89.560 198.360 99.400 198.680 ; 
                RECT 435.680 198.360 440.400 198.680 ; 
                RECT 2.880 199.720 15.760 200.040 ; 
                RECT 20.880 199.720 59.280 200.040 ; 
                RECT 62.360 199.720 75.600 200.040 ; 
                RECT 89.560 199.720 99.400 200.040 ; 
                RECT 435.680 199.720 440.400 200.040 ; 
                RECT 2.880 201.080 15.080 201.400 ; 
                RECT 20.880 201.080 59.280 201.400 ; 
                RECT 62.360 201.080 75.600 201.400 ; 
                RECT 89.560 201.080 99.400 201.400 ; 
                RECT 435.680 201.080 440.400 201.400 ; 
                RECT 2.880 202.440 59.280 202.760 ; 
                RECT 63.040 202.440 75.600 202.760 ; 
                RECT 89.560 202.440 99.400 202.760 ; 
                RECT 435.680 202.440 440.400 202.760 ; 
                RECT 2.880 203.800 14.400 204.120 ; 
                RECT 20.880 203.800 99.400 204.120 ; 
                RECT 435.680 203.800 440.400 204.120 ; 
                RECT 2.880 205.160 13.720 205.480 ; 
                RECT 20.880 205.160 34.120 205.480 ; 
                RECT 41.960 205.160 75.600 205.480 ; 
                RECT 89.560 205.160 99.400 205.480 ; 
                RECT 435.680 205.160 440.400 205.480 ; 
                RECT 2.880 206.520 75.600 206.840 ; 
                RECT 89.560 206.520 99.400 206.840 ; 
                RECT 435.680 206.520 440.400 206.840 ; 
                RECT 2.880 207.880 13.040 208.200 ; 
                RECT 20.880 207.880 34.120 208.200 ; 
                RECT 40.600 207.880 75.600 208.200 ; 
                RECT 89.560 207.880 99.400 208.200 ; 
                RECT 435.680 207.880 440.400 208.200 ; 
                RECT 2.880 209.240 12.360 209.560 ; 
                RECT 20.880 209.240 34.120 209.560 ; 
                RECT 39.920 209.240 75.600 209.560 ; 
                RECT 89.560 209.240 99.400 209.560 ; 
                RECT 435.680 209.240 440.400 209.560 ; 
                RECT 2.880 210.600 11.680 210.920 ; 
                RECT 20.880 210.600 34.120 210.920 ; 
                RECT 39.240 210.600 75.600 210.920 ; 
                RECT 85.480 210.600 99.400 210.920 ; 
                RECT 435.680 210.600 440.400 210.920 ; 
                RECT 2.880 211.960 11.000 212.280 ; 
                RECT 20.880 211.960 80.360 212.280 ; 
                RECT 89.560 211.960 99.400 212.280 ; 
                RECT 435.680 211.960 440.400 212.280 ; 
                RECT 2.880 213.320 75.600 213.640 ; 
                RECT 89.560 213.320 99.400 213.640 ; 
                RECT 435.680 213.320 440.400 213.640 ; 
                RECT 2.880 214.680 10.320 215.000 ; 
                RECT 20.880 214.680 34.120 215.000 ; 
                RECT 37.880 214.680 75.600 215.000 ; 
                RECT 89.560 214.680 99.400 215.000 ; 
                RECT 435.680 214.680 440.400 215.000 ; 
                RECT 2.880 216.040 9.640 216.360 ; 
                RECT 20.880 216.040 75.600 216.360 ; 
                RECT 89.560 216.040 99.400 216.360 ; 
                RECT 435.680 216.040 440.400 216.360 ; 
                RECT 2.880 217.400 75.600 217.720 ; 
                RECT 89.560 217.400 99.400 217.720 ; 
                RECT 435.680 217.400 440.400 217.720 ; 
                RECT 2.880 218.760 75.600 219.080 ; 
                RECT 86.160 218.760 99.400 219.080 ; 
                RECT 435.680 218.760 440.400 219.080 ; 
                RECT 2.880 220.120 75.600 220.440 ; 
                RECT 89.560 220.120 99.400 220.440 ; 
                RECT 435.680 220.120 440.400 220.440 ; 
                RECT 2.880 221.480 75.600 221.800 ; 
                RECT 89.560 221.480 99.400 221.800 ; 
                RECT 435.680 221.480 440.400 221.800 ; 
                RECT 2.880 222.840 75.600 223.160 ; 
                RECT 89.560 222.840 99.400 223.160 ; 
                RECT 435.680 222.840 440.400 223.160 ; 
                RECT 2.880 224.200 75.600 224.520 ; 
                RECT 89.560 224.200 99.400 224.520 ; 
                RECT 435.680 224.200 440.400 224.520 ; 
                RECT 2.880 225.560 75.600 225.880 ; 
                RECT 89.560 225.560 99.400 225.880 ; 
                RECT 435.680 225.560 440.400 225.880 ; 
                RECT 2.880 226.920 75.600 227.240 ; 
                RECT 86.840 226.920 99.400 227.240 ; 
                RECT 435.680 226.920 440.400 227.240 ; 
                RECT 2.880 228.280 75.600 228.600 ; 
                RECT 89.560 228.280 99.400 228.600 ; 
                RECT 435.680 228.280 440.400 228.600 ; 
                RECT 2.880 229.640 75.600 229.960 ; 
                RECT 89.560 229.640 99.400 229.960 ; 
                RECT 435.680 229.640 440.400 229.960 ; 
                RECT 2.880 231.000 75.600 231.320 ; 
                RECT 89.560 231.000 99.400 231.320 ; 
                RECT 435.680 231.000 440.400 231.320 ; 
                RECT 2.880 232.360 75.600 232.680 ; 
                RECT 89.560 232.360 99.400 232.680 ; 
                RECT 435.680 232.360 440.400 232.680 ; 
                RECT 2.880 233.720 75.600 234.040 ; 
                RECT 89.560 233.720 99.400 234.040 ; 
                RECT 435.680 233.720 440.400 234.040 ; 
                RECT 2.880 235.080 99.400 235.400 ; 
                RECT 435.680 235.080 440.400 235.400 ; 
                RECT 2.880 236.440 75.600 236.760 ; 
                RECT 89.560 236.440 99.400 236.760 ; 
                RECT 435.680 236.440 440.400 236.760 ; 
                RECT 2.880 237.800 75.600 238.120 ; 
                RECT 89.560 237.800 99.400 238.120 ; 
                RECT 435.680 237.800 440.400 238.120 ; 
                RECT 2.880 239.160 75.600 239.480 ; 
                RECT 89.560 239.160 99.400 239.480 ; 
                RECT 435.680 239.160 440.400 239.480 ; 
                RECT 2.880 240.520 75.600 240.840 ; 
                RECT 89.560 240.520 99.400 240.840 ; 
                RECT 435.680 240.520 440.400 240.840 ; 
                RECT 2.880 241.880 75.600 242.200 ; 
                RECT 89.560 241.880 99.400 242.200 ; 
                RECT 435.680 241.880 440.400 242.200 ; 
                RECT 2.880 243.240 99.400 243.560 ; 
                RECT 435.680 243.240 440.400 243.560 ; 
                RECT 2.880 244.600 77.640 244.920 ; 
                RECT 89.560 244.600 99.400 244.920 ; 
                RECT 435.680 244.600 440.400 244.920 ; 
                RECT 2.880 245.960 77.640 246.280 ; 
                RECT 89.560 245.960 99.400 246.280 ; 
                RECT 435.680 245.960 440.400 246.280 ; 
                RECT 2.880 247.320 77.640 247.640 ; 
                RECT 89.560 247.320 99.400 247.640 ; 
                RECT 435.680 247.320 440.400 247.640 ; 
                RECT 2.880 248.680 81.720 249.000 ; 
                RECT 89.560 248.680 99.400 249.000 ; 
                RECT 435.680 248.680 440.400 249.000 ; 
                RECT 2.880 250.040 77.640 250.360 ; 
                RECT 89.560 250.040 99.400 250.360 ; 
                RECT 435.680 250.040 440.400 250.360 ; 
                RECT 2.880 251.400 38.880 251.720 ; 
                RECT 64.400 251.400 99.400 251.720 ; 
                RECT 435.680 251.400 440.400 251.720 ; 
                RECT 2.880 252.760 37.520 253.080 ; 
                RECT 63.720 252.760 75.600 253.080 ; 
                RECT 89.560 252.760 99.400 253.080 ; 
                RECT 435.680 252.760 440.400 253.080 ; 
                RECT 2.880 254.120 36.160 254.440 ; 
                RECT 63.040 254.120 75.600 254.440 ; 
                RECT 89.560 254.120 99.400 254.440 ; 
                RECT 435.680 254.120 440.400 254.440 ; 
                RECT 2.880 255.480 77.640 255.800 ; 
                RECT 89.560 255.480 99.400 255.800 ; 
                RECT 435.680 255.480 440.400 255.800 ; 
                RECT 2.880 256.840 75.600 257.160 ; 
                RECT 89.560 256.840 99.400 257.160 ; 
                RECT 435.680 256.840 440.400 257.160 ; 
                RECT 2.880 258.200 75.600 258.520 ; 
                RECT 78.000 258.200 99.400 258.520 ; 
                RECT 435.680 258.200 440.400 258.520 ; 
                RECT 2.880 259.560 83.760 259.880 ; 
                RECT 89.560 259.560 99.400 259.880 ; 
                RECT 435.680 259.560 440.400 259.880 ; 
                RECT 2.880 260.920 75.600 261.240 ; 
                RECT 89.560 260.920 99.400 261.240 ; 
                RECT 435.680 260.920 440.400 261.240 ; 
                RECT 2.880 262.280 75.600 262.600 ; 
                RECT 89.560 262.280 99.400 262.600 ; 
                RECT 435.680 262.280 440.400 262.600 ; 
                RECT 2.880 263.640 75.600 263.960 ; 
                RECT 89.560 263.640 99.400 263.960 ; 
                RECT 435.680 263.640 440.400 263.960 ; 
                RECT 2.880 265.000 75.600 265.320 ; 
                RECT 89.560 265.000 99.400 265.320 ; 
                RECT 435.680 265.000 440.400 265.320 ; 
                RECT 2.880 266.360 75.600 266.680 ; 
                RECT 78.680 266.360 99.400 266.680 ; 
                RECT 435.680 266.360 440.400 266.680 ; 
                RECT 2.880 267.720 85.800 268.040 ; 
                RECT 89.560 267.720 99.400 268.040 ; 
                RECT 435.680 267.720 440.400 268.040 ; 
                RECT 2.880 269.080 75.600 269.400 ; 
                RECT 89.560 269.080 99.400 269.400 ; 
                RECT 435.680 269.080 440.400 269.400 ; 
                RECT 2.880 270.440 75.600 270.760 ; 
                RECT 89.560 270.440 99.400 270.760 ; 
                RECT 435.680 270.440 440.400 270.760 ; 
                RECT 2.880 271.800 75.600 272.120 ; 
                RECT 89.560 271.800 99.400 272.120 ; 
                RECT 435.680 271.800 440.400 272.120 ; 
                RECT 2.880 273.160 75.600 273.480 ; 
                RECT 89.560 273.160 99.400 273.480 ; 
                RECT 435.680 273.160 440.400 273.480 ; 
                RECT 2.880 274.520 99.400 274.840 ; 
                RECT 435.680 274.520 440.400 274.840 ; 
                RECT 2.880 275.880 77.640 276.200 ; 
                RECT 89.560 275.880 99.400 276.200 ; 
                RECT 435.680 275.880 440.400 276.200 ; 
                RECT 2.880 277.240 75.600 277.560 ; 
                RECT 89.560 277.240 99.400 277.560 ; 
                RECT 435.680 277.240 440.400 277.560 ; 
                RECT 2.880 278.600 75.600 278.920 ; 
                RECT 89.560 278.600 99.400 278.920 ; 
                RECT 435.680 278.600 440.400 278.920 ; 
                RECT 2.880 279.960 75.600 280.280 ; 
                RECT 89.560 279.960 99.400 280.280 ; 
                RECT 435.680 279.960 440.400 280.280 ; 
                RECT 2.880 281.320 75.600 281.640 ; 
                RECT 89.560 281.320 99.400 281.640 ; 
                RECT 435.680 281.320 440.400 281.640 ; 
                RECT 2.880 282.680 99.400 283.000 ; 
                RECT 435.680 282.680 440.400 283.000 ; 
                RECT 2.880 284.040 77.640 284.360 ; 
                RECT 89.560 284.040 99.400 284.360 ; 
                RECT 435.680 284.040 440.400 284.360 ; 
                RECT 2.880 285.400 75.600 285.720 ; 
                RECT 89.560 285.400 99.400 285.720 ; 
                RECT 435.680 285.400 440.400 285.720 ; 
                RECT 2.880 286.760 75.600 287.080 ; 
                RECT 89.560 286.760 99.400 287.080 ; 
                RECT 435.680 286.760 440.400 287.080 ; 
                RECT 2.880 288.120 75.600 288.440 ; 
                RECT 89.560 288.120 99.400 288.440 ; 
                RECT 435.680 288.120 440.400 288.440 ; 
                RECT 2.880 289.480 75.600 289.800 ; 
                RECT 89.560 289.480 99.400 289.800 ; 
                RECT 435.680 289.480 440.400 289.800 ; 
                RECT 2.880 290.840 99.400 291.160 ; 
                RECT 435.680 290.840 440.400 291.160 ; 
                RECT 2.880 292.200 75.600 292.520 ; 
                RECT 89.560 292.200 99.400 292.520 ; 
                RECT 435.680 292.200 440.400 292.520 ; 
                RECT 2.880 293.560 75.600 293.880 ; 
                RECT 89.560 293.560 99.400 293.880 ; 
                RECT 435.680 293.560 440.400 293.880 ; 
                RECT 2.880 294.920 77.640 295.240 ; 
                RECT 89.560 294.920 99.400 295.240 ; 
                RECT 435.680 294.920 440.400 295.240 ; 
                RECT 2.880 296.280 75.600 296.600 ; 
                RECT 89.560 296.280 99.400 296.600 ; 
                RECT 435.680 296.280 440.400 296.600 ; 
                RECT 2.880 297.640 75.600 297.960 ; 
                RECT 80.720 297.640 99.400 297.960 ; 
                RECT 435.680 297.640 440.400 297.960 ; 
                RECT 2.880 299.000 85.800 299.320 ; 
                RECT 89.560 299.000 99.400 299.320 ; 
                RECT 435.680 299.000 440.400 299.320 ; 
                RECT 2.880 300.360 75.600 300.680 ; 
                RECT 89.560 300.360 99.400 300.680 ; 
                RECT 435.680 300.360 440.400 300.680 ; 
                RECT 2.880 301.720 75.600 302.040 ; 
                RECT 89.560 301.720 99.400 302.040 ; 
                RECT 435.680 301.720 440.400 302.040 ; 
                RECT 2.880 303.080 75.600 303.400 ; 
                RECT 89.560 303.080 99.400 303.400 ; 
                RECT 435.680 303.080 440.400 303.400 ; 
                RECT 2.880 304.440 75.600 304.760 ; 
                RECT 89.560 304.440 99.400 304.760 ; 
                RECT 435.680 304.440 440.400 304.760 ; 
                RECT 2.880 305.800 75.600 306.120 ; 
                RECT 80.720 305.800 99.400 306.120 ; 
                RECT 435.680 305.800 440.400 306.120 ; 
                RECT 2.880 307.160 80.360 307.480 ; 
                RECT 89.560 307.160 99.400 307.480 ; 
                RECT 435.680 307.160 440.400 307.480 ; 
                RECT 2.880 308.520 75.600 308.840 ; 
                RECT 89.560 308.520 99.400 308.840 ; 
                RECT 435.680 308.520 440.400 308.840 ; 
                RECT 2.880 309.880 75.600 310.200 ; 
                RECT 89.560 309.880 99.400 310.200 ; 
                RECT 435.680 309.880 440.400 310.200 ; 
                RECT 2.880 311.240 75.600 311.560 ; 
                RECT 89.560 311.240 99.400 311.560 ; 
                RECT 435.680 311.240 440.400 311.560 ; 
                RECT 2.880 312.600 75.600 312.920 ; 
                RECT 89.560 312.600 99.400 312.920 ; 
                RECT 435.680 312.600 440.400 312.920 ; 
                RECT 2.880 313.960 99.400 314.280 ; 
                RECT 435.680 313.960 440.400 314.280 ; 
                RECT 2.880 315.320 78.320 315.640 ; 
                RECT 89.560 315.320 99.400 315.640 ; 
                RECT 435.680 315.320 440.400 315.640 ; 
                RECT 2.880 316.680 82.400 317.000 ; 
                RECT 89.560 316.680 99.400 317.000 ; 
                RECT 435.680 316.680 440.400 317.000 ; 
                RECT 2.880 318.040 83.080 318.360 ; 
                RECT 89.560 318.040 99.400 318.360 ; 
                RECT 435.680 318.040 440.400 318.360 ; 
                RECT 2.880 319.400 78.320 319.720 ; 
                RECT 89.560 319.400 99.400 319.720 ; 
                RECT 435.680 319.400 440.400 319.720 ; 
                RECT 2.880 320.760 78.320 321.080 ; 
                RECT 89.560 320.760 99.400 321.080 ; 
                RECT 435.680 320.760 440.400 321.080 ; 
                RECT 2.880 322.120 99.400 322.440 ; 
                RECT 435.680 322.120 440.400 322.440 ; 
                RECT 2.880 323.480 78.320 323.800 ; 
                RECT 89.560 323.480 99.400 323.800 ; 
                RECT 435.680 323.480 440.400 323.800 ; 
                RECT 2.880 324.840 78.320 325.160 ; 
                RECT 89.560 324.840 99.400 325.160 ; 
                RECT 435.680 324.840 440.400 325.160 ; 
                RECT 2.880 326.200 78.320 326.520 ; 
                RECT 89.560 326.200 99.400 326.520 ; 
                RECT 435.680 326.200 440.400 326.520 ; 
                RECT 2.880 327.560 85.800 327.880 ; 
                RECT 89.560 327.560 99.400 327.880 ; 
                RECT 435.680 327.560 440.400 327.880 ; 
                RECT 2.880 328.920 78.320 329.240 ; 
                RECT 89.560 328.920 99.400 329.240 ; 
                RECT 435.680 328.920 440.400 329.240 ; 
                RECT 2.880 330.280 99.400 330.600 ; 
                RECT 435.680 330.280 440.400 330.600 ; 
                RECT 2.880 331.640 78.320 331.960 ; 
                RECT 89.560 331.640 99.400 331.960 ; 
                RECT 435.680 331.640 440.400 331.960 ; 
                RECT 2.880 333.000 78.320 333.320 ; 
                RECT 89.560 333.000 99.400 333.320 ; 
                RECT 435.680 333.000 440.400 333.320 ; 
                RECT 2.880 334.360 78.320 334.680 ; 
                RECT 89.560 334.360 99.400 334.680 ; 
                RECT 435.680 334.360 440.400 334.680 ; 
                RECT 2.880 335.720 78.320 336.040 ; 
                RECT 89.560 335.720 99.400 336.040 ; 
                RECT 435.680 335.720 440.400 336.040 ; 
                RECT 2.880 337.080 99.400 337.400 ; 
                RECT 435.680 337.080 440.400 337.400 ; 
                RECT 2.880 338.440 80.360 338.760 ; 
                RECT 89.560 338.440 99.400 338.760 ; 
                RECT 435.680 338.440 440.400 338.760 ; 
                RECT 2.880 339.800 79.000 340.120 ; 
                RECT 89.560 339.800 99.400 340.120 ; 
                RECT 435.680 339.800 440.400 340.120 ; 
                RECT 2.880 341.160 79.000 341.480 ; 
                RECT 89.560 341.160 99.400 341.480 ; 
                RECT 435.680 341.160 440.400 341.480 ; 
                RECT 2.880 342.520 79.000 342.840 ; 
                RECT 89.560 342.520 99.400 342.840 ; 
                RECT 435.680 342.520 440.400 342.840 ; 
                RECT 2.880 343.880 79.000 344.200 ; 
                RECT 89.560 343.880 99.400 344.200 ; 
                RECT 435.680 343.880 440.400 344.200 ; 
                RECT 2.880 345.240 99.400 345.560 ; 
                RECT 435.680 345.240 440.400 345.560 ; 
                RECT 2.880 346.600 82.400 346.920 ; 
                RECT 89.560 346.600 99.400 346.920 ; 
                RECT 435.680 346.600 440.400 346.920 ; 
                RECT 2.880 347.960 79.000 348.280 ; 
                RECT 89.560 347.960 99.400 348.280 ; 
                RECT 435.680 347.960 440.400 348.280 ; 
                RECT 2.880 349.320 79.000 349.640 ; 
                RECT 89.560 349.320 99.400 349.640 ; 
                RECT 435.680 349.320 440.400 349.640 ; 
                RECT 2.880 350.680 79.000 351.000 ; 
                RECT 89.560 350.680 99.400 351.000 ; 
                RECT 435.680 350.680 440.400 351.000 ; 
                RECT 2.880 352.040 79.000 352.360 ; 
                RECT 89.560 352.040 99.400 352.360 ; 
                RECT 435.680 352.040 440.400 352.360 ; 
                RECT 2.880 353.400 99.400 353.720 ; 
                RECT 435.680 353.400 440.400 353.720 ; 
                RECT 2.880 354.760 79.000 355.080 ; 
                RECT 89.560 354.760 99.400 355.080 ; 
                RECT 435.680 354.760 440.400 355.080 ; 
                RECT 2.880 356.120 84.440 356.440 ; 
                RECT 89.560 356.120 99.400 356.440 ; 
                RECT 435.680 356.120 440.400 356.440 ; 
                RECT 2.880 357.480 79.000 357.800 ; 
                RECT 89.560 357.480 99.400 357.800 ; 
                RECT 435.680 357.480 440.400 357.800 ; 
                RECT 2.880 358.840 79.000 359.160 ; 
                RECT 89.560 358.840 99.400 359.160 ; 
                RECT 435.680 358.840 440.400 359.160 ; 
                RECT 2.880 360.200 79.000 360.520 ; 
                RECT 89.560 360.200 99.400 360.520 ; 
                RECT 435.680 360.200 440.400 360.520 ; 
                RECT 2.880 361.560 99.400 361.880 ; 
                RECT 435.680 361.560 440.400 361.880 ; 
                RECT 2.880 362.920 79.000 363.240 ; 
                RECT 89.560 362.920 99.400 363.240 ; 
                RECT 435.680 362.920 440.400 363.240 ; 
                RECT 2.880 364.280 79.000 364.600 ; 
                RECT 89.560 364.280 99.400 364.600 ; 
                RECT 435.680 364.280 440.400 364.600 ; 
                RECT 2.880 365.640 87.160 365.960 ; 
                RECT 89.560 365.640 99.400 365.960 ; 
                RECT 435.680 365.640 440.400 365.960 ; 
                RECT 2.880 367.000 87.160 367.320 ; 
                RECT 89.560 367.000 99.400 367.320 ; 
                RECT 435.680 367.000 440.400 367.320 ; 
                RECT 2.880 368.360 79.000 368.680 ; 
                RECT 89.560 368.360 99.400 368.680 ; 
                RECT 435.680 368.360 440.400 368.680 ; 
                RECT 2.880 369.720 99.400 370.040 ; 
                RECT 435.680 369.720 440.400 370.040 ; 
                RECT 2.880 371.080 79.000 371.400 ; 
                RECT 89.560 371.080 99.400 371.400 ; 
                RECT 435.680 371.080 440.400 371.400 ; 
                RECT 2.880 372.440 79.000 372.760 ; 
                RECT 89.560 372.440 99.400 372.760 ; 
                RECT 435.680 372.440 440.400 372.760 ; 
                RECT 2.880 373.800 79.000 374.120 ; 
                RECT 89.560 373.800 99.400 374.120 ; 
                RECT 435.680 373.800 440.400 374.120 ; 
                RECT 2.880 375.160 81.720 375.480 ; 
                RECT 89.560 375.160 99.400 375.480 ; 
                RECT 435.680 375.160 440.400 375.480 ; 
                RECT 2.880 376.520 99.400 376.840 ; 
                RECT 435.680 376.520 440.400 376.840 ; 
                RECT 2.880 377.880 82.400 378.200 ; 
                RECT 89.560 377.880 99.400 378.200 ; 
                RECT 435.680 377.880 440.400 378.200 ; 
                RECT 2.880 379.240 79.000 379.560 ; 
                RECT 89.560 379.240 99.400 379.560 ; 
                RECT 435.680 379.240 440.400 379.560 ; 
                RECT 2.880 380.600 79.000 380.920 ; 
                RECT 89.560 380.600 99.400 380.920 ; 
                RECT 435.680 380.600 440.400 380.920 ; 
                RECT 2.880 381.960 79.000 382.280 ; 
                RECT 89.560 381.960 99.400 382.280 ; 
                RECT 435.680 381.960 440.400 382.280 ; 
                RECT 2.880 383.320 79.000 383.640 ; 
                RECT 89.560 383.320 99.400 383.640 ; 
                RECT 435.680 383.320 440.400 383.640 ; 
                RECT 2.880 384.680 99.400 385.000 ; 
                RECT 435.680 384.680 440.400 385.000 ; 
                RECT 2.880 386.040 83.760 386.360 ; 
                RECT 89.560 386.040 99.400 386.360 ; 
                RECT 435.680 386.040 440.400 386.360 ; 
                RECT 2.880 387.400 79.000 387.720 ; 
                RECT 89.560 387.400 99.400 387.720 ; 
                RECT 435.680 387.400 440.400 387.720 ; 
                RECT 2.880 388.760 79.000 389.080 ; 
                RECT 89.560 388.760 99.400 389.080 ; 
                RECT 435.680 388.760 440.400 389.080 ; 
                RECT 2.880 390.120 79.000 390.440 ; 
                RECT 89.560 390.120 99.400 390.440 ; 
                RECT 435.680 390.120 440.400 390.440 ; 
                RECT 2.880 391.480 79.000 391.800 ; 
                RECT 89.560 391.480 99.400 391.800 ; 
                RECT 435.680 391.480 440.400 391.800 ; 
                RECT 2.880 392.840 99.400 393.160 ; 
                RECT 435.680 392.840 440.400 393.160 ; 
                RECT 2.880 394.200 79.000 394.520 ; 
                RECT 89.560 394.200 99.400 394.520 ; 
                RECT 435.680 394.200 440.400 394.520 ; 
                RECT 2.880 395.560 86.480 395.880 ; 
                RECT 89.560 395.560 99.400 395.880 ; 
                RECT 435.680 395.560 440.400 395.880 ; 
                RECT 2.880 396.920 79.000 397.240 ; 
                RECT 89.560 396.920 99.400 397.240 ; 
                RECT 435.680 396.920 440.400 397.240 ; 
                RECT 2.880 398.280 79.000 398.600 ; 
                RECT 89.560 398.280 99.400 398.600 ; 
                RECT 435.680 398.280 440.400 398.600 ; 
                RECT 2.880 399.640 79.000 399.960 ; 
                RECT 89.560 399.640 99.400 399.960 ; 
                RECT 435.680 399.640 440.400 399.960 ; 
                RECT 2.880 401.000 99.400 401.320 ; 
                RECT 435.680 401.000 440.400 401.320 ; 
                RECT 2.880 402.360 79.680 402.680 ; 
                RECT 89.560 402.360 99.400 402.680 ; 
                RECT 435.680 402.360 440.400 402.680 ; 
                RECT 2.880 403.720 79.680 404.040 ; 
                RECT 89.560 403.720 99.400 404.040 ; 
                RECT 435.680 403.720 440.400 404.040 ; 
                RECT 2.880 405.080 81.040 405.400 ; 
                RECT 89.560 405.080 99.400 405.400 ; 
                RECT 435.680 405.080 440.400 405.400 ; 
                RECT 2.880 406.440 79.680 406.760 ; 
                RECT 89.560 406.440 99.400 406.760 ; 
                RECT 435.680 406.440 440.400 406.760 ; 
                RECT 2.880 407.800 79.680 408.120 ; 
                RECT 89.560 407.800 99.400 408.120 ; 
                RECT 435.680 407.800 440.400 408.120 ; 
                RECT 2.880 409.160 99.400 409.480 ; 
                RECT 435.680 409.160 440.400 409.480 ; 
                RECT 2.880 410.520 79.680 410.840 ; 
                RECT 89.560 410.520 99.400 410.840 ; 
                RECT 435.680 410.520 440.400 410.840 ; 
                RECT 2.880 411.880 79.680 412.200 ; 
                RECT 89.560 411.880 99.400 412.200 ; 
                RECT 435.680 411.880 440.400 412.200 ; 
                RECT 2.880 413.240 79.680 413.560 ; 
                RECT 89.560 413.240 99.400 413.560 ; 
                RECT 435.680 413.240 440.400 413.560 ; 
                RECT 2.880 414.600 83.760 414.920 ; 
                RECT 89.560 414.600 99.400 414.920 ; 
                RECT 435.680 414.600 440.400 414.920 ; 
                RECT 2.880 415.960 79.680 416.280 ; 
                RECT 89.560 415.960 99.400 416.280 ; 
                RECT 435.680 415.960 440.400 416.280 ; 
                RECT 2.880 417.320 99.400 417.640 ; 
                RECT 435.680 417.320 440.400 417.640 ; 
                RECT 2.880 418.680 79.680 419.000 ; 
                RECT 89.560 418.680 99.400 419.000 ; 
                RECT 435.680 418.680 440.400 419.000 ; 
                RECT 2.880 420.040 79.680 420.360 ; 
                RECT 89.560 420.040 99.400 420.360 ; 
                RECT 435.680 420.040 440.400 420.360 ; 
                RECT 2.880 421.400 79.680 421.720 ; 
                RECT 89.560 421.400 99.400 421.720 ; 
                RECT 435.680 421.400 440.400 421.720 ; 
                RECT 2.880 422.760 79.680 423.080 ; 
                RECT 89.560 422.760 99.400 423.080 ; 
                RECT 435.680 422.760 440.400 423.080 ; 
                RECT 2.880 424.120 99.400 424.440 ; 
                RECT 435.680 424.120 440.400 424.440 ; 
                RECT 2.880 425.480 85.800 425.800 ; 
                RECT 89.560 425.480 99.400 425.800 ; 
                RECT 435.680 425.480 440.400 425.800 ; 
                RECT 2.880 426.840 79.680 427.160 ; 
                RECT 89.560 426.840 99.400 427.160 ; 
                RECT 435.680 426.840 440.400 427.160 ; 
                RECT 2.880 428.200 79.680 428.520 ; 
                RECT 89.560 428.200 99.400 428.520 ; 
                RECT 435.680 428.200 440.400 428.520 ; 
                RECT 2.880 429.560 79.680 429.880 ; 
                RECT 89.560 429.560 99.400 429.880 ; 
                RECT 435.680 429.560 440.400 429.880 ; 
                RECT 2.880 430.920 79.680 431.240 ; 
                RECT 89.560 430.920 99.400 431.240 ; 
                RECT 435.680 430.920 440.400 431.240 ; 
                RECT 2.880 432.280 99.400 432.600 ; 
                RECT 435.680 432.280 440.400 432.600 ; 
                RECT 2.880 433.640 99.400 433.960 ; 
                RECT 435.680 433.640 440.400 433.960 ; 
                RECT 2.880 435.000 221.120 435.320 ; 
                RECT 435.680 435.000 440.400 435.320 ; 
                RECT 2.880 436.360 221.120 436.680 ; 
                RECT 435.680 436.360 440.400 436.680 ; 
                RECT 2.880 437.720 440.400 438.040 ; 
                RECT 2.880 439.080 440.400 439.400 ; 
                RECT 2.880 440.440 440.400 440.760 ; 
                RECT 2.880 441.800 440.400 442.120 ; 
                RECT 2.880 443.160 440.400 443.480 ; 
                RECT 2.880 2.880 440.400 4.240 ; 
                RECT 2.880 444.480 440.400 445.840 ; 
                RECT 225.260 29.725 231.060 30.845 ; 
                RECT 425.960 29.725 431.760 30.845 ; 
                RECT 225.260 35.515 231.060 36.135 ; 
                RECT 425.960 35.515 431.760 36.135 ; 
                RECT 225.260 40.540 231.060 41.180 ; 
                RECT 425.960 40.540 431.760 41.180 ; 
                RECT 225.260 45.670 231.060 46.320 ; 
                RECT 425.960 45.670 431.760 46.320 ; 
                RECT 225.260 50.885 231.060 51.495 ; 
                RECT 425.960 50.885 431.760 51.495 ; 
                RECT 225.260 55.815 231.060 56.425 ; 
                RECT 425.960 55.815 431.760 56.425 ; 
                RECT 225.260 86.500 431.760 87.300 ; 
                RECT 225.260 142.855 431.760 144.655 ; 
                RECT 225.260 90.185 431.760 93.785 ; 
                RECT 225.260 69.550 431.760 71.350 ; 
                RECT 225.260 81.610 431.760 82.410 ; 
                RECT 225.260 115.645 431.760 115.935 ; 
                RECT 225.260 78.600 431.760 79.400 ; 
                RECT 225.260 83.290 431.760 84.090 ; 
                RECT 225.260 20.355 431.760 22.155 ; 
                RECT 100.285 179.035 101.605 433.415 ; 
                RECT 110.830 179.035 112.750 433.415 ; 
                RECT 128.570 179.035 130.490 433.415 ; 
                RECT 132.410 179.035 134.330 433.415 ; 
                RECT 161.590 179.035 163.510 433.415 ; 
                RECT 165.430 179.035 167.350 433.415 ; 
                RECT 169.270 179.035 171.190 433.415 ; 
                RECT 173.110 179.035 175.030 433.415 ; 
                RECT 149.110 61.485 150.000 114.085 ; 
                RECT 155.870 61.485 156.760 114.085 ; 
                RECT 161.770 61.485 162.660 114.085 ; 
                RECT 168.960 61.485 170.710 114.085 ; 
                RECT 181.885 61.485 183.805 114.085 ; 
                RECT 185.725 61.485 187.645 114.085 ; 
                RECT 161.665 139.540 162.775 172.400 ; 
                RECT 169.180 139.540 170.070 172.400 ; 
                RECT 175.940 139.540 176.830 172.400 ; 
                RECT 182.375 139.540 183.485 172.400 ; 
                RECT 191.525 139.540 193.445 172.400 ; 
                RECT 169.165 126.800 170.275 133.540 ; 
                RECT 177.645 126.800 178.755 133.540 ; 
                RECT 187.870 126.800 189.790 133.540 ; 
                RECT 200.765 51.905 201.875 55.485 ; 
                RECT 26.170 180.100 35.330 180.470 ; 
                RECT 26.170 183.435 35.330 184.325 ; 
                RECT 73.280 165.510 90.520 166.180 ; 
                RECT 73.280 166.840 90.520 168.190 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 443.280 448.720 ; 
        LAYER met2 ;
            RECT 0.000 0.000 443.280 448.720 ; 
    END 
END sram22_512x32m4w8 
END LIBRARY 

