VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_512x64m4w8
    CLASS BLOCK  ;
    FOREIGN sram22_512x64m4w8   ;
    SIZE 805.720 BY 450.080 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 402.310 0.000 402.450 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 408.410 0.000 408.550 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 414.510 0.000 414.650 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 420.610 0.000 420.750 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 426.710 0.000 426.850 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 432.810 0.000 432.950 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 438.910 0.000 439.050 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 445.010 0.000 445.150 0.140 ; 
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 451.110 0.000 451.250 0.140 ; 
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 457.210 0.000 457.350 0.140 ; 
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 463.310 0.000 463.450 0.140 ; 
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 469.410 0.000 469.550 0.140 ; 
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 475.510 0.000 475.650 0.140 ; 
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 481.610 0.000 481.750 0.140 ; 
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 487.710 0.000 487.850 0.140 ; 
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 493.810 0.000 493.950 0.140 ; 
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 499.910 0.000 500.050 0.140 ; 
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 506.010 0.000 506.150 0.140 ; 
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 512.110 0.000 512.250 0.140 ; 
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 518.210 0.000 518.350 0.140 ; 
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 524.310 0.000 524.450 0.140 ; 
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 530.410 0.000 530.550 0.140 ; 
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 536.510 0.000 536.650 0.140 ; 
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 542.610 0.000 542.750 0.140 ; 
        END 
    END dout[23] 
    PIN dout[24] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 548.710 0.000 548.850 0.140 ; 
        END 
    END dout[24] 
    PIN dout[25] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 554.810 0.000 554.950 0.140 ; 
        END 
    END dout[25] 
    PIN dout[26] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 560.910 0.000 561.050 0.140 ; 
        END 
    END dout[26] 
    PIN dout[27] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 567.010 0.000 567.150 0.140 ; 
        END 
    END dout[27] 
    PIN dout[28] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 573.110 0.000 573.250 0.140 ; 
        END 
    END dout[28] 
    PIN dout[29] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 579.210 0.000 579.350 0.140 ; 
        END 
    END dout[29] 
    PIN dout[30] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 585.310 0.000 585.450 0.140 ; 
        END 
    END dout[30] 
    PIN dout[31] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 591.410 0.000 591.550 0.140 ; 
        END 
    END dout[31] 
    PIN dout[32] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 597.510 0.000 597.650 0.140 ; 
        END 
    END dout[32] 
    PIN dout[33] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 603.610 0.000 603.750 0.140 ; 
        END 
    END dout[33] 
    PIN dout[34] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 609.710 0.000 609.850 0.140 ; 
        END 
    END dout[34] 
    PIN dout[35] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 615.810 0.000 615.950 0.140 ; 
        END 
    END dout[35] 
    PIN dout[36] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 621.910 0.000 622.050 0.140 ; 
        END 
    END dout[36] 
    PIN dout[37] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 628.010 0.000 628.150 0.140 ; 
        END 
    END dout[37] 
    PIN dout[38] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 634.110 0.000 634.250 0.140 ; 
        END 
    END dout[38] 
    PIN dout[39] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 640.210 0.000 640.350 0.140 ; 
        END 
    END dout[39] 
    PIN dout[40] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 646.310 0.000 646.450 0.140 ; 
        END 
    END dout[40] 
    PIN dout[41] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 652.410 0.000 652.550 0.140 ; 
        END 
    END dout[41] 
    PIN dout[42] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 658.510 0.000 658.650 0.140 ; 
        END 
    END dout[42] 
    PIN dout[43] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 664.610 0.000 664.750 0.140 ; 
        END 
    END dout[43] 
    PIN dout[44] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 670.710 0.000 670.850 0.140 ; 
        END 
    END dout[44] 
    PIN dout[45] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 676.810 0.000 676.950 0.140 ; 
        END 
    END dout[45] 
    PIN dout[46] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 682.910 0.000 683.050 0.140 ; 
        END 
    END dout[46] 
    PIN dout[47] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 689.010 0.000 689.150 0.140 ; 
        END 
    END dout[47] 
    PIN dout[48] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 695.110 0.000 695.250 0.140 ; 
        END 
    END dout[48] 
    PIN dout[49] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 701.210 0.000 701.350 0.140 ; 
        END 
    END dout[49] 
    PIN dout[50] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 707.310 0.000 707.450 0.140 ; 
        END 
    END dout[50] 
    PIN dout[51] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 713.410 0.000 713.550 0.140 ; 
        END 
    END dout[51] 
    PIN dout[52] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 719.510 0.000 719.650 0.140 ; 
        END 
    END dout[52] 
    PIN dout[53] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 725.610 0.000 725.750 0.140 ; 
        END 
    END dout[53] 
    PIN dout[54] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 731.710 0.000 731.850 0.140 ; 
        END 
    END dout[54] 
    PIN dout[55] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 737.810 0.000 737.950 0.140 ; 
        END 
    END dout[55] 
    PIN dout[56] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 743.910 0.000 744.050 0.140 ; 
        END 
    END dout[56] 
    PIN dout[57] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 750.010 0.000 750.150 0.140 ; 
        END 
    END dout[57] 
    PIN dout[58] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 756.110 0.000 756.250 0.140 ; 
        END 
    END dout[58] 
    PIN dout[59] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 762.210 0.000 762.350 0.140 ; 
        END 
    END dout[59] 
    PIN dout[60] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 768.310 0.000 768.450 0.140 ; 
        END 
    END dout[60] 
    PIN dout[61] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 774.410 0.000 774.550 0.140 ; 
        END 
    END dout[61] 
    PIN dout[62] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 780.510 0.000 780.650 0.140 ; 
        END 
    END dout[62] 
    PIN dout[63] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.891800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 786.610 0.000 786.750 0.140 ; 
        END 
    END dout[63] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 401.890 0.000 402.030 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 407.990 0.000 408.130 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 414.090 0.000 414.230 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 420.190 0.000 420.330 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 426.290 0.000 426.430 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 432.390 0.000 432.530 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 438.490 0.000 438.630 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 444.590 0.000 444.730 0.140 ; 
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 450.690 0.000 450.830 0.140 ; 
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 456.790 0.000 456.930 0.140 ; 
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 462.890 0.000 463.030 0.140 ; 
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 468.990 0.000 469.130 0.140 ; 
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 475.090 0.000 475.230 0.140 ; 
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 481.190 0.000 481.330 0.140 ; 
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 487.290 0.000 487.430 0.140 ; 
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 493.390 0.000 493.530 0.140 ; 
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 499.490 0.000 499.630 0.140 ; 
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 505.590 0.000 505.730 0.140 ; 
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 511.690 0.000 511.830 0.140 ; 
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 517.790 0.000 517.930 0.140 ; 
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 523.890 0.000 524.030 0.140 ; 
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 529.990 0.000 530.130 0.140 ; 
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 536.090 0.000 536.230 0.140 ; 
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 542.190 0.000 542.330 0.140 ; 
        END 
    END din[23] 
    PIN din[24] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 548.290 0.000 548.430 0.140 ; 
        END 
    END din[24] 
    PIN din[25] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 554.390 0.000 554.530 0.140 ; 
        END 
    END din[25] 
    PIN din[26] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 560.490 0.000 560.630 0.140 ; 
        END 
    END din[26] 
    PIN din[27] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 566.590 0.000 566.730 0.140 ; 
        END 
    END din[27] 
    PIN din[28] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 572.690 0.000 572.830 0.140 ; 
        END 
    END din[28] 
    PIN din[29] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 578.790 0.000 578.930 0.140 ; 
        END 
    END din[29] 
    PIN din[30] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 584.890 0.000 585.030 0.140 ; 
        END 
    END din[30] 
    PIN din[31] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 590.990 0.000 591.130 0.140 ; 
        END 
    END din[31] 
    PIN din[32] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 597.090 0.000 597.230 0.140 ; 
        END 
    END din[32] 
    PIN din[33] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 603.190 0.000 603.330 0.140 ; 
        END 
    END din[33] 
    PIN din[34] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 609.290 0.000 609.430 0.140 ; 
        END 
    END din[34] 
    PIN din[35] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 615.390 0.000 615.530 0.140 ; 
        END 
    END din[35] 
    PIN din[36] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 621.490 0.000 621.630 0.140 ; 
        END 
    END din[36] 
    PIN din[37] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 627.590 0.000 627.730 0.140 ; 
        END 
    END din[37] 
    PIN din[38] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 633.690 0.000 633.830 0.140 ; 
        END 
    END din[38] 
    PIN din[39] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 639.790 0.000 639.930 0.140 ; 
        END 
    END din[39] 
    PIN din[40] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 645.890 0.000 646.030 0.140 ; 
        END 
    END din[40] 
    PIN din[41] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 651.990 0.000 652.130 0.140 ; 
        END 
    END din[41] 
    PIN din[42] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 658.090 0.000 658.230 0.140 ; 
        END 
    END din[42] 
    PIN din[43] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 664.190 0.000 664.330 0.140 ; 
        END 
    END din[43] 
    PIN din[44] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 670.290 0.000 670.430 0.140 ; 
        END 
    END din[44] 
    PIN din[45] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 676.390 0.000 676.530 0.140 ; 
        END 
    END din[45] 
    PIN din[46] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 682.490 0.000 682.630 0.140 ; 
        END 
    END din[46] 
    PIN din[47] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 688.590 0.000 688.730 0.140 ; 
        END 
    END din[47] 
    PIN din[48] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 694.690 0.000 694.830 0.140 ; 
        END 
    END din[48] 
    PIN din[49] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 700.790 0.000 700.930 0.140 ; 
        END 
    END din[49] 
    PIN din[50] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 706.890 0.000 707.030 0.140 ; 
        END 
    END din[50] 
    PIN din[51] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 712.990 0.000 713.130 0.140 ; 
        END 
    END din[51] 
    PIN din[52] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 719.090 0.000 719.230 0.140 ; 
        END 
    END din[52] 
    PIN din[53] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 725.190 0.000 725.330 0.140 ; 
        END 
    END din[53] 
    PIN din[54] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 731.290 0.000 731.430 0.140 ; 
        END 
    END din[54] 
    PIN din[55] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 737.390 0.000 737.530 0.140 ; 
        END 
    END din[55] 
    PIN din[56] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 743.490 0.000 743.630 0.140 ; 
        END 
    END din[56] 
    PIN din[57] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 749.590 0.000 749.730 0.140 ; 
        END 
    END din[57] 
    PIN din[58] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 755.690 0.000 755.830 0.140 ; 
        END 
    END din[58] 
    PIN din[59] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 761.790 0.000 761.930 0.140 ; 
        END 
    END din[59] 
    PIN din[60] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 767.890 0.000 768.030 0.140 ; 
        END 
    END din[60] 
    PIN din[61] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 773.990 0.000 774.130 0.140 ; 
        END 
    END din[61] 
    PIN din[62] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 780.090 0.000 780.230 0.140 ; 
        END 
    END din[62] 
    PIN din[63] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.830800 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 9.613400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 786.190 0.000 786.330 0.140 ; 
        END 
    END din[63] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.641200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 401.540 0.000 401.680 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.641200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 450.340 0.000 450.480 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.641200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 499.140 0.000 499.280 0.140 ; 
        END 
    END wmask[2] 
    PIN wmask[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.641200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 547.940 0.000 548.080 0.140 ; 
        END 
    END wmask[3] 
    PIN wmask[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.641200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 596.740 0.000 596.880 0.140 ; 
        END 
    END wmask[4] 
    PIN wmask[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.641200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 645.540 0.000 645.680 0.140 ; 
        END 
    END wmask[5] 
    PIN wmask[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.641200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 694.340 0.000 694.480 0.140 ; 
        END 
    END wmask[6] 
    PIN wmask[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 1.641200 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 743.140 0.000 743.280 0.140 ; 
        END 
    END wmask[7] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 359.520 0.000 359.840 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 353.400 0.000 353.720 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 347.280 0.000 347.600 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 341.160 0.000 341.480 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 335.040 0.000 335.360 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 328.920 0.000 329.240 0.320 ; 
        END 
    END addr[5] 
    PIN addr[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 322.800 0.000 323.120 0.320 ; 
        END 
    END addr[6] 
    PIN addr[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 316.680 0.000 317.000 0.320 ; 
        END 
    END addr[7] 
    PIN addr[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 310.560 0.000 310.880 0.320 ; 
        END 
    END addr[8] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 371.760 0.000 372.080 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.063100 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 365.640 0.000 365.960 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 41.571000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 374.480 0.000 374.800 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 45.477000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 375.160 0.000 375.480 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 401.320 6.240 ; 
                RECT 787.240 5.920 805.560 6.240 ; 
                RECT 0.160 7.280 805.560 7.600 ; 
                RECT 0.160 8.640 805.560 8.960 ; 
                RECT 0.160 10.000 374.120 10.320 ; 
                RECT 796.080 10.000 805.560 10.320 ; 
                RECT 0.160 11.360 391.120 11.680 ; 
                RECT 796.080 11.360 805.560 11.680 ; 
                RECT 0.160 12.720 391.120 13.040 ; 
                RECT 796.080 12.720 805.560 13.040 ; 
                RECT 0.160 14.080 391.120 14.400 ; 
                RECT 796.080 14.080 805.560 14.400 ; 
                RECT 0.160 15.440 391.120 15.760 ; 
                RECT 796.080 15.440 805.560 15.760 ; 
                RECT 0.160 16.800 391.120 17.120 ; 
                RECT 796.080 16.800 805.560 17.120 ; 
                RECT 0.160 18.160 391.120 18.480 ; 
                RECT 796.080 18.160 805.560 18.480 ; 
                RECT 0.160 19.520 391.120 19.840 ; 
                RECT 796.080 19.520 805.560 19.840 ; 
                RECT 0.160 20.880 306.800 21.200 ; 
                RECT 375.840 20.880 391.120 21.200 ; 
                RECT 796.080 20.880 805.560 21.200 ; 
                RECT 0.160 22.240 391.120 22.560 ; 
                RECT 796.080 22.240 805.560 22.560 ; 
                RECT 0.160 23.600 391.120 23.920 ; 
                RECT 796.080 23.600 805.560 23.920 ; 
                RECT 0.160 24.960 306.800 25.280 ; 
                RECT 375.160 24.960 391.120 25.280 ; 
                RECT 796.080 24.960 805.560 25.280 ; 
                RECT 0.160 26.320 391.120 26.640 ; 
                RECT 796.080 26.320 805.560 26.640 ; 
                RECT 0.160 27.680 390.440 28.000 ; 
                RECT 796.080 27.680 805.560 28.000 ; 
                RECT 0.160 29.040 391.120 29.360 ; 
                RECT 796.080 29.040 805.560 29.360 ; 
                RECT 0.160 30.400 391.120 30.720 ; 
                RECT 796.080 30.400 805.560 30.720 ; 
                RECT 0.160 31.760 391.120 32.080 ; 
                RECT 796.080 31.760 805.560 32.080 ; 
                RECT 0.160 33.120 391.120 33.440 ; 
                RECT 796.080 33.120 805.560 33.440 ; 
                RECT 0.160 34.480 391.120 34.800 ; 
                RECT 796.080 34.480 805.560 34.800 ; 
                RECT 0.160 35.840 391.120 36.160 ; 
                RECT 796.080 35.840 805.560 36.160 ; 
                RECT 0.160 37.200 391.120 37.520 ; 
                RECT 796.080 37.200 805.560 37.520 ; 
                RECT 0.160 38.560 391.120 38.880 ; 
                RECT 796.080 38.560 805.560 38.880 ; 
                RECT 0.160 39.920 391.120 40.240 ; 
                RECT 796.080 39.920 805.560 40.240 ; 
                RECT 0.160 41.280 391.120 41.600 ; 
                RECT 796.080 41.280 805.560 41.600 ; 
                RECT 0.160 42.640 276.880 42.960 ; 
                RECT 352.720 42.640 391.120 42.960 ; 
                RECT 796.080 42.640 805.560 42.960 ; 
                RECT 0.160 44.000 275.520 44.320 ; 
                RECT 358.840 44.000 391.120 44.320 ; 
                RECT 796.080 44.000 805.560 44.320 ; 
                RECT 0.160 45.360 255.800 45.680 ; 
                RECT 375.840 45.360 391.120 45.680 ; 
                RECT 796.080 45.360 805.560 45.680 ; 
                RECT 0.160 46.720 255.120 47.040 ; 
                RECT 371.760 46.720 391.120 47.040 ; 
                RECT 796.080 46.720 805.560 47.040 ; 
                RECT 0.160 48.080 391.120 48.400 ; 
                RECT 796.080 48.080 805.560 48.400 ; 
                RECT 0.160 49.440 391.120 49.760 ; 
                RECT 796.080 49.440 805.560 49.760 ; 
                RECT 0.160 50.800 368.000 51.120 ; 
                RECT 373.800 50.800 391.120 51.120 ; 
                RECT 796.080 50.800 805.560 51.120 ; 
                RECT 0.160 52.160 368.000 52.480 ; 
                RECT 796.080 52.160 805.560 52.480 ; 
                RECT 0.160 53.520 368.000 53.840 ; 
                RECT 796.080 53.520 805.560 53.840 ; 
                RECT 0.160 54.880 274.160 55.200 ; 
                RECT 365.640 54.880 368.000 55.200 ; 
                RECT 373.800 54.880 391.120 55.200 ; 
                RECT 796.080 54.880 805.560 55.200 ; 
                RECT 0.160 56.240 391.120 56.560 ; 
                RECT 796.080 56.240 805.560 56.560 ; 
                RECT 0.160 57.600 391.120 57.920 ; 
                RECT 796.080 57.600 805.560 57.920 ; 
                RECT 0.160 58.960 391.120 59.280 ; 
                RECT 796.080 58.960 805.560 59.280 ; 
                RECT 0.160 60.320 391.120 60.640 ; 
                RECT 796.080 60.320 805.560 60.640 ; 
                RECT 0.160 61.680 275.520 62.000 ; 
                RECT 281.320 61.680 286.400 62.000 ; 
                RECT 373.120 61.680 391.120 62.000 ; 
                RECT 796.080 61.680 805.560 62.000 ; 
                RECT 0.160 63.040 276.880 63.360 ; 
                RECT 279.960 63.040 286.400 63.360 ; 
                RECT 383.320 63.040 391.120 63.360 ; 
                RECT 796.080 63.040 805.560 63.360 ; 
                RECT 0.160 64.400 286.400 64.720 ; 
                RECT 373.120 64.400 391.120 64.720 ; 
                RECT 796.080 64.400 805.560 64.720 ; 
                RECT 0.160 65.760 286.400 66.080 ; 
                RECT 381.960 65.760 391.120 66.080 ; 
                RECT 796.080 65.760 805.560 66.080 ; 
                RECT 0.160 67.120 286.400 67.440 ; 
                RECT 383.320 67.120 391.120 67.440 ; 
                RECT 796.080 67.120 805.560 67.440 ; 
                RECT 0.160 68.480 286.400 68.800 ; 
                RECT 383.320 68.480 391.120 68.800 ; 
                RECT 796.080 68.480 805.560 68.800 ; 
                RECT 0.160 69.840 286.400 70.160 ; 
                RECT 381.960 69.840 391.120 70.160 ; 
                RECT 796.080 69.840 805.560 70.160 ; 
                RECT 0.160 71.200 251.040 71.520 ; 
                RECT 262.280 71.200 286.400 71.520 ; 
                RECT 383.320 71.200 391.120 71.520 ; 
                RECT 796.080 71.200 805.560 71.520 ; 
                RECT 0.160 72.560 252.400 72.880 ; 
                RECT 258.200 72.560 266.000 72.880 ; 
                RECT 268.400 72.560 286.400 72.880 ; 
                RECT 381.960 72.560 391.120 72.880 ; 
                RECT 796.080 72.560 805.560 72.880 ; 
                RECT 0.160 73.920 253.760 74.240 ; 
                RECT 257.520 73.920 286.400 74.240 ; 
                RECT 383.320 73.920 391.120 74.240 ; 
                RECT 796.080 73.920 805.560 74.240 ; 
                RECT 0.160 75.280 260.560 75.600 ; 
                RECT 267.720 75.280 286.400 75.600 ; 
                RECT 386.040 75.280 391.120 75.600 ; 
                RECT 796.080 75.280 805.560 75.600 ; 
                RECT 0.160 76.640 255.800 76.960 ; 
                RECT 269.080 76.640 286.400 76.960 ; 
                RECT 384.680 76.640 391.120 76.960 ; 
                RECT 796.080 76.640 805.560 76.960 ; 
                RECT 0.160 78.000 253.080 78.320 ; 
                RECT 262.280 78.000 286.400 78.320 ; 
                RECT 386.040 78.000 391.120 78.320 ; 
                RECT 796.080 78.000 805.560 78.320 ; 
                RECT 0.160 79.360 286.400 79.680 ; 
                RECT 373.120 79.360 391.120 79.680 ; 
                RECT 796.080 79.360 805.560 79.680 ; 
                RECT 0.160 80.720 252.400 81.040 ; 
                RECT 255.480 80.720 286.400 81.040 ; 
                RECT 386.040 80.720 391.120 81.040 ; 
                RECT 796.080 80.720 805.560 81.040 ; 
                RECT 0.160 82.080 250.360 82.400 ; 
                RECT 268.400 82.080 286.400 82.400 ; 
                RECT 386.040 82.080 391.120 82.400 ; 
                RECT 796.080 82.080 805.560 82.400 ; 
                RECT 0.160 83.440 259.200 83.760 ; 
                RECT 262.280 83.440 286.400 83.760 ; 
                RECT 373.120 83.440 391.120 83.760 ; 
                RECT 796.080 83.440 805.560 83.760 ; 
                RECT 0.160 84.800 286.400 85.120 ; 
                RECT 384.680 84.800 391.120 85.120 ; 
                RECT 796.080 84.800 805.560 85.120 ; 
                RECT 0.160 86.160 260.560 86.480 ; 
                RECT 268.400 86.160 286.400 86.480 ; 
                RECT 386.040 86.160 391.120 86.480 ; 
                RECT 796.080 86.160 805.560 86.480 ; 
                RECT 0.160 87.520 257.160 87.840 ; 
                RECT 262.280 87.520 286.400 87.840 ; 
                RECT 373.120 87.520 391.120 87.840 ; 
                RECT 796.080 87.520 805.560 87.840 ; 
                RECT 0.160 88.880 259.200 89.200 ; 
                RECT 262.280 88.880 286.400 89.200 ; 
                RECT 388.760 88.880 391.120 89.200 ; 
                RECT 796.080 88.880 805.560 89.200 ; 
                RECT 0.160 90.240 286.400 90.560 ; 
                RECT 388.760 90.240 391.120 90.560 ; 
                RECT 796.080 90.240 805.560 90.560 ; 
                RECT 0.160 91.600 251.040 91.920 ; 
                RECT 273.840 91.600 286.400 91.920 ; 
                RECT 387.400 91.600 391.120 91.920 ; 
                RECT 796.080 91.600 805.560 91.920 ; 
                RECT 0.160 92.960 269.400 93.280 ; 
                RECT 275.200 92.960 286.400 93.280 ; 
                RECT 388.760 92.960 391.120 93.280 ; 
                RECT 796.080 92.960 805.560 93.280 ; 
                RECT 0.160 94.320 259.200 94.640 ; 
                RECT 262.280 94.320 272.120 94.640 ; 
                RECT 275.880 94.320 286.400 94.640 ; 
                RECT 388.760 94.320 391.120 94.640 ; 
                RECT 796.080 94.320 805.560 94.640 ; 
                RECT 0.160 95.680 251.040 96.000 ; 
                RECT 265.000 95.680 286.400 96.000 ; 
                RECT 387.400 95.680 391.120 96.000 ; 
                RECT 796.080 95.680 805.560 96.000 ; 
                RECT 0.160 97.040 259.880 97.360 ; 
                RECT 268.400 97.040 286.400 97.360 ; 
                RECT 388.760 97.040 391.120 97.360 ; 
                RECT 796.080 97.040 805.560 97.360 ; 
                RECT 0.160 98.400 257.840 98.720 ; 
                RECT 261.600 98.400 286.400 98.720 ; 
                RECT 387.400 98.400 391.120 98.720 ; 
                RECT 796.080 98.400 805.560 98.720 ; 
                RECT 0.160 99.760 260.560 100.080 ; 
                RECT 269.080 99.760 286.400 100.080 ; 
                RECT 388.760 99.760 391.120 100.080 ; 
                RECT 796.080 99.760 805.560 100.080 ; 
                RECT 0.160 101.120 286.400 101.440 ; 
                RECT 796.080 101.120 805.560 101.440 ; 
                RECT 0.160 102.480 253.760 102.800 ; 
                RECT 256.160 102.480 286.400 102.800 ; 
                RECT 796.080 102.480 805.560 102.800 ; 
                RECT 0.160 103.840 253.080 104.160 ; 
                RECT 262.280 103.840 286.400 104.160 ; 
                RECT 796.080 103.840 805.560 104.160 ; 
                RECT 0.160 105.200 286.400 105.520 ; 
                RECT 373.120 105.200 391.120 105.520 ; 
                RECT 796.080 105.200 805.560 105.520 ; 
                RECT 0.160 106.560 259.200 106.880 ; 
                RECT 261.600 106.560 286.400 106.880 ; 
                RECT 796.080 106.560 805.560 106.880 ; 
                RECT 0.160 107.920 252.400 108.240 ; 
                RECT 258.200 107.920 260.560 108.240 ; 
                RECT 262.280 107.920 286.400 108.240 ; 
                RECT 796.080 107.920 805.560 108.240 ; 
                RECT 0.160 109.280 256.480 109.600 ; 
                RECT 267.720 109.280 286.400 109.600 ; 
                RECT 373.120 109.280 391.120 109.600 ; 
                RECT 796.080 109.280 805.560 109.600 ; 
                RECT 0.160 110.640 259.200 110.960 ; 
                RECT 261.600 110.640 286.400 110.960 ; 
                RECT 796.080 110.640 805.560 110.960 ; 
                RECT 0.160 112.000 254.440 112.320 ; 
                RECT 262.280 112.000 286.400 112.320 ; 
                RECT 796.080 112.000 805.560 112.320 ; 
                RECT 0.160 113.360 259.880 113.680 ; 
                RECT 262.280 113.360 286.400 113.680 ; 
                RECT 373.120 113.360 391.120 113.680 ; 
                RECT 796.080 113.360 805.560 113.680 ; 
                RECT 0.160 114.720 251.040 115.040 ; 
                RECT 258.200 114.720 391.120 115.040 ; 
                RECT 796.080 114.720 805.560 115.040 ; 
                RECT 0.160 116.080 250.360 116.400 ; 
                RECT 268.400 116.080 391.120 116.400 ; 
                RECT 796.080 116.080 805.560 116.400 ; 
                RECT 0.160 117.440 247.640 117.760 ; 
                RECT 260.920 117.440 377.520 117.760 ; 
                RECT 796.080 117.440 805.560 117.760 ; 
                RECT 0.160 118.800 251.040 119.120 ; 
                RECT 265.000 118.800 388.400 119.120 ; 
                RECT 796.080 118.800 805.560 119.120 ; 
                RECT 0.160 120.160 266.680 120.480 ; 
                RECT 268.400 120.160 385.680 120.480 ; 
                RECT 796.080 120.160 805.560 120.480 ; 
                RECT 0.160 121.520 380.240 121.840 ; 
                RECT 796.080 121.520 805.560 121.840 ; 
                RECT 0.160 122.880 229.280 123.200 ; 
                RECT 248.000 122.880 263.280 123.200 ; 
                RECT 271.120 122.880 380.240 123.200 ; 
                RECT 796.080 122.880 805.560 123.200 ; 
                RECT 0.160 124.240 229.280 124.560 ; 
                RECT 248.000 124.240 391.120 124.560 ; 
                RECT 796.080 124.240 805.560 124.560 ; 
                RECT 0.160 125.600 229.280 125.920 ; 
                RECT 248.000 125.600 391.120 125.920 ; 
                RECT 796.080 125.600 805.560 125.920 ; 
                RECT 0.160 126.960 229.280 127.280 ; 
                RECT 248.000 126.960 253.080 127.280 ; 
                RECT 256.160 126.960 391.120 127.280 ; 
                RECT 796.080 126.960 805.560 127.280 ; 
                RECT 0.160 128.320 229.280 128.640 ; 
                RECT 248.000 128.320 251.040 128.640 ; 
                RECT 254.800 128.320 274.840 128.640 ; 
                RECT 317.360 128.320 320.400 128.640 ; 
                RECT 373.120 128.320 391.120 128.640 ; 
                RECT 796.080 128.320 805.560 128.640 ; 
                RECT 0.160 129.680 229.280 130.000 ; 
                RECT 248.000 129.680 320.400 130.000 ; 
                RECT 373.120 129.680 391.120 130.000 ; 
                RECT 796.080 129.680 805.560 130.000 ; 
                RECT 0.160 131.040 229.280 131.360 ; 
                RECT 248.000 131.040 320.400 131.360 ; 
                RECT 373.120 131.040 391.120 131.360 ; 
                RECT 796.080 131.040 805.560 131.360 ; 
                RECT 0.160 132.400 229.280 132.720 ; 
                RECT 248.000 132.400 256.480 132.720 ; 
                RECT 268.400 132.400 320.400 132.720 ; 
                RECT 373.120 132.400 391.120 132.720 ; 
                RECT 796.080 132.400 805.560 132.720 ; 
                RECT 0.160 133.760 229.280 134.080 ; 
                RECT 248.000 133.760 320.400 134.080 ; 
                RECT 373.120 133.760 391.120 134.080 ; 
                RECT 796.080 133.760 805.560 134.080 ; 
                RECT 0.160 135.120 229.280 135.440 ; 
                RECT 248.000 135.120 320.400 135.440 ; 
                RECT 373.120 135.120 391.120 135.440 ; 
                RECT 796.080 135.120 805.560 135.440 ; 
                RECT 0.160 136.480 229.280 136.800 ; 
                RECT 248.000 136.480 391.120 136.800 ; 
                RECT 796.080 136.480 805.560 136.800 ; 
                RECT 0.160 137.840 229.280 138.160 ; 
                RECT 248.000 137.840 253.080 138.160 ; 
                RECT 258.200 137.840 391.120 138.160 ; 
                RECT 796.080 137.840 805.560 138.160 ; 
                RECT 0.160 139.200 229.280 139.520 ; 
                RECT 248.000 139.200 391.120 139.520 ; 
                RECT 796.080 139.200 805.560 139.520 ; 
                RECT 0.160 140.560 229.280 140.880 ; 
                RECT 248.000 140.560 266.680 140.880 ; 
                RECT 269.080 140.560 310.880 140.880 ; 
                RECT 373.120 140.560 391.120 140.880 ; 
                RECT 796.080 140.560 805.560 140.880 ; 
                RECT 0.160 141.920 229.280 142.240 ; 
                RECT 248.680 141.920 310.880 142.240 ; 
                RECT 373.120 141.920 391.120 142.240 ; 
                RECT 796.080 141.920 805.560 142.240 ; 
                RECT 0.160 143.280 229.280 143.600 ; 
                RECT 248.000 143.280 310.880 143.600 ; 
                RECT 373.120 143.280 391.120 143.600 ; 
                RECT 796.080 143.280 805.560 143.600 ; 
                RECT 0.160 144.640 229.280 144.960 ; 
                RECT 248.000 144.640 252.400 144.960 ; 
                RECT 255.480 144.640 310.880 144.960 ; 
                RECT 373.120 144.640 391.120 144.960 ; 
                RECT 796.080 144.640 805.560 144.960 ; 
                RECT 0.160 146.000 229.280 146.320 ; 
                RECT 248.000 146.000 310.880 146.320 ; 
                RECT 373.120 146.000 391.120 146.320 ; 
                RECT 796.080 146.000 805.560 146.320 ; 
                RECT 0.160 147.360 229.280 147.680 ; 
                RECT 248.000 147.360 310.880 147.680 ; 
                RECT 373.120 147.360 391.120 147.680 ; 
                RECT 796.080 147.360 805.560 147.680 ; 
                RECT 0.160 148.720 229.280 149.040 ; 
                RECT 248.000 148.720 259.200 149.040 ; 
                RECT 268.400 148.720 310.880 149.040 ; 
                RECT 373.120 148.720 381.600 149.040 ; 
                RECT 796.080 148.720 805.560 149.040 ; 
                RECT 0.160 150.080 229.280 150.400 ; 
                RECT 248.000 150.080 310.880 150.400 ; 
                RECT 373.120 150.080 381.600 150.400 ; 
                RECT 796.080 150.080 805.560 150.400 ; 
                RECT 0.160 151.440 229.280 151.760 ; 
                RECT 248.000 151.440 255.800 151.760 ; 
                RECT 258.200 151.440 310.880 151.760 ; 
                RECT 373.120 151.440 384.320 151.760 ; 
                RECT 796.080 151.440 805.560 151.760 ; 
                RECT 0.160 152.800 229.280 153.120 ; 
                RECT 248.000 152.800 310.880 153.120 ; 
                RECT 373.120 152.800 387.040 153.120 ; 
                RECT 796.080 152.800 805.560 153.120 ; 
                RECT 0.160 154.160 229.280 154.480 ; 
                RECT 248.000 154.160 310.880 154.480 ; 
                RECT 796.080 154.160 805.560 154.480 ; 
                RECT 0.160 155.520 229.280 155.840 ; 
                RECT 248.000 155.520 310.880 155.840 ; 
                RECT 796.080 155.520 805.560 155.840 ; 
                RECT 0.160 156.880 229.280 157.200 ; 
                RECT 248.000 156.880 310.880 157.200 ; 
                RECT 373.120 156.880 391.120 157.200 ; 
                RECT 796.080 156.880 805.560 157.200 ; 
                RECT 0.160 158.240 229.280 158.560 ; 
                RECT 248.000 158.240 310.880 158.560 ; 
                RECT 373.120 158.240 391.120 158.560 ; 
                RECT 796.080 158.240 805.560 158.560 ; 
                RECT 0.160 159.600 229.280 159.920 ; 
                RECT 248.000 159.600 310.880 159.920 ; 
                RECT 373.120 159.600 391.120 159.920 ; 
                RECT 796.080 159.600 805.560 159.920 ; 
                RECT 0.160 160.960 229.280 161.280 ; 
                RECT 248.000 160.960 310.880 161.280 ; 
                RECT 373.120 160.960 391.120 161.280 ; 
                RECT 796.080 160.960 805.560 161.280 ; 
                RECT 0.160 162.320 229.280 162.640 ; 
                RECT 248.000 162.320 310.880 162.640 ; 
                RECT 373.120 162.320 391.120 162.640 ; 
                RECT 796.080 162.320 805.560 162.640 ; 
                RECT 0.160 163.680 254.440 164.000 ; 
                RECT 258.200 163.680 310.880 164.000 ; 
                RECT 373.120 163.680 391.120 164.000 ; 
                RECT 796.080 163.680 805.560 164.000 ; 
                RECT 0.160 165.040 310.880 165.360 ; 
                RECT 373.120 165.040 391.120 165.360 ; 
                RECT 796.080 165.040 805.560 165.360 ; 
                RECT 0.160 166.400 210.920 166.720 ; 
                RECT 229.640 166.400 310.880 166.720 ; 
                RECT 373.120 166.400 391.120 166.720 ; 
                RECT 796.080 166.400 805.560 166.720 ; 
                RECT 0.160 167.760 210.920 168.080 ; 
                RECT 229.640 167.760 256.480 168.080 ; 
                RECT 262.280 167.760 310.880 168.080 ; 
                RECT 373.120 167.760 391.120 168.080 ; 
                RECT 796.080 167.760 805.560 168.080 ; 
                RECT 0.160 169.120 210.920 169.440 ; 
                RECT 229.640 169.120 235.400 169.440 ; 
                RECT 242.560 169.120 310.880 169.440 ; 
                RECT 373.120 169.120 391.120 169.440 ; 
                RECT 796.080 169.120 805.560 169.440 ; 
                RECT 0.160 170.480 210.920 170.800 ; 
                RECT 247.320 170.480 310.880 170.800 ; 
                RECT 796.080 170.480 805.560 170.800 ; 
                RECT 0.160 171.840 210.920 172.160 ; 
                RECT 229.640 171.840 310.880 172.160 ; 
                RECT 796.080 171.840 805.560 172.160 ; 
                RECT 0.160 173.200 208.200 173.520 ; 
                RECT 242.560 173.200 251.040 173.520 ; 
                RECT 260.920 173.200 310.880 173.520 ; 
                RECT 373.120 173.200 391.120 173.520 ; 
                RECT 796.080 173.200 805.560 173.520 ; 
                RECT 0.160 174.560 235.400 174.880 ; 
                RECT 255.480 174.560 805.560 174.880 ; 
                RECT 0.160 175.920 32.080 176.240 ; 
                RECT 254.800 175.920 805.560 176.240 ; 
                RECT 0.160 177.280 388.400 177.600 ; 
                RECT 798.120 177.280 805.560 177.600 ; 
                RECT 0.160 178.640 388.400 178.960 ; 
                RECT 798.120 178.640 805.560 178.960 ; 
                RECT 0.160 180.000 27.320 180.320 ; 
                RECT 33.800 180.000 99.400 180.320 ; 
                RECT 798.120 180.000 805.560 180.320 ; 
                RECT 0.160 181.360 25.280 181.680 ; 
                RECT 35.840 181.360 36.840 181.680 ; 
                RECT 48.760 181.360 99.400 181.680 ; 
                RECT 798.120 181.360 805.560 181.680 ; 
                RECT 0.160 182.720 25.280 183.040 ; 
                RECT 35.840 182.720 38.200 183.040 ; 
                RECT 47.400 182.720 59.280 183.040 ; 
                RECT 61.000 182.720 75.600 183.040 ; 
                RECT 89.560 182.720 99.400 183.040 ; 
                RECT 798.120 182.720 805.560 183.040 ; 
                RECT 0.160 184.080 59.280 184.400 ; 
                RECT 61.000 184.080 75.600 184.400 ; 
                RECT 89.560 184.080 99.400 184.400 ; 
                RECT 798.120 184.080 805.560 184.400 ; 
                RECT 0.160 185.440 25.280 185.760 ; 
                RECT 35.840 185.440 59.280 185.760 ; 
                RECT 63.720 185.440 75.600 185.760 ; 
                RECT 89.560 185.440 99.400 185.760 ; 
                RECT 798.120 185.440 805.560 185.760 ; 
                RECT 0.160 186.800 25.280 187.120 ; 
                RECT 35.840 186.800 59.280 187.120 ; 
                RECT 64.400 186.800 75.600 187.120 ; 
                RECT 89.560 186.800 99.400 187.120 ; 
                RECT 798.120 186.800 805.560 187.120 ; 
                RECT 0.160 188.160 25.280 188.480 ; 
                RECT 35.840 188.160 59.280 188.480 ; 
                RECT 65.080 188.160 75.600 188.480 ; 
                RECT 89.560 188.160 99.400 188.480 ; 
                RECT 798.120 188.160 805.560 188.480 ; 
                RECT 0.160 189.520 25.280 189.840 ; 
                RECT 35.840 189.520 99.400 189.840 ; 
                RECT 798.120 189.520 805.560 189.840 ; 
                RECT 0.160 190.880 75.600 191.200 ; 
                RECT 89.560 190.880 99.400 191.200 ; 
                RECT 798.120 190.880 805.560 191.200 ; 
                RECT 0.160 192.240 75.600 192.560 ; 
                RECT 89.560 192.240 99.400 192.560 ; 
                RECT 798.120 192.240 805.560 192.560 ; 
                RECT 0.160 193.600 18.480 193.920 ; 
                RECT 20.880 193.600 75.600 193.920 ; 
                RECT 89.560 193.600 99.400 193.920 ; 
                RECT 798.120 193.600 805.560 193.920 ; 
                RECT 0.160 194.960 17.800 195.280 ; 
                RECT 20.880 194.960 75.600 195.280 ; 
                RECT 89.560 194.960 99.400 195.280 ; 
                RECT 798.120 194.960 805.560 195.280 ; 
                RECT 0.160 196.320 38.880 196.640 ; 
                RECT 48.760 196.320 75.600 196.640 ; 
                RECT 83.440 196.320 99.400 196.640 ; 
                RECT 798.120 196.320 805.560 196.640 ; 
                RECT 0.160 197.680 17.120 198.000 ; 
                RECT 20.880 197.680 34.120 198.000 ; 
                RECT 48.080 197.680 83.760 198.000 ; 
                RECT 89.560 197.680 99.400 198.000 ; 
                RECT 798.120 197.680 805.560 198.000 ; 
                RECT 0.160 199.040 16.440 199.360 ; 
                RECT 20.880 199.040 34.120 199.360 ; 
                RECT 39.240 199.040 59.280 199.360 ; 
                RECT 61.680 199.040 75.600 199.360 ; 
                RECT 89.560 199.040 99.400 199.360 ; 
                RECT 798.120 199.040 805.560 199.360 ; 
                RECT 0.160 200.400 59.280 200.720 ; 
                RECT 62.360 200.400 75.600 200.720 ; 
                RECT 89.560 200.400 99.400 200.720 ; 
                RECT 798.120 200.400 805.560 200.720 ; 
                RECT 0.160 201.760 15.760 202.080 ; 
                RECT 20.880 201.760 34.120 202.080 ; 
                RECT 39.920 201.760 59.280 202.080 ; 
                RECT 62.360 201.760 75.600 202.080 ; 
                RECT 89.560 201.760 99.400 202.080 ; 
                RECT 798.120 201.760 805.560 202.080 ; 
                RECT 0.160 203.120 15.080 203.440 ; 
                RECT 20.880 203.120 34.120 203.440 ; 
                RECT 40.600 203.120 59.280 203.440 ; 
                RECT 61.000 203.120 75.600 203.440 ; 
                RECT 89.560 203.120 99.400 203.440 ; 
                RECT 798.120 203.120 805.560 203.440 ; 
                RECT 0.160 204.480 14.400 204.800 ; 
                RECT 20.880 204.480 34.120 204.800 ; 
                RECT 41.280 204.480 59.280 204.800 ; 
                RECT 63.040 204.480 75.600 204.800 ; 
                RECT 84.120 204.480 99.400 204.800 ; 
                RECT 798.120 204.480 805.560 204.800 ; 
                RECT 0.160 205.840 13.720 206.160 ; 
                RECT 20.880 205.840 75.600 206.160 ; 
                RECT 89.560 205.840 99.400 206.160 ; 
                RECT 798.120 205.840 805.560 206.160 ; 
                RECT 0.160 207.200 75.600 207.520 ; 
                RECT 89.560 207.200 99.400 207.520 ; 
                RECT 798.120 207.200 805.560 207.520 ; 
                RECT 0.160 208.560 13.040 208.880 ; 
                RECT 20.880 208.560 75.600 208.880 ; 
                RECT 89.560 208.560 99.400 208.880 ; 
                RECT 798.120 208.560 805.560 208.880 ; 
                RECT 0.160 209.920 12.360 210.240 ; 
                RECT 20.880 209.920 75.600 210.240 ; 
                RECT 89.560 209.920 99.400 210.240 ; 
                RECT 798.120 209.920 805.560 210.240 ; 
                RECT 0.160 211.280 11.680 211.600 ; 
                RECT 20.880 211.280 75.600 211.600 ; 
                RECT 89.560 211.280 99.400 211.600 ; 
                RECT 798.120 211.280 805.560 211.600 ; 
                RECT 0.160 212.640 99.400 212.960 ; 
                RECT 798.120 212.640 805.560 212.960 ; 
                RECT 0.160 214.000 11.000 214.320 ; 
                RECT 20.880 214.000 34.120 214.320 ; 
                RECT 38.560 214.000 75.600 214.320 ; 
                RECT 89.560 214.000 99.400 214.320 ; 
                RECT 798.120 214.000 805.560 214.320 ; 
                RECT 0.160 215.360 10.320 215.680 ; 
                RECT 20.880 215.360 75.600 215.680 ; 
                RECT 89.560 215.360 99.400 215.680 ; 
                RECT 798.120 215.360 805.560 215.680 ; 
                RECT 0.160 216.720 75.600 217.040 ; 
                RECT 89.560 216.720 99.400 217.040 ; 
                RECT 798.120 216.720 805.560 217.040 ; 
                RECT 0.160 218.080 9.640 218.400 ; 
                RECT 20.880 218.080 34.120 218.400 ; 
                RECT 37.200 218.080 75.600 218.400 ; 
                RECT 89.560 218.080 99.400 218.400 ; 
                RECT 798.120 218.080 805.560 218.400 ; 
                RECT 0.160 219.440 75.600 219.760 ; 
                RECT 89.560 219.440 99.400 219.760 ; 
                RECT 798.120 219.440 805.560 219.760 ; 
                RECT 0.160 220.800 99.400 221.120 ; 
                RECT 798.120 220.800 805.560 221.120 ; 
                RECT 0.160 222.160 75.600 222.480 ; 
                RECT 89.560 222.160 99.400 222.480 ; 
                RECT 798.120 222.160 805.560 222.480 ; 
                RECT 0.160 223.520 75.600 223.840 ; 
                RECT 89.560 223.520 99.400 223.840 ; 
                RECT 798.120 223.520 805.560 223.840 ; 
                RECT 0.160 224.880 75.600 225.200 ; 
                RECT 89.560 224.880 99.400 225.200 ; 
                RECT 798.120 224.880 805.560 225.200 ; 
                RECT 0.160 226.240 75.600 226.560 ; 
                RECT 89.560 226.240 99.400 226.560 ; 
                RECT 798.120 226.240 805.560 226.560 ; 
                RECT 0.160 227.600 75.600 227.920 ; 
                RECT 89.560 227.600 99.400 227.920 ; 
                RECT 798.120 227.600 805.560 227.920 ; 
                RECT 0.160 228.960 99.400 229.280 ; 
                RECT 798.120 228.960 805.560 229.280 ; 
                RECT 0.160 230.320 75.600 230.640 ; 
                RECT 89.560 230.320 99.400 230.640 ; 
                RECT 798.120 230.320 805.560 230.640 ; 
                RECT 0.160 231.680 75.600 232.000 ; 
                RECT 89.560 231.680 99.400 232.000 ; 
                RECT 798.120 231.680 805.560 232.000 ; 
                RECT 0.160 233.040 75.600 233.360 ; 
                RECT 89.560 233.040 99.400 233.360 ; 
                RECT 798.120 233.040 805.560 233.360 ; 
                RECT 0.160 234.400 75.600 234.720 ; 
                RECT 89.560 234.400 99.400 234.720 ; 
                RECT 798.120 234.400 805.560 234.720 ; 
                RECT 0.160 235.760 75.600 236.080 ; 
                RECT 88.200 235.760 99.400 236.080 ; 
                RECT 798.120 235.760 805.560 236.080 ; 
                RECT 0.160 237.120 85.800 237.440 ; 
                RECT 89.560 237.120 99.400 237.440 ; 
                RECT 798.120 237.120 805.560 237.440 ; 
                RECT 0.160 238.480 75.600 238.800 ; 
                RECT 89.560 238.480 99.400 238.800 ; 
                RECT 798.120 238.480 805.560 238.800 ; 
                RECT 0.160 239.840 75.600 240.160 ; 
                RECT 89.560 239.840 99.400 240.160 ; 
                RECT 798.120 239.840 805.560 240.160 ; 
                RECT 0.160 241.200 75.600 241.520 ; 
                RECT 89.560 241.200 99.400 241.520 ; 
                RECT 798.120 241.200 805.560 241.520 ; 
                RECT 0.160 242.560 75.600 242.880 ; 
                RECT 89.560 242.560 99.400 242.880 ; 
                RECT 798.120 242.560 805.560 242.880 ; 
                RECT 0.160 243.920 75.600 244.240 ; 
                RECT 88.880 243.920 99.400 244.240 ; 
                RECT 798.120 243.920 805.560 244.240 ; 
                RECT 0.160 245.280 80.360 245.600 ; 
                RECT 89.560 245.280 99.400 245.600 ; 
                RECT 798.120 245.280 805.560 245.600 ; 
                RECT 0.160 246.640 77.640 246.960 ; 
                RECT 89.560 246.640 99.400 246.960 ; 
                RECT 798.120 246.640 805.560 246.960 ; 
                RECT 0.160 248.000 77.640 248.320 ; 
                RECT 89.560 248.000 99.400 248.320 ; 
                RECT 798.120 248.000 805.560 248.320 ; 
                RECT 0.160 249.360 77.640 249.680 ; 
                RECT 89.560 249.360 99.400 249.680 ; 
                RECT 798.120 249.360 805.560 249.680 ; 
                RECT 0.160 250.720 77.640 251.040 ; 
                RECT 89.560 250.720 99.400 251.040 ; 
                RECT 798.120 250.720 805.560 251.040 ; 
                RECT 0.160 252.080 39.560 252.400 ; 
                RECT 65.080 252.080 99.400 252.400 ; 
                RECT 798.120 252.080 805.560 252.400 ; 
                RECT 0.160 253.440 38.200 253.760 ; 
                RECT 64.400 253.440 77.640 253.760 ; 
                RECT 89.560 253.440 99.400 253.760 ; 
                RECT 798.120 253.440 805.560 253.760 ; 
                RECT 0.160 254.800 36.840 255.120 ; 
                RECT 63.040 254.800 75.600 255.120 ; 
                RECT 89.560 254.800 99.400 255.120 ; 
                RECT 798.120 254.800 805.560 255.120 ; 
                RECT 0.160 256.160 75.600 256.480 ; 
                RECT 89.560 256.160 99.400 256.480 ; 
                RECT 798.120 256.160 805.560 256.480 ; 
                RECT 0.160 257.520 75.600 257.840 ; 
                RECT 89.560 257.520 99.400 257.840 ; 
                RECT 798.120 257.520 805.560 257.840 ; 
                RECT 0.160 258.880 75.600 259.200 ; 
                RECT 89.560 258.880 99.400 259.200 ; 
                RECT 798.120 258.880 805.560 259.200 ; 
                RECT 0.160 260.240 99.400 260.560 ; 
                RECT 798.120 260.240 805.560 260.560 ; 
                RECT 0.160 261.600 77.640 261.920 ; 
                RECT 89.560 261.600 99.400 261.920 ; 
                RECT 798.120 261.600 805.560 261.920 ; 
                RECT 0.160 262.960 75.600 263.280 ; 
                RECT 89.560 262.960 99.400 263.280 ; 
                RECT 798.120 262.960 805.560 263.280 ; 
                RECT 0.160 264.320 75.600 264.640 ; 
                RECT 89.560 264.320 99.400 264.640 ; 
                RECT 798.120 264.320 805.560 264.640 ; 
                RECT 0.160 265.680 75.600 266.000 ; 
                RECT 89.560 265.680 99.400 266.000 ; 
                RECT 798.120 265.680 805.560 266.000 ; 
                RECT 0.160 267.040 75.600 267.360 ; 
                RECT 89.560 267.040 99.400 267.360 ; 
                RECT 798.120 267.040 805.560 267.360 ; 
                RECT 0.160 268.400 99.400 268.720 ; 
                RECT 798.120 268.400 805.560 268.720 ; 
                RECT 0.160 269.760 75.600 270.080 ; 
                RECT 89.560 269.760 99.400 270.080 ; 
                RECT 798.120 269.760 805.560 270.080 ; 
                RECT 0.160 271.120 75.600 271.440 ; 
                RECT 89.560 271.120 99.400 271.440 ; 
                RECT 798.120 271.120 805.560 271.440 ; 
                RECT 0.160 272.480 75.600 272.800 ; 
                RECT 89.560 272.480 99.400 272.800 ; 
                RECT 798.120 272.480 805.560 272.800 ; 
                RECT 0.160 273.840 75.600 274.160 ; 
                RECT 89.560 273.840 99.400 274.160 ; 
                RECT 798.120 273.840 805.560 274.160 ; 
                RECT 0.160 275.200 75.600 275.520 ; 
                RECT 79.360 275.200 99.400 275.520 ; 
                RECT 798.120 275.200 805.560 275.520 ; 
                RECT 0.160 276.560 80.360 276.880 ; 
                RECT 89.560 276.560 99.400 276.880 ; 
                RECT 798.120 276.560 805.560 276.880 ; 
                RECT 0.160 277.920 75.600 278.240 ; 
                RECT 89.560 277.920 99.400 278.240 ; 
                RECT 798.120 277.920 805.560 278.240 ; 
                RECT 0.160 279.280 75.600 279.600 ; 
                RECT 89.560 279.280 99.400 279.600 ; 
                RECT 798.120 279.280 805.560 279.600 ; 
                RECT 0.160 280.640 77.640 280.960 ; 
                RECT 89.560 280.640 99.400 280.960 ; 
                RECT 798.120 280.640 805.560 280.960 ; 
                RECT 0.160 282.000 75.600 282.320 ; 
                RECT 89.560 282.000 99.400 282.320 ; 
                RECT 798.120 282.000 805.560 282.320 ; 
                RECT 0.160 283.360 75.600 283.680 ; 
                RECT 79.360 283.360 99.400 283.680 ; 
                RECT 798.120 283.360 805.560 283.680 ; 
                RECT 0.160 284.720 82.400 285.040 ; 
                RECT 89.560 284.720 99.400 285.040 ; 
                RECT 798.120 284.720 805.560 285.040 ; 
                RECT 0.160 286.080 75.600 286.400 ; 
                RECT 89.560 286.080 99.400 286.400 ; 
                RECT 798.120 286.080 805.560 286.400 ; 
                RECT 0.160 287.440 75.600 287.760 ; 
                RECT 89.560 287.440 99.400 287.760 ; 
                RECT 798.120 287.440 805.560 287.760 ; 
                RECT 0.160 288.800 75.600 289.120 ; 
                RECT 89.560 288.800 99.400 289.120 ; 
                RECT 798.120 288.800 805.560 289.120 ; 
                RECT 0.160 290.160 75.600 290.480 ; 
                RECT 89.560 290.160 99.400 290.480 ; 
                RECT 798.120 290.160 805.560 290.480 ; 
                RECT 0.160 291.520 99.400 291.840 ; 
                RECT 798.120 291.520 805.560 291.840 ; 
                RECT 0.160 292.880 77.640 293.200 ; 
                RECT 89.560 292.880 99.400 293.200 ; 
                RECT 798.120 292.880 805.560 293.200 ; 
                RECT 0.160 294.240 75.600 294.560 ; 
                RECT 89.560 294.240 99.400 294.560 ; 
                RECT 798.120 294.240 805.560 294.560 ; 
                RECT 0.160 295.600 75.600 295.920 ; 
                RECT 89.560 295.600 99.400 295.920 ; 
                RECT 798.120 295.600 805.560 295.920 ; 
                RECT 0.160 296.960 75.600 297.280 ; 
                RECT 89.560 296.960 99.400 297.280 ; 
                RECT 798.120 296.960 805.560 297.280 ; 
                RECT 0.160 298.320 75.600 298.640 ; 
                RECT 89.560 298.320 99.400 298.640 ; 
                RECT 798.120 298.320 805.560 298.640 ; 
                RECT 0.160 299.680 99.400 300.000 ; 
                RECT 798.120 299.680 805.560 300.000 ; 
                RECT 0.160 301.040 77.640 301.360 ; 
                RECT 89.560 301.040 99.400 301.360 ; 
                RECT 798.120 301.040 805.560 301.360 ; 
                RECT 0.160 302.400 75.600 302.720 ; 
                RECT 89.560 302.400 99.400 302.720 ; 
                RECT 798.120 302.400 805.560 302.720 ; 
                RECT 0.160 303.760 75.600 304.080 ; 
                RECT 89.560 303.760 99.400 304.080 ; 
                RECT 798.120 303.760 805.560 304.080 ; 
                RECT 0.160 305.120 75.600 305.440 ; 
                RECT 89.560 305.120 99.400 305.440 ; 
                RECT 798.120 305.120 805.560 305.440 ; 
                RECT 0.160 306.480 75.600 306.800 ; 
                RECT 89.560 306.480 99.400 306.800 ; 
                RECT 798.120 306.480 805.560 306.800 ; 
                RECT 0.160 307.840 99.400 308.160 ; 
                RECT 798.120 307.840 805.560 308.160 ; 
                RECT 0.160 309.200 75.600 309.520 ; 
                RECT 89.560 309.200 99.400 309.520 ; 
                RECT 798.120 309.200 805.560 309.520 ; 
                RECT 0.160 310.560 75.600 310.880 ; 
                RECT 89.560 310.560 99.400 310.880 ; 
                RECT 798.120 310.560 805.560 310.880 ; 
                RECT 0.160 311.920 75.600 312.240 ; 
                RECT 89.560 311.920 99.400 312.240 ; 
                RECT 798.120 311.920 805.560 312.240 ; 
                RECT 0.160 313.280 75.600 313.600 ; 
                RECT 89.560 313.280 99.400 313.600 ; 
                RECT 798.120 313.280 805.560 313.600 ; 
                RECT 0.160 314.640 75.600 314.960 ; 
                RECT 81.400 314.640 99.400 314.960 ; 
                RECT 798.120 314.640 805.560 314.960 ; 
                RECT 0.160 316.000 99.400 316.320 ; 
                RECT 798.120 316.000 805.560 316.320 ; 
                RECT 0.160 317.360 78.320 317.680 ; 
                RECT 89.560 317.360 99.400 317.680 ; 
                RECT 798.120 317.360 805.560 317.680 ; 
                RECT 0.160 318.720 78.320 319.040 ; 
                RECT 89.560 318.720 99.400 319.040 ; 
                RECT 798.120 318.720 805.560 319.040 ; 
                RECT 0.160 320.080 78.320 320.400 ; 
                RECT 89.560 320.080 99.400 320.400 ; 
                RECT 798.120 320.080 805.560 320.400 ; 
                RECT 0.160 321.440 78.320 321.760 ; 
                RECT 89.560 321.440 99.400 321.760 ; 
                RECT 798.120 321.440 805.560 321.760 ; 
                RECT 0.160 322.800 99.400 323.120 ; 
                RECT 798.120 322.800 805.560 323.120 ; 
                RECT 0.160 324.160 83.760 324.480 ; 
                RECT 89.560 324.160 99.400 324.480 ; 
                RECT 798.120 324.160 805.560 324.480 ; 
                RECT 0.160 325.520 78.320 325.840 ; 
                RECT 89.560 325.520 99.400 325.840 ; 
                RECT 798.120 325.520 805.560 325.840 ; 
                RECT 0.160 326.880 78.320 327.200 ; 
                RECT 89.560 326.880 99.400 327.200 ; 
                RECT 798.120 326.880 805.560 327.200 ; 
                RECT 0.160 328.240 78.320 328.560 ; 
                RECT 89.560 328.240 99.400 328.560 ; 
                RECT 798.120 328.240 805.560 328.560 ; 
                RECT 0.160 329.600 78.320 329.920 ; 
                RECT 89.560 329.600 99.400 329.920 ; 
                RECT 798.120 329.600 805.560 329.920 ; 
                RECT 0.160 330.960 99.400 331.280 ; 
                RECT 798.120 330.960 805.560 331.280 ; 
                RECT 0.160 332.320 78.320 332.640 ; 
                RECT 89.560 332.320 99.400 332.640 ; 
                RECT 798.120 332.320 805.560 332.640 ; 
                RECT 0.160 333.680 86.480 334.000 ; 
                RECT 89.560 333.680 99.400 334.000 ; 
                RECT 798.120 333.680 805.560 334.000 ; 
                RECT 0.160 335.040 78.320 335.360 ; 
                RECT 89.560 335.040 99.400 335.360 ; 
                RECT 798.120 335.040 805.560 335.360 ; 
                RECT 0.160 336.400 78.320 336.720 ; 
                RECT 89.560 336.400 99.400 336.720 ; 
                RECT 798.120 336.400 805.560 336.720 ; 
                RECT 0.160 337.760 78.320 338.080 ; 
                RECT 89.560 337.760 99.400 338.080 ; 
                RECT 798.120 337.760 805.560 338.080 ; 
                RECT 0.160 339.120 99.400 339.440 ; 
                RECT 798.120 339.120 805.560 339.440 ; 
                RECT 0.160 340.480 79.000 340.800 ; 
                RECT 89.560 340.480 99.400 340.800 ; 
                RECT 798.120 340.480 805.560 340.800 ; 
                RECT 0.160 341.840 79.000 342.160 ; 
                RECT 89.560 341.840 99.400 342.160 ; 
                RECT 798.120 341.840 805.560 342.160 ; 
                RECT 0.160 343.200 81.040 343.520 ; 
                RECT 89.560 343.200 99.400 343.520 ; 
                RECT 798.120 343.200 805.560 343.520 ; 
                RECT 0.160 344.560 79.000 344.880 ; 
                RECT 89.560 344.560 99.400 344.880 ; 
                RECT 798.120 344.560 805.560 344.880 ; 
                RECT 0.160 345.920 79.000 346.240 ; 
                RECT 89.560 345.920 99.400 346.240 ; 
                RECT 798.120 345.920 805.560 346.240 ; 
                RECT 0.160 347.280 99.400 347.600 ; 
                RECT 798.120 347.280 805.560 347.600 ; 
                RECT 0.160 348.640 79.000 348.960 ; 
                RECT 89.560 348.640 99.400 348.960 ; 
                RECT 798.120 348.640 805.560 348.960 ; 
                RECT 0.160 350.000 79.000 350.320 ; 
                RECT 89.560 350.000 99.400 350.320 ; 
                RECT 798.120 350.000 805.560 350.320 ; 
                RECT 0.160 351.360 79.000 351.680 ; 
                RECT 89.560 351.360 99.400 351.680 ; 
                RECT 798.120 351.360 805.560 351.680 ; 
                RECT 0.160 352.720 83.760 353.040 ; 
                RECT 89.560 352.720 99.400 353.040 ; 
                RECT 798.120 352.720 805.560 353.040 ; 
                RECT 0.160 354.080 79.000 354.400 ; 
                RECT 89.560 354.080 99.400 354.400 ; 
                RECT 798.120 354.080 805.560 354.400 ; 
                RECT 0.160 355.440 99.400 355.760 ; 
                RECT 798.120 355.440 805.560 355.760 ; 
                RECT 0.160 356.800 79.000 357.120 ; 
                RECT 89.560 356.800 99.400 357.120 ; 
                RECT 798.120 356.800 805.560 357.120 ; 
                RECT 0.160 358.160 79.000 358.480 ; 
                RECT 89.560 358.160 99.400 358.480 ; 
                RECT 798.120 358.160 805.560 358.480 ; 
                RECT 0.160 359.520 79.000 359.840 ; 
                RECT 89.560 359.520 99.400 359.840 ; 
                RECT 798.120 359.520 805.560 359.840 ; 
                RECT 0.160 360.880 79.000 361.200 ; 
                RECT 89.560 360.880 99.400 361.200 ; 
                RECT 798.120 360.880 805.560 361.200 ; 
                RECT 0.160 362.240 99.400 362.560 ; 
                RECT 798.120 362.240 805.560 362.560 ; 
                RECT 0.160 363.600 85.800 363.920 ; 
                RECT 89.560 363.600 99.400 363.920 ; 
                RECT 798.120 363.600 805.560 363.920 ; 
                RECT 0.160 364.960 79.000 365.280 ; 
                RECT 89.560 364.960 99.400 365.280 ; 
                RECT 798.120 364.960 805.560 365.280 ; 
                RECT 0.160 366.320 79.000 366.640 ; 
                RECT 89.560 366.320 99.400 366.640 ; 
                RECT 798.120 366.320 805.560 366.640 ; 
                RECT 0.160 367.680 79.000 368.000 ; 
                RECT 89.560 367.680 99.400 368.000 ; 
                RECT 798.120 367.680 805.560 368.000 ; 
                RECT 0.160 369.040 79.000 369.360 ; 
                RECT 89.560 369.040 99.400 369.360 ; 
                RECT 798.120 369.040 805.560 369.360 ; 
                RECT 0.160 370.400 99.400 370.720 ; 
                RECT 798.120 370.400 805.560 370.720 ; 
                RECT 0.160 371.760 80.360 372.080 ; 
                RECT 89.560 371.760 99.400 372.080 ; 
                RECT 798.120 371.760 805.560 372.080 ; 
                RECT 0.160 373.120 81.040 373.440 ; 
                RECT 89.560 373.120 99.400 373.440 ; 
                RECT 798.120 373.120 805.560 373.440 ; 
                RECT 0.160 374.480 79.000 374.800 ; 
                RECT 89.560 374.480 99.400 374.800 ; 
                RECT 798.120 374.480 805.560 374.800 ; 
                RECT 0.160 375.840 79.000 376.160 ; 
                RECT 89.560 375.840 99.400 376.160 ; 
                RECT 798.120 375.840 805.560 376.160 ; 
                RECT 0.160 377.200 79.000 377.520 ; 
                RECT 89.560 377.200 99.400 377.520 ; 
                RECT 798.120 377.200 805.560 377.520 ; 
                RECT 0.160 378.560 99.400 378.880 ; 
                RECT 798.120 378.560 805.560 378.880 ; 
                RECT 0.160 379.920 79.000 380.240 ; 
                RECT 89.560 379.920 99.400 380.240 ; 
                RECT 798.120 379.920 805.560 380.240 ; 
                RECT 0.160 381.280 79.000 381.600 ; 
                RECT 89.560 381.280 99.400 381.600 ; 
                RECT 798.120 381.280 805.560 381.600 ; 
                RECT 0.160 382.640 83.080 382.960 ; 
                RECT 89.560 382.640 99.400 382.960 ; 
                RECT 798.120 382.640 805.560 382.960 ; 
                RECT 0.160 384.000 79.000 384.320 ; 
                RECT 89.560 384.000 99.400 384.320 ; 
                RECT 798.120 384.000 805.560 384.320 ; 
                RECT 0.160 385.360 79.000 385.680 ; 
                RECT 89.560 385.360 99.400 385.680 ; 
                RECT 798.120 385.360 805.560 385.680 ; 
                RECT 0.160 386.720 99.400 387.040 ; 
                RECT 798.120 386.720 805.560 387.040 ; 
                RECT 0.160 388.080 79.000 388.400 ; 
                RECT 89.560 388.080 99.400 388.400 ; 
                RECT 798.120 388.080 805.560 388.400 ; 
                RECT 0.160 389.440 79.000 389.760 ; 
                RECT 89.560 389.440 99.400 389.760 ; 
                RECT 798.120 389.440 805.560 389.760 ; 
                RECT 0.160 390.800 79.000 391.120 ; 
                RECT 89.560 390.800 99.400 391.120 ; 
                RECT 798.120 390.800 805.560 391.120 ; 
                RECT 0.160 392.160 85.800 392.480 ; 
                RECT 89.560 392.160 99.400 392.480 ; 
                RECT 798.120 392.160 805.560 392.480 ; 
                RECT 0.160 393.520 79.000 393.840 ; 
                RECT 89.560 393.520 99.400 393.840 ; 
                RECT 798.120 393.520 805.560 393.840 ; 
                RECT 0.160 394.880 99.400 395.200 ; 
                RECT 798.120 394.880 805.560 395.200 ; 
                RECT 0.160 396.240 79.000 396.560 ; 
                RECT 89.560 396.240 99.400 396.560 ; 
                RECT 798.120 396.240 805.560 396.560 ; 
                RECT 0.160 397.600 79.000 397.920 ; 
                RECT 89.560 397.600 99.400 397.920 ; 
                RECT 798.120 397.600 805.560 397.920 ; 
                RECT 0.160 398.960 79.000 399.280 ; 
                RECT 89.560 398.960 99.400 399.280 ; 
                RECT 798.120 398.960 805.560 399.280 ; 
                RECT 0.160 400.320 79.000 400.640 ; 
                RECT 89.560 400.320 99.400 400.640 ; 
                RECT 798.120 400.320 805.560 400.640 ; 
                RECT 0.160 401.680 99.400 402.000 ; 
                RECT 798.120 401.680 805.560 402.000 ; 
                RECT 0.160 403.040 80.360 403.360 ; 
                RECT 89.560 403.040 99.400 403.360 ; 
                RECT 798.120 403.040 805.560 403.360 ; 
                RECT 0.160 404.400 79.680 404.720 ; 
                RECT 89.560 404.400 99.400 404.720 ; 
                RECT 798.120 404.400 805.560 404.720 ; 
                RECT 0.160 405.760 79.680 406.080 ; 
                RECT 89.560 405.760 99.400 406.080 ; 
                RECT 798.120 405.760 805.560 406.080 ; 
                RECT 0.160 407.120 79.680 407.440 ; 
                RECT 89.560 407.120 99.400 407.440 ; 
                RECT 798.120 407.120 805.560 407.440 ; 
                RECT 0.160 408.480 79.680 408.800 ; 
                RECT 89.560 408.480 99.400 408.800 ; 
                RECT 798.120 408.480 805.560 408.800 ; 
                RECT 0.160 409.840 99.400 410.160 ; 
                RECT 798.120 409.840 805.560 410.160 ; 
                RECT 0.160 411.200 82.400 411.520 ; 
                RECT 89.560 411.200 99.400 411.520 ; 
                RECT 798.120 411.200 805.560 411.520 ; 
                RECT 0.160 412.560 79.680 412.880 ; 
                RECT 89.560 412.560 99.400 412.880 ; 
                RECT 798.120 412.560 805.560 412.880 ; 
                RECT 0.160 413.920 79.680 414.240 ; 
                RECT 89.560 413.920 99.400 414.240 ; 
                RECT 798.120 413.920 805.560 414.240 ; 
                RECT 0.160 415.280 79.680 415.600 ; 
                RECT 89.560 415.280 99.400 415.600 ; 
                RECT 798.120 415.280 805.560 415.600 ; 
                RECT 0.160 416.640 79.680 416.960 ; 
                RECT 89.560 416.640 99.400 416.960 ; 
                RECT 798.120 416.640 805.560 416.960 ; 
                RECT 0.160 418.000 99.400 418.320 ; 
                RECT 798.120 418.000 805.560 418.320 ; 
                RECT 0.160 419.360 79.680 419.680 ; 
                RECT 89.560 419.360 99.400 419.680 ; 
                RECT 798.120 419.360 805.560 419.680 ; 
                RECT 0.160 420.720 84.440 421.040 ; 
                RECT 89.560 420.720 99.400 421.040 ; 
                RECT 798.120 420.720 805.560 421.040 ; 
                RECT 0.160 422.080 85.120 422.400 ; 
                RECT 89.560 422.080 99.400 422.400 ; 
                RECT 798.120 422.080 805.560 422.400 ; 
                RECT 0.160 423.440 79.680 423.760 ; 
                RECT 89.560 423.440 99.400 423.760 ; 
                RECT 798.120 423.440 805.560 423.760 ; 
                RECT 0.160 424.800 79.680 425.120 ; 
                RECT 89.560 424.800 99.400 425.120 ; 
                RECT 798.120 424.800 805.560 425.120 ; 
                RECT 0.160 426.160 99.400 426.480 ; 
                RECT 798.120 426.160 805.560 426.480 ; 
                RECT 0.160 427.520 79.680 427.840 ; 
                RECT 89.560 427.520 99.400 427.840 ; 
                RECT 798.120 427.520 805.560 427.840 ; 
                RECT 0.160 428.880 79.680 429.200 ; 
                RECT 89.560 428.880 99.400 429.200 ; 
                RECT 798.120 428.880 805.560 429.200 ; 
                RECT 0.160 430.240 87.160 430.560 ; 
                RECT 89.560 430.240 99.400 430.560 ; 
                RECT 798.120 430.240 805.560 430.560 ; 
                RECT 0.160 431.600 87.160 431.920 ; 
                RECT 89.560 431.600 99.400 431.920 ; 
                RECT 798.120 431.600 805.560 431.920 ; 
                RECT 0.160 432.960 79.680 433.280 ; 
                RECT 89.560 432.960 99.400 433.280 ; 
                RECT 798.120 432.960 805.560 433.280 ; 
                RECT 0.160 434.320 99.400 434.640 ; 
                RECT 798.120 434.320 805.560 434.640 ; 
                RECT 0.160 435.680 388.400 436.000 ; 
                RECT 798.120 435.680 805.560 436.000 ; 
                RECT 0.160 437.040 388.400 437.360 ; 
                RECT 798.120 437.040 805.560 437.360 ; 
                RECT 0.160 438.400 388.400 438.720 ; 
                RECT 798.120 438.400 805.560 438.720 ; 
                RECT 0.160 439.760 805.560 440.080 ; 
                RECT 0.160 441.120 805.560 441.440 ; 
                RECT 0.160 442.480 805.560 442.800 ; 
                RECT 0.160 443.840 805.560 444.160 ; 
                RECT 0.160 0.160 805.560 1.520 ; 
                RECT 0.160 448.560 805.560 449.920 ; 
                RECT 392.540 32.220 398.340 33.590 ; 
                RECT 788.440 32.220 794.240 33.590 ; 
                RECT 392.540 37.255 398.340 38.615 ; 
                RECT 788.440 37.255 794.240 38.615 ; 
                RECT 392.540 42.320 398.340 43.720 ; 
                RECT 788.440 42.320 794.240 43.720 ; 
                RECT 392.540 47.495 398.340 48.935 ; 
                RECT 788.440 47.495 794.240 48.935 ; 
                RECT 392.540 52.590 398.340 53.920 ; 
                RECT 788.440 52.590 794.240 53.920 ; 
                RECT 392.540 57.520 398.340 58.850 ; 
                RECT 788.440 57.520 794.240 58.850 ; 
                RECT 392.540 80.140 794.240 80.940 ; 
                RECT 392.540 77.130 794.240 77.930 ; 
                RECT 392.540 102.935 794.240 103.225 ; 
                RECT 392.540 95.555 794.240 99.155 ; 
                RECT 392.540 163.165 794.240 166.765 ; 
                RECT 392.540 65.660 794.240 67.460 ; 
                RECT 392.540 85.030 794.240 85.830 ; 
                RECT 392.540 129.975 794.240 131.775 ; 
                RECT 392.540 16.465 794.240 18.265 ; 
                RECT 103.590 180.395 105.510 434.775 ; 
                RECT 113.805 180.395 115.725 434.775 ; 
                RECT 117.645 180.395 119.565 434.775 ; 
                RECT 130.055 180.395 131.975 434.775 ; 
                RECT 133.895 180.395 135.815 434.775 ; 
                RECT 137.735 180.395 139.655 434.775 ; 
                RECT 141.575 180.395 143.495 434.775 ; 
                RECT 159.220 180.395 161.140 434.775 ; 
                RECT 163.060 180.395 164.980 434.775 ; 
                RECT 166.900 180.395 168.820 434.775 ; 
                RECT 170.740 180.395 172.660 434.775 ; 
                RECT 174.580 180.395 176.500 434.775 ; 
                RECT 178.420 180.395 180.340 434.775 ; 
                RECT 182.260 180.395 184.180 434.775 ; 
                RECT 209.070 180.395 210.990 434.775 ; 
                RECT 212.910 180.395 214.830 434.775 ; 
                RECT 216.750 180.395 218.670 434.775 ; 
                RECT 220.590 180.395 222.510 434.775 ; 
                RECT 224.430 180.395 226.350 434.775 ; 
                RECT 228.270 180.395 230.190 434.775 ; 
                RECT 232.110 180.395 234.030 434.775 ; 
                RECT 235.950 180.395 237.870 434.775 ; 
                RECT 239.790 180.395 241.710 434.775 ; 
                RECT 243.630 180.395 245.550 434.775 ; 
                RECT 247.470 180.395 249.390 434.775 ; 
                RECT 251.310 180.395 253.230 434.775 ; 
                RECT 255.150 180.395 257.070 434.775 ; 
                RECT 298.970 180.395 300.890 434.775 ; 
                RECT 302.810 180.395 304.730 434.775 ; 
                RECT 306.650 180.395 308.570 434.775 ; 
                RECT 310.490 180.395 312.410 434.775 ; 
                RECT 314.330 180.395 316.250 434.775 ; 
                RECT 318.170 180.395 320.090 434.775 ; 
                RECT 322.010 180.395 323.930 434.775 ; 
                RECT 325.850 180.395 327.770 434.775 ; 
                RECT 329.690 180.395 331.610 434.775 ; 
                RECT 333.530 180.395 335.450 434.775 ; 
                RECT 337.370 180.395 339.290 434.775 ; 
                RECT 341.210 180.395 343.130 434.775 ; 
                RECT 345.050 180.395 346.970 434.775 ; 
                RECT 348.890 180.395 350.810 434.775 ; 
                RECT 352.730 180.395 354.650 434.775 ; 
                RECT 356.570 180.395 358.490 434.775 ; 
                RECT 360.410 180.395 362.330 434.775 ; 
                RECT 364.250 180.395 366.170 434.775 ; 
                RECT 368.090 180.395 370.010 434.775 ; 
                RECT 371.930 180.395 373.850 434.775 ; 
                RECT 375.770 180.395 377.690 434.775 ; 
                RECT 379.610 180.395 381.530 434.775 ; 
                RECT 383.450 180.395 385.370 434.775 ; 
                RECT 290.580 61.335 292.500 113.935 ; 
                RECT 297.555 61.335 299.475 113.935 ; 
                RECT 305.390 61.335 307.310 113.935 ; 
                RECT 316.695 61.335 318.615 113.935 ; 
                RECT 320.535 61.335 322.455 113.935 ; 
                RECT 324.375 61.335 326.295 113.935 ; 
                RECT 343.525 61.335 345.445 113.935 ; 
                RECT 347.365 61.335 349.285 113.935 ; 
                RECT 351.205 61.335 353.125 113.935 ; 
                RECT 355.045 61.335 356.965 113.935 ; 
                RECT 358.885 61.335 360.805 113.935 ; 
                RECT 362.725 61.335 364.645 113.935 ; 
                RECT 366.565 61.335 368.485 113.935 ; 
                RECT 370.405 61.335 372.325 113.935 ; 
                RECT 315.500 140.900 317.420 173.760 ; 
                RECT 322.905 140.900 324.825 173.760 ; 
                RECT 329.535 140.900 331.285 173.760 ; 
                RECT 339.005 140.900 340.925 173.760 ; 
                RECT 355.070 140.900 356.990 173.760 ; 
                RECT 358.910 140.900 360.830 173.760 ; 
                RECT 362.750 140.900 364.670 173.760 ; 
                RECT 366.590 140.900 368.510 173.760 ; 
                RECT 370.430 140.900 372.350 173.760 ; 
                RECT 323.515 128.160 325.265 134.900 ; 
                RECT 332.985 128.160 334.905 134.900 ; 
                RECT 351.000 128.160 352.920 134.900 ; 
                RECT 354.840 128.160 356.760 134.900 ; 
                RECT 358.680 128.160 360.600 134.900 ; 
                RECT 362.520 128.160 364.440 134.900 ; 
                RECT 366.360 128.160 368.280 134.900 ; 
                RECT 370.200 128.160 372.120 134.900 ; 
                RECT 371.435 50.175 373.185 55.335 ; 
                RECT 26.230 182.665 35.390 183.415 ; 
                RECT 26.230 187.420 35.390 189.340 ; 
                RECT 230.680 170.375 246.720 171.225 ; 
                RECT 211.480 170.715 228.720 172.745 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 401.320 5.560 ; 
                RECT 787.240 5.240 802.840 5.560 ; 
                RECT 2.880 6.600 802.840 6.920 ; 
                RECT 2.880 7.960 802.840 8.280 ; 
                RECT 2.880 9.320 374.800 9.640 ; 
                RECT 396.920 9.320 802.840 9.640 ; 
                RECT 2.880 10.680 391.120 11.000 ; 
                RECT 796.080 10.680 802.840 11.000 ; 
                RECT 2.880 12.040 391.120 12.360 ; 
                RECT 796.080 12.040 802.840 12.360 ; 
                RECT 2.880 13.400 391.120 13.720 ; 
                RECT 796.080 13.400 802.840 13.720 ; 
                RECT 2.880 14.760 391.120 15.080 ; 
                RECT 796.080 14.760 802.840 15.080 ; 
                RECT 2.880 16.120 391.120 16.440 ; 
                RECT 796.080 16.120 802.840 16.440 ; 
                RECT 2.880 17.480 391.120 17.800 ; 
                RECT 796.080 17.480 802.840 17.800 ; 
                RECT 2.880 18.840 391.120 19.160 ; 
                RECT 796.080 18.840 802.840 19.160 ; 
                RECT 2.880 20.200 306.800 20.520 ; 
                RECT 375.840 20.200 391.120 20.520 ; 
                RECT 796.080 20.200 802.840 20.520 ; 
                RECT 2.880 21.560 391.120 21.880 ; 
                RECT 796.080 21.560 802.840 21.880 ; 
                RECT 2.880 22.920 391.120 23.240 ; 
                RECT 796.080 22.920 802.840 23.240 ; 
                RECT 2.880 24.280 306.800 24.600 ; 
                RECT 375.160 24.280 391.120 24.600 ; 
                RECT 796.080 24.280 802.840 24.600 ; 
                RECT 2.880 25.640 391.120 25.960 ; 
                RECT 796.080 25.640 802.840 25.960 ; 
                RECT 2.880 27.000 391.120 27.320 ; 
                RECT 796.080 27.000 802.840 27.320 ; 
                RECT 2.880 28.360 390.440 28.680 ; 
                RECT 796.080 28.360 802.840 28.680 ; 
                RECT 2.880 29.720 391.120 30.040 ; 
                RECT 796.080 29.720 802.840 30.040 ; 
                RECT 2.880 31.080 391.120 31.400 ; 
                RECT 796.080 31.080 802.840 31.400 ; 
                RECT 2.880 32.440 391.120 32.760 ; 
                RECT 796.080 32.440 802.840 32.760 ; 
                RECT 2.880 33.800 391.120 34.120 ; 
                RECT 796.080 33.800 802.840 34.120 ; 
                RECT 2.880 35.160 391.120 35.480 ; 
                RECT 796.080 35.160 802.840 35.480 ; 
                RECT 2.880 36.520 391.120 36.840 ; 
                RECT 796.080 36.520 802.840 36.840 ; 
                RECT 2.880 37.880 391.120 38.200 ; 
                RECT 796.080 37.880 802.840 38.200 ; 
                RECT 2.880 39.240 391.120 39.560 ; 
                RECT 796.080 39.240 802.840 39.560 ; 
                RECT 2.880 40.600 391.120 40.920 ; 
                RECT 796.080 40.600 802.840 40.920 ; 
                RECT 2.880 41.960 277.560 42.280 ; 
                RECT 354.080 41.960 391.120 42.280 ; 
                RECT 796.080 41.960 802.840 42.280 ; 
                RECT 2.880 43.320 276.200 43.640 ; 
                RECT 360.200 43.320 391.120 43.640 ; 
                RECT 796.080 43.320 802.840 43.640 ; 
                RECT 2.880 44.680 253.080 45.000 ; 
                RECT 375.160 44.680 391.120 45.000 ; 
                RECT 796.080 44.680 802.840 45.000 ; 
                RECT 2.880 46.040 253.760 46.360 ; 
                RECT 365.640 46.040 391.120 46.360 ; 
                RECT 796.080 46.040 802.840 46.360 ; 
                RECT 2.880 47.400 391.120 47.720 ; 
                RECT 796.080 47.400 802.840 47.720 ; 
                RECT 2.880 48.760 391.120 49.080 ; 
                RECT 796.080 48.760 802.840 49.080 ; 
                RECT 2.880 50.120 368.000 50.440 ; 
                RECT 373.800 50.120 391.120 50.440 ; 
                RECT 796.080 50.120 802.840 50.440 ; 
                RECT 2.880 51.480 368.000 51.800 ; 
                RECT 796.080 51.480 802.840 51.800 ; 
                RECT 2.880 52.840 368.000 53.160 ; 
                RECT 796.080 52.840 802.840 53.160 ; 
                RECT 2.880 54.200 368.000 54.520 ; 
                RECT 373.800 54.200 391.120 54.520 ; 
                RECT 796.080 54.200 802.840 54.520 ; 
                RECT 2.880 55.560 368.000 55.880 ; 
                RECT 373.800 55.560 391.120 55.880 ; 
                RECT 796.080 55.560 802.840 55.880 ; 
                RECT 2.880 56.920 391.120 57.240 ; 
                RECT 796.080 56.920 802.840 57.240 ; 
                RECT 2.880 58.280 391.120 58.600 ; 
                RECT 796.080 58.280 802.840 58.600 ; 
                RECT 2.880 59.640 391.120 59.960 ; 
                RECT 796.080 59.640 802.840 59.960 ; 
                RECT 2.880 61.000 286.400 61.320 ; 
                RECT 373.120 61.000 391.120 61.320 ; 
                RECT 796.080 61.000 802.840 61.320 ; 
                RECT 2.880 62.360 276.200 62.680 ; 
                RECT 280.640 62.360 286.400 62.680 ; 
                RECT 373.120 62.360 391.120 62.680 ; 
                RECT 796.080 62.360 802.840 62.680 ; 
                RECT 2.880 63.720 277.560 64.040 ; 
                RECT 279.960 63.720 286.400 64.040 ; 
                RECT 383.320 63.720 391.120 64.040 ; 
                RECT 796.080 63.720 802.840 64.040 ; 
                RECT 2.880 65.080 286.400 65.400 ; 
                RECT 383.320 65.080 391.120 65.400 ; 
                RECT 796.080 65.080 802.840 65.400 ; 
                RECT 2.880 66.440 286.400 66.760 ; 
                RECT 383.320 66.440 391.120 66.760 ; 
                RECT 796.080 66.440 802.840 66.760 ; 
                RECT 2.880 67.800 286.400 68.120 ; 
                RECT 381.960 67.800 391.120 68.120 ; 
                RECT 796.080 67.800 802.840 68.120 ; 
                RECT 2.880 69.160 286.400 69.480 ; 
                RECT 383.320 69.160 391.120 69.480 ; 
                RECT 796.080 69.160 802.840 69.480 ; 
                RECT 2.880 70.520 251.040 70.840 ; 
                RECT 262.280 70.520 286.400 70.840 ; 
                RECT 373.120 70.520 391.120 70.840 ; 
                RECT 796.080 70.520 802.840 70.840 ; 
                RECT 2.880 71.880 252.400 72.200 ; 
                RECT 256.160 71.880 286.400 72.200 ; 
                RECT 383.320 71.880 391.120 72.200 ; 
                RECT 796.080 71.880 802.840 72.200 ; 
                RECT 2.880 73.240 253.760 73.560 ; 
                RECT 258.200 73.240 266.000 73.560 ; 
                RECT 268.400 73.240 286.400 73.560 ; 
                RECT 383.320 73.240 391.120 73.560 ; 
                RECT 796.080 73.240 802.840 73.560 ; 
                RECT 2.880 74.600 286.400 74.920 ; 
                RECT 381.960 74.600 391.120 74.920 ; 
                RECT 796.080 74.600 802.840 74.920 ; 
                RECT 2.880 75.960 260.560 76.280 ; 
                RECT 269.080 75.960 286.400 76.280 ; 
                RECT 386.040 75.960 391.120 76.280 ; 
                RECT 796.080 75.960 802.840 76.280 ; 
                RECT 2.880 77.320 253.080 77.640 ; 
                RECT 262.280 77.320 286.400 77.640 ; 
                RECT 386.040 77.320 391.120 77.640 ; 
                RECT 796.080 77.320 802.840 77.640 ; 
                RECT 2.880 78.680 256.480 79.000 ; 
                RECT 261.600 78.680 286.400 79.000 ; 
                RECT 373.120 78.680 391.120 79.000 ; 
                RECT 796.080 78.680 802.840 79.000 ; 
                RECT 2.880 80.040 286.400 80.360 ; 
                RECT 386.040 80.040 391.120 80.360 ; 
                RECT 796.080 80.040 802.840 80.360 ; 
                RECT 2.880 81.400 250.360 81.720 ; 
                RECT 262.280 81.400 286.400 81.720 ; 
                RECT 384.680 81.400 391.120 81.720 ; 
                RECT 796.080 81.400 802.840 81.720 ; 
                RECT 2.880 82.760 260.560 83.080 ; 
                RECT 268.400 82.760 286.400 83.080 ; 
                RECT 386.040 82.760 391.120 83.080 ; 
                RECT 796.080 82.760 802.840 83.080 ; 
                RECT 2.880 84.120 259.200 84.440 ; 
                RECT 262.280 84.120 286.400 84.440 ; 
                RECT 386.040 84.120 391.120 84.440 ; 
                RECT 796.080 84.120 802.840 84.440 ; 
                RECT 2.880 85.480 286.400 85.800 ; 
                RECT 386.040 85.480 391.120 85.800 ; 
                RECT 796.080 85.480 802.840 85.800 ; 
                RECT 2.880 86.840 260.560 87.160 ; 
                RECT 268.400 86.840 286.400 87.160 ; 
                RECT 384.680 86.840 391.120 87.160 ; 
                RECT 796.080 86.840 802.840 87.160 ; 
                RECT 2.880 88.200 257.160 88.520 ; 
                RECT 262.280 88.200 286.400 88.520 ; 
                RECT 373.120 88.200 391.120 88.520 ; 
                RECT 796.080 88.200 802.840 88.520 ; 
                RECT 2.880 89.560 259.200 89.880 ; 
                RECT 262.280 89.560 286.400 89.880 ; 
                RECT 388.760 89.560 391.120 89.880 ; 
                RECT 796.080 89.560 802.840 89.880 ; 
                RECT 2.880 90.920 263.280 91.240 ; 
                RECT 273.840 90.920 286.400 91.240 ; 
                RECT 388.760 90.920 391.120 91.240 ; 
                RECT 796.080 90.920 802.840 91.240 ; 
                RECT 2.880 92.280 251.040 92.600 ; 
                RECT 268.400 92.280 286.400 92.600 ; 
                RECT 388.760 92.280 391.120 92.600 ; 
                RECT 796.080 92.280 802.840 92.600 ; 
                RECT 2.880 93.640 259.200 93.960 ; 
                RECT 262.280 93.640 269.400 93.960 ; 
                RECT 275.200 93.640 286.400 93.960 ; 
                RECT 387.400 93.640 391.120 93.960 ; 
                RECT 796.080 93.640 802.840 93.960 ; 
                RECT 2.880 95.000 272.120 95.320 ; 
                RECT 275.880 95.000 286.400 95.320 ; 
                RECT 388.760 95.000 391.120 95.320 ; 
                RECT 796.080 95.000 802.840 95.320 ; 
                RECT 2.880 96.360 251.040 96.680 ; 
                RECT 265.000 96.360 286.400 96.680 ; 
                RECT 373.120 96.360 391.120 96.680 ; 
                RECT 796.080 96.360 802.840 96.680 ; 
                RECT 2.880 97.720 259.880 98.040 ; 
                RECT 268.400 97.720 286.400 98.040 ; 
                RECT 388.760 97.720 391.120 98.040 ; 
                RECT 796.080 97.720 802.840 98.040 ; 
                RECT 2.880 99.080 257.840 99.400 ; 
                RECT 269.080 99.080 286.400 99.400 ; 
                RECT 388.760 99.080 391.120 99.400 ; 
                RECT 796.080 99.080 802.840 99.400 ; 
                RECT 2.880 100.440 286.400 100.760 ; 
                RECT 387.400 100.440 391.120 100.760 ; 
                RECT 796.080 100.440 802.840 100.760 ; 
                RECT 2.880 101.800 253.760 102.120 ; 
                RECT 256.160 101.800 286.400 102.120 ; 
                RECT 796.080 101.800 802.840 102.120 ; 
                RECT 2.880 103.160 253.080 103.480 ; 
                RECT 262.280 103.160 286.400 103.480 ; 
                RECT 796.080 103.160 802.840 103.480 ; 
                RECT 2.880 104.520 255.800 104.840 ; 
                RECT 259.560 104.520 286.400 104.840 ; 
                RECT 373.120 104.520 391.120 104.840 ; 
                RECT 796.080 104.520 802.840 104.840 ; 
                RECT 2.880 105.880 286.400 106.200 ; 
                RECT 796.080 105.880 802.840 106.200 ; 
                RECT 2.880 107.240 259.200 107.560 ; 
                RECT 261.600 107.240 286.400 107.560 ; 
                RECT 796.080 107.240 802.840 107.560 ; 
                RECT 2.880 108.600 252.400 108.920 ; 
                RECT 267.720 108.600 286.400 108.920 ; 
                RECT 796.080 108.600 802.840 108.920 ; 
                RECT 2.880 109.960 259.200 110.280 ; 
                RECT 261.600 109.960 286.400 110.280 ; 
                RECT 796.080 109.960 802.840 110.280 ; 
                RECT 2.880 111.320 286.400 111.640 ; 
                RECT 796.080 111.320 802.840 111.640 ; 
                RECT 2.880 112.680 254.440 113.000 ; 
                RECT 262.280 112.680 286.400 113.000 ; 
                RECT 796.080 112.680 802.840 113.000 ; 
                RECT 2.880 114.040 251.040 114.360 ; 
                RECT 262.280 114.040 286.400 114.360 ; 
                RECT 373.120 114.040 391.120 114.360 ; 
                RECT 796.080 114.040 802.840 114.360 ; 
                RECT 2.880 115.400 391.120 115.720 ; 
                RECT 796.080 115.400 802.840 115.720 ; 
                RECT 2.880 116.760 250.360 117.080 ; 
                RECT 268.400 116.760 377.520 117.080 ; 
                RECT 796.080 116.760 802.840 117.080 ; 
                RECT 2.880 118.120 247.640 118.440 ; 
                RECT 260.920 118.120 388.400 118.440 ; 
                RECT 796.080 118.120 802.840 118.440 ; 
                RECT 2.880 119.480 251.040 119.800 ; 
                RECT 265.000 119.480 385.680 119.800 ; 
                RECT 796.080 119.480 802.840 119.800 ; 
                RECT 2.880 120.840 266.680 121.160 ; 
                RECT 268.400 120.840 382.960 121.160 ; 
                RECT 796.080 120.840 802.840 121.160 ; 
                RECT 2.880 122.200 380.240 122.520 ; 
                RECT 796.080 122.200 802.840 122.520 ; 
                RECT 2.880 123.560 229.280 123.880 ; 
                RECT 248.000 123.560 263.280 123.880 ; 
                RECT 271.120 123.560 391.120 123.880 ; 
                RECT 796.080 123.560 802.840 123.880 ; 
                RECT 2.880 124.920 229.280 125.240 ; 
                RECT 248.000 124.920 391.120 125.240 ; 
                RECT 796.080 124.920 802.840 125.240 ; 
                RECT 2.880 126.280 229.280 126.600 ; 
                RECT 248.000 126.280 391.120 126.600 ; 
                RECT 796.080 126.280 802.840 126.600 ; 
                RECT 2.880 127.640 229.280 127.960 ; 
                RECT 248.000 127.640 253.080 127.960 ; 
                RECT 256.160 127.640 320.400 127.960 ; 
                RECT 373.120 127.640 391.120 127.960 ; 
                RECT 796.080 127.640 802.840 127.960 ; 
                RECT 2.880 129.000 229.280 129.320 ; 
                RECT 248.000 129.000 251.040 129.320 ; 
                RECT 254.800 129.000 320.400 129.320 ; 
                RECT 373.120 129.000 391.120 129.320 ; 
                RECT 796.080 129.000 802.840 129.320 ; 
                RECT 2.880 130.360 229.280 130.680 ; 
                RECT 248.000 130.360 320.400 130.680 ; 
                RECT 373.120 130.360 391.120 130.680 ; 
                RECT 796.080 130.360 802.840 130.680 ; 
                RECT 2.880 131.720 229.280 132.040 ; 
                RECT 248.000 131.720 256.480 132.040 ; 
                RECT 268.400 131.720 320.400 132.040 ; 
                RECT 373.120 131.720 391.120 132.040 ; 
                RECT 796.080 131.720 802.840 132.040 ; 
                RECT 2.880 133.080 229.280 133.400 ; 
                RECT 248.000 133.080 320.400 133.400 ; 
                RECT 373.120 133.080 391.120 133.400 ; 
                RECT 796.080 133.080 802.840 133.400 ; 
                RECT 2.880 134.440 229.280 134.760 ; 
                RECT 248.000 134.440 320.400 134.760 ; 
                RECT 373.120 134.440 391.120 134.760 ; 
                RECT 796.080 134.440 802.840 134.760 ; 
                RECT 2.880 135.800 229.280 136.120 ; 
                RECT 248.000 135.800 391.120 136.120 ; 
                RECT 796.080 135.800 802.840 136.120 ; 
                RECT 2.880 137.160 229.280 137.480 ; 
                RECT 248.000 137.160 253.080 137.480 ; 
                RECT 258.200 137.160 391.120 137.480 ; 
                RECT 796.080 137.160 802.840 137.480 ; 
                RECT 2.880 138.520 229.280 138.840 ; 
                RECT 248.000 138.520 391.120 138.840 ; 
                RECT 796.080 138.520 802.840 138.840 ; 
                RECT 2.880 139.880 229.280 140.200 ; 
                RECT 248.000 139.880 266.680 140.200 ; 
                RECT 269.080 139.880 391.120 140.200 ; 
                RECT 796.080 139.880 802.840 140.200 ; 
                RECT 2.880 141.240 229.280 141.560 ; 
                RECT 248.680 141.240 310.880 141.560 ; 
                RECT 373.120 141.240 391.120 141.560 ; 
                RECT 796.080 141.240 802.840 141.560 ; 
                RECT 2.880 142.600 229.280 142.920 ; 
                RECT 248.000 142.600 310.880 142.920 ; 
                RECT 373.120 142.600 391.120 142.920 ; 
                RECT 796.080 142.600 802.840 142.920 ; 
                RECT 2.880 143.960 229.280 144.280 ; 
                RECT 248.000 143.960 252.400 144.280 ; 
                RECT 255.480 143.960 310.880 144.280 ; 
                RECT 373.120 143.960 391.120 144.280 ; 
                RECT 796.080 143.960 802.840 144.280 ; 
                RECT 2.880 145.320 229.280 145.640 ; 
                RECT 248.000 145.320 310.880 145.640 ; 
                RECT 373.120 145.320 391.120 145.640 ; 
                RECT 796.080 145.320 802.840 145.640 ; 
                RECT 2.880 146.680 229.280 147.000 ; 
                RECT 248.000 146.680 310.880 147.000 ; 
                RECT 373.120 146.680 391.120 147.000 ; 
                RECT 796.080 146.680 802.840 147.000 ; 
                RECT 2.880 148.040 229.280 148.360 ; 
                RECT 248.000 148.040 310.880 148.360 ; 
                RECT 373.120 148.040 391.120 148.360 ; 
                RECT 796.080 148.040 802.840 148.360 ; 
                RECT 2.880 149.400 229.280 149.720 ; 
                RECT 248.000 149.400 259.200 149.720 ; 
                RECT 268.400 149.400 310.880 149.720 ; 
                RECT 373.120 149.400 381.600 149.720 ; 
                RECT 796.080 149.400 802.840 149.720 ; 
                RECT 2.880 150.760 229.280 151.080 ; 
                RECT 248.000 150.760 310.880 151.080 ; 
                RECT 373.120 150.760 384.320 151.080 ; 
                RECT 796.080 150.760 802.840 151.080 ; 
                RECT 2.880 152.120 229.280 152.440 ; 
                RECT 248.000 152.120 255.800 152.440 ; 
                RECT 258.200 152.120 310.880 152.440 ; 
                RECT 373.120 152.120 387.040 152.440 ; 
                RECT 796.080 152.120 802.840 152.440 ; 
                RECT 2.880 153.480 229.280 153.800 ; 
                RECT 248.000 153.480 310.880 153.800 ; 
                RECT 373.120 153.480 389.760 153.800 ; 
                RECT 796.080 153.480 802.840 153.800 ; 
                RECT 2.880 154.840 229.280 155.160 ; 
                RECT 248.000 154.840 310.880 155.160 ; 
                RECT 796.080 154.840 802.840 155.160 ; 
                RECT 2.880 156.200 229.280 156.520 ; 
                RECT 248.000 156.200 310.880 156.520 ; 
                RECT 796.080 156.200 802.840 156.520 ; 
                RECT 2.880 157.560 229.280 157.880 ; 
                RECT 248.000 157.560 310.880 157.880 ; 
                RECT 373.120 157.560 391.120 157.880 ; 
                RECT 796.080 157.560 802.840 157.880 ; 
                RECT 2.880 158.920 229.280 159.240 ; 
                RECT 248.000 158.920 310.880 159.240 ; 
                RECT 373.120 158.920 391.120 159.240 ; 
                RECT 796.080 158.920 802.840 159.240 ; 
                RECT 2.880 160.280 229.280 160.600 ; 
                RECT 248.000 160.280 310.880 160.600 ; 
                RECT 373.120 160.280 391.120 160.600 ; 
                RECT 796.080 160.280 802.840 160.600 ; 
                RECT 2.880 161.640 229.280 161.960 ; 
                RECT 248.000 161.640 310.880 161.960 ; 
                RECT 373.120 161.640 391.120 161.960 ; 
                RECT 796.080 161.640 802.840 161.960 ; 
                RECT 2.880 163.000 254.440 163.320 ; 
                RECT 258.200 163.000 310.880 163.320 ; 
                RECT 373.120 163.000 391.120 163.320 ; 
                RECT 796.080 163.000 802.840 163.320 ; 
                RECT 2.880 164.360 310.880 164.680 ; 
                RECT 373.120 164.360 391.120 164.680 ; 
                RECT 796.080 164.360 802.840 164.680 ; 
                RECT 2.880 165.720 310.880 166.040 ; 
                RECT 373.120 165.720 391.120 166.040 ; 
                RECT 796.080 165.720 802.840 166.040 ; 
                RECT 2.880 167.080 210.920 167.400 ; 
                RECT 229.640 167.080 256.480 167.400 ; 
                RECT 262.280 167.080 310.880 167.400 ; 
                RECT 373.120 167.080 391.120 167.400 ; 
                RECT 796.080 167.080 802.840 167.400 ; 
                RECT 2.880 168.440 210.920 168.760 ; 
                RECT 229.640 168.440 235.400 168.760 ; 
                RECT 242.560 168.440 310.880 168.760 ; 
                RECT 373.120 168.440 391.120 168.760 ; 
                RECT 796.080 168.440 802.840 168.760 ; 
                RECT 2.880 169.800 210.920 170.120 ; 
                RECT 247.320 169.800 310.880 170.120 ; 
                RECT 373.120 169.800 391.120 170.120 ; 
                RECT 796.080 169.800 802.840 170.120 ; 
                RECT 2.880 171.160 210.920 171.480 ; 
                RECT 247.320 171.160 310.880 171.480 ; 
                RECT 796.080 171.160 802.840 171.480 ; 
                RECT 2.880 172.520 210.920 172.840 ; 
                RECT 229.640 172.520 235.400 172.840 ; 
                RECT 242.560 172.520 251.040 172.840 ; 
                RECT 260.920 172.520 310.880 172.840 ; 
                RECT 796.080 172.520 802.840 172.840 ; 
                RECT 2.880 173.880 208.200 174.200 ; 
                RECT 241.880 173.880 310.880 174.200 ; 
                RECT 373.120 173.880 802.840 174.200 ; 
                RECT 2.880 175.240 241.520 175.560 ; 
                RECT 308.520 175.240 802.840 175.560 ; 
                RECT 2.880 176.600 388.400 176.920 ; 
                RECT 798.120 176.600 802.840 176.920 ; 
                RECT 2.880 177.960 388.400 178.280 ; 
                RECT 798.120 177.960 802.840 178.280 ; 
                RECT 2.880 179.320 388.400 179.640 ; 
                RECT 798.120 179.320 802.840 179.640 ; 
                RECT 2.880 180.680 27.320 181.000 ; 
                RECT 33.800 180.680 36.160 181.000 ; 
                RECT 48.760 180.680 99.400 181.000 ; 
                RECT 798.120 180.680 802.840 181.000 ; 
                RECT 2.880 182.040 25.280 182.360 ; 
                RECT 48.080 182.040 59.280 182.360 ; 
                RECT 61.000 182.040 75.600 182.360 ; 
                RECT 89.560 182.040 99.400 182.360 ; 
                RECT 798.120 182.040 802.840 182.360 ; 
                RECT 2.880 183.400 25.280 183.720 ; 
                RECT 35.840 183.400 59.280 183.720 ; 
                RECT 63.720 183.400 75.600 183.720 ; 
                RECT 89.560 183.400 99.400 183.720 ; 
                RECT 798.120 183.400 802.840 183.720 ; 
                RECT 2.880 184.760 25.280 185.080 ; 
                RECT 35.840 184.760 59.280 185.080 ; 
                RECT 63.720 184.760 75.600 185.080 ; 
                RECT 89.560 184.760 99.400 185.080 ; 
                RECT 798.120 184.760 802.840 185.080 ; 
                RECT 2.880 186.120 59.280 186.440 ; 
                RECT 64.400 186.120 75.600 186.440 ; 
                RECT 89.560 186.120 99.400 186.440 ; 
                RECT 798.120 186.120 802.840 186.440 ; 
                RECT 2.880 187.480 25.280 187.800 ; 
                RECT 35.840 187.480 59.280 187.800 ; 
                RECT 61.000 187.480 75.600 187.800 ; 
                RECT 89.560 187.480 99.400 187.800 ; 
                RECT 798.120 187.480 802.840 187.800 ; 
                RECT 2.880 188.840 25.280 189.160 ; 
                RECT 35.840 188.840 99.400 189.160 ; 
                RECT 798.120 188.840 802.840 189.160 ; 
                RECT 2.880 190.200 75.600 190.520 ; 
                RECT 89.560 190.200 99.400 190.520 ; 
                RECT 798.120 190.200 802.840 190.520 ; 
                RECT 2.880 191.560 75.600 191.880 ; 
                RECT 89.560 191.560 99.400 191.880 ; 
                RECT 798.120 191.560 802.840 191.880 ; 
                RECT 2.880 192.920 75.600 193.240 ; 
                RECT 89.560 192.920 99.400 193.240 ; 
                RECT 798.120 192.920 802.840 193.240 ; 
                RECT 2.880 194.280 18.480 194.600 ; 
                RECT 20.880 194.280 34.120 194.600 ; 
                RECT 37.200 194.280 75.600 194.600 ; 
                RECT 89.560 194.280 99.400 194.600 ; 
                RECT 798.120 194.280 802.840 194.600 ; 
                RECT 2.880 195.640 17.800 195.960 ; 
                RECT 20.880 195.640 34.120 195.960 ; 
                RECT 37.880 195.640 75.600 195.960 ; 
                RECT 89.560 195.640 99.400 195.960 ; 
                RECT 798.120 195.640 802.840 195.960 ; 
                RECT 2.880 197.000 17.120 197.320 ; 
                RECT 20.880 197.000 39.560 197.320 ; 
                RECT 48.760 197.000 99.400 197.320 ; 
                RECT 798.120 197.000 802.840 197.320 ; 
                RECT 2.880 198.360 16.440 198.680 ; 
                RECT 20.880 198.360 40.920 198.680 ; 
                RECT 47.400 198.360 59.280 198.680 ; 
                RECT 61.000 198.360 75.600 198.680 ; 
                RECT 89.560 198.360 99.400 198.680 ; 
                RECT 798.120 198.360 802.840 198.680 ; 
                RECT 2.880 199.720 59.280 200.040 ; 
                RECT 61.680 199.720 75.600 200.040 ; 
                RECT 89.560 199.720 99.400 200.040 ; 
                RECT 798.120 199.720 802.840 200.040 ; 
                RECT 2.880 201.080 15.760 201.400 ; 
                RECT 20.880 201.080 59.280 201.400 ; 
                RECT 62.360 201.080 75.600 201.400 ; 
                RECT 89.560 201.080 99.400 201.400 ; 
                RECT 798.120 201.080 802.840 201.400 ; 
                RECT 2.880 202.440 15.080 202.760 ; 
                RECT 20.880 202.440 59.280 202.760 ; 
                RECT 62.360 202.440 75.600 202.760 ; 
                RECT 89.560 202.440 99.400 202.760 ; 
                RECT 798.120 202.440 802.840 202.760 ; 
                RECT 2.880 203.800 59.280 204.120 ; 
                RECT 63.040 203.800 75.600 204.120 ; 
                RECT 89.560 203.800 99.400 204.120 ; 
                RECT 798.120 203.800 802.840 204.120 ; 
                RECT 2.880 205.160 14.400 205.480 ; 
                RECT 20.880 205.160 99.400 205.480 ; 
                RECT 798.120 205.160 802.840 205.480 ; 
                RECT 2.880 206.520 13.720 206.840 ; 
                RECT 20.880 206.520 34.120 206.840 ; 
                RECT 41.960 206.520 75.600 206.840 ; 
                RECT 89.560 206.520 99.400 206.840 ; 
                RECT 798.120 206.520 802.840 206.840 ; 
                RECT 2.880 207.880 75.600 208.200 ; 
                RECT 89.560 207.880 99.400 208.200 ; 
                RECT 798.120 207.880 802.840 208.200 ; 
                RECT 2.880 209.240 13.040 209.560 ; 
                RECT 20.880 209.240 34.120 209.560 ; 
                RECT 40.600 209.240 75.600 209.560 ; 
                RECT 89.560 209.240 99.400 209.560 ; 
                RECT 798.120 209.240 802.840 209.560 ; 
                RECT 2.880 210.600 12.360 210.920 ; 
                RECT 20.880 210.600 34.120 210.920 ; 
                RECT 39.920 210.600 75.600 210.920 ; 
                RECT 89.560 210.600 99.400 210.920 ; 
                RECT 798.120 210.600 802.840 210.920 ; 
                RECT 2.880 211.960 11.680 212.280 ; 
                RECT 20.880 211.960 34.120 212.280 ; 
                RECT 39.240 211.960 75.600 212.280 ; 
                RECT 85.480 211.960 99.400 212.280 ; 
                RECT 798.120 211.960 802.840 212.280 ; 
                RECT 2.880 213.320 11.000 213.640 ; 
                RECT 20.880 213.320 80.360 213.640 ; 
                RECT 89.560 213.320 99.400 213.640 ; 
                RECT 798.120 213.320 802.840 213.640 ; 
                RECT 2.880 214.680 75.600 215.000 ; 
                RECT 89.560 214.680 99.400 215.000 ; 
                RECT 798.120 214.680 802.840 215.000 ; 
                RECT 2.880 216.040 10.320 216.360 ; 
                RECT 20.880 216.040 34.120 216.360 ; 
                RECT 37.880 216.040 75.600 216.360 ; 
                RECT 89.560 216.040 99.400 216.360 ; 
                RECT 798.120 216.040 802.840 216.360 ; 
                RECT 2.880 217.400 9.640 217.720 ; 
                RECT 20.880 217.400 75.600 217.720 ; 
                RECT 89.560 217.400 99.400 217.720 ; 
                RECT 798.120 217.400 802.840 217.720 ; 
                RECT 2.880 218.760 75.600 219.080 ; 
                RECT 89.560 218.760 99.400 219.080 ; 
                RECT 798.120 218.760 802.840 219.080 ; 
                RECT 2.880 220.120 75.600 220.440 ; 
                RECT 86.160 220.120 99.400 220.440 ; 
                RECT 798.120 220.120 802.840 220.440 ; 
                RECT 2.880 221.480 75.600 221.800 ; 
                RECT 89.560 221.480 99.400 221.800 ; 
                RECT 798.120 221.480 802.840 221.800 ; 
                RECT 2.880 222.840 75.600 223.160 ; 
                RECT 89.560 222.840 99.400 223.160 ; 
                RECT 798.120 222.840 802.840 223.160 ; 
                RECT 2.880 224.200 75.600 224.520 ; 
                RECT 89.560 224.200 99.400 224.520 ; 
                RECT 798.120 224.200 802.840 224.520 ; 
                RECT 2.880 225.560 75.600 225.880 ; 
                RECT 89.560 225.560 99.400 225.880 ; 
                RECT 798.120 225.560 802.840 225.880 ; 
                RECT 2.880 226.920 75.600 227.240 ; 
                RECT 89.560 226.920 99.400 227.240 ; 
                RECT 798.120 226.920 802.840 227.240 ; 
                RECT 2.880 228.280 75.600 228.600 ; 
                RECT 87.520 228.280 99.400 228.600 ; 
                RECT 798.120 228.280 802.840 228.600 ; 
                RECT 2.880 229.640 75.600 229.960 ; 
                RECT 89.560 229.640 99.400 229.960 ; 
                RECT 798.120 229.640 802.840 229.960 ; 
                RECT 2.880 231.000 75.600 231.320 ; 
                RECT 89.560 231.000 99.400 231.320 ; 
                RECT 798.120 231.000 802.840 231.320 ; 
                RECT 2.880 232.360 75.600 232.680 ; 
                RECT 89.560 232.360 99.400 232.680 ; 
                RECT 798.120 232.360 802.840 232.680 ; 
                RECT 2.880 233.720 75.600 234.040 ; 
                RECT 89.560 233.720 99.400 234.040 ; 
                RECT 798.120 233.720 802.840 234.040 ; 
                RECT 2.880 235.080 75.600 235.400 ; 
                RECT 89.560 235.080 99.400 235.400 ; 
                RECT 798.120 235.080 802.840 235.400 ; 
                RECT 2.880 236.440 99.400 236.760 ; 
                RECT 798.120 236.440 802.840 236.760 ; 
                RECT 2.880 237.800 75.600 238.120 ; 
                RECT 89.560 237.800 99.400 238.120 ; 
                RECT 798.120 237.800 802.840 238.120 ; 
                RECT 2.880 239.160 75.600 239.480 ; 
                RECT 89.560 239.160 99.400 239.480 ; 
                RECT 798.120 239.160 802.840 239.480 ; 
                RECT 2.880 240.520 75.600 240.840 ; 
                RECT 89.560 240.520 99.400 240.840 ; 
                RECT 798.120 240.520 802.840 240.840 ; 
                RECT 2.880 241.880 75.600 242.200 ; 
                RECT 89.560 241.880 99.400 242.200 ; 
                RECT 798.120 241.880 802.840 242.200 ; 
                RECT 2.880 243.240 75.600 243.560 ; 
                RECT 89.560 243.240 99.400 243.560 ; 
                RECT 798.120 243.240 802.840 243.560 ; 
                RECT 2.880 244.600 99.400 244.920 ; 
                RECT 798.120 244.600 802.840 244.920 ; 
                RECT 2.880 245.960 77.640 246.280 ; 
                RECT 89.560 245.960 99.400 246.280 ; 
                RECT 798.120 245.960 802.840 246.280 ; 
                RECT 2.880 247.320 77.640 247.640 ; 
                RECT 89.560 247.320 99.400 247.640 ; 
                RECT 798.120 247.320 802.840 247.640 ; 
                RECT 2.880 248.680 77.640 249.000 ; 
                RECT 89.560 248.680 99.400 249.000 ; 
                RECT 798.120 248.680 802.840 249.000 ; 
                RECT 2.880 250.040 81.720 250.360 ; 
                RECT 89.560 250.040 99.400 250.360 ; 
                RECT 798.120 250.040 802.840 250.360 ; 
                RECT 2.880 251.400 77.640 251.720 ; 
                RECT 89.560 251.400 99.400 251.720 ; 
                RECT 798.120 251.400 802.840 251.720 ; 
                RECT 2.880 252.760 38.880 253.080 ; 
                RECT 65.080 252.760 99.400 253.080 ; 
                RECT 798.120 252.760 802.840 253.080 ; 
                RECT 2.880 254.120 37.520 254.440 ; 
                RECT 63.720 254.120 75.600 254.440 ; 
                RECT 89.560 254.120 99.400 254.440 ; 
                RECT 798.120 254.120 802.840 254.440 ; 
                RECT 2.880 255.480 36.160 255.800 ; 
                RECT 63.040 255.480 75.600 255.800 ; 
                RECT 89.560 255.480 99.400 255.800 ; 
                RECT 798.120 255.480 802.840 255.800 ; 
                RECT 2.880 256.840 77.640 257.160 ; 
                RECT 89.560 256.840 99.400 257.160 ; 
                RECT 798.120 256.840 802.840 257.160 ; 
                RECT 2.880 258.200 75.600 258.520 ; 
                RECT 89.560 258.200 99.400 258.520 ; 
                RECT 798.120 258.200 802.840 258.520 ; 
                RECT 2.880 259.560 75.600 259.880 ; 
                RECT 78.000 259.560 99.400 259.880 ; 
                RECT 798.120 259.560 802.840 259.880 ; 
                RECT 2.880 260.920 83.760 261.240 ; 
                RECT 89.560 260.920 99.400 261.240 ; 
                RECT 798.120 260.920 802.840 261.240 ; 
                RECT 2.880 262.280 75.600 262.600 ; 
                RECT 89.560 262.280 99.400 262.600 ; 
                RECT 798.120 262.280 802.840 262.600 ; 
                RECT 2.880 263.640 75.600 263.960 ; 
                RECT 89.560 263.640 99.400 263.960 ; 
                RECT 798.120 263.640 802.840 263.960 ; 
                RECT 2.880 265.000 75.600 265.320 ; 
                RECT 89.560 265.000 99.400 265.320 ; 
                RECT 798.120 265.000 802.840 265.320 ; 
                RECT 2.880 266.360 75.600 266.680 ; 
                RECT 89.560 266.360 99.400 266.680 ; 
                RECT 798.120 266.360 802.840 266.680 ; 
                RECT 2.880 267.720 75.600 268.040 ; 
                RECT 78.680 267.720 99.400 268.040 ; 
                RECT 798.120 267.720 802.840 268.040 ; 
                RECT 2.880 269.080 85.800 269.400 ; 
                RECT 89.560 269.080 99.400 269.400 ; 
                RECT 798.120 269.080 802.840 269.400 ; 
                RECT 2.880 270.440 75.600 270.760 ; 
                RECT 89.560 270.440 99.400 270.760 ; 
                RECT 798.120 270.440 802.840 270.760 ; 
                RECT 2.880 271.800 75.600 272.120 ; 
                RECT 89.560 271.800 99.400 272.120 ; 
                RECT 798.120 271.800 802.840 272.120 ; 
                RECT 2.880 273.160 75.600 273.480 ; 
                RECT 89.560 273.160 99.400 273.480 ; 
                RECT 798.120 273.160 802.840 273.480 ; 
                RECT 2.880 274.520 75.600 274.840 ; 
                RECT 89.560 274.520 99.400 274.840 ; 
                RECT 798.120 274.520 802.840 274.840 ; 
                RECT 2.880 275.880 99.400 276.200 ; 
                RECT 798.120 275.880 802.840 276.200 ; 
                RECT 2.880 277.240 77.640 277.560 ; 
                RECT 89.560 277.240 99.400 277.560 ; 
                RECT 798.120 277.240 802.840 277.560 ; 
                RECT 2.880 278.600 75.600 278.920 ; 
                RECT 89.560 278.600 99.400 278.920 ; 
                RECT 798.120 278.600 802.840 278.920 ; 
                RECT 2.880 279.960 75.600 280.280 ; 
                RECT 89.560 279.960 99.400 280.280 ; 
                RECT 798.120 279.960 802.840 280.280 ; 
                RECT 2.880 281.320 75.600 281.640 ; 
                RECT 89.560 281.320 99.400 281.640 ; 
                RECT 798.120 281.320 802.840 281.640 ; 
                RECT 2.880 282.680 75.600 283.000 ; 
                RECT 89.560 282.680 99.400 283.000 ; 
                RECT 798.120 282.680 802.840 283.000 ; 
                RECT 2.880 284.040 99.400 284.360 ; 
                RECT 798.120 284.040 802.840 284.360 ; 
                RECT 2.880 285.400 77.640 285.720 ; 
                RECT 89.560 285.400 99.400 285.720 ; 
                RECT 798.120 285.400 802.840 285.720 ; 
                RECT 2.880 286.760 75.600 287.080 ; 
                RECT 89.560 286.760 99.400 287.080 ; 
                RECT 798.120 286.760 802.840 287.080 ; 
                RECT 2.880 288.120 75.600 288.440 ; 
                RECT 89.560 288.120 99.400 288.440 ; 
                RECT 798.120 288.120 802.840 288.440 ; 
                RECT 2.880 289.480 75.600 289.800 ; 
                RECT 89.560 289.480 99.400 289.800 ; 
                RECT 798.120 289.480 802.840 289.800 ; 
                RECT 2.880 290.840 75.600 291.160 ; 
                RECT 89.560 290.840 99.400 291.160 ; 
                RECT 798.120 290.840 802.840 291.160 ; 
                RECT 2.880 292.200 99.400 292.520 ; 
                RECT 798.120 292.200 802.840 292.520 ; 
                RECT 2.880 293.560 75.600 293.880 ; 
                RECT 89.560 293.560 99.400 293.880 ; 
                RECT 798.120 293.560 802.840 293.880 ; 
                RECT 2.880 294.920 75.600 295.240 ; 
                RECT 89.560 294.920 99.400 295.240 ; 
                RECT 798.120 294.920 802.840 295.240 ; 
                RECT 2.880 296.280 77.640 296.600 ; 
                RECT 89.560 296.280 99.400 296.600 ; 
                RECT 798.120 296.280 802.840 296.600 ; 
                RECT 2.880 297.640 75.600 297.960 ; 
                RECT 89.560 297.640 99.400 297.960 ; 
                RECT 798.120 297.640 802.840 297.960 ; 
                RECT 2.880 299.000 75.600 299.320 ; 
                RECT 80.720 299.000 99.400 299.320 ; 
                RECT 798.120 299.000 802.840 299.320 ; 
                RECT 2.880 300.360 85.800 300.680 ; 
                RECT 89.560 300.360 99.400 300.680 ; 
                RECT 798.120 300.360 802.840 300.680 ; 
                RECT 2.880 301.720 75.600 302.040 ; 
                RECT 89.560 301.720 99.400 302.040 ; 
                RECT 798.120 301.720 802.840 302.040 ; 
                RECT 2.880 303.080 75.600 303.400 ; 
                RECT 89.560 303.080 99.400 303.400 ; 
                RECT 798.120 303.080 802.840 303.400 ; 
                RECT 2.880 304.440 75.600 304.760 ; 
                RECT 89.560 304.440 99.400 304.760 ; 
                RECT 798.120 304.440 802.840 304.760 ; 
                RECT 2.880 305.800 75.600 306.120 ; 
                RECT 89.560 305.800 99.400 306.120 ; 
                RECT 798.120 305.800 802.840 306.120 ; 
                RECT 2.880 307.160 75.600 307.480 ; 
                RECT 80.720 307.160 99.400 307.480 ; 
                RECT 798.120 307.160 802.840 307.480 ; 
                RECT 2.880 308.520 80.360 308.840 ; 
                RECT 89.560 308.520 99.400 308.840 ; 
                RECT 798.120 308.520 802.840 308.840 ; 
                RECT 2.880 309.880 75.600 310.200 ; 
                RECT 89.560 309.880 99.400 310.200 ; 
                RECT 798.120 309.880 802.840 310.200 ; 
                RECT 2.880 311.240 75.600 311.560 ; 
                RECT 89.560 311.240 99.400 311.560 ; 
                RECT 798.120 311.240 802.840 311.560 ; 
                RECT 2.880 312.600 75.600 312.920 ; 
                RECT 89.560 312.600 99.400 312.920 ; 
                RECT 798.120 312.600 802.840 312.920 ; 
                RECT 2.880 313.960 75.600 314.280 ; 
                RECT 89.560 313.960 99.400 314.280 ; 
                RECT 798.120 313.960 802.840 314.280 ; 
                RECT 2.880 315.320 99.400 315.640 ; 
                RECT 798.120 315.320 802.840 315.640 ; 
                RECT 2.880 316.680 78.320 317.000 ; 
                RECT 89.560 316.680 99.400 317.000 ; 
                RECT 798.120 316.680 802.840 317.000 ; 
                RECT 2.880 318.040 82.400 318.360 ; 
                RECT 89.560 318.040 99.400 318.360 ; 
                RECT 798.120 318.040 802.840 318.360 ; 
                RECT 2.880 319.400 83.080 319.720 ; 
                RECT 89.560 319.400 99.400 319.720 ; 
                RECT 798.120 319.400 802.840 319.720 ; 
                RECT 2.880 320.760 78.320 321.080 ; 
                RECT 89.560 320.760 99.400 321.080 ; 
                RECT 798.120 320.760 802.840 321.080 ; 
                RECT 2.880 322.120 78.320 322.440 ; 
                RECT 89.560 322.120 99.400 322.440 ; 
                RECT 798.120 322.120 802.840 322.440 ; 
                RECT 2.880 323.480 99.400 323.800 ; 
                RECT 798.120 323.480 802.840 323.800 ; 
                RECT 2.880 324.840 78.320 325.160 ; 
                RECT 89.560 324.840 99.400 325.160 ; 
                RECT 798.120 324.840 802.840 325.160 ; 
                RECT 2.880 326.200 78.320 326.520 ; 
                RECT 89.560 326.200 99.400 326.520 ; 
                RECT 798.120 326.200 802.840 326.520 ; 
                RECT 2.880 327.560 78.320 327.880 ; 
                RECT 89.560 327.560 99.400 327.880 ; 
                RECT 798.120 327.560 802.840 327.880 ; 
                RECT 2.880 328.920 85.800 329.240 ; 
                RECT 89.560 328.920 99.400 329.240 ; 
                RECT 798.120 328.920 802.840 329.240 ; 
                RECT 2.880 330.280 78.320 330.600 ; 
                RECT 89.560 330.280 99.400 330.600 ; 
                RECT 798.120 330.280 802.840 330.600 ; 
                RECT 2.880 331.640 99.400 331.960 ; 
                RECT 798.120 331.640 802.840 331.960 ; 
                RECT 2.880 333.000 78.320 333.320 ; 
                RECT 89.560 333.000 99.400 333.320 ; 
                RECT 798.120 333.000 802.840 333.320 ; 
                RECT 2.880 334.360 78.320 334.680 ; 
                RECT 89.560 334.360 99.400 334.680 ; 
                RECT 798.120 334.360 802.840 334.680 ; 
                RECT 2.880 335.720 78.320 336.040 ; 
                RECT 89.560 335.720 99.400 336.040 ; 
                RECT 798.120 335.720 802.840 336.040 ; 
                RECT 2.880 337.080 78.320 337.400 ; 
                RECT 89.560 337.080 99.400 337.400 ; 
                RECT 798.120 337.080 802.840 337.400 ; 
                RECT 2.880 338.440 99.400 338.760 ; 
                RECT 798.120 338.440 802.840 338.760 ; 
                RECT 2.880 339.800 80.360 340.120 ; 
                RECT 89.560 339.800 99.400 340.120 ; 
                RECT 798.120 339.800 802.840 340.120 ; 
                RECT 2.880 341.160 79.000 341.480 ; 
                RECT 89.560 341.160 99.400 341.480 ; 
                RECT 798.120 341.160 802.840 341.480 ; 
                RECT 2.880 342.520 79.000 342.840 ; 
                RECT 89.560 342.520 99.400 342.840 ; 
                RECT 798.120 342.520 802.840 342.840 ; 
                RECT 2.880 343.880 79.000 344.200 ; 
                RECT 89.560 343.880 99.400 344.200 ; 
                RECT 798.120 343.880 802.840 344.200 ; 
                RECT 2.880 345.240 79.000 345.560 ; 
                RECT 89.560 345.240 99.400 345.560 ; 
                RECT 798.120 345.240 802.840 345.560 ; 
                RECT 2.880 346.600 99.400 346.920 ; 
                RECT 798.120 346.600 802.840 346.920 ; 
                RECT 2.880 347.960 82.400 348.280 ; 
                RECT 89.560 347.960 99.400 348.280 ; 
                RECT 798.120 347.960 802.840 348.280 ; 
                RECT 2.880 349.320 79.000 349.640 ; 
                RECT 89.560 349.320 99.400 349.640 ; 
                RECT 798.120 349.320 802.840 349.640 ; 
                RECT 2.880 350.680 79.000 351.000 ; 
                RECT 89.560 350.680 99.400 351.000 ; 
                RECT 798.120 350.680 802.840 351.000 ; 
                RECT 2.880 352.040 79.000 352.360 ; 
                RECT 89.560 352.040 99.400 352.360 ; 
                RECT 798.120 352.040 802.840 352.360 ; 
                RECT 2.880 353.400 79.000 353.720 ; 
                RECT 89.560 353.400 99.400 353.720 ; 
                RECT 798.120 353.400 802.840 353.720 ; 
                RECT 2.880 354.760 99.400 355.080 ; 
                RECT 798.120 354.760 802.840 355.080 ; 
                RECT 2.880 356.120 79.000 356.440 ; 
                RECT 89.560 356.120 99.400 356.440 ; 
                RECT 798.120 356.120 802.840 356.440 ; 
                RECT 2.880 357.480 84.440 357.800 ; 
                RECT 89.560 357.480 99.400 357.800 ; 
                RECT 798.120 357.480 802.840 357.800 ; 
                RECT 2.880 358.840 79.000 359.160 ; 
                RECT 89.560 358.840 99.400 359.160 ; 
                RECT 798.120 358.840 802.840 359.160 ; 
                RECT 2.880 360.200 79.000 360.520 ; 
                RECT 89.560 360.200 99.400 360.520 ; 
                RECT 798.120 360.200 802.840 360.520 ; 
                RECT 2.880 361.560 79.000 361.880 ; 
                RECT 89.560 361.560 99.400 361.880 ; 
                RECT 798.120 361.560 802.840 361.880 ; 
                RECT 2.880 362.920 99.400 363.240 ; 
                RECT 798.120 362.920 802.840 363.240 ; 
                RECT 2.880 364.280 79.000 364.600 ; 
                RECT 89.560 364.280 99.400 364.600 ; 
                RECT 798.120 364.280 802.840 364.600 ; 
                RECT 2.880 365.640 79.000 365.960 ; 
                RECT 89.560 365.640 99.400 365.960 ; 
                RECT 798.120 365.640 802.840 365.960 ; 
                RECT 2.880 367.000 87.160 367.320 ; 
                RECT 89.560 367.000 99.400 367.320 ; 
                RECT 798.120 367.000 802.840 367.320 ; 
                RECT 2.880 368.360 87.160 368.680 ; 
                RECT 89.560 368.360 99.400 368.680 ; 
                RECT 798.120 368.360 802.840 368.680 ; 
                RECT 2.880 369.720 79.000 370.040 ; 
                RECT 89.560 369.720 99.400 370.040 ; 
                RECT 798.120 369.720 802.840 370.040 ; 
                RECT 2.880 371.080 99.400 371.400 ; 
                RECT 798.120 371.080 802.840 371.400 ; 
                RECT 2.880 372.440 79.000 372.760 ; 
                RECT 89.560 372.440 99.400 372.760 ; 
                RECT 798.120 372.440 802.840 372.760 ; 
                RECT 2.880 373.800 79.000 374.120 ; 
                RECT 89.560 373.800 99.400 374.120 ; 
                RECT 798.120 373.800 802.840 374.120 ; 
                RECT 2.880 375.160 79.000 375.480 ; 
                RECT 89.560 375.160 99.400 375.480 ; 
                RECT 798.120 375.160 802.840 375.480 ; 
                RECT 2.880 376.520 81.720 376.840 ; 
                RECT 89.560 376.520 99.400 376.840 ; 
                RECT 798.120 376.520 802.840 376.840 ; 
                RECT 2.880 377.880 99.400 378.200 ; 
                RECT 798.120 377.880 802.840 378.200 ; 
                RECT 2.880 379.240 82.400 379.560 ; 
                RECT 89.560 379.240 99.400 379.560 ; 
                RECT 798.120 379.240 802.840 379.560 ; 
                RECT 2.880 380.600 79.000 380.920 ; 
                RECT 89.560 380.600 99.400 380.920 ; 
                RECT 798.120 380.600 802.840 380.920 ; 
                RECT 2.880 381.960 79.000 382.280 ; 
                RECT 89.560 381.960 99.400 382.280 ; 
                RECT 798.120 381.960 802.840 382.280 ; 
                RECT 2.880 383.320 79.000 383.640 ; 
                RECT 89.560 383.320 99.400 383.640 ; 
                RECT 798.120 383.320 802.840 383.640 ; 
                RECT 2.880 384.680 79.000 385.000 ; 
                RECT 89.560 384.680 99.400 385.000 ; 
                RECT 798.120 384.680 802.840 385.000 ; 
                RECT 2.880 386.040 99.400 386.360 ; 
                RECT 798.120 386.040 802.840 386.360 ; 
                RECT 2.880 387.400 83.760 387.720 ; 
                RECT 89.560 387.400 99.400 387.720 ; 
                RECT 798.120 387.400 802.840 387.720 ; 
                RECT 2.880 388.760 79.000 389.080 ; 
                RECT 89.560 388.760 99.400 389.080 ; 
                RECT 798.120 388.760 802.840 389.080 ; 
                RECT 2.880 390.120 79.000 390.440 ; 
                RECT 89.560 390.120 99.400 390.440 ; 
                RECT 798.120 390.120 802.840 390.440 ; 
                RECT 2.880 391.480 79.000 391.800 ; 
                RECT 89.560 391.480 99.400 391.800 ; 
                RECT 798.120 391.480 802.840 391.800 ; 
                RECT 2.880 392.840 79.000 393.160 ; 
                RECT 89.560 392.840 99.400 393.160 ; 
                RECT 798.120 392.840 802.840 393.160 ; 
                RECT 2.880 394.200 99.400 394.520 ; 
                RECT 798.120 394.200 802.840 394.520 ; 
                RECT 2.880 395.560 79.000 395.880 ; 
                RECT 89.560 395.560 99.400 395.880 ; 
                RECT 798.120 395.560 802.840 395.880 ; 
                RECT 2.880 396.920 86.480 397.240 ; 
                RECT 89.560 396.920 99.400 397.240 ; 
                RECT 798.120 396.920 802.840 397.240 ; 
                RECT 2.880 398.280 79.000 398.600 ; 
                RECT 89.560 398.280 99.400 398.600 ; 
                RECT 798.120 398.280 802.840 398.600 ; 
                RECT 2.880 399.640 79.000 399.960 ; 
                RECT 89.560 399.640 99.400 399.960 ; 
                RECT 798.120 399.640 802.840 399.960 ; 
                RECT 2.880 401.000 79.000 401.320 ; 
                RECT 89.560 401.000 99.400 401.320 ; 
                RECT 798.120 401.000 802.840 401.320 ; 
                RECT 2.880 402.360 99.400 402.680 ; 
                RECT 798.120 402.360 802.840 402.680 ; 
                RECT 2.880 403.720 79.680 404.040 ; 
                RECT 89.560 403.720 99.400 404.040 ; 
                RECT 798.120 403.720 802.840 404.040 ; 
                RECT 2.880 405.080 79.680 405.400 ; 
                RECT 89.560 405.080 99.400 405.400 ; 
                RECT 798.120 405.080 802.840 405.400 ; 
                RECT 2.880 406.440 81.040 406.760 ; 
                RECT 89.560 406.440 99.400 406.760 ; 
                RECT 798.120 406.440 802.840 406.760 ; 
                RECT 2.880 407.800 79.680 408.120 ; 
                RECT 89.560 407.800 99.400 408.120 ; 
                RECT 798.120 407.800 802.840 408.120 ; 
                RECT 2.880 409.160 79.680 409.480 ; 
                RECT 89.560 409.160 99.400 409.480 ; 
                RECT 798.120 409.160 802.840 409.480 ; 
                RECT 2.880 410.520 99.400 410.840 ; 
                RECT 798.120 410.520 802.840 410.840 ; 
                RECT 2.880 411.880 79.680 412.200 ; 
                RECT 89.560 411.880 99.400 412.200 ; 
                RECT 798.120 411.880 802.840 412.200 ; 
                RECT 2.880 413.240 79.680 413.560 ; 
                RECT 89.560 413.240 99.400 413.560 ; 
                RECT 798.120 413.240 802.840 413.560 ; 
                RECT 2.880 414.600 79.680 414.920 ; 
                RECT 89.560 414.600 99.400 414.920 ; 
                RECT 798.120 414.600 802.840 414.920 ; 
                RECT 2.880 415.960 83.760 416.280 ; 
                RECT 89.560 415.960 99.400 416.280 ; 
                RECT 798.120 415.960 802.840 416.280 ; 
                RECT 2.880 417.320 79.680 417.640 ; 
                RECT 89.560 417.320 99.400 417.640 ; 
                RECT 798.120 417.320 802.840 417.640 ; 
                RECT 2.880 418.680 99.400 419.000 ; 
                RECT 798.120 418.680 802.840 419.000 ; 
                RECT 2.880 420.040 79.680 420.360 ; 
                RECT 89.560 420.040 99.400 420.360 ; 
                RECT 798.120 420.040 802.840 420.360 ; 
                RECT 2.880 421.400 79.680 421.720 ; 
                RECT 89.560 421.400 99.400 421.720 ; 
                RECT 798.120 421.400 802.840 421.720 ; 
                RECT 2.880 422.760 79.680 423.080 ; 
                RECT 89.560 422.760 99.400 423.080 ; 
                RECT 798.120 422.760 802.840 423.080 ; 
                RECT 2.880 424.120 79.680 424.440 ; 
                RECT 89.560 424.120 99.400 424.440 ; 
                RECT 798.120 424.120 802.840 424.440 ; 
                RECT 2.880 425.480 99.400 425.800 ; 
                RECT 798.120 425.480 802.840 425.800 ; 
                RECT 2.880 426.840 85.800 427.160 ; 
                RECT 89.560 426.840 99.400 427.160 ; 
                RECT 798.120 426.840 802.840 427.160 ; 
                RECT 2.880 428.200 79.680 428.520 ; 
                RECT 89.560 428.200 99.400 428.520 ; 
                RECT 798.120 428.200 802.840 428.520 ; 
                RECT 2.880 429.560 79.680 429.880 ; 
                RECT 89.560 429.560 99.400 429.880 ; 
                RECT 798.120 429.560 802.840 429.880 ; 
                RECT 2.880 430.920 79.680 431.240 ; 
                RECT 89.560 430.920 99.400 431.240 ; 
                RECT 798.120 430.920 802.840 431.240 ; 
                RECT 2.880 432.280 79.680 432.600 ; 
                RECT 89.560 432.280 99.400 432.600 ; 
                RECT 798.120 432.280 802.840 432.600 ; 
                RECT 2.880 433.640 99.400 433.960 ; 
                RECT 798.120 433.640 802.840 433.960 ; 
                RECT 2.880 435.000 99.400 435.320 ; 
                RECT 798.120 435.000 802.840 435.320 ; 
                RECT 2.880 436.360 388.400 436.680 ; 
                RECT 798.120 436.360 802.840 436.680 ; 
                RECT 2.880 437.720 388.400 438.040 ; 
                RECT 798.120 437.720 802.840 438.040 ; 
                RECT 2.880 439.080 802.840 439.400 ; 
                RECT 2.880 440.440 802.840 440.760 ; 
                RECT 2.880 441.800 802.840 442.120 ; 
                RECT 2.880 443.160 802.840 443.480 ; 
                RECT 2.880 444.520 802.840 444.840 ; 
                RECT 2.880 2.880 802.840 4.240 ; 
                RECT 2.880 445.840 802.840 447.200 ; 
                RECT 392.540 29.575 398.340 30.695 ; 
                RECT 788.440 29.575 794.240 30.695 ; 
                RECT 392.540 35.365 398.340 35.985 ; 
                RECT 788.440 35.365 794.240 35.985 ; 
                RECT 392.540 40.390 398.340 41.030 ; 
                RECT 788.440 40.390 794.240 41.030 ; 
                RECT 392.540 45.520 398.340 46.170 ; 
                RECT 788.440 45.520 794.240 46.170 ; 
                RECT 392.540 50.735 398.340 51.345 ; 
                RECT 788.440 50.735 794.240 51.345 ; 
                RECT 392.540 55.665 398.340 56.275 ; 
                RECT 788.440 55.665 794.240 56.275 ; 
                RECT 392.540 86.350 794.240 87.150 ; 
                RECT 392.540 69.400 794.240 71.200 ; 
                RECT 392.540 90.035 794.240 93.635 ; 
                RECT 392.540 83.140 794.240 83.940 ; 
                RECT 392.540 78.450 794.240 79.250 ; 
                RECT 392.540 115.495 794.240 115.785 ; 
                RECT 392.540 81.460 794.240 82.260 ; 
                RECT 392.540 142.705 794.240 144.505 ; 
                RECT 392.540 20.205 794.240 22.005 ; 
                RECT 99.995 180.395 101.105 434.775 ; 
                RECT 108.930 180.395 110.850 434.775 ; 
                RECT 124.290 180.395 126.210 434.775 ; 
                RECT 146.560 180.395 148.480 434.775 ; 
                RECT 150.400 180.395 152.320 434.775 ; 
                RECT 154.240 180.395 156.160 434.775 ; 
                RECT 188.395 180.395 190.315 434.775 ; 
                RECT 192.235 180.395 194.155 434.775 ; 
                RECT 196.075 180.395 197.995 434.775 ; 
                RECT 199.915 180.395 201.835 434.775 ; 
                RECT 203.755 180.395 205.675 434.775 ; 
                RECT 261.435 180.395 263.355 434.775 ; 
                RECT 265.275 180.395 267.195 434.775 ; 
                RECT 269.115 180.395 271.035 434.775 ; 
                RECT 272.955 180.395 274.875 434.775 ; 
                RECT 276.795 180.395 278.715 434.775 ; 
                RECT 280.635 180.395 282.555 434.775 ; 
                RECT 284.475 180.395 286.395 434.775 ; 
                RECT 288.315 180.395 290.235 434.775 ; 
                RECT 292.155 180.395 294.075 434.775 ; 
                RECT 287.415 61.335 288.525 113.935 ; 
                RECT 294.930 61.335 295.820 113.935 ; 
                RECT 301.795 61.335 302.905 113.935 ; 
                RECT 311.375 61.335 313.295 113.935 ; 
                RECT 330.205 61.335 332.125 113.935 ; 
                RECT 334.045 61.335 335.965 113.935 ; 
                RECT 337.885 61.335 339.805 113.935 ; 
                RECT 311.905 140.900 313.015 173.760 ; 
                RECT 320.280 140.900 321.170 173.760 ; 
                RECT 327.040 140.900 327.930 173.760 ; 
                RECT 333.690 140.900 335.230 173.760 ; 
                RECT 345.865 140.900 347.785 173.760 ; 
                RECT 349.705 140.900 351.625 173.760 ; 
                RECT 321.020 128.160 321.910 134.900 ; 
                RECT 327.670 128.160 329.210 134.900 ; 
                RECT 340.705 128.160 342.625 134.900 ; 
                RECT 344.545 128.160 346.465 134.900 ; 
                RECT 368.940 50.175 369.830 55.335 ; 
                RECT 26.230 181.460 35.390 181.830 ; 
                RECT 26.230 184.795 35.390 185.685 ; 
                RECT 211.480 166.870 228.720 167.540 ; 
                RECT 211.480 168.200 228.720 169.550 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 805.720 450.080 ; 
        LAYER met2 ;
            RECT 0.000 0.000 805.720 450.080 ; 
    END 
END sram22_512x64m4w8 
END LIBRARY 

