VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram22_64x4m4w2
  CLASS BLOCK ;
  ORIGIN 61.96 159.085 ;
  FOREIGN sram22_64x4m4w2 -61.96 -159.085 ;
  SIZE 104.105 BY 205.29 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 20.96 -94.075 21.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 44.8 21.925 45.93 ;
        RECT 21.595 39.955 21.925 40.285 ;
        RECT 21.595 38.595 21.925 38.925 ;
        RECT 21.6 37.92 21.92 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 -96.045 21.925 -95.715 ;
        RECT 21.595 -97.405 21.925 -97.075 ;
        RECT 21.595 -98.765 21.925 -98.435 ;
        RECT 21.595 -100.125 21.925 -99.795 ;
        RECT 21.595 -101.485 21.925 -101.155 ;
        RECT 21.595 -102.845 21.925 -102.515 ;
        RECT 21.595 -104.205 21.925 -103.875 ;
        RECT 21.595 -105.565 21.925 -105.235 ;
        RECT 21.595 -106.925 21.925 -106.595 ;
        RECT 21.595 -108.285 21.925 -107.955 ;
        RECT 21.595 -109.645 21.925 -109.315 ;
        RECT 21.595 -111.005 21.925 -110.675 ;
        RECT 21.595 -112.365 21.925 -112.035 ;
        RECT 21.595 -113.725 21.925 -113.395 ;
        RECT 21.595 -115.085 21.925 -114.755 ;
        RECT 21.595 -116.445 21.925 -116.115 ;
        RECT 21.595 -117.805 21.925 -117.475 ;
        RECT 21.595 -119.165 21.925 -118.835 ;
        RECT 21.595 -120.525 21.925 -120.195 ;
        RECT 21.595 -121.885 21.925 -121.555 ;
        RECT 21.595 -123.245 21.925 -122.915 ;
        RECT 21.595 -124.605 21.925 -124.275 ;
        RECT 21.595 -125.965 21.925 -125.635 ;
        RECT 21.595 -127.325 21.925 -126.995 ;
        RECT 21.595 -128.685 21.925 -128.355 ;
        RECT 21.595 -130.045 21.925 -129.715 ;
        RECT 21.595 -131.405 21.925 -131.075 ;
        RECT 21.595 -132.765 21.925 -132.435 ;
        RECT 21.595 -134.125 21.925 -133.795 ;
        RECT 21.595 -135.485 21.925 -135.155 ;
        RECT 21.595 -136.845 21.925 -136.515 ;
        RECT 21.595 -138.205 21.925 -137.875 ;
        RECT 21.595 -139.565 21.925 -139.235 ;
        RECT 21.595 -140.925 21.925 -140.595 ;
        RECT 21.595 -142.285 21.925 -141.955 ;
        RECT 21.595 -143.645 21.925 -143.315 ;
        RECT 21.595 -145.005 21.925 -144.675 ;
        RECT 21.595 -146.365 21.925 -146.035 ;
        RECT 21.595 -147.725 21.925 -147.395 ;
        RECT 21.595 -149.085 21.925 -148.755 ;
        RECT 21.595 -150.445 21.925 -150.115 ;
        RECT 21.595 -151.805 21.925 -151.475 ;
        RECT 21.595 -153.165 21.925 -152.835 ;
        RECT 21.595 -158.81 21.925 -157.68 ;
        RECT 21.6 -158.925 21.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 44.8 23.285 45.93 ;
        RECT 22.955 39.955 23.285 40.285 ;
        RECT 22.955 38.595 23.285 38.925 ;
        RECT 22.96 37.92 23.28 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 -0.845 23.285 -0.515 ;
        RECT 22.955 -2.205 23.285 -1.875 ;
        RECT 22.955 -3.565 23.285 -3.235 ;
        RECT 22.96 -3.565 23.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 44.8 24.645 45.93 ;
        RECT 24.315 39.955 24.645 40.285 ;
        RECT 24.315 38.595 24.645 38.925 ;
        RECT 24.32 37.92 24.64 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 -0.845 24.645 -0.515 ;
        RECT 24.315 -2.205 24.645 -1.875 ;
        RECT 24.315 -3.565 24.645 -3.235 ;
        RECT 24.32 -3.565 24.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 44.8 26.005 45.93 ;
        RECT 25.675 39.955 26.005 40.285 ;
        RECT 25.675 38.595 26.005 38.925 ;
        RECT 25.68 37.92 26 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 -0.845 26.005 -0.515 ;
        RECT 25.675 -2.205 26.005 -1.875 ;
        RECT 25.675 -3.565 26.005 -3.235 ;
        RECT 25.68 -3.565 26 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 -91.965 26.005 -91.635 ;
        RECT 25.675 -93.325 26.005 -92.995 ;
        RECT 25.675 -94.685 26.005 -94.355 ;
        RECT 25.675 -96.045 26.005 -95.715 ;
        RECT 25.675 -97.405 26.005 -97.075 ;
        RECT 25.675 -98.765 26.005 -98.435 ;
        RECT 25.675 -100.125 26.005 -99.795 ;
        RECT 25.675 -101.485 26.005 -101.155 ;
        RECT 25.675 -102.845 26.005 -102.515 ;
        RECT 25.675 -104.205 26.005 -103.875 ;
        RECT 25.675 -105.565 26.005 -105.235 ;
        RECT 25.675 -106.925 26.005 -106.595 ;
        RECT 25.675 -108.285 26.005 -107.955 ;
        RECT 25.675 -109.645 26.005 -109.315 ;
        RECT 25.675 -111.005 26.005 -110.675 ;
        RECT 25.675 -112.365 26.005 -112.035 ;
        RECT 25.675 -113.725 26.005 -113.395 ;
        RECT 25.675 -115.085 26.005 -114.755 ;
        RECT 25.675 -116.445 26.005 -116.115 ;
        RECT 25.675 -117.805 26.005 -117.475 ;
        RECT 25.675 -119.165 26.005 -118.835 ;
        RECT 25.675 -120.525 26.005 -120.195 ;
        RECT 25.675 -121.885 26.005 -121.555 ;
        RECT 25.675 -123.245 26.005 -122.915 ;
        RECT 25.675 -124.605 26.005 -124.275 ;
        RECT 25.675 -125.965 26.005 -125.635 ;
        RECT 25.675 -127.325 26.005 -126.995 ;
        RECT 25.675 -128.685 26.005 -128.355 ;
        RECT 25.675 -130.045 26.005 -129.715 ;
        RECT 25.675 -131.405 26.005 -131.075 ;
        RECT 25.675 -132.765 26.005 -132.435 ;
        RECT 25.675 -134.125 26.005 -133.795 ;
        RECT 25.675 -135.485 26.005 -135.155 ;
        RECT 25.675 -136.845 26.005 -136.515 ;
        RECT 25.675 -138.205 26.005 -137.875 ;
        RECT 25.675 -139.565 26.005 -139.235 ;
        RECT 25.675 -140.925 26.005 -140.595 ;
        RECT 25.675 -142.285 26.005 -141.955 ;
        RECT 25.675 -143.645 26.005 -143.315 ;
        RECT 25.675 -145.005 26.005 -144.675 ;
        RECT 25.675 -146.365 26.005 -146.035 ;
        RECT 25.675 -147.725 26.005 -147.395 ;
        RECT 25.675 -149.085 26.005 -148.755 ;
        RECT 25.675 -150.445 26.005 -150.115 ;
        RECT 25.675 -151.805 26.005 -151.475 ;
        RECT 25.675 -153.165 26.005 -152.835 ;
        RECT 25.675 -158.81 26.005 -157.68 ;
        RECT 25.68 -158.925 26 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 44.8 27.365 45.93 ;
        RECT 27.035 39.955 27.365 40.285 ;
        RECT 27.035 38.595 27.365 38.925 ;
        RECT 27.04 37.92 27.36 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 -96.045 27.365 -95.715 ;
        RECT 27.035 -97.405 27.365 -97.075 ;
        RECT 27.035 -98.765 27.365 -98.435 ;
        RECT 27.035 -100.125 27.365 -99.795 ;
        RECT 27.035 -101.485 27.365 -101.155 ;
        RECT 27.035 -102.845 27.365 -102.515 ;
        RECT 27.035 -104.205 27.365 -103.875 ;
        RECT 27.035 -105.565 27.365 -105.235 ;
        RECT 27.035 -106.925 27.365 -106.595 ;
        RECT 27.035 -108.285 27.365 -107.955 ;
        RECT 27.035 -109.645 27.365 -109.315 ;
        RECT 27.035 -111.005 27.365 -110.675 ;
        RECT 27.035 -112.365 27.365 -112.035 ;
        RECT 27.035 -113.725 27.365 -113.395 ;
        RECT 27.035 -115.085 27.365 -114.755 ;
        RECT 27.035 -116.445 27.365 -116.115 ;
        RECT 27.035 -117.805 27.365 -117.475 ;
        RECT 27.035 -119.165 27.365 -118.835 ;
        RECT 27.035 -120.525 27.365 -120.195 ;
        RECT 27.035 -121.885 27.365 -121.555 ;
        RECT 27.035 -123.245 27.365 -122.915 ;
        RECT 27.035 -124.605 27.365 -124.275 ;
        RECT 27.035 -125.965 27.365 -125.635 ;
        RECT 27.035 -127.325 27.365 -126.995 ;
        RECT 27.035 -128.685 27.365 -128.355 ;
        RECT 27.035 -130.045 27.365 -129.715 ;
        RECT 27.035 -131.405 27.365 -131.075 ;
        RECT 27.035 -132.765 27.365 -132.435 ;
        RECT 27.035 -134.125 27.365 -133.795 ;
        RECT 27.035 -135.485 27.365 -135.155 ;
        RECT 27.035 -136.845 27.365 -136.515 ;
        RECT 27.035 -138.205 27.365 -137.875 ;
        RECT 27.035 -139.565 27.365 -139.235 ;
        RECT 27.035 -140.925 27.365 -140.595 ;
        RECT 27.035 -142.285 27.365 -141.955 ;
        RECT 27.035 -143.645 27.365 -143.315 ;
        RECT 27.035 -145.005 27.365 -144.675 ;
        RECT 27.035 -146.365 27.365 -146.035 ;
        RECT 27.035 -147.725 27.365 -147.395 ;
        RECT 27.035 -149.085 27.365 -148.755 ;
        RECT 27.035 -150.445 27.365 -150.115 ;
        RECT 27.035 -151.805 27.365 -151.475 ;
        RECT 27.035 -153.165 27.365 -152.835 ;
        RECT 27.035 -158.81 27.365 -157.68 ;
        RECT 27.04 -158.925 27.36 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.71 -94.075 28.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 44.8 28.725 45.93 ;
        RECT 28.395 39.955 28.725 40.285 ;
        RECT 28.395 38.595 28.725 38.925 ;
        RECT 28.4 37.92 28.72 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 -0.845 28.725 -0.515 ;
        RECT 28.395 -2.205 28.725 -1.875 ;
        RECT 28.395 -3.565 28.725 -3.235 ;
        RECT 28.4 -3.565 28.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 -91.965 28.725 -91.635 ;
        RECT 28.395 -93.325 28.725 -92.995 ;
        RECT 28.395 -94.685 28.725 -94.355 ;
        RECT 28.395 -96.045 28.725 -95.715 ;
        RECT 28.395 -97.405 28.725 -97.075 ;
        RECT 28.395 -98.765 28.725 -98.435 ;
        RECT 28.395 -100.125 28.725 -99.795 ;
        RECT 28.395 -101.485 28.725 -101.155 ;
        RECT 28.395 -102.845 28.725 -102.515 ;
        RECT 28.395 -104.205 28.725 -103.875 ;
        RECT 28.395 -105.565 28.725 -105.235 ;
        RECT 28.395 -106.925 28.725 -106.595 ;
        RECT 28.395 -108.285 28.725 -107.955 ;
        RECT 28.395 -109.645 28.725 -109.315 ;
        RECT 28.395 -111.005 28.725 -110.675 ;
        RECT 28.395 -112.365 28.725 -112.035 ;
        RECT 28.395 -113.725 28.725 -113.395 ;
        RECT 28.395 -115.085 28.725 -114.755 ;
        RECT 28.395 -116.445 28.725 -116.115 ;
        RECT 28.395 -117.805 28.725 -117.475 ;
        RECT 28.395 -119.165 28.725 -118.835 ;
        RECT 28.395 -120.525 28.725 -120.195 ;
        RECT 28.395 -121.885 28.725 -121.555 ;
        RECT 28.395 -123.245 28.725 -122.915 ;
        RECT 28.395 -124.605 28.725 -124.275 ;
        RECT 28.395 -125.965 28.725 -125.635 ;
        RECT 28.395 -127.325 28.725 -126.995 ;
        RECT 28.395 -128.685 28.725 -128.355 ;
        RECT 28.395 -130.045 28.725 -129.715 ;
        RECT 28.395 -131.405 28.725 -131.075 ;
        RECT 28.395 -132.765 28.725 -132.435 ;
        RECT 28.395 -134.125 28.725 -133.795 ;
        RECT 28.395 -135.485 28.725 -135.155 ;
        RECT 28.395 -136.845 28.725 -136.515 ;
        RECT 28.395 -138.205 28.725 -137.875 ;
        RECT 28.395 -139.565 28.725 -139.235 ;
        RECT 28.395 -140.925 28.725 -140.595 ;
        RECT 28.395 -142.285 28.725 -141.955 ;
        RECT 28.395 -143.645 28.725 -143.315 ;
        RECT 28.395 -145.005 28.725 -144.675 ;
        RECT 28.395 -146.365 28.725 -146.035 ;
        RECT 28.395 -147.725 28.725 -147.395 ;
        RECT 28.395 -149.085 28.725 -148.755 ;
        RECT 28.395 -150.445 28.725 -150.115 ;
        RECT 28.395 -151.805 28.725 -151.475 ;
        RECT 28.395 -153.165 28.725 -152.835 ;
        RECT 28.395 -158.81 28.725 -157.68 ;
        RECT 28.4 -158.925 28.72 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 44.8 30.085 45.93 ;
        RECT 29.755 39.955 30.085 40.285 ;
        RECT 29.755 38.595 30.085 38.925 ;
        RECT 29.76 37.92 30.08 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 -0.845 30.085 -0.515 ;
        RECT 29.755 -2.205 30.085 -1.875 ;
        RECT 29.755 -3.565 30.085 -3.235 ;
        RECT 29.76 -3.565 30.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 -91.965 30.085 -91.635 ;
        RECT 29.755 -93.325 30.085 -92.995 ;
        RECT 29.755 -94.685 30.085 -94.355 ;
        RECT 29.755 -96.045 30.085 -95.715 ;
        RECT 29.755 -97.405 30.085 -97.075 ;
        RECT 29.755 -98.765 30.085 -98.435 ;
        RECT 29.755 -100.125 30.085 -99.795 ;
        RECT 29.755 -101.485 30.085 -101.155 ;
        RECT 29.755 -102.845 30.085 -102.515 ;
        RECT 29.755 -104.205 30.085 -103.875 ;
        RECT 29.755 -105.565 30.085 -105.235 ;
        RECT 29.755 -106.925 30.085 -106.595 ;
        RECT 29.755 -108.285 30.085 -107.955 ;
        RECT 29.755 -109.645 30.085 -109.315 ;
        RECT 29.755 -111.005 30.085 -110.675 ;
        RECT 29.755 -112.365 30.085 -112.035 ;
        RECT 29.755 -113.725 30.085 -113.395 ;
        RECT 29.755 -115.085 30.085 -114.755 ;
        RECT 29.755 -116.445 30.085 -116.115 ;
        RECT 29.755 -117.805 30.085 -117.475 ;
        RECT 29.755 -119.165 30.085 -118.835 ;
        RECT 29.755 -120.525 30.085 -120.195 ;
        RECT 29.755 -121.885 30.085 -121.555 ;
        RECT 29.755 -123.245 30.085 -122.915 ;
        RECT 29.755 -124.605 30.085 -124.275 ;
        RECT 29.755 -125.965 30.085 -125.635 ;
        RECT 29.755 -127.325 30.085 -126.995 ;
        RECT 29.755 -128.685 30.085 -128.355 ;
        RECT 29.755 -130.045 30.085 -129.715 ;
        RECT 29.755 -131.405 30.085 -131.075 ;
        RECT 29.755 -132.765 30.085 -132.435 ;
        RECT 29.755 -134.125 30.085 -133.795 ;
        RECT 29.755 -135.485 30.085 -135.155 ;
        RECT 29.755 -136.845 30.085 -136.515 ;
        RECT 29.755 -138.205 30.085 -137.875 ;
        RECT 29.755 -139.565 30.085 -139.235 ;
        RECT 29.755 -140.925 30.085 -140.595 ;
        RECT 29.755 -142.285 30.085 -141.955 ;
        RECT 29.755 -143.645 30.085 -143.315 ;
        RECT 29.755 -145.005 30.085 -144.675 ;
        RECT 29.755 -146.365 30.085 -146.035 ;
        RECT 29.755 -147.725 30.085 -147.395 ;
        RECT 29.755 -149.085 30.085 -148.755 ;
        RECT 29.755 -150.445 30.085 -150.115 ;
        RECT 29.755 -151.805 30.085 -151.475 ;
        RECT 29.755 -153.165 30.085 -152.835 ;
        RECT 29.755 -158.81 30.085 -157.68 ;
        RECT 29.76 -158.925 30.08 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 44.8 31.445 45.93 ;
        RECT 31.115 39.955 31.445 40.285 ;
        RECT 31.115 38.595 31.445 38.925 ;
        RECT 31.115 36.09 31.445 36.42 ;
        RECT 31.115 33.915 31.445 34.245 ;
        RECT 31.115 32.335 31.445 32.665 ;
        RECT 31.115 31.485 31.445 31.815 ;
        RECT 31.115 29.175 31.445 29.505 ;
        RECT 31.115 28.325 31.445 28.655 ;
        RECT 31.115 26.015 31.445 26.345 ;
        RECT 31.115 25.165 31.445 25.495 ;
        RECT 31.115 22.855 31.445 23.185 ;
        RECT 31.115 22.005 31.445 22.335 ;
        RECT 31.115 19.695 31.445 20.025 ;
        RECT 31.115 18.115 31.445 18.445 ;
        RECT 31.115 17.265 31.445 17.595 ;
        RECT 31.115 14.955 31.445 15.285 ;
        RECT 31.115 14.105 31.445 14.435 ;
        RECT 31.115 11.795 31.445 12.125 ;
        RECT 31.115 10.945 31.445 11.275 ;
        RECT 31.115 8.635 31.445 8.965 ;
        RECT 31.115 7.785 31.445 8.115 ;
        RECT 31.115 5.475 31.445 5.805 ;
        RECT 31.115 3.895 31.445 4.225 ;
        RECT 31.115 3.045 31.445 3.375 ;
        RECT 31.115 0.87 31.445 1.2 ;
        RECT 31.115 -0.845 31.445 -0.515 ;
        RECT 31.115 -2.205 31.445 -1.875 ;
        RECT 31.115 -3.565 31.445 -3.235 ;
        RECT 31.115 -4.925 31.445 -4.595 ;
        RECT 31.115 -6.285 31.445 -5.955 ;
        RECT 31.115 -7.645 31.445 -7.315 ;
        RECT 31.115 -9.005 31.445 -8.675 ;
        RECT 31.115 -10.365 31.445 -10.035 ;
        RECT 31.115 -11.725 31.445 -11.395 ;
        RECT 31.115 -13.085 31.445 -12.755 ;
        RECT 31.115 -14.445 31.445 -14.115 ;
        RECT 31.115 -15.805 31.445 -15.475 ;
        RECT 31.115 -17.165 31.445 -16.835 ;
        RECT 31.115 -18.525 31.445 -18.195 ;
        RECT 31.115 -19.885 31.445 -19.555 ;
        RECT 31.115 -21.245 31.445 -20.915 ;
        RECT 31.115 -22.605 31.445 -22.275 ;
        RECT 31.115 -23.965 31.445 -23.635 ;
        RECT 31.115 -25.325 31.445 -24.995 ;
        RECT 31.115 -26.685 31.445 -26.355 ;
        RECT 31.115 -28.045 31.445 -27.715 ;
        RECT 31.115 -29.405 31.445 -29.075 ;
        RECT 31.115 -30.765 31.445 -30.435 ;
        RECT 31.115 -32.125 31.445 -31.795 ;
        RECT 31.115 -33.485 31.445 -33.155 ;
        RECT 31.115 -34.845 31.445 -34.515 ;
        RECT 31.115 -36.205 31.445 -35.875 ;
        RECT 31.115 -37.565 31.445 -37.235 ;
        RECT 31.115 -38.925 31.445 -38.595 ;
        RECT 31.115 -40.285 31.445 -39.955 ;
        RECT 31.115 -41.645 31.445 -41.315 ;
        RECT 31.115 -43.005 31.445 -42.675 ;
        RECT 31.115 -44.365 31.445 -44.035 ;
        RECT 31.115 -45.725 31.445 -45.395 ;
        RECT 31.115 -47.085 31.445 -46.755 ;
        RECT 31.115 -48.445 31.445 -48.115 ;
        RECT 31.115 -49.805 31.445 -49.475 ;
        RECT 31.115 -51.165 31.445 -50.835 ;
        RECT 31.115 -52.525 31.445 -52.195 ;
        RECT 31.115 -53.885 31.445 -53.555 ;
        RECT 31.115 -55.245 31.445 -54.915 ;
        RECT 31.115 -56.605 31.445 -56.275 ;
        RECT 31.115 -57.965 31.445 -57.635 ;
        RECT 31.115 -59.325 31.445 -58.995 ;
        RECT 31.115 -60.685 31.445 -60.355 ;
        RECT 31.115 -62.045 31.445 -61.715 ;
        RECT 31.115 -63.405 31.445 -63.075 ;
        RECT 31.115 -64.765 31.445 -64.435 ;
        RECT 31.115 -66.125 31.445 -65.795 ;
        RECT 31.115 -67.485 31.445 -67.155 ;
        RECT 31.115 -68.845 31.445 -68.515 ;
        RECT 31.115 -70.205 31.445 -69.875 ;
        RECT 31.115 -71.565 31.445 -71.235 ;
        RECT 31.115 -72.925 31.445 -72.595 ;
        RECT 31.115 -74.285 31.445 -73.955 ;
        RECT 31.115 -75.645 31.445 -75.315 ;
        RECT 31.115 -77.005 31.445 -76.675 ;
        RECT 31.115 -78.365 31.445 -78.035 ;
        RECT 31.115 -79.725 31.445 -79.395 ;
        RECT 31.115 -81.085 31.445 -80.755 ;
        RECT 31.115 -82.445 31.445 -82.115 ;
        RECT 31.115 -83.805 31.445 -83.475 ;
        RECT 31.115 -85.165 31.445 -84.835 ;
        RECT 31.115 -86.525 31.445 -86.195 ;
        RECT 31.115 -87.885 31.445 -87.555 ;
        RECT 31.115 -89.245 31.445 -88.915 ;
        RECT 31.115 -90.605 31.445 -90.275 ;
        RECT 31.115 -91.965 31.445 -91.635 ;
        RECT 31.115 -93.325 31.445 -92.995 ;
        RECT 31.115 -94.685 31.445 -94.355 ;
        RECT 31.115 -96.045 31.445 -95.715 ;
        RECT 31.115 -97.405 31.445 -97.075 ;
        RECT 31.115 -98.765 31.445 -98.435 ;
        RECT 31.115 -100.125 31.445 -99.795 ;
        RECT 31.115 -101.485 31.445 -101.155 ;
        RECT 31.115 -102.845 31.445 -102.515 ;
        RECT 31.115 -104.205 31.445 -103.875 ;
        RECT 31.115 -105.565 31.445 -105.235 ;
        RECT 31.115 -106.925 31.445 -106.595 ;
        RECT 31.115 -108.285 31.445 -107.955 ;
        RECT 31.115 -109.645 31.445 -109.315 ;
        RECT 31.115 -111.005 31.445 -110.675 ;
        RECT 31.115 -112.365 31.445 -112.035 ;
        RECT 31.115 -113.725 31.445 -113.395 ;
        RECT 31.115 -115.085 31.445 -114.755 ;
        RECT 31.115 -116.445 31.445 -116.115 ;
        RECT 31.115 -117.805 31.445 -117.475 ;
        RECT 31.115 -119.165 31.445 -118.835 ;
        RECT 31.115 -120.525 31.445 -120.195 ;
        RECT 31.115 -121.885 31.445 -121.555 ;
        RECT 31.115 -123.245 31.445 -122.915 ;
        RECT 31.115 -124.605 31.445 -124.275 ;
        RECT 31.115 -125.965 31.445 -125.635 ;
        RECT 31.115 -127.325 31.445 -126.995 ;
        RECT 31.115 -128.685 31.445 -128.355 ;
        RECT 31.115 -130.045 31.445 -129.715 ;
        RECT 31.115 -131.405 31.445 -131.075 ;
        RECT 31.115 -132.765 31.445 -132.435 ;
        RECT 31.115 -134.125 31.445 -133.795 ;
        RECT 31.115 -135.485 31.445 -135.155 ;
        RECT 31.115 -136.845 31.445 -136.515 ;
        RECT 31.115 -138.205 31.445 -137.875 ;
        RECT 31.115 -139.565 31.445 -139.235 ;
        RECT 31.115 -140.925 31.445 -140.595 ;
        RECT 31.115 -142.285 31.445 -141.955 ;
        RECT 31.115 -143.645 31.445 -143.315 ;
        RECT 31.115 -145.005 31.445 -144.675 ;
        RECT 31.115 -146.365 31.445 -146.035 ;
        RECT 31.115 -147.725 31.445 -147.395 ;
        RECT 31.115 -149.085 31.445 -148.755 ;
        RECT 31.115 -150.445 31.445 -150.115 ;
        RECT 31.115 -151.805 31.445 -151.475 ;
        RECT 31.115 -153.165 31.445 -152.835 ;
        RECT 31.115 -158.81 31.445 -157.68 ;
        RECT 31.12 -158.925 31.44 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 44.8 32.805 45.93 ;
        RECT 32.475 39.955 32.805 40.285 ;
        RECT 32.475 38.595 32.805 38.925 ;
        RECT 32.475 36.09 32.805 36.42 ;
        RECT 32.475 33.915 32.805 34.245 ;
        RECT 32.475 32.335 32.805 32.665 ;
        RECT 32.475 31.485 32.805 31.815 ;
        RECT 32.475 29.175 32.805 29.505 ;
        RECT 32.475 28.325 32.805 28.655 ;
        RECT 32.475 26.015 32.805 26.345 ;
        RECT 32.475 25.165 32.805 25.495 ;
        RECT 32.475 22.855 32.805 23.185 ;
        RECT 32.475 22.005 32.805 22.335 ;
        RECT 32.475 19.695 32.805 20.025 ;
        RECT 32.475 18.115 32.805 18.445 ;
        RECT 32.475 17.265 32.805 17.595 ;
        RECT 32.475 14.955 32.805 15.285 ;
        RECT 32.475 14.105 32.805 14.435 ;
        RECT 32.475 11.795 32.805 12.125 ;
        RECT 32.475 10.945 32.805 11.275 ;
        RECT 32.475 8.635 32.805 8.965 ;
        RECT 32.475 7.785 32.805 8.115 ;
        RECT 32.475 5.475 32.805 5.805 ;
        RECT 32.475 3.895 32.805 4.225 ;
        RECT 32.475 3.045 32.805 3.375 ;
        RECT 32.475 0.87 32.805 1.2 ;
        RECT 32.475 -0.845 32.805 -0.515 ;
        RECT 32.475 -2.205 32.805 -1.875 ;
        RECT 32.475 -3.565 32.805 -3.235 ;
        RECT 32.475 -4.925 32.805 -4.595 ;
        RECT 32.475 -6.285 32.805 -5.955 ;
        RECT 32.475 -7.645 32.805 -7.315 ;
        RECT 32.475 -9.005 32.805 -8.675 ;
        RECT 32.475 -10.365 32.805 -10.035 ;
        RECT 32.475 -11.725 32.805 -11.395 ;
        RECT 32.475 -13.085 32.805 -12.755 ;
        RECT 32.475 -14.445 32.805 -14.115 ;
        RECT 32.475 -15.805 32.805 -15.475 ;
        RECT 32.475 -17.165 32.805 -16.835 ;
        RECT 32.475 -18.525 32.805 -18.195 ;
        RECT 32.475 -19.885 32.805 -19.555 ;
        RECT 32.475 -21.245 32.805 -20.915 ;
        RECT 32.475 -22.605 32.805 -22.275 ;
        RECT 32.475 -23.965 32.805 -23.635 ;
        RECT 32.475 -25.325 32.805 -24.995 ;
        RECT 32.475 -26.685 32.805 -26.355 ;
        RECT 32.475 -28.045 32.805 -27.715 ;
        RECT 32.475 -29.405 32.805 -29.075 ;
        RECT 32.475 -30.765 32.805 -30.435 ;
        RECT 32.475 -32.125 32.805 -31.795 ;
        RECT 32.475 -33.485 32.805 -33.155 ;
        RECT 32.475 -34.845 32.805 -34.515 ;
        RECT 32.475 -36.205 32.805 -35.875 ;
        RECT 32.475 -37.565 32.805 -37.235 ;
        RECT 32.475 -38.925 32.805 -38.595 ;
        RECT 32.475 -40.285 32.805 -39.955 ;
        RECT 32.475 -41.645 32.805 -41.315 ;
        RECT 32.475 -43.005 32.805 -42.675 ;
        RECT 32.475 -44.365 32.805 -44.035 ;
        RECT 32.475 -45.725 32.805 -45.395 ;
        RECT 32.475 -47.085 32.805 -46.755 ;
        RECT 32.475 -48.445 32.805 -48.115 ;
        RECT 32.475 -49.805 32.805 -49.475 ;
        RECT 32.475 -51.165 32.805 -50.835 ;
        RECT 32.475 -52.525 32.805 -52.195 ;
        RECT 32.475 -53.885 32.805 -53.555 ;
        RECT 32.475 -55.245 32.805 -54.915 ;
        RECT 32.475 -56.605 32.805 -56.275 ;
        RECT 32.475 -57.965 32.805 -57.635 ;
        RECT 32.475 -59.325 32.805 -58.995 ;
        RECT 32.475 -60.685 32.805 -60.355 ;
        RECT 32.475 -62.045 32.805 -61.715 ;
        RECT 32.475 -63.405 32.805 -63.075 ;
        RECT 32.475 -64.765 32.805 -64.435 ;
        RECT 32.475 -66.125 32.805 -65.795 ;
        RECT 32.475 -67.485 32.805 -67.155 ;
        RECT 32.475 -68.845 32.805 -68.515 ;
        RECT 32.475 -70.205 32.805 -69.875 ;
        RECT 32.475 -71.565 32.805 -71.235 ;
        RECT 32.475 -72.925 32.805 -72.595 ;
        RECT 32.475 -74.285 32.805 -73.955 ;
        RECT 32.475 -75.645 32.805 -75.315 ;
        RECT 32.475 -77.005 32.805 -76.675 ;
        RECT 32.475 -78.365 32.805 -78.035 ;
        RECT 32.475 -79.725 32.805 -79.395 ;
        RECT 32.475 -81.085 32.805 -80.755 ;
        RECT 32.475 -82.445 32.805 -82.115 ;
        RECT 32.475 -83.805 32.805 -83.475 ;
        RECT 32.475 -85.165 32.805 -84.835 ;
        RECT 32.475 -86.525 32.805 -86.195 ;
        RECT 32.475 -87.885 32.805 -87.555 ;
        RECT 32.475 -89.245 32.805 -88.915 ;
        RECT 32.475 -90.605 32.805 -90.275 ;
        RECT 32.475 -91.965 32.805 -91.635 ;
        RECT 32.475 -93.325 32.805 -92.995 ;
        RECT 32.475 -94.685 32.805 -94.355 ;
        RECT 32.475 -96.045 32.805 -95.715 ;
        RECT 32.475 -97.405 32.805 -97.075 ;
        RECT 32.475 -98.765 32.805 -98.435 ;
        RECT 32.475 -100.125 32.805 -99.795 ;
        RECT 32.475 -101.485 32.805 -101.155 ;
        RECT 32.475 -102.845 32.805 -102.515 ;
        RECT 32.475 -104.205 32.805 -103.875 ;
        RECT 32.475 -105.565 32.805 -105.235 ;
        RECT 32.475 -106.925 32.805 -106.595 ;
        RECT 32.475 -108.285 32.805 -107.955 ;
        RECT 32.475 -109.645 32.805 -109.315 ;
        RECT 32.475 -111.005 32.805 -110.675 ;
        RECT 32.475 -112.365 32.805 -112.035 ;
        RECT 32.475 -113.725 32.805 -113.395 ;
        RECT 32.475 -115.085 32.805 -114.755 ;
        RECT 32.475 -116.445 32.805 -116.115 ;
        RECT 32.475 -117.805 32.805 -117.475 ;
        RECT 32.475 -119.165 32.805 -118.835 ;
        RECT 32.475 -120.525 32.805 -120.195 ;
        RECT 32.475 -121.885 32.805 -121.555 ;
        RECT 32.475 -123.245 32.805 -122.915 ;
        RECT 32.475 -124.605 32.805 -124.275 ;
        RECT 32.475 -125.965 32.805 -125.635 ;
        RECT 32.475 -127.325 32.805 -126.995 ;
        RECT 32.475 -128.685 32.805 -128.355 ;
        RECT 32.475 -130.045 32.805 -129.715 ;
        RECT 32.475 -131.405 32.805 -131.075 ;
        RECT 32.475 -132.765 32.805 -132.435 ;
        RECT 32.475 -134.125 32.805 -133.795 ;
        RECT 32.475 -135.485 32.805 -135.155 ;
        RECT 32.475 -136.845 32.805 -136.515 ;
        RECT 32.475 -138.205 32.805 -137.875 ;
        RECT 32.475 -139.565 32.805 -139.235 ;
        RECT 32.475 -140.925 32.805 -140.595 ;
        RECT 32.475 -142.285 32.805 -141.955 ;
        RECT 32.475 -143.645 32.805 -143.315 ;
        RECT 32.475 -145.005 32.805 -144.675 ;
        RECT 32.475 -146.365 32.805 -146.035 ;
        RECT 32.475 -147.725 32.805 -147.395 ;
        RECT 32.475 -149.085 32.805 -148.755 ;
        RECT 32.475 -150.445 32.805 -150.115 ;
        RECT 32.475 -151.805 32.805 -151.475 ;
        RECT 32.475 -153.165 32.805 -152.835 ;
        RECT 32.475 -158.81 32.805 -157.68 ;
        RECT 32.48 -158.925 32.8 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 44.8 34.165 45.93 ;
        RECT 33.835 39.955 34.165 40.285 ;
        RECT 33.835 38.595 34.165 38.925 ;
        RECT 33.835 36.09 34.165 36.42 ;
        RECT 33.835 33.915 34.165 34.245 ;
        RECT 33.835 32.335 34.165 32.665 ;
        RECT 33.835 31.485 34.165 31.815 ;
        RECT 33.835 29.175 34.165 29.505 ;
        RECT 33.835 28.325 34.165 28.655 ;
        RECT 33.835 26.015 34.165 26.345 ;
        RECT 33.835 25.165 34.165 25.495 ;
        RECT 33.835 22.855 34.165 23.185 ;
        RECT 33.835 22.005 34.165 22.335 ;
        RECT 33.835 19.695 34.165 20.025 ;
        RECT 33.835 18.115 34.165 18.445 ;
        RECT 33.835 17.265 34.165 17.595 ;
        RECT 33.835 14.955 34.165 15.285 ;
        RECT 33.835 14.105 34.165 14.435 ;
        RECT 33.835 11.795 34.165 12.125 ;
        RECT 33.835 10.945 34.165 11.275 ;
        RECT 33.835 8.635 34.165 8.965 ;
        RECT 33.835 7.785 34.165 8.115 ;
        RECT 33.835 5.475 34.165 5.805 ;
        RECT 33.835 3.895 34.165 4.225 ;
        RECT 33.835 3.045 34.165 3.375 ;
        RECT 33.835 0.87 34.165 1.2 ;
        RECT 33.835 -0.845 34.165 -0.515 ;
        RECT 33.835 -2.205 34.165 -1.875 ;
        RECT 33.835 -3.565 34.165 -3.235 ;
        RECT 33.835 -4.925 34.165 -4.595 ;
        RECT 33.835 -6.285 34.165 -5.955 ;
        RECT 33.835 -7.645 34.165 -7.315 ;
        RECT 33.835 -9.005 34.165 -8.675 ;
        RECT 33.835 -10.365 34.165 -10.035 ;
        RECT 33.835 -11.725 34.165 -11.395 ;
        RECT 33.835 -13.085 34.165 -12.755 ;
        RECT 33.835 -14.445 34.165 -14.115 ;
        RECT 33.835 -15.805 34.165 -15.475 ;
        RECT 33.835 -17.165 34.165 -16.835 ;
        RECT 33.835 -18.525 34.165 -18.195 ;
        RECT 33.835 -19.885 34.165 -19.555 ;
        RECT 33.835 -21.245 34.165 -20.915 ;
        RECT 33.835 -22.605 34.165 -22.275 ;
        RECT 33.835 -23.965 34.165 -23.635 ;
        RECT 33.835 -25.325 34.165 -24.995 ;
        RECT 33.835 -26.685 34.165 -26.355 ;
        RECT 33.835 -28.045 34.165 -27.715 ;
        RECT 33.835 -29.405 34.165 -29.075 ;
        RECT 33.835 -30.765 34.165 -30.435 ;
        RECT 33.835 -32.125 34.165 -31.795 ;
        RECT 33.835 -33.485 34.165 -33.155 ;
        RECT 33.835 -34.845 34.165 -34.515 ;
        RECT 33.835 -36.205 34.165 -35.875 ;
        RECT 33.835 -37.565 34.165 -37.235 ;
        RECT 33.835 -38.925 34.165 -38.595 ;
        RECT 33.835 -40.285 34.165 -39.955 ;
        RECT 33.835 -41.645 34.165 -41.315 ;
        RECT 33.835 -43.005 34.165 -42.675 ;
        RECT 33.835 -44.365 34.165 -44.035 ;
        RECT 33.835 -45.725 34.165 -45.395 ;
        RECT 33.835 -47.085 34.165 -46.755 ;
        RECT 33.835 -48.445 34.165 -48.115 ;
        RECT 33.835 -49.805 34.165 -49.475 ;
        RECT 33.835 -51.165 34.165 -50.835 ;
        RECT 33.835 -52.525 34.165 -52.195 ;
        RECT 33.835 -53.885 34.165 -53.555 ;
        RECT 33.835 -55.245 34.165 -54.915 ;
        RECT 33.835 -56.605 34.165 -56.275 ;
        RECT 33.835 -57.965 34.165 -57.635 ;
        RECT 33.835 -59.325 34.165 -58.995 ;
        RECT 33.835 -60.685 34.165 -60.355 ;
        RECT 33.835 -62.045 34.165 -61.715 ;
        RECT 33.835 -63.405 34.165 -63.075 ;
        RECT 33.835 -64.765 34.165 -64.435 ;
        RECT 33.835 -66.125 34.165 -65.795 ;
        RECT 33.835 -67.485 34.165 -67.155 ;
        RECT 33.835 -68.845 34.165 -68.515 ;
        RECT 33.835 -70.205 34.165 -69.875 ;
        RECT 33.835 -71.565 34.165 -71.235 ;
        RECT 33.835 -72.925 34.165 -72.595 ;
        RECT 33.835 -74.285 34.165 -73.955 ;
        RECT 33.835 -75.645 34.165 -75.315 ;
        RECT 33.835 -77.005 34.165 -76.675 ;
        RECT 33.835 -78.365 34.165 -78.035 ;
        RECT 33.835 -79.725 34.165 -79.395 ;
        RECT 33.835 -81.085 34.165 -80.755 ;
        RECT 33.835 -82.445 34.165 -82.115 ;
        RECT 33.835 -83.805 34.165 -83.475 ;
        RECT 33.835 -85.165 34.165 -84.835 ;
        RECT 33.835 -86.525 34.165 -86.195 ;
        RECT 33.835 -87.885 34.165 -87.555 ;
        RECT 33.835 -89.245 34.165 -88.915 ;
        RECT 33.835 -90.605 34.165 -90.275 ;
        RECT 33.835 -91.965 34.165 -91.635 ;
        RECT 33.835 -93.325 34.165 -92.995 ;
        RECT 33.835 -94.685 34.165 -94.355 ;
        RECT 33.835 -96.045 34.165 -95.715 ;
        RECT 33.835 -97.405 34.165 -97.075 ;
        RECT 33.835 -98.765 34.165 -98.435 ;
        RECT 33.835 -100.125 34.165 -99.795 ;
        RECT 33.835 -101.485 34.165 -101.155 ;
        RECT 33.835 -102.845 34.165 -102.515 ;
        RECT 33.835 -104.205 34.165 -103.875 ;
        RECT 33.835 -105.565 34.165 -105.235 ;
        RECT 33.835 -106.925 34.165 -106.595 ;
        RECT 33.835 -108.285 34.165 -107.955 ;
        RECT 33.835 -109.645 34.165 -109.315 ;
        RECT 33.835 -111.005 34.165 -110.675 ;
        RECT 33.835 -112.365 34.165 -112.035 ;
        RECT 33.835 -113.725 34.165 -113.395 ;
        RECT 33.835 -115.085 34.165 -114.755 ;
        RECT 33.835 -116.445 34.165 -116.115 ;
        RECT 33.835 -117.805 34.165 -117.475 ;
        RECT 33.835 -119.165 34.165 -118.835 ;
        RECT 33.835 -120.525 34.165 -120.195 ;
        RECT 33.835 -121.885 34.165 -121.555 ;
        RECT 33.835 -123.245 34.165 -122.915 ;
        RECT 33.835 -124.605 34.165 -124.275 ;
        RECT 33.835 -125.965 34.165 -125.635 ;
        RECT 33.835 -127.325 34.165 -126.995 ;
        RECT 33.835 -128.685 34.165 -128.355 ;
        RECT 33.835 -130.045 34.165 -129.715 ;
        RECT 33.835 -131.405 34.165 -131.075 ;
        RECT 33.835 -132.765 34.165 -132.435 ;
        RECT 33.835 -134.125 34.165 -133.795 ;
        RECT 33.835 -135.485 34.165 -135.155 ;
        RECT 33.835 -136.845 34.165 -136.515 ;
        RECT 33.835 -138.205 34.165 -137.875 ;
        RECT 33.835 -139.565 34.165 -139.235 ;
        RECT 33.835 -140.925 34.165 -140.595 ;
        RECT 33.835 -142.285 34.165 -141.955 ;
        RECT 33.835 -143.645 34.165 -143.315 ;
        RECT 33.835 -145.005 34.165 -144.675 ;
        RECT 33.835 -146.365 34.165 -146.035 ;
        RECT 33.835 -147.725 34.165 -147.395 ;
        RECT 33.835 -149.085 34.165 -148.755 ;
        RECT 33.835 -150.445 34.165 -150.115 ;
        RECT 33.835 -151.805 34.165 -151.475 ;
        RECT 33.835 -153.165 34.165 -152.835 ;
        RECT 33.835 -158.81 34.165 -157.68 ;
        RECT 33.84 -158.925 34.16 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 44.8 35.525 45.93 ;
        RECT 35.195 39.955 35.525 40.285 ;
        RECT 35.195 38.595 35.525 38.925 ;
        RECT 35.195 36.09 35.525 36.42 ;
        RECT 35.195 33.915 35.525 34.245 ;
        RECT 35.195 32.335 35.525 32.665 ;
        RECT 35.195 31.485 35.525 31.815 ;
        RECT 35.195 29.175 35.525 29.505 ;
        RECT 35.195 28.325 35.525 28.655 ;
        RECT 35.195 26.015 35.525 26.345 ;
        RECT 35.195 25.165 35.525 25.495 ;
        RECT 35.195 22.855 35.525 23.185 ;
        RECT 35.195 22.005 35.525 22.335 ;
        RECT 35.195 19.695 35.525 20.025 ;
        RECT 35.195 18.115 35.525 18.445 ;
        RECT 35.195 17.265 35.525 17.595 ;
        RECT 35.195 14.955 35.525 15.285 ;
        RECT 35.195 14.105 35.525 14.435 ;
        RECT 35.195 11.795 35.525 12.125 ;
        RECT 35.195 10.945 35.525 11.275 ;
        RECT 35.195 8.635 35.525 8.965 ;
        RECT 35.195 7.785 35.525 8.115 ;
        RECT 35.195 5.475 35.525 5.805 ;
        RECT 35.195 3.895 35.525 4.225 ;
        RECT 35.195 3.045 35.525 3.375 ;
        RECT 35.195 0.87 35.525 1.2 ;
        RECT 35.195 -0.845 35.525 -0.515 ;
        RECT 35.195 -2.205 35.525 -1.875 ;
        RECT 35.195 -3.565 35.525 -3.235 ;
        RECT 35.195 -4.925 35.525 -4.595 ;
        RECT 35.195 -6.285 35.525 -5.955 ;
        RECT 35.195 -7.645 35.525 -7.315 ;
        RECT 35.195 -9.005 35.525 -8.675 ;
        RECT 35.195 -10.365 35.525 -10.035 ;
        RECT 35.195 -11.725 35.525 -11.395 ;
        RECT 35.195 -13.085 35.525 -12.755 ;
        RECT 35.195 -14.445 35.525 -14.115 ;
        RECT 35.195 -15.805 35.525 -15.475 ;
        RECT 35.195 -17.165 35.525 -16.835 ;
        RECT 35.195 -18.525 35.525 -18.195 ;
        RECT 35.195 -19.885 35.525 -19.555 ;
        RECT 35.195 -21.245 35.525 -20.915 ;
        RECT 35.195 -22.605 35.525 -22.275 ;
        RECT 35.195 -23.965 35.525 -23.635 ;
        RECT 35.195 -25.325 35.525 -24.995 ;
        RECT 35.195 -26.685 35.525 -26.355 ;
        RECT 35.195 -28.045 35.525 -27.715 ;
        RECT 35.195 -29.405 35.525 -29.075 ;
        RECT 35.195 -30.765 35.525 -30.435 ;
        RECT 35.195 -32.125 35.525 -31.795 ;
        RECT 35.195 -33.485 35.525 -33.155 ;
        RECT 35.195 -34.845 35.525 -34.515 ;
        RECT 35.195 -36.205 35.525 -35.875 ;
        RECT 35.195 -37.565 35.525 -37.235 ;
        RECT 35.195 -38.925 35.525 -38.595 ;
        RECT 35.195 -40.285 35.525 -39.955 ;
        RECT 35.195 -41.645 35.525 -41.315 ;
        RECT 35.195 -43.005 35.525 -42.675 ;
        RECT 35.195 -44.365 35.525 -44.035 ;
        RECT 35.195 -45.725 35.525 -45.395 ;
        RECT 35.195 -47.085 35.525 -46.755 ;
        RECT 35.195 -48.445 35.525 -48.115 ;
        RECT 35.195 -49.805 35.525 -49.475 ;
        RECT 35.195 -51.165 35.525 -50.835 ;
        RECT 35.195 -52.525 35.525 -52.195 ;
        RECT 35.195 -53.885 35.525 -53.555 ;
        RECT 35.195 -55.245 35.525 -54.915 ;
        RECT 35.195 -56.605 35.525 -56.275 ;
        RECT 35.195 -57.965 35.525 -57.635 ;
        RECT 35.195 -59.325 35.525 -58.995 ;
        RECT 35.195 -60.685 35.525 -60.355 ;
        RECT 35.195 -62.045 35.525 -61.715 ;
        RECT 35.195 -63.405 35.525 -63.075 ;
        RECT 35.195 -64.765 35.525 -64.435 ;
        RECT 35.195 -66.125 35.525 -65.795 ;
        RECT 35.195 -67.485 35.525 -67.155 ;
        RECT 35.195 -68.845 35.525 -68.515 ;
        RECT 35.195 -70.205 35.525 -69.875 ;
        RECT 35.195 -71.565 35.525 -71.235 ;
        RECT 35.195 -72.925 35.525 -72.595 ;
        RECT 35.195 -74.285 35.525 -73.955 ;
        RECT 35.195 -75.645 35.525 -75.315 ;
        RECT 35.195 -77.005 35.525 -76.675 ;
        RECT 35.195 -78.365 35.525 -78.035 ;
        RECT 35.195 -79.725 35.525 -79.395 ;
        RECT 35.195 -81.085 35.525 -80.755 ;
        RECT 35.195 -82.445 35.525 -82.115 ;
        RECT 35.195 -83.805 35.525 -83.475 ;
        RECT 35.195 -85.165 35.525 -84.835 ;
        RECT 35.195 -86.525 35.525 -86.195 ;
        RECT 35.195 -87.885 35.525 -87.555 ;
        RECT 35.195 -89.245 35.525 -88.915 ;
        RECT 35.195 -90.605 35.525 -90.275 ;
        RECT 35.195 -91.965 35.525 -91.635 ;
        RECT 35.195 -93.325 35.525 -92.995 ;
        RECT 35.195 -94.685 35.525 -94.355 ;
        RECT 35.195 -96.045 35.525 -95.715 ;
        RECT 35.195 -97.405 35.525 -97.075 ;
        RECT 35.195 -98.765 35.525 -98.435 ;
        RECT 35.195 -100.125 35.525 -99.795 ;
        RECT 35.195 -101.485 35.525 -101.155 ;
        RECT 35.195 -102.845 35.525 -102.515 ;
        RECT 35.195 -104.205 35.525 -103.875 ;
        RECT 35.195 -105.565 35.525 -105.235 ;
        RECT 35.195 -106.925 35.525 -106.595 ;
        RECT 35.195 -108.285 35.525 -107.955 ;
        RECT 35.195 -109.645 35.525 -109.315 ;
        RECT 35.195 -111.005 35.525 -110.675 ;
        RECT 35.195 -112.365 35.525 -112.035 ;
        RECT 35.195 -113.725 35.525 -113.395 ;
        RECT 35.195 -115.085 35.525 -114.755 ;
        RECT 35.195 -116.445 35.525 -116.115 ;
        RECT 35.195 -117.805 35.525 -117.475 ;
        RECT 35.195 -119.165 35.525 -118.835 ;
        RECT 35.195 -120.525 35.525 -120.195 ;
        RECT 35.195 -121.885 35.525 -121.555 ;
        RECT 35.195 -123.245 35.525 -122.915 ;
        RECT 35.195 -124.605 35.525 -124.275 ;
        RECT 35.195 -125.965 35.525 -125.635 ;
        RECT 35.195 -127.325 35.525 -126.995 ;
        RECT 35.195 -128.685 35.525 -128.355 ;
        RECT 35.195 -130.045 35.525 -129.715 ;
        RECT 35.195 -131.405 35.525 -131.075 ;
        RECT 35.195 -132.765 35.525 -132.435 ;
        RECT 35.195 -134.125 35.525 -133.795 ;
        RECT 35.195 -135.485 35.525 -135.155 ;
        RECT 35.195 -136.845 35.525 -136.515 ;
        RECT 35.195 -138.205 35.525 -137.875 ;
        RECT 35.195 -139.565 35.525 -139.235 ;
        RECT 35.195 -140.925 35.525 -140.595 ;
        RECT 35.195 -142.285 35.525 -141.955 ;
        RECT 35.195 -143.645 35.525 -143.315 ;
        RECT 35.195 -145.005 35.525 -144.675 ;
        RECT 35.195 -146.365 35.525 -146.035 ;
        RECT 35.195 -147.725 35.525 -147.395 ;
        RECT 35.195 -149.085 35.525 -148.755 ;
        RECT 35.195 -150.445 35.525 -150.115 ;
        RECT 35.195 -151.805 35.525 -151.475 ;
        RECT 35.195 -153.165 35.525 -152.835 ;
        RECT 35.195 -158.81 35.525 -157.68 ;
        RECT 35.2 -158.925 35.52 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.555 44.8 36.885 45.93 ;
        RECT 36.555 39.955 36.885 40.285 ;
        RECT 36.555 38.595 36.885 38.925 ;
        RECT 36.555 -0.845 36.885 -0.515 ;
        RECT 36.555 -2.205 36.885 -1.875 ;
        RECT 36.555 -3.565 36.885 -3.235 ;
        RECT 36.555 -4.925 36.885 -4.595 ;
        RECT 36.555 -6.285 36.885 -5.955 ;
        RECT 36.555 -7.645 36.885 -7.315 ;
        RECT 36.555 -9.005 36.885 -8.675 ;
        RECT 36.555 -10.365 36.885 -10.035 ;
        RECT 36.555 -11.725 36.885 -11.395 ;
        RECT 36.555 -13.085 36.885 -12.755 ;
        RECT 36.555 -14.445 36.885 -14.115 ;
        RECT 36.555 -15.805 36.885 -15.475 ;
        RECT 36.555 -17.165 36.885 -16.835 ;
        RECT 36.555 -18.525 36.885 -18.195 ;
        RECT 36.555 -19.885 36.885 -19.555 ;
        RECT 36.555 -21.245 36.885 -20.915 ;
        RECT 36.555 -22.605 36.885 -22.275 ;
        RECT 36.555 -23.965 36.885 -23.635 ;
        RECT 36.555 -25.325 36.885 -24.995 ;
        RECT 36.555 -26.685 36.885 -26.355 ;
        RECT 36.555 -28.045 36.885 -27.715 ;
        RECT 36.555 -29.405 36.885 -29.075 ;
        RECT 36.555 -30.765 36.885 -30.435 ;
        RECT 36.555 -32.125 36.885 -31.795 ;
        RECT 36.555 -33.485 36.885 -33.155 ;
        RECT 36.555 -34.845 36.885 -34.515 ;
        RECT 36.555 -36.205 36.885 -35.875 ;
        RECT 36.555 -37.565 36.885 -37.235 ;
        RECT 36.555 -38.925 36.885 -38.595 ;
        RECT 36.555 -40.285 36.885 -39.955 ;
        RECT 36.555 -41.645 36.885 -41.315 ;
        RECT 36.555 -43.005 36.885 -42.675 ;
        RECT 36.555 -44.365 36.885 -44.035 ;
        RECT 36.555 -45.725 36.885 -45.395 ;
        RECT 36.555 -47.085 36.885 -46.755 ;
        RECT 36.555 -48.445 36.885 -48.115 ;
        RECT 36.555 -49.805 36.885 -49.475 ;
        RECT 36.555 -51.165 36.885 -50.835 ;
        RECT 36.555 -52.525 36.885 -52.195 ;
        RECT 36.555 -53.885 36.885 -53.555 ;
        RECT 36.555 -55.245 36.885 -54.915 ;
        RECT 36.555 -56.605 36.885 -56.275 ;
        RECT 36.555 -57.965 36.885 -57.635 ;
        RECT 36.555 -59.325 36.885 -58.995 ;
        RECT 36.555 -60.685 36.885 -60.355 ;
        RECT 36.555 -62.045 36.885 -61.715 ;
        RECT 36.555 -63.405 36.885 -63.075 ;
        RECT 36.555 -64.765 36.885 -64.435 ;
        RECT 36.555 -66.125 36.885 -65.795 ;
        RECT 36.555 -67.485 36.885 -67.155 ;
        RECT 36.555 -68.845 36.885 -68.515 ;
        RECT 36.555 -70.205 36.885 -69.875 ;
        RECT 36.555 -71.565 36.885 -71.235 ;
        RECT 36.555 -72.925 36.885 -72.595 ;
        RECT 36.555 -74.285 36.885 -73.955 ;
        RECT 36.555 -75.645 36.885 -75.315 ;
        RECT 36.555 -77.005 36.885 -76.675 ;
        RECT 36.555 -78.365 36.885 -78.035 ;
        RECT 36.555 -79.725 36.885 -79.395 ;
        RECT 36.555 -81.085 36.885 -80.755 ;
        RECT 36.555 -82.445 36.885 -82.115 ;
        RECT 36.555 -83.805 36.885 -83.475 ;
        RECT 36.555 -85.165 36.885 -84.835 ;
        RECT 36.555 -86.525 36.885 -86.195 ;
        RECT 36.555 -87.885 36.885 -87.555 ;
        RECT 36.555 -89.245 36.885 -88.915 ;
        RECT 36.555 -90.605 36.885 -90.275 ;
        RECT 36.555 -91.965 36.885 -91.635 ;
        RECT 36.555 -93.325 36.885 -92.995 ;
        RECT 36.555 -94.685 36.885 -94.355 ;
        RECT 36.555 -96.045 36.885 -95.715 ;
        RECT 36.555 -97.405 36.885 -97.075 ;
        RECT 36.555 -98.765 36.885 -98.435 ;
        RECT 36.555 -100.125 36.885 -99.795 ;
        RECT 36.555 -101.485 36.885 -101.155 ;
        RECT 36.555 -102.845 36.885 -102.515 ;
        RECT 36.555 -104.205 36.885 -103.875 ;
        RECT 36.555 -105.565 36.885 -105.235 ;
        RECT 36.555 -106.925 36.885 -106.595 ;
        RECT 36.555 -108.285 36.885 -107.955 ;
        RECT 36.555 -109.645 36.885 -109.315 ;
        RECT 36.555 -111.005 36.885 -110.675 ;
        RECT 36.555 -112.365 36.885 -112.035 ;
        RECT 36.555 -113.725 36.885 -113.395 ;
        RECT 36.555 -115.085 36.885 -114.755 ;
        RECT 36.555 -116.445 36.885 -116.115 ;
        RECT 36.555 -117.805 36.885 -117.475 ;
        RECT 36.555 -119.165 36.885 -118.835 ;
        RECT 36.555 -120.525 36.885 -120.195 ;
        RECT 36.555 -121.885 36.885 -121.555 ;
        RECT 36.555 -123.245 36.885 -122.915 ;
        RECT 36.555 -124.605 36.885 -124.275 ;
        RECT 36.555 -125.965 36.885 -125.635 ;
        RECT 36.555 -127.325 36.885 -126.995 ;
        RECT 36.555 -128.685 36.885 -128.355 ;
        RECT 36.555 -130.045 36.885 -129.715 ;
        RECT 36.555 -131.405 36.885 -131.075 ;
        RECT 36.555 -132.765 36.885 -132.435 ;
        RECT 36.555 -134.125 36.885 -133.795 ;
        RECT 36.555 -135.485 36.885 -135.155 ;
        RECT 36.555 -136.845 36.885 -136.515 ;
        RECT 36.555 -138.205 36.885 -137.875 ;
        RECT 36.555 -139.565 36.885 -139.235 ;
        RECT 36.555 -140.925 36.885 -140.595 ;
        RECT 36.555 -142.285 36.885 -141.955 ;
        RECT 36.555 -143.645 36.885 -143.315 ;
        RECT 36.555 -145.005 36.885 -144.675 ;
        RECT 36.555 -146.365 36.885 -146.035 ;
        RECT 36.555 -147.725 36.885 -147.395 ;
        RECT 36.555 -149.085 36.885 -148.755 ;
        RECT 36.555 -150.445 36.885 -150.115 ;
        RECT 36.555 -151.805 36.885 -151.475 ;
        RECT 36.555 -153.165 36.885 -152.835 ;
        RECT 36.555 -158.81 36.885 -157.68 ;
        RECT 36.56 -158.925 36.88 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.605 44.8 -5.275 45.93 ;
        RECT -5.605 39.955 -5.275 40.285 ;
        RECT -5.605 38.595 -5.275 38.925 ;
        RECT -5.605 36.09 -5.275 36.42 ;
        RECT -5.605 33.915 -5.275 34.245 ;
        RECT -5.605 32.335 -5.275 32.665 ;
        RECT -5.605 31.485 -5.275 31.815 ;
        RECT -5.605 29.175 -5.275 29.505 ;
        RECT -5.605 28.325 -5.275 28.655 ;
        RECT -5.605 26.015 -5.275 26.345 ;
        RECT -5.605 25.165 -5.275 25.495 ;
        RECT -5.605 22.855 -5.275 23.185 ;
        RECT -5.605 22.005 -5.275 22.335 ;
        RECT -5.605 19.695 -5.275 20.025 ;
        RECT -5.605 18.115 -5.275 18.445 ;
        RECT -5.605 17.265 -5.275 17.595 ;
        RECT -5.605 14.955 -5.275 15.285 ;
        RECT -5.605 14.105 -5.275 14.435 ;
        RECT -5.605 11.795 -5.275 12.125 ;
        RECT -5.605 10.945 -5.275 11.275 ;
        RECT -5.605 8.635 -5.275 8.965 ;
        RECT -5.605 7.785 -5.275 8.115 ;
        RECT -5.605 5.475 -5.275 5.805 ;
        RECT -5.605 3.895 -5.275 4.225 ;
        RECT -5.605 3.045 -5.275 3.375 ;
        RECT -5.605 0.87 -5.275 1.2 ;
        RECT -5.605 -0.845 -5.275 -0.515 ;
        RECT -5.605 -2.205 -5.275 -1.875 ;
        RECT -5.605 -3.565 -5.275 -3.235 ;
        RECT -5.605 -4.925 -5.275 -4.595 ;
        RECT -5.605 -6.285 -5.275 -5.955 ;
        RECT -5.605 -7.645 -5.275 -7.315 ;
        RECT -5.605 -9.005 -5.275 -8.675 ;
        RECT -5.605 -10.365 -5.275 -10.035 ;
        RECT -5.605 -11.725 -5.275 -11.395 ;
        RECT -5.605 -13.085 -5.275 -12.755 ;
        RECT -5.605 -14.445 -5.275 -14.115 ;
        RECT -5.605 -15.805 -5.275 -15.475 ;
        RECT -5.605 -17.165 -5.275 -16.835 ;
        RECT -5.605 -21.245 -5.275 -20.915 ;
        RECT -5.605 -22.605 -5.275 -22.275 ;
        RECT -5.605 -23.965 -5.275 -23.635 ;
        RECT -5.605 -25.325 -5.275 -24.995 ;
        RECT -5.605 -26.685 -5.275 -26.355 ;
        RECT -5.605 -28.045 -5.275 -27.715 ;
        RECT -5.605 -29.405 -5.275 -29.075 ;
        RECT -5.605 -30.765 -5.275 -30.435 ;
        RECT -5.605 -32.125 -5.275 -31.795 ;
        RECT -5.605 -33.485 -5.275 -33.155 ;
        RECT -5.605 -36.205 -5.275 -35.875 ;
        RECT -5.605 -37.565 -5.275 -37.235 ;
        RECT -5.605 -38.925 -5.275 -38.595 ;
        RECT -5.605 -40.285 -5.275 -39.955 ;
        RECT -5.605 -43.005 -5.275 -42.675 ;
        RECT -5.605 -45.725 -5.275 -45.395 ;
        RECT -5.605 -47.085 -5.275 -46.755 ;
        RECT -5.605 -48.445 -5.275 -48.115 ;
        RECT -5.605 -49.805 -5.275 -49.475 ;
        RECT -5.605 -51.165 -5.275 -50.835 ;
        RECT -5.605 -52.525 -5.275 -52.195 ;
        RECT -5.605 -53.885 -5.275 -53.555 ;
        RECT -5.605 -55.245 -5.275 -54.915 ;
        RECT -5.605 -56.605 -5.275 -56.275 ;
        RECT -5.605 -57.965 -5.275 -57.635 ;
        RECT -5.605 -59.325 -5.275 -58.995 ;
        RECT -5.605 -60.685 -5.275 -60.355 ;
        RECT -5.605 -62.045 -5.275 -61.715 ;
        RECT -5.605 -63.405 -5.275 -63.075 ;
        RECT -5.605 -64.765 -5.275 -64.435 ;
        RECT -5.605 -66.125 -5.275 -65.795 ;
        RECT -5.605 -67.485 -5.275 -67.155 ;
        RECT -5.605 -68.845 -5.275 -68.515 ;
        RECT -5.605 -70.205 -5.275 -69.875 ;
        RECT -5.605 -71.565 -5.275 -71.235 ;
        RECT -5.605 -72.925 -5.275 -72.595 ;
        RECT -5.605 -74.285 -5.275 -73.955 ;
        RECT -5.605 -75.645 -5.275 -75.315 ;
        RECT -5.605 -77.005 -5.275 -76.675 ;
        RECT -5.605 -78.365 -5.275 -78.035 ;
        RECT -5.605 -79.725 -5.275 -79.395 ;
        RECT -5.605 -81.085 -5.275 -80.755 ;
        RECT -5.605 -82.445 -5.275 -82.115 ;
        RECT -5.605 -83.805 -5.275 -83.475 ;
        RECT -5.605 -85.165 -5.275 -84.835 ;
        RECT -5.605 -87.885 -5.275 -87.555 ;
        RECT -5.605 -89.245 -5.275 -88.915 ;
        RECT -5.605 -90.605 -5.275 -90.275 ;
        RECT -5.605 -91.965 -5.275 -91.635 ;
        RECT -5.605 -93.325 -5.275 -92.995 ;
        RECT -5.605 -94.685 -5.275 -94.355 ;
        RECT -5.605 -96.045 -5.275 -95.715 ;
        RECT -5.605 -97.405 -5.275 -97.075 ;
        RECT -5.605 -98.765 -5.275 -98.435 ;
        RECT -5.605 -100.125 -5.275 -99.795 ;
        RECT -5.605 -101.485 -5.275 -101.155 ;
        RECT -5.605 -102.845 -5.275 -102.515 ;
        RECT -5.605 -104.205 -5.275 -103.875 ;
        RECT -5.605 -105.565 -5.275 -105.235 ;
        RECT -5.605 -106.925 -5.275 -106.595 ;
        RECT -5.605 -108.285 -5.275 -107.955 ;
        RECT -5.605 -109.645 -5.275 -109.315 ;
        RECT -5.605 -111.005 -5.275 -110.675 ;
        RECT -5.605 -112.365 -5.275 -112.035 ;
        RECT -5.605 -113.725 -5.275 -113.395 ;
        RECT -5.605 -115.085 -5.275 -114.755 ;
        RECT -5.605 -116.445 -5.275 -116.115 ;
        RECT -5.605 -117.805 -5.275 -117.475 ;
        RECT -5.605 -119.165 -5.275 -118.835 ;
        RECT -5.605 -120.525 -5.275 -120.195 ;
        RECT -5.605 -121.885 -5.275 -121.555 ;
        RECT -5.605 -123.245 -5.275 -122.915 ;
        RECT -5.605 -124.605 -5.275 -124.275 ;
        RECT -5.605 -125.965 -5.275 -125.635 ;
        RECT -5.605 -127.325 -5.275 -126.995 ;
        RECT -5.605 -128.685 -5.275 -128.355 ;
        RECT -5.605 -130.045 -5.275 -129.715 ;
        RECT -5.605 -131.405 -5.275 -131.075 ;
        RECT -5.605 -132.765 -5.275 -132.435 ;
        RECT -5.605 -134.125 -5.275 -133.795 ;
        RECT -5.605 -135.485 -5.275 -135.155 ;
        RECT -5.605 -136.845 -5.275 -136.515 ;
        RECT -5.605 -138.205 -5.275 -137.875 ;
        RECT -5.605 -139.565 -5.275 -139.235 ;
        RECT -5.605 -140.925 -5.275 -140.595 ;
        RECT -5.605 -142.285 -5.275 -141.955 ;
        RECT -5.605 -143.645 -5.275 -143.315 ;
        RECT -5.605 -145.005 -5.275 -144.675 ;
        RECT -5.605 -146.365 -5.275 -146.035 ;
        RECT -5.605 -147.725 -5.275 -147.395 ;
        RECT -5.605 -149.085 -5.275 -148.755 ;
        RECT -5.605 -150.445 -5.275 -150.115 ;
        RECT -5.605 -151.805 -5.275 -151.475 ;
        RECT -5.605 -153.165 -5.275 -152.835 ;
        RECT -5.605 -158.81 -5.275 -157.68 ;
        RECT -5.6 -158.925 -5.28 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.245 44.8 -3.915 45.93 ;
        RECT -4.245 39.955 -3.915 40.285 ;
        RECT -4.245 38.595 -3.915 38.925 ;
        RECT -4.245 36.09 -3.915 36.42 ;
        RECT -4.245 33.915 -3.915 34.245 ;
        RECT -4.245 32.335 -3.915 32.665 ;
        RECT -4.245 31.485 -3.915 31.815 ;
        RECT -4.245 29.175 -3.915 29.505 ;
        RECT -4.245 28.325 -3.915 28.655 ;
        RECT -4.245 26.015 -3.915 26.345 ;
        RECT -4.245 25.165 -3.915 25.495 ;
        RECT -4.245 22.855 -3.915 23.185 ;
        RECT -4.245 22.005 -3.915 22.335 ;
        RECT -4.245 19.695 -3.915 20.025 ;
        RECT -4.245 18.115 -3.915 18.445 ;
        RECT -4.245 17.265 -3.915 17.595 ;
        RECT -4.245 14.955 -3.915 15.285 ;
        RECT -4.245 14.105 -3.915 14.435 ;
        RECT -4.245 11.795 -3.915 12.125 ;
        RECT -4.245 10.945 -3.915 11.275 ;
        RECT -4.245 8.635 -3.915 8.965 ;
        RECT -4.245 7.785 -3.915 8.115 ;
        RECT -4.245 5.475 -3.915 5.805 ;
        RECT -4.245 3.895 -3.915 4.225 ;
        RECT -4.245 3.045 -3.915 3.375 ;
        RECT -4.245 0.87 -3.915 1.2 ;
        RECT -4.245 -0.845 -3.915 -0.515 ;
        RECT -4.245 -2.205 -3.915 -1.875 ;
        RECT -4.245 -3.565 -3.915 -3.235 ;
        RECT -4.245 -4.925 -3.915 -4.595 ;
        RECT -4.245 -6.285 -3.915 -5.955 ;
        RECT -4.245 -7.645 -3.915 -7.315 ;
        RECT -4.245 -9.005 -3.915 -8.675 ;
        RECT -4.245 -10.365 -3.915 -10.035 ;
        RECT -4.245 -11.725 -3.915 -11.395 ;
        RECT -4.245 -13.085 -3.915 -12.755 ;
        RECT -4.245 -14.445 -3.915 -14.115 ;
        RECT -4.245 -15.805 -3.915 -15.475 ;
        RECT -4.245 -17.165 -3.915 -16.835 ;
        RECT -4.245 -21.245 -3.915 -20.915 ;
        RECT -4.245 -22.605 -3.915 -22.275 ;
        RECT -4.245 -23.965 -3.915 -23.635 ;
        RECT -4.245 -25.325 -3.915 -24.995 ;
        RECT -4.245 -26.685 -3.915 -26.355 ;
        RECT -4.245 -28.045 -3.915 -27.715 ;
        RECT -4.245 -29.405 -3.915 -29.075 ;
        RECT -4.245 -30.765 -3.915 -30.435 ;
        RECT -4.245 -32.125 -3.915 -31.795 ;
        RECT -4.245 -33.485 -3.915 -33.155 ;
        RECT -4.245 -36.205 -3.915 -35.875 ;
        RECT -4.245 -37.565 -3.915 -37.235 ;
        RECT -4.245 -38.925 -3.915 -38.595 ;
        RECT -4.245 -40.285 -3.915 -39.955 ;
        RECT -4.245 -43.005 -3.915 -42.675 ;
        RECT -4.245 -45.725 -3.915 -45.395 ;
        RECT -4.245 -47.085 -3.915 -46.755 ;
        RECT -4.245 -48.445 -3.915 -48.115 ;
        RECT -4.245 -49.805 -3.915 -49.475 ;
        RECT -4.245 -51.165 -3.915 -50.835 ;
        RECT -4.245 -52.525 -3.915 -52.195 ;
        RECT -4.245 -53.885 -3.915 -53.555 ;
        RECT -4.245 -55.245 -3.915 -54.915 ;
        RECT -4.245 -56.605 -3.915 -56.275 ;
        RECT -4.245 -57.965 -3.915 -57.635 ;
        RECT -4.245 -59.325 -3.915 -58.995 ;
        RECT -4.245 -60.685 -3.915 -60.355 ;
        RECT -4.245 -62.045 -3.915 -61.715 ;
        RECT -4.245 -63.405 -3.915 -63.075 ;
        RECT -4.245 -64.765 -3.915 -64.435 ;
        RECT -4.245 -66.125 -3.915 -65.795 ;
        RECT -4.245 -67.485 -3.915 -67.155 ;
        RECT -4.245 -68.845 -3.915 -68.515 ;
        RECT -4.245 -70.205 -3.915 -69.875 ;
        RECT -4.245 -71.565 -3.915 -71.235 ;
        RECT -4.245 -72.925 -3.915 -72.595 ;
        RECT -4.245 -74.285 -3.915 -73.955 ;
        RECT -4.245 -75.645 -3.915 -75.315 ;
        RECT -4.245 -77.005 -3.915 -76.675 ;
        RECT -4.245 -78.365 -3.915 -78.035 ;
        RECT -4.245 -79.725 -3.915 -79.395 ;
        RECT -4.245 -81.085 -3.915 -80.755 ;
        RECT -4.245 -82.445 -3.915 -82.115 ;
        RECT -4.245 -83.805 -3.915 -83.475 ;
        RECT -4.245 -85.165 -3.915 -84.835 ;
        RECT -4.245 -87.885 -3.915 -87.555 ;
        RECT -4.245 -89.245 -3.915 -88.915 ;
        RECT -4.245 -90.605 -3.915 -90.275 ;
        RECT -4.245 -91.965 -3.915 -91.635 ;
        RECT -4.245 -93.325 -3.915 -92.995 ;
        RECT -4.245 -94.685 -3.915 -94.355 ;
        RECT -4.245 -96.045 -3.915 -95.715 ;
        RECT -4.245 -97.405 -3.915 -97.075 ;
        RECT -4.245 -98.765 -3.915 -98.435 ;
        RECT -4.245 -100.125 -3.915 -99.795 ;
        RECT -4.245 -101.485 -3.915 -101.155 ;
        RECT -4.245 -102.845 -3.915 -102.515 ;
        RECT -4.245 -104.205 -3.915 -103.875 ;
        RECT -4.245 -105.565 -3.915 -105.235 ;
        RECT -4.245 -106.925 -3.915 -106.595 ;
        RECT -4.245 -108.285 -3.915 -107.955 ;
        RECT -4.245 -109.645 -3.915 -109.315 ;
        RECT -4.245 -111.005 -3.915 -110.675 ;
        RECT -4.245 -112.365 -3.915 -112.035 ;
        RECT -4.245 -113.725 -3.915 -113.395 ;
        RECT -4.245 -115.085 -3.915 -114.755 ;
        RECT -4.245 -116.445 -3.915 -116.115 ;
        RECT -4.245 -117.805 -3.915 -117.475 ;
        RECT -4.245 -119.165 -3.915 -118.835 ;
        RECT -4.245 -120.525 -3.915 -120.195 ;
        RECT -4.245 -121.885 -3.915 -121.555 ;
        RECT -4.245 -123.245 -3.915 -122.915 ;
        RECT -4.245 -124.605 -3.915 -124.275 ;
        RECT -4.245 -125.965 -3.915 -125.635 ;
        RECT -4.245 -127.325 -3.915 -126.995 ;
        RECT -4.245 -128.685 -3.915 -128.355 ;
        RECT -4.245 -130.045 -3.915 -129.715 ;
        RECT -4.245 -131.405 -3.915 -131.075 ;
        RECT -4.245 -132.765 -3.915 -132.435 ;
        RECT -4.245 -134.125 -3.915 -133.795 ;
        RECT -4.245 -135.485 -3.915 -135.155 ;
        RECT -4.245 -136.845 -3.915 -136.515 ;
        RECT -4.245 -138.205 -3.915 -137.875 ;
        RECT -4.245 -139.565 -3.915 -139.235 ;
        RECT -4.245 -140.925 -3.915 -140.595 ;
        RECT -4.245 -142.285 -3.915 -141.955 ;
        RECT -4.245 -143.645 -3.915 -143.315 ;
        RECT -4.245 -145.005 -3.915 -144.675 ;
        RECT -4.245 -146.365 -3.915 -146.035 ;
        RECT -4.245 -147.725 -3.915 -147.395 ;
        RECT -4.245 -149.085 -3.915 -148.755 ;
        RECT -4.245 -150.445 -3.915 -150.115 ;
        RECT -4.245 -151.805 -3.915 -151.475 ;
        RECT -4.245 -153.165 -3.915 -152.835 ;
        RECT -4.245 -158.81 -3.915 -157.68 ;
        RECT -4.24 -158.925 -3.92 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.885 44.8 -2.555 45.93 ;
        RECT -2.885 39.955 -2.555 40.285 ;
        RECT -2.885 38.595 -2.555 38.925 ;
        RECT -2.885 36.09 -2.555 36.42 ;
        RECT -2.885 33.915 -2.555 34.245 ;
        RECT -2.885 32.335 -2.555 32.665 ;
        RECT -2.885 31.485 -2.555 31.815 ;
        RECT -2.885 29.175 -2.555 29.505 ;
        RECT -2.885 28.325 -2.555 28.655 ;
        RECT -2.885 26.015 -2.555 26.345 ;
        RECT -2.885 25.165 -2.555 25.495 ;
        RECT -2.885 22.855 -2.555 23.185 ;
        RECT -2.885 22.005 -2.555 22.335 ;
        RECT -2.885 19.695 -2.555 20.025 ;
        RECT -2.885 18.115 -2.555 18.445 ;
        RECT -2.885 17.265 -2.555 17.595 ;
        RECT -2.885 14.955 -2.555 15.285 ;
        RECT -2.885 14.105 -2.555 14.435 ;
        RECT -2.885 11.795 -2.555 12.125 ;
        RECT -2.885 10.945 -2.555 11.275 ;
        RECT -2.885 8.635 -2.555 8.965 ;
        RECT -2.885 7.785 -2.555 8.115 ;
        RECT -2.885 5.475 -2.555 5.805 ;
        RECT -2.885 3.895 -2.555 4.225 ;
        RECT -2.885 3.045 -2.555 3.375 ;
        RECT -2.885 0.87 -2.555 1.2 ;
        RECT -2.885 -0.845 -2.555 -0.515 ;
        RECT -2.885 -2.205 -2.555 -1.875 ;
        RECT -2.885 -3.565 -2.555 -3.235 ;
        RECT -2.885 -4.925 -2.555 -4.595 ;
        RECT -2.885 -6.285 -2.555 -5.955 ;
        RECT -2.885 -7.645 -2.555 -7.315 ;
        RECT -2.885 -9.005 -2.555 -8.675 ;
        RECT -2.885 -10.365 -2.555 -10.035 ;
        RECT -2.885 -11.725 -2.555 -11.395 ;
        RECT -2.885 -13.085 -2.555 -12.755 ;
        RECT -2.885 -14.445 -2.555 -14.115 ;
        RECT -2.885 -15.805 -2.555 -15.475 ;
        RECT -2.885 -17.165 -2.555 -16.835 ;
        RECT -2.885 -21.245 -2.555 -20.915 ;
        RECT -2.885 -22.605 -2.555 -22.275 ;
        RECT -2.885 -23.965 -2.555 -23.635 ;
        RECT -2.885 -25.325 -2.555 -24.995 ;
        RECT -2.885 -26.685 -2.555 -26.355 ;
        RECT -2.885 -28.045 -2.555 -27.715 ;
        RECT -2.885 -29.405 -2.555 -29.075 ;
        RECT -2.885 -30.765 -2.555 -30.435 ;
        RECT -2.885 -32.125 -2.555 -31.795 ;
        RECT -2.885 -33.485 -2.555 -33.155 ;
        RECT -2.885 -36.205 -2.555 -35.875 ;
        RECT -2.885 -37.565 -2.555 -37.235 ;
        RECT -2.885 -38.925 -2.555 -38.595 ;
        RECT -2.885 -40.285 -2.555 -39.955 ;
        RECT -2.885 -43.005 -2.555 -42.675 ;
        RECT -2.885 -45.725 -2.555 -45.395 ;
        RECT -2.885 -47.085 -2.555 -46.755 ;
        RECT -2.885 -48.445 -2.555 -48.115 ;
        RECT -2.885 -49.805 -2.555 -49.475 ;
        RECT -2.885 -51.165 -2.555 -50.835 ;
        RECT -2.885 -52.525 -2.555 -52.195 ;
        RECT -2.885 -53.885 -2.555 -53.555 ;
        RECT -2.885 -55.245 -2.555 -54.915 ;
        RECT -2.885 -56.605 -2.555 -56.275 ;
        RECT -2.885 -57.965 -2.555 -57.635 ;
        RECT -2.885 -59.325 -2.555 -58.995 ;
        RECT -2.885 -60.685 -2.555 -60.355 ;
        RECT -2.885 -62.045 -2.555 -61.715 ;
        RECT -2.885 -63.405 -2.555 -63.075 ;
        RECT -2.885 -64.765 -2.555 -64.435 ;
        RECT -2.885 -66.125 -2.555 -65.795 ;
        RECT -2.885 -67.485 -2.555 -67.155 ;
        RECT -2.885 -68.845 -2.555 -68.515 ;
        RECT -2.885 -70.205 -2.555 -69.875 ;
        RECT -2.885 -71.565 -2.555 -71.235 ;
        RECT -2.885 -72.925 -2.555 -72.595 ;
        RECT -2.885 -74.285 -2.555 -73.955 ;
        RECT -2.885 -75.645 -2.555 -75.315 ;
        RECT -2.885 -77.005 -2.555 -76.675 ;
        RECT -2.885 -78.365 -2.555 -78.035 ;
        RECT -2.885 -79.725 -2.555 -79.395 ;
        RECT -2.885 -81.085 -2.555 -80.755 ;
        RECT -2.885 -82.445 -2.555 -82.115 ;
        RECT -2.885 -83.805 -2.555 -83.475 ;
        RECT -2.885 -85.165 -2.555 -84.835 ;
        RECT -2.885 -87.885 -2.555 -87.555 ;
        RECT -2.885 -89.245 -2.555 -88.915 ;
        RECT -2.885 -90.605 -2.555 -90.275 ;
        RECT -2.885 -91.965 -2.555 -91.635 ;
        RECT -2.885 -93.325 -2.555 -92.995 ;
        RECT -2.885 -94.685 -2.555 -94.355 ;
        RECT -2.885 -96.045 -2.555 -95.715 ;
        RECT -2.885 -97.405 -2.555 -97.075 ;
        RECT -2.885 -98.765 -2.555 -98.435 ;
        RECT -2.885 -100.125 -2.555 -99.795 ;
        RECT -2.885 -101.485 -2.555 -101.155 ;
        RECT -2.885 -102.845 -2.555 -102.515 ;
        RECT -2.885 -104.205 -2.555 -103.875 ;
        RECT -2.885 -105.565 -2.555 -105.235 ;
        RECT -2.885 -106.925 -2.555 -106.595 ;
        RECT -2.885 -108.285 -2.555 -107.955 ;
        RECT -2.885 -109.645 -2.555 -109.315 ;
        RECT -2.885 -111.005 -2.555 -110.675 ;
        RECT -2.885 -112.365 -2.555 -112.035 ;
        RECT -2.885 -113.725 -2.555 -113.395 ;
        RECT -2.885 -115.085 -2.555 -114.755 ;
        RECT -2.885 -116.445 -2.555 -116.115 ;
        RECT -2.885 -117.805 -2.555 -117.475 ;
        RECT -2.885 -119.165 -2.555 -118.835 ;
        RECT -2.885 -120.525 -2.555 -120.195 ;
        RECT -2.885 -121.885 -2.555 -121.555 ;
        RECT -2.885 -123.245 -2.555 -122.915 ;
        RECT -2.885 -124.605 -2.555 -124.275 ;
        RECT -2.885 -125.965 -2.555 -125.635 ;
        RECT -2.885 -127.325 -2.555 -126.995 ;
        RECT -2.885 -128.685 -2.555 -128.355 ;
        RECT -2.885 -130.045 -2.555 -129.715 ;
        RECT -2.885 -131.405 -2.555 -131.075 ;
        RECT -2.885 -132.765 -2.555 -132.435 ;
        RECT -2.885 -134.125 -2.555 -133.795 ;
        RECT -2.885 -135.485 -2.555 -135.155 ;
        RECT -2.885 -136.845 -2.555 -136.515 ;
        RECT -2.885 -138.205 -2.555 -137.875 ;
        RECT -2.885 -139.565 -2.555 -139.235 ;
        RECT -2.885 -140.925 -2.555 -140.595 ;
        RECT -2.885 -142.285 -2.555 -141.955 ;
        RECT -2.885 -143.645 -2.555 -143.315 ;
        RECT -2.885 -145.005 -2.555 -144.675 ;
        RECT -2.885 -146.365 -2.555 -146.035 ;
        RECT -2.885 -147.725 -2.555 -147.395 ;
        RECT -2.885 -149.085 -2.555 -148.755 ;
        RECT -2.885 -150.445 -2.555 -150.115 ;
        RECT -2.885 -151.805 -2.555 -151.475 ;
        RECT -2.885 -153.165 -2.555 -152.835 ;
        RECT -2.885 -158.81 -2.555 -157.68 ;
        RECT -2.88 -158.925 -2.56 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 44.8 -1.195 45.93 ;
        RECT -1.525 39.955 -1.195 40.285 ;
        RECT -1.525 38.595 -1.195 38.925 ;
        RECT -1.525 36.09 -1.195 36.42 ;
        RECT -1.525 33.915 -1.195 34.245 ;
        RECT -1.525 32.335 -1.195 32.665 ;
        RECT -1.525 31.485 -1.195 31.815 ;
        RECT -1.525 29.175 -1.195 29.505 ;
        RECT -1.525 28.325 -1.195 28.655 ;
        RECT -1.525 26.015 -1.195 26.345 ;
        RECT -1.525 25.165 -1.195 25.495 ;
        RECT -1.525 22.855 -1.195 23.185 ;
        RECT -1.525 22.005 -1.195 22.335 ;
        RECT -1.525 19.695 -1.195 20.025 ;
        RECT -1.525 18.115 -1.195 18.445 ;
        RECT -1.525 17.265 -1.195 17.595 ;
        RECT -1.525 14.955 -1.195 15.285 ;
        RECT -1.525 14.105 -1.195 14.435 ;
        RECT -1.525 11.795 -1.195 12.125 ;
        RECT -1.525 10.945 -1.195 11.275 ;
        RECT -1.525 8.635 -1.195 8.965 ;
        RECT -1.525 7.785 -1.195 8.115 ;
        RECT -1.525 5.475 -1.195 5.805 ;
        RECT -1.525 3.895 -1.195 4.225 ;
        RECT -1.525 3.045 -1.195 3.375 ;
        RECT -1.525 0.87 -1.195 1.2 ;
        RECT -1.525 -0.845 -1.195 -0.515 ;
        RECT -1.525 -2.205 -1.195 -1.875 ;
        RECT -1.525 -3.565 -1.195 -3.235 ;
        RECT -1.525 -4.925 -1.195 -4.595 ;
        RECT -1.525 -6.285 -1.195 -5.955 ;
        RECT -1.525 -7.645 -1.195 -7.315 ;
        RECT -1.525 -9.005 -1.195 -8.675 ;
        RECT -1.525 -10.365 -1.195 -10.035 ;
        RECT -1.525 -11.725 -1.195 -11.395 ;
        RECT -1.525 -13.085 -1.195 -12.755 ;
        RECT -1.525 -14.445 -1.195 -14.115 ;
        RECT -1.525 -15.805 -1.195 -15.475 ;
        RECT -1.525 -17.165 -1.195 -16.835 ;
        RECT -1.525 -21.245 -1.195 -20.915 ;
        RECT -1.525 -22.605 -1.195 -22.275 ;
        RECT -1.525 -23.965 -1.195 -23.635 ;
        RECT -1.525 -25.325 -1.195 -24.995 ;
        RECT -1.525 -26.685 -1.195 -26.355 ;
        RECT -1.525 -28.045 -1.195 -27.715 ;
        RECT -1.525 -29.405 -1.195 -29.075 ;
        RECT -1.525 -30.765 -1.195 -30.435 ;
        RECT -1.525 -32.125 -1.195 -31.795 ;
        RECT -1.525 -33.485 -1.195 -33.155 ;
        RECT -1.525 -36.205 -1.195 -35.875 ;
        RECT -1.525 -37.565 -1.195 -37.235 ;
        RECT -1.525 -38.925 -1.195 -38.595 ;
        RECT -1.525 -40.285 -1.195 -39.955 ;
        RECT -1.525 -43.005 -1.195 -42.675 ;
        RECT -1.525 -45.725 -1.195 -45.395 ;
        RECT -1.525 -47.085 -1.195 -46.755 ;
        RECT -1.525 -48.445 -1.195 -48.115 ;
        RECT -1.525 -49.805 -1.195 -49.475 ;
        RECT -1.525 -51.165 -1.195 -50.835 ;
        RECT -1.525 -52.525 -1.195 -52.195 ;
        RECT -1.525 -53.885 -1.195 -53.555 ;
        RECT -1.525 -55.245 -1.195 -54.915 ;
        RECT -1.525 -56.605 -1.195 -56.275 ;
        RECT -1.525 -57.965 -1.195 -57.635 ;
        RECT -1.525 -59.325 -1.195 -58.995 ;
        RECT -1.525 -60.685 -1.195 -60.355 ;
        RECT -1.525 -62.045 -1.195 -61.715 ;
        RECT -1.525 -63.405 -1.195 -63.075 ;
        RECT -1.525 -64.765 -1.195 -64.435 ;
        RECT -1.525 -66.125 -1.195 -65.795 ;
        RECT -1.525 -67.485 -1.195 -67.155 ;
        RECT -1.525 -68.845 -1.195 -68.515 ;
        RECT -1.525 -70.205 -1.195 -69.875 ;
        RECT -1.525 -71.565 -1.195 -71.235 ;
        RECT -1.525 -72.925 -1.195 -72.595 ;
        RECT -1.525 -74.285 -1.195 -73.955 ;
        RECT -1.525 -75.645 -1.195 -75.315 ;
        RECT -1.525 -77.005 -1.195 -76.675 ;
        RECT -1.525 -78.365 -1.195 -78.035 ;
        RECT -1.525 -79.725 -1.195 -79.395 ;
        RECT -1.525 -81.085 -1.195 -80.755 ;
        RECT -1.525 -82.445 -1.195 -82.115 ;
        RECT -1.525 -83.805 -1.195 -83.475 ;
        RECT -1.525 -85.165 -1.195 -84.835 ;
        RECT -1.525 -87.885 -1.195 -87.555 ;
        RECT -1.525 -89.245 -1.195 -88.915 ;
        RECT -1.525 -90.605 -1.195 -90.275 ;
        RECT -1.525 -91.965 -1.195 -91.635 ;
        RECT -1.525 -93.325 -1.195 -92.995 ;
        RECT -1.525 -94.685 -1.195 -94.355 ;
        RECT -1.525 -96.045 -1.195 -95.715 ;
        RECT -1.525 -97.405 -1.195 -97.075 ;
        RECT -1.525 -98.765 -1.195 -98.435 ;
        RECT -1.525 -100.125 -1.195 -99.795 ;
        RECT -1.525 -101.485 -1.195 -101.155 ;
        RECT -1.525 -102.845 -1.195 -102.515 ;
        RECT -1.525 -104.205 -1.195 -103.875 ;
        RECT -1.525 -105.565 -1.195 -105.235 ;
        RECT -1.525 -106.925 -1.195 -106.595 ;
        RECT -1.525 -108.285 -1.195 -107.955 ;
        RECT -1.525 -109.645 -1.195 -109.315 ;
        RECT -1.525 -111.005 -1.195 -110.675 ;
        RECT -1.525 -112.365 -1.195 -112.035 ;
        RECT -1.525 -113.725 -1.195 -113.395 ;
        RECT -1.525 -115.085 -1.195 -114.755 ;
        RECT -1.525 -116.445 -1.195 -116.115 ;
        RECT -1.525 -117.805 -1.195 -117.475 ;
        RECT -1.525 -119.165 -1.195 -118.835 ;
        RECT -1.525 -120.525 -1.195 -120.195 ;
        RECT -1.525 -121.885 -1.195 -121.555 ;
        RECT -1.525 -123.245 -1.195 -122.915 ;
        RECT -1.525 -124.605 -1.195 -124.275 ;
        RECT -1.525 -125.965 -1.195 -125.635 ;
        RECT -1.525 -127.325 -1.195 -126.995 ;
        RECT -1.525 -128.685 -1.195 -128.355 ;
        RECT -1.525 -130.045 -1.195 -129.715 ;
        RECT -1.525 -131.405 -1.195 -131.075 ;
        RECT -1.525 -132.765 -1.195 -132.435 ;
        RECT -1.525 -134.125 -1.195 -133.795 ;
        RECT -1.525 -135.485 -1.195 -135.155 ;
        RECT -1.525 -136.845 -1.195 -136.515 ;
        RECT -1.525 -138.205 -1.195 -137.875 ;
        RECT -1.525 -139.565 -1.195 -139.235 ;
        RECT -1.525 -140.925 -1.195 -140.595 ;
        RECT -1.525 -142.285 -1.195 -141.955 ;
        RECT -1.525 -143.645 -1.195 -143.315 ;
        RECT -1.525 -145.005 -1.195 -144.675 ;
        RECT -1.525 -146.365 -1.195 -146.035 ;
        RECT -1.525 -147.725 -1.195 -147.395 ;
        RECT -1.525 -149.085 -1.195 -148.755 ;
        RECT -1.525 -150.445 -1.195 -150.115 ;
        RECT -1.525 -151.805 -1.195 -151.475 ;
        RECT -1.525 -153.165 -1.195 -152.835 ;
        RECT -1.525 -158.81 -1.195 -157.68 ;
        RECT -1.52 -158.925 -1.2 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 44.8 0.165 45.93 ;
        RECT -0.165 39.955 0.165 40.285 ;
        RECT -0.165 38.595 0.165 38.925 ;
        RECT -0.16 37.92 0.16 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 -0.845 0.165 -0.515 ;
        RECT -0.165 -2.205 0.165 -1.875 ;
        RECT -0.165 -3.565 0.165 -3.235 ;
        RECT -0.16 -3.565 0.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 -91.965 0.165 -91.635 ;
        RECT -0.165 -93.325 0.165 -92.995 ;
        RECT -0.165 -94.685 0.165 -94.355 ;
        RECT -0.165 -96.045 0.165 -95.715 ;
        RECT -0.165 -97.405 0.165 -97.075 ;
        RECT -0.165 -98.765 0.165 -98.435 ;
        RECT -0.165 -100.125 0.165 -99.795 ;
        RECT -0.165 -101.485 0.165 -101.155 ;
        RECT -0.165 -102.845 0.165 -102.515 ;
        RECT -0.165 -104.205 0.165 -103.875 ;
        RECT -0.165 -105.565 0.165 -105.235 ;
        RECT -0.165 -106.925 0.165 -106.595 ;
        RECT -0.165 -108.285 0.165 -107.955 ;
        RECT -0.165 -109.645 0.165 -109.315 ;
        RECT -0.165 -111.005 0.165 -110.675 ;
        RECT -0.165 -112.365 0.165 -112.035 ;
        RECT -0.165 -113.725 0.165 -113.395 ;
        RECT -0.165 -115.085 0.165 -114.755 ;
        RECT -0.165 -116.445 0.165 -116.115 ;
        RECT -0.165 -117.805 0.165 -117.475 ;
        RECT -0.165 -119.165 0.165 -118.835 ;
        RECT -0.165 -120.525 0.165 -120.195 ;
        RECT -0.165 -121.885 0.165 -121.555 ;
        RECT -0.165 -123.245 0.165 -122.915 ;
        RECT -0.165 -124.605 0.165 -124.275 ;
        RECT -0.165 -125.965 0.165 -125.635 ;
        RECT -0.165 -127.325 0.165 -126.995 ;
        RECT -0.165 -128.685 0.165 -128.355 ;
        RECT -0.165 -130.045 0.165 -129.715 ;
        RECT -0.165 -131.405 0.165 -131.075 ;
        RECT -0.165 -132.765 0.165 -132.435 ;
        RECT -0.165 -134.125 0.165 -133.795 ;
        RECT -0.165 -135.485 0.165 -135.155 ;
        RECT -0.165 -136.845 0.165 -136.515 ;
        RECT -0.165 -138.205 0.165 -137.875 ;
        RECT -0.165 -139.565 0.165 -139.235 ;
        RECT -0.165 -140.925 0.165 -140.595 ;
        RECT -0.165 -142.285 0.165 -141.955 ;
        RECT -0.165 -143.645 0.165 -143.315 ;
        RECT -0.165 -145.005 0.165 -144.675 ;
        RECT -0.165 -146.365 0.165 -146.035 ;
        RECT -0.165 -147.725 0.165 -147.395 ;
        RECT -0.165 -149.085 0.165 -148.755 ;
        RECT -0.165 -150.445 0.165 -150.115 ;
        RECT -0.165 -151.805 0.165 -151.475 ;
        RECT -0.165 -153.165 0.165 -152.835 ;
        RECT -0.165 -158.81 0.165 -157.68 ;
        RECT -0.16 -158.925 0.16 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 44.8 1.525 45.93 ;
        RECT 1.195 39.955 1.525 40.285 ;
        RECT 1.195 38.595 1.525 38.925 ;
        RECT 1.2 37.92 1.52 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 -0.845 1.525 -0.515 ;
        RECT 1.195 -2.205 1.525 -1.875 ;
        RECT 1.195 -3.565 1.525 -3.235 ;
        RECT 1.2 -3.565 1.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 -91.965 1.525 -91.635 ;
        RECT 1.195 -93.325 1.525 -92.995 ;
        RECT 1.195 -94.685 1.525 -94.355 ;
        RECT 1.195 -96.045 1.525 -95.715 ;
        RECT 1.195 -97.405 1.525 -97.075 ;
        RECT 1.195 -98.765 1.525 -98.435 ;
        RECT 1.195 -100.125 1.525 -99.795 ;
        RECT 1.195 -101.485 1.525 -101.155 ;
        RECT 1.195 -102.845 1.525 -102.515 ;
        RECT 1.195 -104.205 1.525 -103.875 ;
        RECT 1.195 -105.565 1.525 -105.235 ;
        RECT 1.195 -106.925 1.525 -106.595 ;
        RECT 1.195 -108.285 1.525 -107.955 ;
        RECT 1.195 -109.645 1.525 -109.315 ;
        RECT 1.195 -111.005 1.525 -110.675 ;
        RECT 1.195 -112.365 1.525 -112.035 ;
        RECT 1.195 -113.725 1.525 -113.395 ;
        RECT 1.195 -115.085 1.525 -114.755 ;
        RECT 1.195 -116.445 1.525 -116.115 ;
        RECT 1.195 -117.805 1.525 -117.475 ;
        RECT 1.195 -119.165 1.525 -118.835 ;
        RECT 1.195 -120.525 1.525 -120.195 ;
        RECT 1.195 -121.885 1.525 -121.555 ;
        RECT 1.195 -123.245 1.525 -122.915 ;
        RECT 1.195 -124.605 1.525 -124.275 ;
        RECT 1.195 -125.965 1.525 -125.635 ;
        RECT 1.195 -127.325 1.525 -126.995 ;
        RECT 1.195 -128.685 1.525 -128.355 ;
        RECT 1.195 -130.045 1.525 -129.715 ;
        RECT 1.195 -131.405 1.525 -131.075 ;
        RECT 1.195 -132.765 1.525 -132.435 ;
        RECT 1.195 -134.125 1.525 -133.795 ;
        RECT 1.195 -135.485 1.525 -135.155 ;
        RECT 1.195 -136.845 1.525 -136.515 ;
        RECT 1.195 -138.205 1.525 -137.875 ;
        RECT 1.195 -139.565 1.525 -139.235 ;
        RECT 1.195 -140.925 1.525 -140.595 ;
        RECT 1.195 -142.285 1.525 -141.955 ;
        RECT 1.195 -143.645 1.525 -143.315 ;
        RECT 1.195 -145.005 1.525 -144.675 ;
        RECT 1.195 -146.365 1.525 -146.035 ;
        RECT 1.195 -147.725 1.525 -147.395 ;
        RECT 1.195 -149.085 1.525 -148.755 ;
        RECT 1.195 -150.445 1.525 -150.115 ;
        RECT 1.195 -151.805 1.525 -151.475 ;
        RECT 1.195 -153.165 1.525 -152.835 ;
        RECT 1.195 -158.81 1.525 -157.68 ;
        RECT 1.2 -158.925 1.52 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 44.8 2.885 45.93 ;
        RECT 2.555 39.955 2.885 40.285 ;
        RECT 2.555 38.595 2.885 38.925 ;
        RECT 2.56 37.92 2.88 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 -96.045 2.885 -95.715 ;
        RECT 2.555 -97.405 2.885 -97.075 ;
        RECT 2.555 -98.765 2.885 -98.435 ;
        RECT 2.555 -100.125 2.885 -99.795 ;
        RECT 2.555 -101.485 2.885 -101.155 ;
        RECT 2.555 -102.845 2.885 -102.515 ;
        RECT 2.555 -104.205 2.885 -103.875 ;
        RECT 2.555 -105.565 2.885 -105.235 ;
        RECT 2.555 -106.925 2.885 -106.595 ;
        RECT 2.555 -108.285 2.885 -107.955 ;
        RECT 2.555 -109.645 2.885 -109.315 ;
        RECT 2.555 -111.005 2.885 -110.675 ;
        RECT 2.555 -112.365 2.885 -112.035 ;
        RECT 2.555 -113.725 2.885 -113.395 ;
        RECT 2.555 -115.085 2.885 -114.755 ;
        RECT 2.555 -116.445 2.885 -116.115 ;
        RECT 2.555 -117.805 2.885 -117.475 ;
        RECT 2.555 -119.165 2.885 -118.835 ;
        RECT 2.555 -120.525 2.885 -120.195 ;
        RECT 2.555 -121.885 2.885 -121.555 ;
        RECT 2.555 -123.245 2.885 -122.915 ;
        RECT 2.555 -124.605 2.885 -124.275 ;
        RECT 2.555 -125.965 2.885 -125.635 ;
        RECT 2.555 -127.325 2.885 -126.995 ;
        RECT 2.555 -128.685 2.885 -128.355 ;
        RECT 2.555 -130.045 2.885 -129.715 ;
        RECT 2.555 -131.405 2.885 -131.075 ;
        RECT 2.555 -132.765 2.885 -132.435 ;
        RECT 2.555 -134.125 2.885 -133.795 ;
        RECT 2.555 -135.485 2.885 -135.155 ;
        RECT 2.555 -136.845 2.885 -136.515 ;
        RECT 2.555 -138.205 2.885 -137.875 ;
        RECT 2.555 -139.565 2.885 -139.235 ;
        RECT 2.555 -140.925 2.885 -140.595 ;
        RECT 2.555 -142.285 2.885 -141.955 ;
        RECT 2.555 -143.645 2.885 -143.315 ;
        RECT 2.555 -145.005 2.885 -144.675 ;
        RECT 2.555 -146.365 2.885 -146.035 ;
        RECT 2.555 -147.725 2.885 -147.395 ;
        RECT 2.555 -149.085 2.885 -148.755 ;
        RECT 2.555 -150.445 2.885 -150.115 ;
        RECT 2.555 -151.805 2.885 -151.475 ;
        RECT 2.555 -153.165 2.885 -152.835 ;
        RECT 2.555 -158.81 2.885 -157.68 ;
        RECT 2.56 -158.925 2.88 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.66 -94.075 2.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.915 44.8 4.245 45.93 ;
        RECT 3.915 39.955 4.245 40.285 ;
        RECT 3.915 38.595 4.245 38.925 ;
        RECT 3.92 37.92 4.24 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 44.8 5.605 45.93 ;
        RECT 5.275 39.955 5.605 40.285 ;
        RECT 5.275 38.595 5.605 38.925 ;
        RECT 5.28 37.92 5.6 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 -0.845 5.605 -0.515 ;
        RECT 5.275 -2.205 5.605 -1.875 ;
        RECT 5.275 -3.565 5.605 -3.235 ;
        RECT 5.28 -3.565 5.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 44.8 6.965 45.93 ;
        RECT 6.635 39.955 6.965 40.285 ;
        RECT 6.635 38.595 6.965 38.925 ;
        RECT 6.64 37.92 6.96 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 -0.845 6.965 -0.515 ;
        RECT 6.635 -2.205 6.965 -1.875 ;
        RECT 6.635 -3.565 6.965 -3.235 ;
        RECT 6.64 -3.565 6.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 44.8 8.325 45.93 ;
        RECT 7.995 39.955 8.325 40.285 ;
        RECT 7.995 38.595 8.325 38.925 ;
        RECT 8 37.92 8.32 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 -0.845 8.325 -0.515 ;
        RECT 7.995 -2.205 8.325 -1.875 ;
        RECT 7.995 -3.565 8.325 -3.235 ;
        RECT 8 -3.565 8.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 -91.965 8.325 -91.635 ;
        RECT 7.995 -93.325 8.325 -92.995 ;
        RECT 7.995 -94.685 8.325 -94.355 ;
        RECT 7.995 -96.045 8.325 -95.715 ;
        RECT 7.995 -97.405 8.325 -97.075 ;
        RECT 7.995 -98.765 8.325 -98.435 ;
        RECT 7.995 -100.125 8.325 -99.795 ;
        RECT 7.995 -101.485 8.325 -101.155 ;
        RECT 7.995 -102.845 8.325 -102.515 ;
        RECT 7.995 -104.205 8.325 -103.875 ;
        RECT 7.995 -105.565 8.325 -105.235 ;
        RECT 7.995 -106.925 8.325 -106.595 ;
        RECT 7.995 -108.285 8.325 -107.955 ;
        RECT 7.995 -109.645 8.325 -109.315 ;
        RECT 7.995 -111.005 8.325 -110.675 ;
        RECT 7.995 -112.365 8.325 -112.035 ;
        RECT 7.995 -113.725 8.325 -113.395 ;
        RECT 7.995 -115.085 8.325 -114.755 ;
        RECT 7.995 -116.445 8.325 -116.115 ;
        RECT 7.995 -117.805 8.325 -117.475 ;
        RECT 7.995 -119.165 8.325 -118.835 ;
        RECT 7.995 -120.525 8.325 -120.195 ;
        RECT 7.995 -121.885 8.325 -121.555 ;
        RECT 7.995 -123.245 8.325 -122.915 ;
        RECT 7.995 -124.605 8.325 -124.275 ;
        RECT 7.995 -125.965 8.325 -125.635 ;
        RECT 7.995 -127.325 8.325 -126.995 ;
        RECT 7.995 -128.685 8.325 -128.355 ;
        RECT 7.995 -130.045 8.325 -129.715 ;
        RECT 7.995 -131.405 8.325 -131.075 ;
        RECT 7.995 -132.765 8.325 -132.435 ;
        RECT 7.995 -134.125 8.325 -133.795 ;
        RECT 7.995 -135.485 8.325 -135.155 ;
        RECT 7.995 -136.845 8.325 -136.515 ;
        RECT 7.995 -138.205 8.325 -137.875 ;
        RECT 7.995 -139.565 8.325 -139.235 ;
        RECT 7.995 -140.925 8.325 -140.595 ;
        RECT 7.995 -142.285 8.325 -141.955 ;
        RECT 7.995 -143.645 8.325 -143.315 ;
        RECT 7.995 -145.005 8.325 -144.675 ;
        RECT 7.995 -146.365 8.325 -146.035 ;
        RECT 7.995 -147.725 8.325 -147.395 ;
        RECT 7.995 -149.085 8.325 -148.755 ;
        RECT 7.995 -150.445 8.325 -150.115 ;
        RECT 7.995 -151.805 8.325 -151.475 ;
        RECT 7.995 -153.165 8.325 -152.835 ;
        RECT 7.995 -158.81 8.325 -157.68 ;
        RECT 8 -158.925 8.32 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.76 -94.075 9.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 44.8 9.685 45.93 ;
        RECT 9.355 39.955 9.685 40.285 ;
        RECT 9.355 38.595 9.685 38.925 ;
        RECT 9.36 37.92 9.68 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 -96.045 9.685 -95.715 ;
        RECT 9.355 -97.405 9.685 -97.075 ;
        RECT 9.355 -98.765 9.685 -98.435 ;
        RECT 9.355 -100.125 9.685 -99.795 ;
        RECT 9.355 -101.485 9.685 -101.155 ;
        RECT 9.355 -102.845 9.685 -102.515 ;
        RECT 9.355 -104.205 9.685 -103.875 ;
        RECT 9.355 -105.565 9.685 -105.235 ;
        RECT 9.355 -106.925 9.685 -106.595 ;
        RECT 9.355 -108.285 9.685 -107.955 ;
        RECT 9.355 -109.645 9.685 -109.315 ;
        RECT 9.355 -111.005 9.685 -110.675 ;
        RECT 9.355 -112.365 9.685 -112.035 ;
        RECT 9.355 -113.725 9.685 -113.395 ;
        RECT 9.355 -115.085 9.685 -114.755 ;
        RECT 9.355 -116.445 9.685 -116.115 ;
        RECT 9.355 -117.805 9.685 -117.475 ;
        RECT 9.355 -119.165 9.685 -118.835 ;
        RECT 9.355 -120.525 9.685 -120.195 ;
        RECT 9.355 -121.885 9.685 -121.555 ;
        RECT 9.355 -123.245 9.685 -122.915 ;
        RECT 9.355 -124.605 9.685 -124.275 ;
        RECT 9.355 -125.965 9.685 -125.635 ;
        RECT 9.355 -127.325 9.685 -126.995 ;
        RECT 9.355 -128.685 9.685 -128.355 ;
        RECT 9.355 -130.045 9.685 -129.715 ;
        RECT 9.355 -131.405 9.685 -131.075 ;
        RECT 9.355 -132.765 9.685 -132.435 ;
        RECT 9.355 -134.125 9.685 -133.795 ;
        RECT 9.355 -135.485 9.685 -135.155 ;
        RECT 9.355 -136.845 9.685 -136.515 ;
        RECT 9.355 -138.205 9.685 -137.875 ;
        RECT 9.355 -139.565 9.685 -139.235 ;
        RECT 9.355 -140.925 9.685 -140.595 ;
        RECT 9.355 -142.285 9.685 -141.955 ;
        RECT 9.355 -143.645 9.685 -143.315 ;
        RECT 9.355 -145.005 9.685 -144.675 ;
        RECT 9.355 -146.365 9.685 -146.035 ;
        RECT 9.355 -147.725 9.685 -147.395 ;
        RECT 9.355 -149.085 9.685 -148.755 ;
        RECT 9.355 -150.445 9.685 -150.115 ;
        RECT 9.355 -151.805 9.685 -151.475 ;
        RECT 9.355 -153.165 9.685 -152.835 ;
        RECT 9.355 -158.81 9.685 -157.68 ;
        RECT 9.36 -158.925 9.68 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 44.8 11.045 45.93 ;
        RECT 10.715 39.955 11.045 40.285 ;
        RECT 10.715 38.595 11.045 38.925 ;
        RECT 10.72 37.92 11.04 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 -0.845 11.045 -0.515 ;
        RECT 10.715 -2.205 11.045 -1.875 ;
        RECT 10.715 -3.565 11.045 -3.235 ;
        RECT 10.72 -3.565 11.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 44.8 12.405 45.93 ;
        RECT 12.075 39.955 12.405 40.285 ;
        RECT 12.075 38.595 12.405 38.925 ;
        RECT 12.08 37.92 12.4 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 -0.845 12.405 -0.515 ;
        RECT 12.075 -2.205 12.405 -1.875 ;
        RECT 12.075 -3.565 12.405 -3.235 ;
        RECT 12.08 -3.565 12.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 44.8 13.765 45.93 ;
        RECT 13.435 39.955 13.765 40.285 ;
        RECT 13.435 38.595 13.765 38.925 ;
        RECT 13.44 37.92 13.76 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 -0.845 13.765 -0.515 ;
        RECT 13.435 -2.205 13.765 -1.875 ;
        RECT 13.435 -3.565 13.765 -3.235 ;
        RECT 13.44 -3.565 13.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 -91.965 13.765 -91.635 ;
        RECT 13.435 -93.325 13.765 -92.995 ;
        RECT 13.435 -94.685 13.765 -94.355 ;
        RECT 13.435 -96.045 13.765 -95.715 ;
        RECT 13.435 -97.405 13.765 -97.075 ;
        RECT 13.435 -98.765 13.765 -98.435 ;
        RECT 13.435 -100.125 13.765 -99.795 ;
        RECT 13.435 -101.485 13.765 -101.155 ;
        RECT 13.435 -102.845 13.765 -102.515 ;
        RECT 13.435 -104.205 13.765 -103.875 ;
        RECT 13.435 -105.565 13.765 -105.235 ;
        RECT 13.435 -106.925 13.765 -106.595 ;
        RECT 13.435 -108.285 13.765 -107.955 ;
        RECT 13.435 -109.645 13.765 -109.315 ;
        RECT 13.435 -111.005 13.765 -110.675 ;
        RECT 13.435 -112.365 13.765 -112.035 ;
        RECT 13.435 -113.725 13.765 -113.395 ;
        RECT 13.435 -115.085 13.765 -114.755 ;
        RECT 13.435 -116.445 13.765 -116.115 ;
        RECT 13.435 -117.805 13.765 -117.475 ;
        RECT 13.435 -119.165 13.765 -118.835 ;
        RECT 13.435 -120.525 13.765 -120.195 ;
        RECT 13.435 -121.885 13.765 -121.555 ;
        RECT 13.435 -123.245 13.765 -122.915 ;
        RECT 13.435 -124.605 13.765 -124.275 ;
        RECT 13.435 -125.965 13.765 -125.635 ;
        RECT 13.435 -127.325 13.765 -126.995 ;
        RECT 13.435 -128.685 13.765 -128.355 ;
        RECT 13.435 -130.045 13.765 -129.715 ;
        RECT 13.435 -131.405 13.765 -131.075 ;
        RECT 13.435 -132.765 13.765 -132.435 ;
        RECT 13.435 -134.125 13.765 -133.795 ;
        RECT 13.435 -135.485 13.765 -135.155 ;
        RECT 13.435 -136.845 13.765 -136.515 ;
        RECT 13.435 -138.205 13.765 -137.875 ;
        RECT 13.435 -139.565 13.765 -139.235 ;
        RECT 13.435 -140.925 13.765 -140.595 ;
        RECT 13.435 -142.285 13.765 -141.955 ;
        RECT 13.435 -143.645 13.765 -143.315 ;
        RECT 13.435 -145.005 13.765 -144.675 ;
        RECT 13.435 -146.365 13.765 -146.035 ;
        RECT 13.435 -147.725 13.765 -147.395 ;
        RECT 13.435 -149.085 13.765 -148.755 ;
        RECT 13.435 -150.445 13.765 -150.115 ;
        RECT 13.435 -151.805 13.765 -151.475 ;
        RECT 13.435 -153.165 13.765 -152.835 ;
        RECT 13.435 -158.81 13.765 -157.68 ;
        RECT 13.44 -158.925 13.76 -90.96 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 44.8 15.125 45.93 ;
        RECT 14.795 39.955 15.125 40.285 ;
        RECT 14.795 38.595 15.125 38.925 ;
        RECT 14.8 37.92 15.12 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 -96.045 15.125 -95.715 ;
        RECT 14.795 -97.405 15.125 -97.075 ;
        RECT 14.795 -98.765 15.125 -98.435 ;
        RECT 14.795 -100.125 15.125 -99.795 ;
        RECT 14.795 -101.485 15.125 -101.155 ;
        RECT 14.795 -102.845 15.125 -102.515 ;
        RECT 14.795 -104.205 15.125 -103.875 ;
        RECT 14.795 -105.565 15.125 -105.235 ;
        RECT 14.795 -106.925 15.125 -106.595 ;
        RECT 14.795 -108.285 15.125 -107.955 ;
        RECT 14.795 -109.645 15.125 -109.315 ;
        RECT 14.795 -111.005 15.125 -110.675 ;
        RECT 14.795 -112.365 15.125 -112.035 ;
        RECT 14.795 -113.725 15.125 -113.395 ;
        RECT 14.795 -115.085 15.125 -114.755 ;
        RECT 14.795 -116.445 15.125 -116.115 ;
        RECT 14.795 -117.805 15.125 -117.475 ;
        RECT 14.795 -119.165 15.125 -118.835 ;
        RECT 14.795 -120.525 15.125 -120.195 ;
        RECT 14.795 -121.885 15.125 -121.555 ;
        RECT 14.795 -123.245 15.125 -122.915 ;
        RECT 14.795 -124.605 15.125 -124.275 ;
        RECT 14.795 -125.965 15.125 -125.635 ;
        RECT 14.795 -127.325 15.125 -126.995 ;
        RECT 14.795 -128.685 15.125 -128.355 ;
        RECT 14.795 -130.045 15.125 -129.715 ;
        RECT 14.795 -131.405 15.125 -131.075 ;
        RECT 14.795 -132.765 15.125 -132.435 ;
        RECT 14.795 -134.125 15.125 -133.795 ;
        RECT 14.795 -135.485 15.125 -135.155 ;
        RECT 14.795 -136.845 15.125 -136.515 ;
        RECT 14.795 -138.205 15.125 -137.875 ;
        RECT 14.795 -139.565 15.125 -139.235 ;
        RECT 14.795 -140.925 15.125 -140.595 ;
        RECT 14.795 -142.285 15.125 -141.955 ;
        RECT 14.795 -143.645 15.125 -143.315 ;
        RECT 14.795 -145.005 15.125 -144.675 ;
        RECT 14.795 -146.365 15.125 -146.035 ;
        RECT 14.795 -147.725 15.125 -147.395 ;
        RECT 14.795 -149.085 15.125 -148.755 ;
        RECT 14.795 -150.445 15.125 -150.115 ;
        RECT 14.795 -151.805 15.125 -151.475 ;
        RECT 14.795 -153.165 15.125 -152.835 ;
        RECT 14.795 -158.81 15.125 -157.68 ;
        RECT 14.8 -158.925 15.12 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.86 -94.075 15.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.155 44.8 16.485 45.93 ;
        RECT 16.155 39.955 16.485 40.285 ;
        RECT 16.155 38.595 16.485 38.925 ;
        RECT 16.16 37.92 16.48 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 44.8 17.845 45.93 ;
        RECT 17.515 39.955 17.845 40.285 ;
        RECT 17.515 38.595 17.845 38.925 ;
        RECT 17.52 37.92 17.84 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 -0.845 17.845 -0.515 ;
        RECT 17.515 -2.205 17.845 -1.875 ;
        RECT 17.515 -3.565 17.845 -3.235 ;
        RECT 17.52 -3.565 17.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 44.8 19.205 45.93 ;
        RECT 18.875 39.955 19.205 40.285 ;
        RECT 18.875 38.595 19.205 38.925 ;
        RECT 18.88 37.92 19.2 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 -0.845 19.205 -0.515 ;
        RECT 18.875 -2.205 19.205 -1.875 ;
        RECT 18.875 -3.565 19.205 -3.235 ;
        RECT 18.88 -3.565 19.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 44.8 20.565 45.93 ;
        RECT 20.235 39.955 20.565 40.285 ;
        RECT 20.235 38.595 20.565 38.925 ;
        RECT 20.24 37.92 20.56 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 -0.845 20.565 -0.515 ;
        RECT 20.235 -2.205 20.565 -1.875 ;
        RECT 20.235 -3.565 20.565 -3.235 ;
        RECT 20.24 -3.565 20.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 -138.205 20.565 -137.875 ;
        RECT 20.235 -139.565 20.565 -139.235 ;
        RECT 20.235 -140.925 20.565 -140.595 ;
        RECT 20.235 -142.285 20.565 -141.955 ;
        RECT 20.235 -143.645 20.565 -143.315 ;
        RECT 20.235 -145.005 20.565 -144.675 ;
        RECT 20.235 -146.365 20.565 -146.035 ;
        RECT 20.235 -147.725 20.565 -147.395 ;
        RECT 20.235 -149.085 20.565 -148.755 ;
        RECT 20.235 -150.445 20.565 -150.115 ;
        RECT 20.235 -151.805 20.565 -151.475 ;
        RECT 20.235 -153.165 20.565 -152.835 ;
        RECT 20.235 -158.81 20.565 -157.68 ;
        RECT 20.24 -158.925 20.56 -90.96 ;
        RECT 20.235 -91.965 20.565 -91.635 ;
        RECT 20.235 -93.325 20.565 -92.995 ;
        RECT 20.235 -94.685 20.565 -94.355 ;
        RECT 20.235 -96.045 20.565 -95.715 ;
        RECT 20.235 -97.405 20.565 -97.075 ;
        RECT 20.235 -98.765 20.565 -98.435 ;
        RECT 20.235 -100.125 20.565 -99.795 ;
        RECT 20.235 -101.485 20.565 -101.155 ;
        RECT 20.235 -102.845 20.565 -102.515 ;
        RECT 20.235 -104.205 20.565 -103.875 ;
        RECT 20.235 -105.565 20.565 -105.235 ;
        RECT 20.235 -106.925 20.565 -106.595 ;
        RECT 20.235 -108.285 20.565 -107.955 ;
        RECT 20.235 -109.645 20.565 -109.315 ;
        RECT 20.235 -111.005 20.565 -110.675 ;
        RECT 20.235 -112.365 20.565 -112.035 ;
        RECT 20.235 -113.725 20.565 -113.395 ;
        RECT 20.235 -115.085 20.565 -114.755 ;
        RECT 20.235 -116.445 20.565 -116.115 ;
        RECT 20.235 -117.805 20.565 -117.475 ;
        RECT 20.235 -119.165 20.565 -118.835 ;
        RECT 20.235 -120.525 20.565 -120.195 ;
        RECT 20.235 -121.885 20.565 -121.555 ;
        RECT 20.235 -123.245 20.565 -122.915 ;
        RECT 20.235 -124.605 20.565 -124.275 ;
        RECT 20.235 -125.965 20.565 -125.635 ;
        RECT 20.235 -127.325 20.565 -126.995 ;
        RECT 20.235 -128.685 20.565 -128.355 ;
        RECT 20.235 -130.045 20.565 -129.715 ;
        RECT 20.235 -131.405 20.565 -131.075 ;
        RECT 20.235 -132.765 20.565 -132.435 ;
        RECT 20.235 -134.125 20.565 -133.795 ;
        RECT 20.235 -135.485 20.565 -135.155 ;
        RECT 20.235 -136.845 20.565 -136.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 -151.805 -20.235 -151.475 ;
        RECT -20.565 -153.165 -20.235 -152.835 ;
        RECT -20.565 -158.81 -20.235 -157.68 ;
        RECT -20.56 -158.925 -20.24 -147.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 44.8 -18.875 45.93 ;
        RECT -19.205 39.955 -18.875 40.285 ;
        RECT -19.205 38.595 -18.875 38.925 ;
        RECT -19.205 37.235 -18.875 37.565 ;
        RECT -19.205 35.875 -18.875 36.205 ;
        RECT -19.205 34.515 -18.875 34.845 ;
        RECT -19.205 33.155 -18.875 33.485 ;
        RECT -19.205 31.795 -18.875 32.125 ;
        RECT -19.205 30.435 -18.875 30.765 ;
        RECT -19.205 29.075 -18.875 29.405 ;
        RECT -19.205 27.715 -18.875 28.045 ;
        RECT -19.205 26.355 -18.875 26.685 ;
        RECT -19.205 24.995 -18.875 25.325 ;
        RECT -19.205 23.635 -18.875 23.965 ;
        RECT -19.205 22.275 -18.875 22.605 ;
        RECT -19.205 20.915 -18.875 21.245 ;
        RECT -19.205 19.555 -18.875 19.885 ;
        RECT -19.205 18.195 -18.875 18.525 ;
        RECT -19.205 16.835 -18.875 17.165 ;
        RECT -19.205 15.475 -18.875 15.805 ;
        RECT -19.205 14.115 -18.875 14.445 ;
        RECT -19.205 12.755 -18.875 13.085 ;
        RECT -19.205 11.395 -18.875 11.725 ;
        RECT -19.205 10.035 -18.875 10.365 ;
        RECT -19.205 8.675 -18.875 9.005 ;
        RECT -19.205 7.315 -18.875 7.645 ;
        RECT -19.205 5.955 -18.875 6.285 ;
        RECT -19.205 4.595 -18.875 4.925 ;
        RECT -19.205 3.235 -18.875 3.565 ;
        RECT -19.205 1.875 -18.875 2.205 ;
        RECT -19.205 -2.205 -18.875 -1.875 ;
        RECT -19.205 -4.925 -18.875 -4.595 ;
        RECT -19.205 -5.65 -18.875 -5.32 ;
        RECT -19.205 -7.645 -18.875 -7.315 ;
        RECT -19.205 -11.69 -18.875 -11.36 ;
        RECT -19.205 -13.085 -18.875 -12.755 ;
        RECT -19.205 -15.805 -18.875 -15.475 ;
        RECT -19.205 -25.325 -18.875 -24.995 ;
        RECT -19.205 -26.685 -18.875 -26.355 ;
        RECT -19.205 -27.67 -18.875 -27.34 ;
        RECT -19.205 -29.405 -18.875 -29.075 ;
        RECT -19.205 -30.765 -18.875 -30.435 ;
        RECT -19.2 -32.12 -18.88 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 -100.125 -18.875 -99.795 ;
        RECT -19.205 -101.485 -18.875 -101.155 ;
        RECT -19.205 -109.645 -18.875 -109.315 ;
        RECT -19.205 -113.725 -18.875 -113.395 ;
        RECT -19.205 -119.165 -18.875 -118.835 ;
        RECT -19.205 -120.525 -18.875 -120.195 ;
        RECT -19.205 -123.245 -18.875 -122.915 ;
        RECT -19.205 -125.965 -18.875 -125.635 ;
        RECT -19.205 -127.325 -18.875 -126.995 ;
        RECT -19.205 -132.765 -18.875 -132.435 ;
        RECT -19.205 -134.125 -18.875 -133.795 ;
        RECT -19.205 -135.485 -18.875 -135.155 ;
        RECT -19.205 -136.845 -18.875 -136.515 ;
        RECT -19.205 -138.205 -18.875 -137.875 ;
        RECT -19.205 -139.565 -18.875 -139.235 ;
        RECT -19.205 -140.925 -18.875 -140.595 ;
        RECT -19.205 -143.755 -18.875 -143.425 ;
        RECT -19.205 -145.005 -18.875 -144.675 ;
        RECT -19.205 -146.365 -18.875 -146.035 ;
        RECT -19.205 -147.725 -18.875 -147.395 ;
        RECT -19.205 -151.805 -18.875 -151.475 ;
        RECT -19.205 -153.165 -18.875 -152.835 ;
        RECT -19.205 -158.81 -18.875 -157.68 ;
        RECT -19.2 -158.925 -18.88 -96.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.845 44.8 -17.515 45.93 ;
        RECT -17.845 39.955 -17.515 40.285 ;
        RECT -17.845 38.595 -17.515 38.925 ;
        RECT -17.845 37.235 -17.515 37.565 ;
        RECT -17.845 35.875 -17.515 36.205 ;
        RECT -17.845 34.515 -17.515 34.845 ;
        RECT -17.845 33.155 -17.515 33.485 ;
        RECT -17.845 31.795 -17.515 32.125 ;
        RECT -17.845 30.435 -17.515 30.765 ;
        RECT -17.845 29.075 -17.515 29.405 ;
        RECT -17.845 27.715 -17.515 28.045 ;
        RECT -17.845 26.355 -17.515 26.685 ;
        RECT -17.845 24.995 -17.515 25.325 ;
        RECT -17.845 23.635 -17.515 23.965 ;
        RECT -17.845 22.275 -17.515 22.605 ;
        RECT -17.845 20.915 -17.515 21.245 ;
        RECT -17.845 19.555 -17.515 19.885 ;
        RECT -17.845 18.195 -17.515 18.525 ;
        RECT -17.845 16.835 -17.515 17.165 ;
        RECT -17.845 15.475 -17.515 15.805 ;
        RECT -17.845 14.115 -17.515 14.445 ;
        RECT -17.845 12.755 -17.515 13.085 ;
        RECT -17.845 11.395 -17.515 11.725 ;
        RECT -17.845 10.035 -17.515 10.365 ;
        RECT -17.845 8.675 -17.515 9.005 ;
        RECT -17.845 7.315 -17.515 7.645 ;
        RECT -17.845 5.955 -17.515 6.285 ;
        RECT -17.845 4.595 -17.515 4.925 ;
        RECT -17.845 3.235 -17.515 3.565 ;
        RECT -17.845 1.875 -17.515 2.205 ;
        RECT -17.845 -2.205 -17.515 -1.875 ;
        RECT -17.845 -4.925 -17.515 -4.595 ;
        RECT -17.845 -5.65 -17.515 -5.32 ;
        RECT -17.845 -7.645 -17.515 -7.315 ;
        RECT -17.845 -11.69 -17.515 -11.36 ;
        RECT -17.845 -13.085 -17.515 -12.755 ;
        RECT -17.845 -15.805 -17.515 -15.475 ;
        RECT -17.845 -22.605 -17.515 -22.275 ;
        RECT -17.845 -25.325 -17.515 -24.995 ;
        RECT -17.845 -26.685 -17.515 -26.355 ;
        RECT -17.845 -27.67 -17.515 -27.34 ;
        RECT -17.845 -29.405 -17.515 -29.075 ;
        RECT -17.845 -30.765 -17.515 -30.435 ;
        RECT -17.845 -33.71 -17.515 -33.38 ;
        RECT -17.845 -34.845 -17.515 -34.515 ;
        RECT -17.845 -37.565 -17.515 -37.235 ;
        RECT -17.845 -45.725 -17.515 -45.395 ;
        RECT -17.845 -47.085 -17.515 -46.755 ;
        RECT -17.845 -48.29 -17.515 -47.96 ;
        RECT -17.845 -49.805 -17.515 -49.475 ;
        RECT -17.845 -52.525 -17.515 -52.195 ;
        RECT -17.845 -53.885 -17.515 -53.555 ;
        RECT -17.845 -55.83 -17.515 -55.5 ;
        RECT -17.845 -56.605 -17.515 -56.275 ;
        RECT -17.845 -57.965 -17.515 -57.635 ;
        RECT -17.845 -59.325 -17.515 -58.995 ;
        RECT -17.845 -62.045 -17.515 -61.715 ;
        RECT -17.845 -64.765 -17.515 -64.435 ;
        RECT -17.845 -66.125 -17.515 -65.795 ;
        RECT -17.845 -67.485 -17.515 -67.155 ;
        RECT -17.845 -68.845 -17.515 -68.515 ;
        RECT -17.845 -70.47 -17.515 -70.14 ;
        RECT -17.845 -71.565 -17.515 -71.235 ;
        RECT -17.845 -72.925 -17.515 -72.595 ;
        RECT -17.845 -75.645 -17.515 -75.315 ;
        RECT -17.845 -77.005 -17.515 -76.675 ;
        RECT -17.845 -78.01 -17.515 -77.68 ;
        RECT -17.845 -79.725 -17.515 -79.395 ;
        RECT -17.845 -81.085 -17.515 -80.755 ;
        RECT -17.845 -89.245 -17.515 -88.915 ;
        RECT -17.845 -90.605 -17.515 -90.275 ;
        RECT -17.845 -91.965 -17.515 -91.635 ;
        RECT -17.845 -93.325 -17.515 -92.995 ;
        RECT -17.845 -96.045 -17.515 -95.715 ;
        RECT -17.845 -101.485 -17.515 -101.155 ;
        RECT -17.845 -113.725 -17.515 -113.395 ;
        RECT -17.845 -119.165 -17.515 -118.835 ;
        RECT -17.845 -120.525 -17.515 -120.195 ;
        RECT -17.845 -123.245 -17.515 -122.915 ;
        RECT -17.845 -125.965 -17.515 -125.635 ;
        RECT -17.845 -127.325 -17.515 -126.995 ;
        RECT -17.845 -131.405 -17.515 -131.075 ;
        RECT -17.845 -132.765 -17.515 -132.435 ;
        RECT -17.845 -134.125 -17.515 -133.795 ;
        RECT -17.845 -135.485 -17.515 -135.155 ;
        RECT -17.845 -136.845 -17.515 -136.515 ;
        RECT -17.845 -138.205 -17.515 -137.875 ;
        RECT -17.845 -139.565 -17.515 -139.235 ;
        RECT -17.845 -140.925 -17.515 -140.595 ;
        RECT -17.845 -143.755 -17.515 -143.425 ;
        RECT -17.845 -145.005 -17.515 -144.675 ;
        RECT -17.845 -146.365 -17.515 -146.035 ;
        RECT -17.845 -147.725 -17.515 -147.395 ;
        RECT -17.845 -151.805 -17.515 -151.475 ;
        RECT -17.845 -153.165 -17.515 -152.835 ;
        RECT -17.845 -158.81 -17.515 -157.68 ;
        RECT -17.84 -158.925 -17.52 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 44.8 -16.155 45.93 ;
        RECT -16.485 39.955 -16.155 40.285 ;
        RECT -16.485 38.595 -16.155 38.925 ;
        RECT -16.485 37.235 -16.155 37.565 ;
        RECT -16.485 35.875 -16.155 36.205 ;
        RECT -16.485 34.515 -16.155 34.845 ;
        RECT -16.485 33.155 -16.155 33.485 ;
        RECT -16.485 31.795 -16.155 32.125 ;
        RECT -16.485 30.435 -16.155 30.765 ;
        RECT -16.485 29.075 -16.155 29.405 ;
        RECT -16.485 27.715 -16.155 28.045 ;
        RECT -16.485 26.355 -16.155 26.685 ;
        RECT -16.485 24.995 -16.155 25.325 ;
        RECT -16.485 23.635 -16.155 23.965 ;
        RECT -16.485 22.275 -16.155 22.605 ;
        RECT -16.485 20.915 -16.155 21.245 ;
        RECT -16.485 19.555 -16.155 19.885 ;
        RECT -16.485 18.195 -16.155 18.525 ;
        RECT -16.485 16.835 -16.155 17.165 ;
        RECT -16.485 15.475 -16.155 15.805 ;
        RECT -16.485 14.115 -16.155 14.445 ;
        RECT -16.485 12.755 -16.155 13.085 ;
        RECT -16.485 11.395 -16.155 11.725 ;
        RECT -16.485 10.035 -16.155 10.365 ;
        RECT -16.485 8.675 -16.155 9.005 ;
        RECT -16.485 7.315 -16.155 7.645 ;
        RECT -16.485 5.955 -16.155 6.285 ;
        RECT -16.485 4.595 -16.155 4.925 ;
        RECT -16.485 3.235 -16.155 3.565 ;
        RECT -16.485 1.875 -16.155 2.205 ;
        RECT -16.485 0.515 -16.155 0.845 ;
        RECT -16.485 -2.205 -16.155 -1.875 ;
        RECT -16.485 -4.925 -16.155 -4.595 ;
        RECT -16.485 -5.65 -16.155 -5.32 ;
        RECT -16.485 -7.645 -16.155 -7.315 ;
        RECT -16.485 -11.69 -16.155 -11.36 ;
        RECT -16.485 -13.085 -16.155 -12.755 ;
        RECT -16.485 -15.805 -16.155 -15.475 ;
        RECT -16.48 -17.84 -16.16 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 -22.605 -16.155 -22.275 ;
        RECT -16.485 -25.325 -16.155 -24.995 ;
        RECT -16.485 -26.685 -16.155 -26.355 ;
        RECT -16.485 -27.67 -16.155 -27.34 ;
        RECT -16.485 -29.405 -16.155 -29.075 ;
        RECT -16.485 -30.765 -16.155 -30.435 ;
        RECT -16.485 -33.71 -16.155 -33.38 ;
        RECT -16.485 -34.845 -16.155 -34.515 ;
        RECT -16.485 -37.565 -16.155 -37.235 ;
        RECT -16.48 -39.6 -16.16 -22.275 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 -45.725 -16.155 -45.395 ;
        RECT -16.485 -47.085 -16.155 -46.755 ;
        RECT -16.485 -48.29 -16.155 -47.96 ;
        RECT -16.485 -49.805 -16.155 -49.475 ;
        RECT -16.485 -52.525 -16.155 -52.195 ;
        RECT -16.485 -53.885 -16.155 -53.555 ;
        RECT -16.485 -55.83 -16.155 -55.5 ;
        RECT -16.485 -56.605 -16.155 -56.275 ;
        RECT -16.485 -57.965 -16.155 -57.635 ;
        RECT -16.485 -59.325 -16.155 -58.995 ;
        RECT -16.485 -62.045 -16.155 -61.715 ;
        RECT -16.485 -64.765 -16.155 -64.435 ;
        RECT -16.485 -66.125 -16.155 -65.795 ;
        RECT -16.485 -67.485 -16.155 -67.155 ;
        RECT -16.485 -68.845 -16.155 -68.515 ;
        RECT -16.485 -70.47 -16.155 -70.14 ;
        RECT -16.485 -71.565 -16.155 -71.235 ;
        RECT -16.485 -72.925 -16.155 -72.595 ;
        RECT -16.485 -75.645 -16.155 -75.315 ;
        RECT -16.485 -77.005 -16.155 -76.675 ;
        RECT -16.485 -78.01 -16.155 -77.68 ;
        RECT -16.485 -79.725 -16.155 -79.395 ;
        RECT -16.485 -81.085 -16.155 -80.755 ;
        RECT -16.48 -85.84 -16.16 -44.04 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 -151.805 -16.155 -151.475 ;
        RECT -16.485 -153.165 -16.155 -152.835 ;
        RECT -16.485 -158.81 -16.155 -157.68 ;
        RECT -16.48 -158.925 -16.16 -149.44 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.125 44.8 -14.795 45.93 ;
        RECT -15.125 39.955 -14.795 40.285 ;
        RECT -15.125 38.595 -14.795 38.925 ;
        RECT -15.125 37.235 -14.795 37.565 ;
        RECT -15.125 35.875 -14.795 36.205 ;
        RECT -15.125 34.515 -14.795 34.845 ;
        RECT -15.125 33.155 -14.795 33.485 ;
        RECT -15.125 31.795 -14.795 32.125 ;
        RECT -15.125 30.435 -14.795 30.765 ;
        RECT -15.125 29.075 -14.795 29.405 ;
        RECT -15.125 27.715 -14.795 28.045 ;
        RECT -15.125 26.355 -14.795 26.685 ;
        RECT -15.125 24.995 -14.795 25.325 ;
        RECT -15.125 23.635 -14.795 23.965 ;
        RECT -15.125 22.275 -14.795 22.605 ;
        RECT -15.125 20.915 -14.795 21.245 ;
        RECT -15.125 19.555 -14.795 19.885 ;
        RECT -15.125 18.195 -14.795 18.525 ;
        RECT -15.125 16.835 -14.795 17.165 ;
        RECT -15.125 15.475 -14.795 15.805 ;
        RECT -15.125 14.115 -14.795 14.445 ;
        RECT -15.125 12.755 -14.795 13.085 ;
        RECT -15.125 11.395 -14.795 11.725 ;
        RECT -15.125 10.035 -14.795 10.365 ;
        RECT -15.125 8.675 -14.795 9.005 ;
        RECT -15.125 7.315 -14.795 7.645 ;
        RECT -15.125 5.955 -14.795 6.285 ;
        RECT -15.125 4.595 -14.795 4.925 ;
        RECT -15.125 3.235 -14.795 3.565 ;
        RECT -15.125 1.875 -14.795 2.205 ;
        RECT -15.125 0.515 -14.795 0.845 ;
        RECT -15.125 -2.205 -14.795 -1.875 ;
        RECT -15.125 -4.925 -14.795 -4.595 ;
        RECT -15.125 -5.65 -14.795 -5.32 ;
        RECT -15.125 -7.645 -14.795 -7.315 ;
        RECT -15.125 -11.69 -14.795 -11.36 ;
        RECT -15.125 -13.085 -14.795 -12.755 ;
        RECT -15.125 -15.805 -14.795 -15.475 ;
        RECT -15.12 -17.16 -14.8 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.125 -21.245 -14.795 -20.915 ;
        RECT -15.125 -22.605 -14.795 -22.275 ;
        RECT -15.125 -25.325 -14.795 -24.995 ;
        RECT -15.125 -26.685 -14.795 -26.355 ;
        RECT -15.125 -27.67 -14.795 -27.34 ;
        RECT -15.125 -29.405 -14.795 -29.075 ;
        RECT -15.125 -30.765 -14.795 -30.435 ;
        RECT -15.125 -33.71 -14.795 -33.38 ;
        RECT -15.125 -34.845 -14.795 -34.515 ;
        RECT -15.125 -37.565 -14.795 -37.235 ;
        RECT -15.12 -38.92 -14.8 -20.915 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.125 -43.005 -14.795 -42.675 ;
        RECT -15.125 -45.725 -14.795 -45.395 ;
        RECT -15.125 -47.085 -14.795 -46.755 ;
        RECT -15.125 -48.29 -14.795 -47.96 ;
        RECT -15.125 -49.805 -14.795 -49.475 ;
        RECT -15.125 -52.525 -14.795 -52.195 ;
        RECT -15.125 -53.885 -14.795 -53.555 ;
        RECT -15.125 -55.83 -14.795 -55.5 ;
        RECT -15.125 -56.605 -14.795 -56.275 ;
        RECT -15.125 -57.965 -14.795 -57.635 ;
        RECT -15.125 -59.325 -14.795 -58.995 ;
        RECT -15.125 -62.045 -14.795 -61.715 ;
        RECT -15.125 -64.765 -14.795 -64.435 ;
        RECT -15.125 -66.125 -14.795 -65.795 ;
        RECT -15.125 -67.485 -14.795 -67.155 ;
        RECT -15.125 -68.845 -14.795 -68.515 ;
        RECT -15.125 -70.47 -14.795 -70.14 ;
        RECT -15.125 -71.565 -14.795 -71.235 ;
        RECT -15.125 -72.925 -14.795 -72.595 ;
        RECT -15.125 -75.645 -14.795 -75.315 ;
        RECT -15.125 -77.005 -14.795 -76.675 ;
        RECT -15.125 -78.01 -14.795 -77.68 ;
        RECT -15.125 -79.725 -14.795 -79.395 ;
        RECT -15.125 -81.085 -14.795 -80.755 ;
        RECT -15.12 -84.48 -14.8 -42.675 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.125 -89.245 -14.795 -88.915 ;
        RECT -15.125 -90.605 -14.795 -90.275 ;
        RECT -15.125 -91.965 -14.795 -91.635 ;
        RECT -15.125 -93.325 -14.795 -92.995 ;
        RECT -15.125 -94.685 -14.795 -94.355 ;
        RECT -15.125 -102.845 -14.795 -102.515 ;
        RECT -15.125 -108.285 -14.795 -107.955 ;
        RECT -15.125 -109.645 -14.795 -109.315 ;
        RECT -15.125 -113.725 -14.795 -113.395 ;
        RECT -15.125 -116.445 -14.795 -116.115 ;
        RECT -15.125 -120.525 -14.795 -120.195 ;
        RECT -15.125 -121.885 -14.795 -121.555 ;
        RECT -15.125 -127.325 -14.795 -126.995 ;
        RECT -15.125 -131.405 -14.795 -131.075 ;
        RECT -15.125 -132.765 -14.795 -132.435 ;
        RECT -15.125 -134.125 -14.795 -133.795 ;
        RECT -15.125 -135.485 -14.795 -135.155 ;
        RECT -15.125 -136.845 -14.795 -136.515 ;
        RECT -15.125 -138.205 -14.795 -137.875 ;
        RECT -15.125 -139.565 -14.795 -139.235 ;
        RECT -15.125 -140.925 -14.795 -140.595 ;
        RECT -15.125 -143.755 -14.795 -143.425 ;
        RECT -15.125 -145.005 -14.795 -144.675 ;
        RECT -15.125 -146.365 -14.795 -146.035 ;
        RECT -15.125 -149.085 -14.795 -148.755 ;
        RECT -15.125 -151.805 -14.795 -151.475 ;
        RECT -15.125 -153.165 -14.795 -152.835 ;
        RECT -15.125 -158.81 -14.795 -157.68 ;
        RECT -15.12 -158.925 -14.8 -88.915 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.765 44.8 -13.435 45.93 ;
        RECT -13.765 39.955 -13.435 40.285 ;
        RECT -13.765 38.595 -13.435 38.925 ;
        RECT -13.765 37.235 -13.435 37.565 ;
        RECT -13.765 35.875 -13.435 36.205 ;
        RECT -13.765 34.515 -13.435 34.845 ;
        RECT -13.765 33.155 -13.435 33.485 ;
        RECT -13.765 31.795 -13.435 32.125 ;
        RECT -13.765 30.435 -13.435 30.765 ;
        RECT -13.765 29.075 -13.435 29.405 ;
        RECT -13.765 27.715 -13.435 28.045 ;
        RECT -13.765 26.355 -13.435 26.685 ;
        RECT -13.765 24.995 -13.435 25.325 ;
        RECT -13.765 23.635 -13.435 23.965 ;
        RECT -13.765 22.275 -13.435 22.605 ;
        RECT -13.765 20.915 -13.435 21.245 ;
        RECT -13.765 19.555 -13.435 19.885 ;
        RECT -13.765 18.195 -13.435 18.525 ;
        RECT -13.765 16.835 -13.435 17.165 ;
        RECT -13.765 15.475 -13.435 15.805 ;
        RECT -13.765 14.115 -13.435 14.445 ;
        RECT -13.765 12.755 -13.435 13.085 ;
        RECT -13.765 11.395 -13.435 11.725 ;
        RECT -13.765 10.035 -13.435 10.365 ;
        RECT -13.765 8.675 -13.435 9.005 ;
        RECT -13.765 7.315 -13.435 7.645 ;
        RECT -13.765 5.955 -13.435 6.285 ;
        RECT -13.765 4.595 -13.435 4.925 ;
        RECT -13.765 3.235 -13.435 3.565 ;
        RECT -13.765 1.875 -13.435 2.205 ;
        RECT -13.765 0.515 -13.435 0.845 ;
        RECT -13.765 -2.205 -13.435 -1.875 ;
        RECT -13.765 -4.925 -13.435 -4.595 ;
        RECT -13.765 -5.65 -13.435 -5.32 ;
        RECT -13.765 -7.645 -13.435 -7.315 ;
        RECT -13.765 -11.69 -13.435 -11.36 ;
        RECT -13.765 -13.085 -13.435 -12.755 ;
        RECT -13.765 -15.805 -13.435 -15.475 ;
        RECT -13.76 -19.88 -13.44 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.765 -77.005 -13.435 -76.675 ;
        RECT -13.765 -78.01 -13.435 -77.68 ;
        RECT -13.765 -79.725 -13.435 -79.395 ;
        RECT -13.765 -81.085 -13.435 -80.755 ;
        RECT -13.765 -87.885 -13.435 -87.555 ;
        RECT -13.765 -89.245 -13.435 -88.915 ;
        RECT -13.765 -90.605 -13.435 -90.275 ;
        RECT -13.765 -91.965 -13.435 -91.635 ;
        RECT -13.765 -93.325 -13.435 -92.995 ;
        RECT -13.765 -94.685 -13.435 -94.355 ;
        RECT -13.765 -104.205 -13.435 -103.875 ;
        RECT -13.765 -108.285 -13.435 -107.955 ;
        RECT -13.765 -109.645 -13.435 -109.315 ;
        RECT -13.765 -116.445 -13.435 -116.115 ;
        RECT -13.765 -121.885 -13.435 -121.555 ;
        RECT -13.765 -124.605 -13.435 -124.275 ;
        RECT -13.765 -127.325 -13.435 -126.995 ;
        RECT -13.765 -131.405 -13.435 -131.075 ;
        RECT -13.765 -132.765 -13.435 -132.435 ;
        RECT -13.765 -134.125 -13.435 -133.795 ;
        RECT -13.765 -135.485 -13.435 -135.155 ;
        RECT -13.765 -136.845 -13.435 -136.515 ;
        RECT -13.765 -138.205 -13.435 -137.875 ;
        RECT -13.765 -139.565 -13.435 -139.235 ;
        RECT -13.765 -140.925 -13.435 -140.595 ;
        RECT -13.765 -143.755 -13.435 -143.425 ;
        RECT -13.765 -145.005 -13.435 -144.675 ;
        RECT -13.765 -146.365 -13.435 -146.035 ;
        RECT -13.765 -147.725 -13.435 -147.395 ;
        RECT -13.765 -149.085 -13.435 -148.755 ;
        RECT -13.765 -151.805 -13.435 -151.475 ;
        RECT -13.765 -153.165 -13.435 -152.835 ;
        RECT -13.765 -158.81 -13.435 -157.68 ;
        RECT -13.76 -158.925 -13.44 -76.675 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.405 44.8 -12.075 45.93 ;
        RECT -12.405 39.955 -12.075 40.285 ;
        RECT -12.405 38.595 -12.075 38.925 ;
        RECT -12.405 37.235 -12.075 37.565 ;
        RECT -12.405 35.875 -12.075 36.205 ;
        RECT -12.405 34.515 -12.075 34.845 ;
        RECT -12.405 33.155 -12.075 33.485 ;
        RECT -12.405 31.795 -12.075 32.125 ;
        RECT -12.405 30.435 -12.075 30.765 ;
        RECT -12.405 29.075 -12.075 29.405 ;
        RECT -12.405 27.715 -12.075 28.045 ;
        RECT -12.405 26.355 -12.075 26.685 ;
        RECT -12.405 24.995 -12.075 25.325 ;
        RECT -12.405 23.635 -12.075 23.965 ;
        RECT -12.405 22.275 -12.075 22.605 ;
        RECT -12.405 20.915 -12.075 21.245 ;
        RECT -12.405 19.555 -12.075 19.885 ;
        RECT -12.405 18.195 -12.075 18.525 ;
        RECT -12.405 16.835 -12.075 17.165 ;
        RECT -12.405 15.475 -12.075 15.805 ;
        RECT -12.405 14.115 -12.075 14.445 ;
        RECT -12.405 12.755 -12.075 13.085 ;
        RECT -12.405 11.395 -12.075 11.725 ;
        RECT -12.405 10.035 -12.075 10.365 ;
        RECT -12.405 8.675 -12.075 9.005 ;
        RECT -12.405 7.315 -12.075 7.645 ;
        RECT -12.405 5.955 -12.075 6.285 ;
        RECT -12.405 4.595 -12.075 4.925 ;
        RECT -12.405 3.235 -12.075 3.565 ;
        RECT -12.405 1.875 -12.075 2.205 ;
        RECT -12.405 0.515 -12.075 0.845 ;
        RECT -12.405 -0.845 -12.075 -0.515 ;
        RECT -12.405 -2.205 -12.075 -1.875 ;
        RECT -12.405 -3.565 -12.075 -3.235 ;
        RECT -12.405 -4.925 -12.075 -4.595 ;
        RECT -12.405 -5.65 -12.075 -5.32 ;
        RECT -12.405 -7.645 -12.075 -7.315 ;
        RECT -12.405 -11.69 -12.075 -11.36 ;
        RECT -12.405 -13.085 -12.075 -12.755 ;
        RECT -12.405 -15.805 -12.075 -15.475 ;
        RECT -12.405 -21.245 -12.075 -20.915 ;
        RECT -12.405 -22.605 -12.075 -22.275 ;
        RECT -12.405 -23.965 -12.075 -23.635 ;
        RECT -12.405 -25.325 -12.075 -24.995 ;
        RECT -12.405 -26.685 -12.075 -26.355 ;
        RECT -12.405 -27.67 -12.075 -27.34 ;
        RECT -12.405 -29.405 -12.075 -29.075 ;
        RECT -12.405 -30.765 -12.075 -30.435 ;
        RECT -12.405 -33.71 -12.075 -33.38 ;
        RECT -12.405 -37.565 -12.075 -37.235 ;
        RECT -12.405 -43.005 -12.075 -42.675 ;
        RECT -12.405 -45.725 -12.075 -45.395 ;
        RECT -12.405 -47.085 -12.075 -46.755 ;
        RECT -12.405 -48.29 -12.075 -47.96 ;
        RECT -12.405 -49.805 -12.075 -49.475 ;
        RECT -12.405 -52.525 -12.075 -52.195 ;
        RECT -12.405 -53.885 -12.075 -53.555 ;
        RECT -12.405 -55.83 -12.075 -55.5 ;
        RECT -12.405 -56.605 -12.075 -56.275 ;
        RECT -12.405 -57.965 -12.075 -57.635 ;
        RECT -12.405 -59.325 -12.075 -58.995 ;
        RECT -12.405 -62.045 -12.075 -61.715 ;
        RECT -12.405 -64.765 -12.075 -64.435 ;
        RECT -12.405 -66.125 -12.075 -65.795 ;
        RECT -12.405 -67.485 -12.075 -67.155 ;
        RECT -12.405 -68.845 -12.075 -68.515 ;
        RECT -12.405 -70.47 -12.075 -70.14 ;
        RECT -12.405 -71.565 -12.075 -71.235 ;
        RECT -12.405 -72.925 -12.075 -72.595 ;
        RECT -12.405 -75.645 -12.075 -75.315 ;
        RECT -12.405 -77.005 -12.075 -76.675 ;
        RECT -12.405 -78.01 -12.075 -77.68 ;
        RECT -12.405 -79.725 -12.075 -79.395 ;
        RECT -12.405 -81.085 -12.075 -80.755 ;
        RECT -12.405 -83.805 -12.075 -83.475 ;
        RECT -12.405 -87.885 -12.075 -87.555 ;
        RECT -12.405 -89.245 -12.075 -88.915 ;
        RECT -12.405 -90.605 -12.075 -90.275 ;
        RECT -12.405 -91.965 -12.075 -91.635 ;
        RECT -12.405 -93.325 -12.075 -92.995 ;
        RECT -12.405 -94.685 -12.075 -94.355 ;
        RECT -12.405 -104.205 -12.075 -103.875 ;
        RECT -12.405 -108.285 -12.075 -107.955 ;
        RECT -12.405 -109.645 -12.075 -109.315 ;
        RECT -12.405 -112.365 -12.075 -112.035 ;
        RECT -12.405 -113.725 -12.075 -113.395 ;
        RECT -12.405 -115.085 -12.075 -114.755 ;
        RECT -12.405 -116.445 -12.075 -116.115 ;
        RECT -12.405 -119.165 -12.075 -118.835 ;
        RECT -12.405 -121.885 -12.075 -121.555 ;
        RECT -12.405 -123.245 -12.075 -122.915 ;
        RECT -12.405 -124.605 -12.075 -124.275 ;
        RECT -12.405 -127.325 -12.075 -126.995 ;
        RECT -12.405 -128.685 -12.075 -128.355 ;
        RECT -12.405 -130.045 -12.075 -129.715 ;
        RECT -12.405 -131.405 -12.075 -131.075 ;
        RECT -12.405 -132.765 -12.075 -132.435 ;
        RECT -12.405 -134.125 -12.075 -133.795 ;
        RECT -12.405 -135.485 -12.075 -135.155 ;
        RECT -12.405 -136.845 -12.075 -136.515 ;
        RECT -12.405 -138.205 -12.075 -137.875 ;
        RECT -12.405 -139.565 -12.075 -139.235 ;
        RECT -12.405 -140.925 -12.075 -140.595 ;
        RECT -12.405 -143.755 -12.075 -143.425 ;
        RECT -12.405 -145.005 -12.075 -144.675 ;
        RECT -12.405 -146.365 -12.075 -146.035 ;
        RECT -12.405 -147.725 -12.075 -147.395 ;
        RECT -12.405 -149.085 -12.075 -148.755 ;
        RECT -12.405 -151.805 -12.075 -151.475 ;
        RECT -12.405 -153.165 -12.075 -152.835 ;
        RECT -12.405 -158.81 -12.075 -157.68 ;
        RECT -12.4 -158.925 -12.08 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.045 44.8 -10.715 45.93 ;
        RECT -11.045 39.955 -10.715 40.285 ;
        RECT -11.045 38.595 -10.715 38.925 ;
        RECT -11.045 37.235 -10.715 37.565 ;
        RECT -11.045 35.875 -10.715 36.205 ;
        RECT -11.045 34.515 -10.715 34.845 ;
        RECT -11.045 33.155 -10.715 33.485 ;
        RECT -11.045 31.795 -10.715 32.125 ;
        RECT -11.045 29.075 -10.715 29.405 ;
        RECT -11.045 22.275 -10.715 22.605 ;
        RECT -11.045 19.555 -10.715 19.885 ;
        RECT -11.045 18.195 -10.715 18.525 ;
        RECT -11.045 11.395 -10.715 11.725 ;
        RECT -11.045 4.595 -10.715 4.925 ;
        RECT -11.045 3.235 -10.715 3.565 ;
        RECT -11.045 1.875 -10.715 2.205 ;
        RECT -11.045 0.515 -10.715 0.845 ;
        RECT -11.045 -0.845 -10.715 -0.515 ;
        RECT -11.045 -2.205 -10.715 -1.875 ;
        RECT -11.045 -3.565 -10.715 -3.235 ;
        RECT -11.045 -4.925 -10.715 -4.595 ;
        RECT -11.045 -5.65 -10.715 -5.32 ;
        RECT -11.045 -7.645 -10.715 -7.315 ;
        RECT -11.045 -11.69 -10.715 -11.36 ;
        RECT -11.045 -13.085 -10.715 -12.755 ;
        RECT -11.045 -15.805 -10.715 -15.475 ;
        RECT -11.045 -21.245 -10.715 -20.915 ;
        RECT -11.045 -22.605 -10.715 -22.275 ;
        RECT -11.045 -23.965 -10.715 -23.635 ;
        RECT -11.045 -25.325 -10.715 -24.995 ;
        RECT -11.045 -26.685 -10.715 -26.355 ;
        RECT -11.045 -27.67 -10.715 -27.34 ;
        RECT -11.045 -29.405 -10.715 -29.075 ;
        RECT -11.045 -30.765 -10.715 -30.435 ;
        RECT -11.045 -33.71 -10.715 -33.38 ;
        RECT -11.045 -37.565 -10.715 -37.235 ;
        RECT -11.045 -43.005 -10.715 -42.675 ;
        RECT -11.045 -45.725 -10.715 -45.395 ;
        RECT -11.045 -47.085 -10.715 -46.755 ;
        RECT -11.045 -48.29 -10.715 -47.96 ;
        RECT -11.045 -49.805 -10.715 -49.475 ;
        RECT -11.045 -52.525 -10.715 -52.195 ;
        RECT -11.045 -53.885 -10.715 -53.555 ;
        RECT -11.045 -55.83 -10.715 -55.5 ;
        RECT -11.045 -56.605 -10.715 -56.275 ;
        RECT -11.045 -57.965 -10.715 -57.635 ;
        RECT -11.045 -59.325 -10.715 -58.995 ;
        RECT -11.045 -62.045 -10.715 -61.715 ;
        RECT -11.045 -64.765 -10.715 -64.435 ;
        RECT -11.045 -66.125 -10.715 -65.795 ;
        RECT -11.045 -67.485 -10.715 -67.155 ;
        RECT -11.045 -68.845 -10.715 -68.515 ;
        RECT -11.045 -70.47 -10.715 -70.14 ;
        RECT -11.045 -71.565 -10.715 -71.235 ;
        RECT -11.045 -72.925 -10.715 -72.595 ;
        RECT -11.045 -75.645 -10.715 -75.315 ;
        RECT -11.045 -77.005 -10.715 -76.675 ;
        RECT -11.045 -78.01 -10.715 -77.68 ;
        RECT -11.045 -79.725 -10.715 -79.395 ;
        RECT -11.045 -81.085 -10.715 -80.755 ;
        RECT -11.045 -83.805 -10.715 -83.475 ;
        RECT -11.045 -87.885 -10.715 -87.555 ;
        RECT -11.045 -89.245 -10.715 -88.915 ;
        RECT -11.045 -90.605 -10.715 -90.275 ;
        RECT -11.045 -91.965 -10.715 -91.635 ;
        RECT -11.045 -93.325 -10.715 -92.995 ;
        RECT -11.045 -94.685 -10.715 -94.355 ;
        RECT -11.045 -98.765 -10.715 -98.435 ;
        RECT -11.045 -101.485 -10.715 -101.155 ;
        RECT -11.045 -104.205 -10.715 -103.875 ;
        RECT -11.045 -105.565 -10.715 -105.235 ;
        RECT -11.045 -108.285 -10.715 -107.955 ;
        RECT -11.045 -109.645 -10.715 -109.315 ;
        RECT -11.045 -111.005 -10.715 -110.675 ;
        RECT -11.045 -112.365 -10.715 -112.035 ;
        RECT -11.045 -113.725 -10.715 -113.395 ;
        RECT -11.045 -115.085 -10.715 -114.755 ;
        RECT -11.045 -116.445 -10.715 -116.115 ;
        RECT -11.045 -119.165 -10.715 -118.835 ;
        RECT -11.045 -121.885 -10.715 -121.555 ;
        RECT -11.045 -123.245 -10.715 -122.915 ;
        RECT -11.045 -124.605 -10.715 -124.275 ;
        RECT -11.045 -125.965 -10.715 -125.635 ;
        RECT -11.045 -127.325 -10.715 -126.995 ;
        RECT -11.045 -128.685 -10.715 -128.355 ;
        RECT -11.045 -130.045 -10.715 -129.715 ;
        RECT -11.045 -131.405 -10.715 -131.075 ;
        RECT -11.045 -132.765 -10.715 -132.435 ;
        RECT -11.045 -134.125 -10.715 -133.795 ;
        RECT -11.045 -135.485 -10.715 -135.155 ;
        RECT -11.045 -136.845 -10.715 -136.515 ;
        RECT -11.045 -138.205 -10.715 -137.875 ;
        RECT -11.045 -139.565 -10.715 -139.235 ;
        RECT -11.045 -140.925 -10.715 -140.595 ;
        RECT -11.04 -142.28 -10.72 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.045 -149.085 -10.715 -148.755 ;
        RECT -11.045 -151.805 -10.715 -151.475 ;
        RECT -11.045 -153.165 -10.715 -152.835 ;
        RECT -11.045 -158.81 -10.715 -157.68 ;
        RECT -11.04 -158.925 -10.72 -148.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.685 44.8 -9.355 45.93 ;
        RECT -9.685 39.955 -9.355 40.285 ;
        RECT -9.685 38.595 -9.355 38.925 ;
        RECT -9.685 37.235 -9.355 37.565 ;
        RECT -9.685 35.875 -9.355 36.205 ;
        RECT -9.685 34.515 -9.355 34.845 ;
        RECT -9.685 33.155 -9.355 33.485 ;
        RECT -9.685 31.795 -9.355 32.125 ;
        RECT -9.685 29.075 -9.355 29.405 ;
        RECT -9.685 22.275 -9.355 22.605 ;
        RECT -9.685 19.555 -9.355 19.885 ;
        RECT -9.685 18.195 -9.355 18.525 ;
        RECT -9.685 11.395 -9.355 11.725 ;
        RECT -9.685 4.595 -9.355 4.925 ;
        RECT -9.685 3.235 -9.355 3.565 ;
        RECT -9.685 1.875 -9.355 2.205 ;
        RECT -9.685 0.515 -9.355 0.845 ;
        RECT -9.685 -0.845 -9.355 -0.515 ;
        RECT -9.685 -2.205 -9.355 -1.875 ;
        RECT -9.685 -3.565 -9.355 -3.235 ;
        RECT -9.685 -4.925 -9.355 -4.595 ;
        RECT -9.685 -6.285 -9.355 -5.955 ;
        RECT -9.685 -7.645 -9.355 -7.315 ;
        RECT -9.685 -10.365 -9.355 -10.035 ;
        RECT -9.685 -11.725 -9.355 -11.395 ;
        RECT -9.685 -13.085 -9.355 -12.755 ;
        RECT -9.685 -14.445 -9.355 -14.115 ;
        RECT -9.685 -15.805 -9.355 -15.475 ;
        RECT -9.685 -17.165 -9.355 -16.835 ;
        RECT -9.68 -18.52 -9.36 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.685 -77.005 -9.355 -76.675 ;
        RECT -9.685 -78.365 -9.355 -78.035 ;
        RECT -9.685 -79.725 -9.355 -79.395 ;
        RECT -9.685 -81.085 -9.355 -80.755 ;
        RECT -9.685 -82.445 -9.355 -82.115 ;
        RECT -9.685 -83.805 -9.355 -83.475 ;
        RECT -9.685 -85.165 -9.355 -84.835 ;
        RECT -9.68 -85.84 -9.36 -76.675 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.685 -134.125 -9.355 -133.795 ;
        RECT -9.685 -135.485 -9.355 -135.155 ;
        RECT -9.685 -136.845 -9.355 -136.515 ;
        RECT -9.685 -138.205 -9.355 -137.875 ;
        RECT -9.685 -139.565 -9.355 -139.235 ;
        RECT -9.685 -140.925 -9.355 -140.595 ;
        RECT -9.68 -141.6 -9.36 -133.795 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.325 44.8 -7.995 45.93 ;
        RECT -8.325 39.955 -7.995 40.285 ;
        RECT -8.325 38.595 -7.995 38.925 ;
        RECT -8.325 37.235 -7.995 37.565 ;
        RECT -8.325 35.875 -7.995 36.205 ;
        RECT -8.325 34.515 -7.995 34.845 ;
        RECT -8.325 33.155 -7.995 33.485 ;
        RECT -8.325 31.795 -7.995 32.125 ;
        RECT -8.325 29.075 -7.995 29.405 ;
        RECT -8.325 22.275 -7.995 22.605 ;
        RECT -8.325 19.555 -7.995 19.885 ;
        RECT -8.325 18.195 -7.995 18.525 ;
        RECT -8.325 11.395 -7.995 11.725 ;
        RECT -8.325 4.595 -7.995 4.925 ;
        RECT -8.325 3.235 -7.995 3.565 ;
        RECT -8.325 1.875 -7.995 2.205 ;
        RECT -8.325 0.515 -7.995 0.845 ;
        RECT -8.325 -0.845 -7.995 -0.515 ;
        RECT -8.325 -2.205 -7.995 -1.875 ;
        RECT -8.325 -3.565 -7.995 -3.235 ;
        RECT -8.325 -4.925 -7.995 -4.595 ;
        RECT -8.325 -6.285 -7.995 -5.955 ;
        RECT -8.325 -7.645 -7.995 -7.315 ;
        RECT -8.325 -9.005 -7.995 -8.675 ;
        RECT -8.325 -10.365 -7.995 -10.035 ;
        RECT -8.325 -11.725 -7.995 -11.395 ;
        RECT -8.325 -13.085 -7.995 -12.755 ;
        RECT -8.325 -14.445 -7.995 -14.115 ;
        RECT -8.325 -15.805 -7.995 -15.475 ;
        RECT -8.325 -17.165 -7.995 -16.835 ;
        RECT -8.325 -21.245 -7.995 -20.915 ;
        RECT -8.325 -22.605 -7.995 -22.275 ;
        RECT -8.325 -23.965 -7.995 -23.635 ;
        RECT -8.325 -25.325 -7.995 -24.995 ;
        RECT -8.325 -26.685 -7.995 -26.355 ;
        RECT -8.325 -28.045 -7.995 -27.715 ;
        RECT -8.325 -29.405 -7.995 -29.075 ;
        RECT -8.325 -30.765 -7.995 -30.435 ;
        RECT -8.325 -32.125 -7.995 -31.795 ;
        RECT -8.325 -33.485 -7.995 -33.155 ;
        RECT -8.325 -36.205 -7.995 -35.875 ;
        RECT -8.325 -37.565 -7.995 -37.235 ;
        RECT -8.325 -38.925 -7.995 -38.595 ;
        RECT -8.325 -40.285 -7.995 -39.955 ;
        RECT -8.325 -43.005 -7.995 -42.675 ;
        RECT -8.325 -45.725 -7.995 -45.395 ;
        RECT -8.325 -47.085 -7.995 -46.755 ;
        RECT -8.325 -48.445 -7.995 -48.115 ;
        RECT -8.325 -49.805 -7.995 -49.475 ;
        RECT -8.325 -51.165 -7.995 -50.835 ;
        RECT -8.325 -52.525 -7.995 -52.195 ;
        RECT -8.325 -53.885 -7.995 -53.555 ;
        RECT -8.325 -55.245 -7.995 -54.915 ;
        RECT -8.325 -56.605 -7.995 -56.275 ;
        RECT -8.325 -57.965 -7.995 -57.635 ;
        RECT -8.325 -59.325 -7.995 -58.995 ;
        RECT -8.325 -60.685 -7.995 -60.355 ;
        RECT -8.325 -62.045 -7.995 -61.715 ;
        RECT -8.325 -63.405 -7.995 -63.075 ;
        RECT -8.325 -64.765 -7.995 -64.435 ;
        RECT -8.325 -66.125 -7.995 -65.795 ;
        RECT -8.325 -67.485 -7.995 -67.155 ;
        RECT -8.325 -68.845 -7.995 -68.515 ;
        RECT -8.325 -70.205 -7.995 -69.875 ;
        RECT -8.325 -71.565 -7.995 -71.235 ;
        RECT -8.325 -72.925 -7.995 -72.595 ;
        RECT -8.325 -74.285 -7.995 -73.955 ;
        RECT -8.325 -75.645 -7.995 -75.315 ;
        RECT -8.325 -77.005 -7.995 -76.675 ;
        RECT -8.325 -78.365 -7.995 -78.035 ;
        RECT -8.325 -79.725 -7.995 -79.395 ;
        RECT -8.325 -81.085 -7.995 -80.755 ;
        RECT -8.325 -82.445 -7.995 -82.115 ;
        RECT -8.325 -83.805 -7.995 -83.475 ;
        RECT -8.325 -85.165 -7.995 -84.835 ;
        RECT -8.325 -87.885 -7.995 -87.555 ;
        RECT -8.325 -89.245 -7.995 -88.915 ;
        RECT -8.325 -90.605 -7.995 -90.275 ;
        RECT -8.325 -91.965 -7.995 -91.635 ;
        RECT -8.325 -93.325 -7.995 -92.995 ;
        RECT -8.325 -94.685 -7.995 -94.355 ;
        RECT -8.325 -96.045 -7.995 -95.715 ;
        RECT -8.325 -97.405 -7.995 -97.075 ;
        RECT -8.325 -98.765 -7.995 -98.435 ;
        RECT -8.325 -100.125 -7.995 -99.795 ;
        RECT -8.325 -101.485 -7.995 -101.155 ;
        RECT -8.325 -102.845 -7.995 -102.515 ;
        RECT -8.325 -104.205 -7.995 -103.875 ;
        RECT -8.325 -105.565 -7.995 -105.235 ;
        RECT -8.325 -106.925 -7.995 -106.595 ;
        RECT -8.325 -108.285 -7.995 -107.955 ;
        RECT -8.325 -109.645 -7.995 -109.315 ;
        RECT -8.325 -111.005 -7.995 -110.675 ;
        RECT -8.325 -112.365 -7.995 -112.035 ;
        RECT -8.325 -113.725 -7.995 -113.395 ;
        RECT -8.325 -115.085 -7.995 -114.755 ;
        RECT -8.325 -116.445 -7.995 -116.115 ;
        RECT -8.325 -117.805 -7.995 -117.475 ;
        RECT -8.325 -119.165 -7.995 -118.835 ;
        RECT -8.325 -120.525 -7.995 -120.195 ;
        RECT -8.325 -121.885 -7.995 -121.555 ;
        RECT -8.325 -123.245 -7.995 -122.915 ;
        RECT -8.325 -124.605 -7.995 -124.275 ;
        RECT -8.325 -125.965 -7.995 -125.635 ;
        RECT -8.325 -127.325 -7.995 -126.995 ;
        RECT -8.325 -128.685 -7.995 -128.355 ;
        RECT -8.325 -130.045 -7.995 -129.715 ;
        RECT -8.325 -131.405 -7.995 -131.075 ;
        RECT -8.325 -132.765 -7.995 -132.435 ;
        RECT -8.325 -134.125 -7.995 -133.795 ;
        RECT -8.325 -135.485 -7.995 -135.155 ;
        RECT -8.325 -136.845 -7.995 -136.515 ;
        RECT -8.325 -138.205 -7.995 -137.875 ;
        RECT -8.325 -139.565 -7.995 -139.235 ;
        RECT -8.325 -140.925 -7.995 -140.595 ;
        RECT -8.325 -142.285 -7.995 -141.955 ;
        RECT -8.325 -143.645 -7.995 -143.315 ;
        RECT -8.325 -145.005 -7.995 -144.675 ;
        RECT -8.325 -146.365 -7.995 -146.035 ;
        RECT -8.325 -147.725 -7.995 -147.395 ;
        RECT -8.325 -149.085 -7.995 -148.755 ;
        RECT -8.325 -150.445 -7.995 -150.115 ;
        RECT -8.325 -151.805 -7.995 -151.475 ;
        RECT -8.325 -153.165 -7.995 -152.835 ;
        RECT -8.325 -158.81 -7.995 -157.68 ;
        RECT -8.32 -158.925 -8 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.965 29.075 -6.635 29.405 ;
        RECT -6.965 22.275 -6.635 22.605 ;
        RECT -6.965 19.555 -6.635 19.885 ;
        RECT -6.965 18.195 -6.635 18.525 ;
        RECT -6.965 11.395 -6.635 11.725 ;
        RECT -6.965 4.595 -6.635 4.925 ;
        RECT -6.965 3.235 -6.635 3.565 ;
        RECT -6.965 1.875 -6.635 2.205 ;
        RECT -6.965 0.515 -6.635 0.845 ;
        RECT -6.965 -0.845 -6.635 -0.515 ;
        RECT -6.965 -2.205 -6.635 -1.875 ;
        RECT -6.965 -3.565 -6.635 -3.235 ;
        RECT -6.965 -4.925 -6.635 -4.595 ;
        RECT -6.965 -6.285 -6.635 -5.955 ;
        RECT -6.965 -7.645 -6.635 -7.315 ;
        RECT -6.965 -9.005 -6.635 -8.675 ;
        RECT -6.965 -10.365 -6.635 -10.035 ;
        RECT -6.965 -11.725 -6.635 -11.395 ;
        RECT -6.965 -13.085 -6.635 -12.755 ;
        RECT -6.965 -14.445 -6.635 -14.115 ;
        RECT -6.965 -15.805 -6.635 -15.475 ;
        RECT -6.965 -17.165 -6.635 -16.835 ;
        RECT -6.965 -21.245 -6.635 -20.915 ;
        RECT -6.965 -22.605 -6.635 -22.275 ;
        RECT -6.965 -23.965 -6.635 -23.635 ;
        RECT -6.965 -25.325 -6.635 -24.995 ;
        RECT -6.965 -26.685 -6.635 -26.355 ;
        RECT -6.965 -28.045 -6.635 -27.715 ;
        RECT -6.965 -29.405 -6.635 -29.075 ;
        RECT -6.965 -30.765 -6.635 -30.435 ;
        RECT -6.965 -32.125 -6.635 -31.795 ;
        RECT -6.965 -33.485 -6.635 -33.155 ;
        RECT -6.965 -36.205 -6.635 -35.875 ;
        RECT -6.965 -37.565 -6.635 -37.235 ;
        RECT -6.965 -38.925 -6.635 -38.595 ;
        RECT -6.965 -40.285 -6.635 -39.955 ;
        RECT -6.965 -43.005 -6.635 -42.675 ;
        RECT -6.965 -45.725 -6.635 -45.395 ;
        RECT -6.965 -47.085 -6.635 -46.755 ;
        RECT -6.965 -48.445 -6.635 -48.115 ;
        RECT -6.965 -49.805 -6.635 -49.475 ;
        RECT -6.965 -51.165 -6.635 -50.835 ;
        RECT -6.965 -52.525 -6.635 -52.195 ;
        RECT -6.965 -53.885 -6.635 -53.555 ;
        RECT -6.965 -55.245 -6.635 -54.915 ;
        RECT -6.965 -56.605 -6.635 -56.275 ;
        RECT -6.965 -57.965 -6.635 -57.635 ;
        RECT -6.965 -59.325 -6.635 -58.995 ;
        RECT -6.965 -60.685 -6.635 -60.355 ;
        RECT -6.965 -62.045 -6.635 -61.715 ;
        RECT -6.965 -63.405 -6.635 -63.075 ;
        RECT -6.965 -64.765 -6.635 -64.435 ;
        RECT -6.965 -66.125 -6.635 -65.795 ;
        RECT -6.965 -67.485 -6.635 -67.155 ;
        RECT -6.965 -68.845 -6.635 -68.515 ;
        RECT -6.965 -70.205 -6.635 -69.875 ;
        RECT -6.965 -71.565 -6.635 -71.235 ;
        RECT -6.965 -72.925 -6.635 -72.595 ;
        RECT -6.965 -74.285 -6.635 -73.955 ;
        RECT -6.965 -75.645 -6.635 -75.315 ;
        RECT -6.965 -77.005 -6.635 -76.675 ;
        RECT -6.965 -78.365 -6.635 -78.035 ;
        RECT -6.965 -79.725 -6.635 -79.395 ;
        RECT -6.965 -81.085 -6.635 -80.755 ;
        RECT -6.965 -82.445 -6.635 -82.115 ;
        RECT -6.965 -83.805 -6.635 -83.475 ;
        RECT -6.965 -85.165 -6.635 -84.835 ;
        RECT -6.965 -87.885 -6.635 -87.555 ;
        RECT -6.965 -89.245 -6.635 -88.915 ;
        RECT -6.965 -90.605 -6.635 -90.275 ;
        RECT -6.965 -91.965 -6.635 -91.635 ;
        RECT -6.965 -93.325 -6.635 -92.995 ;
        RECT -6.965 -94.685 -6.635 -94.355 ;
        RECT -6.965 -96.045 -6.635 -95.715 ;
        RECT -6.965 -97.405 -6.635 -97.075 ;
        RECT -6.965 -98.765 -6.635 -98.435 ;
        RECT -6.965 -100.125 -6.635 -99.795 ;
        RECT -6.965 -101.485 -6.635 -101.155 ;
        RECT -6.965 -102.845 -6.635 -102.515 ;
        RECT -6.965 -104.205 -6.635 -103.875 ;
        RECT -6.965 -105.565 -6.635 -105.235 ;
        RECT -6.965 -106.925 -6.635 -106.595 ;
        RECT -6.965 -108.285 -6.635 -107.955 ;
        RECT -6.965 -109.645 -6.635 -109.315 ;
        RECT -6.965 -111.005 -6.635 -110.675 ;
        RECT -6.965 -112.365 -6.635 -112.035 ;
        RECT -6.965 -113.725 -6.635 -113.395 ;
        RECT -6.965 -115.085 -6.635 -114.755 ;
        RECT -6.965 -116.445 -6.635 -116.115 ;
        RECT -6.965 -117.805 -6.635 -117.475 ;
        RECT -6.965 -119.165 -6.635 -118.835 ;
        RECT -6.965 -120.525 -6.635 -120.195 ;
        RECT -6.965 -121.885 -6.635 -121.555 ;
        RECT -6.965 -123.245 -6.635 -122.915 ;
        RECT -6.965 -124.605 -6.635 -124.275 ;
        RECT -6.965 -125.965 -6.635 -125.635 ;
        RECT -6.965 -127.325 -6.635 -126.995 ;
        RECT -6.965 -128.685 -6.635 -128.355 ;
        RECT -6.965 -130.045 -6.635 -129.715 ;
        RECT -6.965 -131.405 -6.635 -131.075 ;
        RECT -6.965 -132.765 -6.635 -132.435 ;
        RECT -6.965 -134.125 -6.635 -133.795 ;
        RECT -6.965 -135.485 -6.635 -135.155 ;
        RECT -6.965 -136.845 -6.635 -136.515 ;
        RECT -6.965 -138.205 -6.635 -137.875 ;
        RECT -6.965 -139.565 -6.635 -139.235 ;
        RECT -6.965 -140.925 -6.635 -140.595 ;
        RECT -6.965 -142.285 -6.635 -141.955 ;
        RECT -6.965 -143.645 -6.635 -143.315 ;
        RECT -6.965 -145.005 -6.635 -144.675 ;
        RECT -6.965 -146.365 -6.635 -146.035 ;
        RECT -6.965 -147.725 -6.635 -147.395 ;
        RECT -6.965 -149.085 -6.635 -148.755 ;
        RECT -6.965 -150.445 -6.635 -150.115 ;
        RECT -6.965 -151.805 -6.635 -151.475 ;
        RECT -6.965 -153.165 -6.635 -152.835 ;
        RECT -6.965 -158.81 -6.635 -157.68 ;
        RECT -6.96 -158.925 -6.64 46.045 ;
        RECT -6.965 44.8 -6.635 45.93 ;
        RECT -6.965 39.955 -6.635 40.285 ;
        RECT -6.965 38.595 -6.635 38.925 ;
        RECT -6.965 37.235 -6.635 37.565 ;
        RECT -6.965 35.875 -6.635 36.205 ;
        RECT -6.965 34.515 -6.635 34.845 ;
        RECT -6.965 33.155 -6.635 33.485 ;
        RECT -6.965 31.795 -6.635 32.125 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.805 -149.085 -32.475 -148.755 ;
        RECT -32.805 -151.805 -32.475 -151.475 ;
        RECT -32.805 -153.165 -32.475 -152.835 ;
        RECT -32.805 -158.81 -32.475 -157.68 ;
        RECT -32.8 -158.925 -32.48 -147.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.445 44.8 -31.115 45.93 ;
        RECT -31.445 39.955 -31.115 40.285 ;
        RECT -31.445 38.595 -31.115 38.925 ;
        RECT -31.445 37.235 -31.115 37.565 ;
        RECT -31.445 35.875 -31.115 36.205 ;
        RECT -31.445 34.515 -31.115 34.845 ;
        RECT -31.445 33.155 -31.115 33.485 ;
        RECT -31.445 31.795 -31.115 32.125 ;
        RECT -31.445 30.435 -31.115 30.765 ;
        RECT -31.445 29.075 -31.115 29.405 ;
        RECT -31.445 27.715 -31.115 28.045 ;
        RECT -31.445 26.355 -31.115 26.685 ;
        RECT -31.445 24.995 -31.115 25.325 ;
        RECT -31.445 23.635 -31.115 23.965 ;
        RECT -31.445 22.275 -31.115 22.605 ;
        RECT -31.445 20.915 -31.115 21.245 ;
        RECT -31.445 19.555 -31.115 19.885 ;
        RECT -31.445 18.195 -31.115 18.525 ;
        RECT -31.445 16.835 -31.115 17.165 ;
        RECT -31.445 15.475 -31.115 15.805 ;
        RECT -31.445 14.115 -31.115 14.445 ;
        RECT -31.445 12.755 -31.115 13.085 ;
        RECT -31.445 11.395 -31.115 11.725 ;
        RECT -31.445 10.035 -31.115 10.365 ;
        RECT -31.445 8.675 -31.115 9.005 ;
        RECT -31.445 7.315 -31.115 7.645 ;
        RECT -31.445 5.955 -31.115 6.285 ;
        RECT -31.445 4.595 -31.115 4.925 ;
        RECT -31.445 3.235 -31.115 3.565 ;
        RECT -31.445 1.875 -31.115 2.205 ;
        RECT -31.445 -2.205 -31.115 -1.875 ;
        RECT -31.445 -4.925 -31.115 -4.595 ;
        RECT -31.445 -6.285 -31.115 -5.955 ;
        RECT -31.445 -7.645 -31.115 -7.315 ;
        RECT -31.445 -10.365 -31.115 -10.035 ;
        RECT -31.445 -11.725 -31.115 -11.395 ;
        RECT -31.445 -13.085 -31.115 -12.755 ;
        RECT -31.445 -14.445 -31.115 -14.115 ;
        RECT -31.445 -15.805 -31.115 -15.475 ;
        RECT -31.445 -17.165 -31.115 -16.835 ;
        RECT -31.445 -18.525 -31.115 -18.195 ;
        RECT -31.445 -25.325 -31.115 -24.995 ;
        RECT -31.445 -26.685 -31.115 -26.355 ;
        RECT -31.445 -28.045 -31.115 -27.715 ;
        RECT -31.445 -29.405 -31.115 -29.075 ;
        RECT -31.445 -30.765 -31.115 -30.435 ;
        RECT -31.445 -32.125 -31.115 -31.795 ;
        RECT -31.445 -33.485 -31.115 -33.155 ;
        RECT -31.445 -34.845 -31.115 -34.515 ;
        RECT -31.445 -36.205 -31.115 -35.875 ;
        RECT -31.445 -37.565 -31.115 -37.235 ;
        RECT -31.445 -38.925 -31.115 -38.595 ;
        RECT -31.445 -40.285 -31.115 -39.955 ;
        RECT -31.445 -43.005 -31.115 -42.675 ;
        RECT -31.445 -44.365 -31.115 -44.035 ;
        RECT -31.445 -45.725 -31.115 -45.395 ;
        RECT -31.445 -47.085 -31.115 -46.755 ;
        RECT -31.445 -48.445 -31.115 -48.115 ;
        RECT -31.445 -49.805 -31.115 -49.475 ;
        RECT -31.445 -51.165 -31.115 -50.835 ;
        RECT -31.445 -52.525 -31.115 -52.195 ;
        RECT -31.445 -53.885 -31.115 -53.555 ;
        RECT -31.445 -55.245 -31.115 -54.915 ;
        RECT -31.445 -56.605 -31.115 -56.275 ;
        RECT -31.445 -57.965 -31.115 -57.635 ;
        RECT -31.445 -59.325 -31.115 -58.995 ;
        RECT -31.445 -60.685 -31.115 -60.355 ;
        RECT -31.445 -62.045 -31.115 -61.715 ;
        RECT -31.445 -63.405 -31.115 -63.075 ;
        RECT -31.445 -64.765 -31.115 -64.435 ;
        RECT -31.445 -65.91 -31.115 -65.58 ;
        RECT -31.445 -67.485 -31.115 -67.155 ;
        RECT -31.445 -68.845 -31.115 -68.515 ;
        RECT -31.445 -70.205 -31.115 -69.875 ;
        RECT -31.445 -71.565 -31.115 -71.235 ;
        RECT -31.445 -72.925 -31.115 -72.595 ;
        RECT -31.445 -75.645 -31.115 -75.315 ;
        RECT -31.445 -76.45 -31.115 -76.12 ;
        RECT -31.445 -78.365 -31.115 -78.035 ;
        RECT -31.445 -79.725 -31.115 -79.395 ;
        RECT -31.445 -81.085 -31.115 -80.755 ;
        RECT -31.445 -83.805 -31.115 -83.475 ;
        RECT -31.445 -85.165 -31.115 -84.835 ;
        RECT -31.445 -87.885 -31.115 -87.555 ;
        RECT -31.445 -89.245 -31.115 -88.915 ;
        RECT -31.445 -90.605 -31.115 -90.275 ;
        RECT -31.445 -91.965 -31.115 -91.635 ;
        RECT -31.445 -93.325 -31.115 -92.995 ;
        RECT -31.445 -94.685 -31.115 -94.355 ;
        RECT -31.445 -96.045 -31.115 -95.715 ;
        RECT -31.445 -97.405 -31.115 -97.075 ;
        RECT -31.445 -98.765 -31.115 -98.435 ;
        RECT -31.445 -100.125 -31.115 -99.795 ;
        RECT -31.445 -101.485 -31.115 -101.155 ;
        RECT -31.445 -102.845 -31.115 -102.515 ;
        RECT -31.445 -104.205 -31.115 -103.875 ;
        RECT -31.445 -108.285 -31.115 -107.955 ;
        RECT -31.445 -109.645 -31.115 -109.315 ;
        RECT -31.445 -111.005 -31.115 -110.675 ;
        RECT -31.445 -113.725 -31.115 -113.395 ;
        RECT -31.445 -116.445 -31.115 -116.115 ;
        RECT -31.445 -117.805 -31.115 -117.475 ;
        RECT -31.445 -119.165 -31.115 -118.835 ;
        RECT -31.445 -120.525 -31.115 -120.195 ;
        RECT -31.445 -121.885 -31.115 -121.555 ;
        RECT -31.445 -123.245 -31.115 -122.915 ;
        RECT -31.445 -125.965 -31.115 -125.635 ;
        RECT -31.445 -127.325 -31.115 -126.995 ;
        RECT -31.445 -131.405 -31.115 -131.075 ;
        RECT -31.445 -132.765 -31.115 -132.435 ;
        RECT -31.445 -134.125 -31.115 -133.795 ;
        RECT -31.445 -135.485 -31.115 -135.155 ;
        RECT -31.445 -136.845 -31.115 -136.515 ;
        RECT -31.445 -138.205 -31.115 -137.875 ;
        RECT -31.445 -139.565 -31.115 -139.235 ;
        RECT -31.445 -140.925 -31.115 -140.595 ;
        RECT -31.445 -143.755 -31.115 -143.425 ;
        RECT -31.445 -145.005 -31.115 -144.675 ;
        RECT -31.445 -146.365 -31.115 -146.035 ;
        RECT -31.445 -147.725 -31.115 -147.395 ;
        RECT -31.445 -149.085 -31.115 -148.755 ;
        RECT -31.445 -151.805 -31.115 -151.475 ;
        RECT -31.445 -153.165 -31.115 -152.835 ;
        RECT -31.445 -158.81 -31.115 -157.68 ;
        RECT -31.44 -158.925 -31.12 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 44.8 -29.755 45.93 ;
        RECT -30.085 39.955 -29.755 40.285 ;
        RECT -30.085 38.595 -29.755 38.925 ;
        RECT -30.085 37.235 -29.755 37.565 ;
        RECT -30.085 35.875 -29.755 36.205 ;
        RECT -30.085 34.515 -29.755 34.845 ;
        RECT -30.085 33.155 -29.755 33.485 ;
        RECT -30.085 31.795 -29.755 32.125 ;
        RECT -30.085 30.435 -29.755 30.765 ;
        RECT -30.085 29.075 -29.755 29.405 ;
        RECT -30.085 27.715 -29.755 28.045 ;
        RECT -30.085 26.355 -29.755 26.685 ;
        RECT -30.085 24.995 -29.755 25.325 ;
        RECT -30.085 23.635 -29.755 23.965 ;
        RECT -30.085 22.275 -29.755 22.605 ;
        RECT -30.085 20.915 -29.755 21.245 ;
        RECT -30.085 19.555 -29.755 19.885 ;
        RECT -30.085 18.195 -29.755 18.525 ;
        RECT -30.085 16.835 -29.755 17.165 ;
        RECT -30.085 15.475 -29.755 15.805 ;
        RECT -30.085 14.115 -29.755 14.445 ;
        RECT -30.085 12.755 -29.755 13.085 ;
        RECT -30.085 11.395 -29.755 11.725 ;
        RECT -30.085 10.035 -29.755 10.365 ;
        RECT -30.085 8.675 -29.755 9.005 ;
        RECT -30.085 7.315 -29.755 7.645 ;
        RECT -30.085 5.955 -29.755 6.285 ;
        RECT -30.085 4.595 -29.755 4.925 ;
        RECT -30.085 3.235 -29.755 3.565 ;
        RECT -30.085 1.875 -29.755 2.205 ;
        RECT -30.085 -2.205 -29.755 -1.875 ;
        RECT -30.085 -4.925 -29.755 -4.595 ;
        RECT -30.085 -6.285 -29.755 -5.955 ;
        RECT -30.085 -7.645 -29.755 -7.315 ;
        RECT -30.085 -10.365 -29.755 -10.035 ;
        RECT -30.085 -11.725 -29.755 -11.395 ;
        RECT -30.085 -13.085 -29.755 -12.755 ;
        RECT -30.085 -14.445 -29.755 -14.115 ;
        RECT -30.085 -15.805 -29.755 -15.475 ;
        RECT -30.085 -17.165 -29.755 -16.835 ;
        RECT -30.085 -18.525 -29.755 -18.195 ;
        RECT -30.085 -25.325 -29.755 -24.995 ;
        RECT -30.085 -26.685 -29.755 -26.355 ;
        RECT -30.085 -28.045 -29.755 -27.715 ;
        RECT -30.085 -29.405 -29.755 -29.075 ;
        RECT -30.085 -30.765 -29.755 -30.435 ;
        RECT -30.085 -32.125 -29.755 -31.795 ;
        RECT -30.085 -33.485 -29.755 -33.155 ;
        RECT -30.085 -34.845 -29.755 -34.515 ;
        RECT -30.085 -36.205 -29.755 -35.875 ;
        RECT -30.085 -37.565 -29.755 -37.235 ;
        RECT -30.085 -38.925 -29.755 -38.595 ;
        RECT -30.085 -40.285 -29.755 -39.955 ;
        RECT -30.085 -44.365 -29.755 -44.035 ;
        RECT -30.085 -45.725 -29.755 -45.395 ;
        RECT -30.085 -47.085 -29.755 -46.755 ;
        RECT -30.085 -48.445 -29.755 -48.115 ;
        RECT -30.085 -49.805 -29.755 -49.475 ;
        RECT -30.085 -51.165 -29.755 -50.835 ;
        RECT -30.085 -52.525 -29.755 -52.195 ;
        RECT -30.085 -53.885 -29.755 -53.555 ;
        RECT -30.085 -55.245 -29.755 -54.915 ;
        RECT -30.085 -56.605 -29.755 -56.275 ;
        RECT -30.085 -57.965 -29.755 -57.635 ;
        RECT -30.085 -59.325 -29.755 -58.995 ;
        RECT -30.085 -60.685 -29.755 -60.355 ;
        RECT -30.085 -62.045 -29.755 -61.715 ;
        RECT -30.085 -63.405 -29.755 -63.075 ;
        RECT -30.085 -64.765 -29.755 -64.435 ;
        RECT -30.085 -65.91 -29.755 -65.58 ;
        RECT -30.085 -67.485 -29.755 -67.155 ;
        RECT -30.085 -68.845 -29.755 -68.515 ;
        RECT -30.085 -70.205 -29.755 -69.875 ;
        RECT -30.085 -71.565 -29.755 -71.235 ;
        RECT -30.085 -72.925 -29.755 -72.595 ;
        RECT -30.085 -75.645 -29.755 -75.315 ;
        RECT -30.085 -76.45 -29.755 -76.12 ;
        RECT -30.085 -78.365 -29.755 -78.035 ;
        RECT -30.085 -79.725 -29.755 -79.395 ;
        RECT -30.085 -81.085 -29.755 -80.755 ;
        RECT -30.085 -83.805 -29.755 -83.475 ;
        RECT -30.085 -85.165 -29.755 -84.835 ;
        RECT -30.08 -87.88 -29.76 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 -151.805 -29.755 -151.475 ;
        RECT -30.085 -153.165 -29.755 -152.835 ;
        RECT -30.085 -158.81 -29.755 -157.68 ;
        RECT -30.08 -158.925 -29.76 -149.44 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.725 44.8 -28.395 45.93 ;
        RECT -28.725 39.955 -28.395 40.285 ;
        RECT -28.725 38.595 -28.395 38.925 ;
        RECT -28.725 37.235 -28.395 37.565 ;
        RECT -28.725 35.875 -28.395 36.205 ;
        RECT -28.725 34.515 -28.395 34.845 ;
        RECT -28.725 33.155 -28.395 33.485 ;
        RECT -28.725 31.795 -28.395 32.125 ;
        RECT -28.725 30.435 -28.395 30.765 ;
        RECT -28.725 29.075 -28.395 29.405 ;
        RECT -28.725 27.715 -28.395 28.045 ;
        RECT -28.725 26.355 -28.395 26.685 ;
        RECT -28.725 24.995 -28.395 25.325 ;
        RECT -28.725 23.635 -28.395 23.965 ;
        RECT -28.725 22.275 -28.395 22.605 ;
        RECT -28.725 20.915 -28.395 21.245 ;
        RECT -28.725 19.555 -28.395 19.885 ;
        RECT -28.725 18.195 -28.395 18.525 ;
        RECT -28.725 16.835 -28.395 17.165 ;
        RECT -28.725 15.475 -28.395 15.805 ;
        RECT -28.725 14.115 -28.395 14.445 ;
        RECT -28.725 12.755 -28.395 13.085 ;
        RECT -28.725 11.395 -28.395 11.725 ;
        RECT -28.725 10.035 -28.395 10.365 ;
        RECT -28.725 8.675 -28.395 9.005 ;
        RECT -28.725 7.315 -28.395 7.645 ;
        RECT -28.725 5.955 -28.395 6.285 ;
        RECT -28.725 4.595 -28.395 4.925 ;
        RECT -28.725 3.235 -28.395 3.565 ;
        RECT -28.725 1.875 -28.395 2.205 ;
        RECT -28.725 -2.205 -28.395 -1.875 ;
        RECT -28.725 -4.925 -28.395 -4.595 ;
        RECT -28.725 -6.285 -28.395 -5.955 ;
        RECT -28.725 -7.645 -28.395 -7.315 ;
        RECT -28.725 -10.365 -28.395 -10.035 ;
        RECT -28.725 -11.725 -28.395 -11.395 ;
        RECT -28.725 -13.085 -28.395 -12.755 ;
        RECT -28.725 -14.445 -28.395 -14.115 ;
        RECT -28.725 -15.805 -28.395 -15.475 ;
        RECT -28.725 -17.165 -28.395 -16.835 ;
        RECT -28.725 -18.525 -28.395 -18.195 ;
        RECT -28.725 -25.325 -28.395 -24.995 ;
        RECT -28.725 -26.685 -28.395 -26.355 ;
        RECT -28.725 -28.045 -28.395 -27.715 ;
        RECT -28.725 -29.405 -28.395 -29.075 ;
        RECT -28.725 -30.765 -28.395 -30.435 ;
        RECT -28.725 -32.125 -28.395 -31.795 ;
        RECT -28.725 -33.485 -28.395 -33.155 ;
        RECT -28.725 -34.845 -28.395 -34.515 ;
        RECT -28.725 -36.205 -28.395 -35.875 ;
        RECT -28.725 -37.565 -28.395 -37.235 ;
        RECT -28.725 -38.925 -28.395 -38.595 ;
        RECT -28.725 -40.285 -28.395 -39.955 ;
        RECT -28.725 -44.365 -28.395 -44.035 ;
        RECT -28.725 -45.725 -28.395 -45.395 ;
        RECT -28.725 -47.085 -28.395 -46.755 ;
        RECT -28.725 -48.445 -28.395 -48.115 ;
        RECT -28.725 -49.805 -28.395 -49.475 ;
        RECT -28.725 -51.165 -28.395 -50.835 ;
        RECT -28.725 -52.525 -28.395 -52.195 ;
        RECT -28.725 -53.885 -28.395 -53.555 ;
        RECT -28.725 -55.245 -28.395 -54.915 ;
        RECT -28.725 -56.605 -28.395 -56.275 ;
        RECT -28.725 -57.965 -28.395 -57.635 ;
        RECT -28.725 -59.325 -28.395 -58.995 ;
        RECT -28.725 -60.685 -28.395 -60.355 ;
        RECT -28.725 -62.045 -28.395 -61.715 ;
        RECT -28.725 -63.405 -28.395 -63.075 ;
        RECT -28.725 -64.765 -28.395 -64.435 ;
        RECT -28.725 -65.91 -28.395 -65.58 ;
        RECT -28.725 -67.485 -28.395 -67.155 ;
        RECT -28.725 -68.845 -28.395 -68.515 ;
        RECT -28.725 -70.205 -28.395 -69.875 ;
        RECT -28.725 -71.565 -28.395 -71.235 ;
        RECT -28.725 -72.925 -28.395 -72.595 ;
        RECT -28.725 -75.645 -28.395 -75.315 ;
        RECT -28.725 -76.45 -28.395 -76.12 ;
        RECT -28.725 -78.365 -28.395 -78.035 ;
        RECT -28.725 -79.725 -28.395 -79.395 ;
        RECT -28.725 -81.085 -28.395 -80.755 ;
        RECT -28.725 -83.805 -28.395 -83.475 ;
        RECT -28.725 -85.165 -28.395 -84.835 ;
        RECT -28.725 -87.885 -28.395 -87.555 ;
        RECT -28.725 -89.245 -28.395 -88.915 ;
        RECT -28.725 -90.605 -28.395 -90.275 ;
        RECT -28.725 -91.965 -28.395 -91.635 ;
        RECT -28.725 -93.325 -28.395 -92.995 ;
        RECT -28.725 -94.685 -28.395 -94.355 ;
        RECT -28.725 -96.045 -28.395 -95.715 ;
        RECT -28.725 -97.405 -28.395 -97.075 ;
        RECT -28.725 -100.125 -28.395 -99.795 ;
        RECT -28.725 -101.485 -28.395 -101.155 ;
        RECT -28.725 -102.845 -28.395 -102.515 ;
        RECT -28.725 -104.205 -28.395 -103.875 ;
        RECT -28.725 -108.285 -28.395 -107.955 ;
        RECT -28.725 -109.645 -28.395 -109.315 ;
        RECT -28.725 -111.005 -28.395 -110.675 ;
        RECT -28.725 -113.725 -28.395 -113.395 ;
        RECT -28.725 -116.445 -28.395 -116.115 ;
        RECT -28.725 -117.805 -28.395 -117.475 ;
        RECT -28.725 -119.165 -28.395 -118.835 ;
        RECT -28.725 -120.525 -28.395 -120.195 ;
        RECT -28.725 -121.885 -28.395 -121.555 ;
        RECT -28.725 -123.245 -28.395 -122.915 ;
        RECT -28.725 -125.965 -28.395 -125.635 ;
        RECT -28.725 -127.325 -28.395 -126.995 ;
        RECT -28.725 -131.405 -28.395 -131.075 ;
        RECT -28.725 -132.765 -28.395 -132.435 ;
        RECT -28.725 -134.125 -28.395 -133.795 ;
        RECT -28.725 -135.485 -28.395 -135.155 ;
        RECT -28.725 -136.845 -28.395 -136.515 ;
        RECT -28.725 -138.205 -28.395 -137.875 ;
        RECT -28.725 -139.565 -28.395 -139.235 ;
        RECT -28.725 -140.925 -28.395 -140.595 ;
        RECT -28.725 -145.005 -28.395 -144.675 ;
        RECT -28.725 -146.365 -28.395 -146.035 ;
        RECT -28.725 -149.085 -28.395 -148.755 ;
        RECT -28.725 -151.805 -28.395 -151.475 ;
        RECT -28.725 -153.165 -28.395 -152.835 ;
        RECT -28.725 -158.81 -28.395 -157.68 ;
        RECT -28.72 -158.925 -28.4 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.365 44.8 -27.035 45.93 ;
        RECT -27.365 39.955 -27.035 40.285 ;
        RECT -27.365 38.595 -27.035 38.925 ;
        RECT -27.365 37.235 -27.035 37.565 ;
        RECT -27.365 35.875 -27.035 36.205 ;
        RECT -27.365 34.515 -27.035 34.845 ;
        RECT -27.365 33.155 -27.035 33.485 ;
        RECT -27.365 31.795 -27.035 32.125 ;
        RECT -27.365 30.435 -27.035 30.765 ;
        RECT -27.365 29.075 -27.035 29.405 ;
        RECT -27.365 27.715 -27.035 28.045 ;
        RECT -27.365 26.355 -27.035 26.685 ;
        RECT -27.365 24.995 -27.035 25.325 ;
        RECT -27.365 23.635 -27.035 23.965 ;
        RECT -27.365 22.275 -27.035 22.605 ;
        RECT -27.365 20.915 -27.035 21.245 ;
        RECT -27.365 19.555 -27.035 19.885 ;
        RECT -27.365 18.195 -27.035 18.525 ;
        RECT -27.365 16.835 -27.035 17.165 ;
        RECT -27.365 15.475 -27.035 15.805 ;
        RECT -27.365 14.115 -27.035 14.445 ;
        RECT -27.365 12.755 -27.035 13.085 ;
        RECT -27.365 11.395 -27.035 11.725 ;
        RECT -27.365 10.035 -27.035 10.365 ;
        RECT -27.365 8.675 -27.035 9.005 ;
        RECT -27.365 7.315 -27.035 7.645 ;
        RECT -27.365 5.955 -27.035 6.285 ;
        RECT -27.365 4.595 -27.035 4.925 ;
        RECT -27.365 3.235 -27.035 3.565 ;
        RECT -27.365 1.875 -27.035 2.205 ;
        RECT -27.365 -2.205 -27.035 -1.875 ;
        RECT -27.365 -4.925 -27.035 -4.595 ;
        RECT -27.365 -6.285 -27.035 -5.955 ;
        RECT -27.365 -7.645 -27.035 -7.315 ;
        RECT -27.365 -10.365 -27.035 -10.035 ;
        RECT -27.365 -11.725 -27.035 -11.395 ;
        RECT -27.365 -13.085 -27.035 -12.755 ;
        RECT -27.365 -14.445 -27.035 -14.115 ;
        RECT -27.365 -15.805 -27.035 -15.475 ;
        RECT -27.365 -17.165 -27.035 -16.835 ;
        RECT -27.365 -18.525 -27.035 -18.195 ;
        RECT -27.365 -25.325 -27.035 -24.995 ;
        RECT -27.365 -26.685 -27.035 -26.355 ;
        RECT -27.365 -28.045 -27.035 -27.715 ;
        RECT -27.365 -29.405 -27.035 -29.075 ;
        RECT -27.365 -30.765 -27.035 -30.435 ;
        RECT -27.365 -32.125 -27.035 -31.795 ;
        RECT -27.365 -33.485 -27.035 -33.155 ;
        RECT -27.365 -34.845 -27.035 -34.515 ;
        RECT -27.365 -36.205 -27.035 -35.875 ;
        RECT -27.365 -37.565 -27.035 -37.235 ;
        RECT -27.365 -38.925 -27.035 -38.595 ;
        RECT -27.365 -40.285 -27.035 -39.955 ;
        RECT -27.365 -44.365 -27.035 -44.035 ;
        RECT -27.365 -45.725 -27.035 -45.395 ;
        RECT -27.365 -47.085 -27.035 -46.755 ;
        RECT -27.365 -48.445 -27.035 -48.115 ;
        RECT -27.365 -49.805 -27.035 -49.475 ;
        RECT -27.365 -51.165 -27.035 -50.835 ;
        RECT -27.365 -52.525 -27.035 -52.195 ;
        RECT -27.365 -53.885 -27.035 -53.555 ;
        RECT -27.365 -55.245 -27.035 -54.915 ;
        RECT -27.365 -56.605 -27.035 -56.275 ;
        RECT -27.365 -57.965 -27.035 -57.635 ;
        RECT -27.365 -59.325 -27.035 -58.995 ;
        RECT -27.365 -60.685 -27.035 -60.355 ;
        RECT -27.365 -62.045 -27.035 -61.715 ;
        RECT -27.365 -63.405 -27.035 -63.075 ;
        RECT -27.365 -64.765 -27.035 -64.435 ;
        RECT -27.365 -65.91 -27.035 -65.58 ;
        RECT -27.365 -67.485 -27.035 -67.155 ;
        RECT -27.365 -68.845 -27.035 -68.515 ;
        RECT -27.365 -70.205 -27.035 -69.875 ;
        RECT -27.365 -71.565 -27.035 -71.235 ;
        RECT -27.365 -72.925 -27.035 -72.595 ;
        RECT -27.365 -75.645 -27.035 -75.315 ;
        RECT -27.365 -76.45 -27.035 -76.12 ;
        RECT -27.365 -78.365 -27.035 -78.035 ;
        RECT -27.365 -79.725 -27.035 -79.395 ;
        RECT -27.365 -81.085 -27.035 -80.755 ;
        RECT -27.365 -83.805 -27.035 -83.475 ;
        RECT -27.365 -85.165 -27.035 -84.835 ;
        RECT -27.365 -87.885 -27.035 -87.555 ;
        RECT -27.365 -89.245 -27.035 -88.915 ;
        RECT -27.365 -90.605 -27.035 -90.275 ;
        RECT -27.365 -91.965 -27.035 -91.635 ;
        RECT -27.365 -93.325 -27.035 -92.995 ;
        RECT -27.365 -94.685 -27.035 -94.355 ;
        RECT -27.365 -96.045 -27.035 -95.715 ;
        RECT -27.365 -97.405 -27.035 -97.075 ;
        RECT -27.365 -100.125 -27.035 -99.795 ;
        RECT -27.365 -101.485 -27.035 -101.155 ;
        RECT -27.365 -102.845 -27.035 -102.515 ;
        RECT -27.365 -104.205 -27.035 -103.875 ;
        RECT -27.365 -108.285 -27.035 -107.955 ;
        RECT -27.365 -109.645 -27.035 -109.315 ;
        RECT -27.365 -111.005 -27.035 -110.675 ;
        RECT -27.365 -113.725 -27.035 -113.395 ;
        RECT -27.365 -116.445 -27.035 -116.115 ;
        RECT -27.365 -117.805 -27.035 -117.475 ;
        RECT -27.365 -119.165 -27.035 -118.835 ;
        RECT -27.365 -120.525 -27.035 -120.195 ;
        RECT -27.365 -121.885 -27.035 -121.555 ;
        RECT -27.365 -123.245 -27.035 -122.915 ;
        RECT -27.365 -125.965 -27.035 -125.635 ;
        RECT -27.365 -127.325 -27.035 -126.995 ;
        RECT -27.365 -131.405 -27.035 -131.075 ;
        RECT -27.365 -132.765 -27.035 -132.435 ;
        RECT -27.365 -134.125 -27.035 -133.795 ;
        RECT -27.365 -135.485 -27.035 -135.155 ;
        RECT -27.365 -136.845 -27.035 -136.515 ;
        RECT -27.365 -138.205 -27.035 -137.875 ;
        RECT -27.365 -139.565 -27.035 -139.235 ;
        RECT -27.365 -140.925 -27.035 -140.595 ;
        RECT -27.365 -143.755 -27.035 -143.425 ;
        RECT -27.365 -145.005 -27.035 -144.675 ;
        RECT -27.365 -146.365 -27.035 -146.035 ;
        RECT -27.365 -149.085 -27.035 -148.755 ;
        RECT -27.365 -151.805 -27.035 -151.475 ;
        RECT -27.365 -153.165 -27.035 -152.835 ;
        RECT -27.365 -158.81 -27.035 -157.68 ;
        RECT -27.36 -158.925 -27.04 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.005 44.8 -25.675 45.93 ;
        RECT -26.005 39.955 -25.675 40.285 ;
        RECT -26.005 38.595 -25.675 38.925 ;
        RECT -26.005 37.235 -25.675 37.565 ;
        RECT -26.005 35.875 -25.675 36.205 ;
        RECT -26.005 34.515 -25.675 34.845 ;
        RECT -26.005 33.155 -25.675 33.485 ;
        RECT -26.005 31.795 -25.675 32.125 ;
        RECT -26.005 30.435 -25.675 30.765 ;
        RECT -26.005 29.075 -25.675 29.405 ;
        RECT -26.005 27.715 -25.675 28.045 ;
        RECT -26.005 26.355 -25.675 26.685 ;
        RECT -26.005 24.995 -25.675 25.325 ;
        RECT -26.005 23.635 -25.675 23.965 ;
        RECT -26.005 22.275 -25.675 22.605 ;
        RECT -26.005 20.915 -25.675 21.245 ;
        RECT -26.005 19.555 -25.675 19.885 ;
        RECT -26.005 18.195 -25.675 18.525 ;
        RECT -26.005 16.835 -25.675 17.165 ;
        RECT -26.005 15.475 -25.675 15.805 ;
        RECT -26.005 14.115 -25.675 14.445 ;
        RECT -26.005 12.755 -25.675 13.085 ;
        RECT -26.005 11.395 -25.675 11.725 ;
        RECT -26.005 10.035 -25.675 10.365 ;
        RECT -26.005 8.675 -25.675 9.005 ;
        RECT -26.005 7.315 -25.675 7.645 ;
        RECT -26.005 5.955 -25.675 6.285 ;
        RECT -26.005 4.595 -25.675 4.925 ;
        RECT -26.005 3.235 -25.675 3.565 ;
        RECT -26.005 1.875 -25.675 2.205 ;
        RECT -26.005 -2.205 -25.675 -1.875 ;
        RECT -26.005 -4.925 -25.675 -4.595 ;
        RECT -26.005 -6.285 -25.675 -5.955 ;
        RECT -26.005 -7.645 -25.675 -7.315 ;
        RECT -26.005 -10.365 -25.675 -10.035 ;
        RECT -26.005 -11.725 -25.675 -11.395 ;
        RECT -26.005 -13.085 -25.675 -12.755 ;
        RECT -26.005 -14.445 -25.675 -14.115 ;
        RECT -26.005 -15.805 -25.675 -15.475 ;
        RECT -26.005 -17.165 -25.675 -16.835 ;
        RECT -26.005 -18.525 -25.675 -18.195 ;
        RECT -26.005 -25.325 -25.675 -24.995 ;
        RECT -26.005 -26.685 -25.675 -26.355 ;
        RECT -26.005 -28.045 -25.675 -27.715 ;
        RECT -26.005 -29.405 -25.675 -29.075 ;
        RECT -26.005 -30.765 -25.675 -30.435 ;
        RECT -26.005 -32.125 -25.675 -31.795 ;
        RECT -26.005 -33.485 -25.675 -33.155 ;
        RECT -26.005 -34.845 -25.675 -34.515 ;
        RECT -26.005 -36.205 -25.675 -35.875 ;
        RECT -26.005 -37.565 -25.675 -37.235 ;
        RECT -26.005 -38.925 -25.675 -38.595 ;
        RECT -26.005 -40.285 -25.675 -39.955 ;
        RECT -26.005 -44.365 -25.675 -44.035 ;
        RECT -26.005 -45.725 -25.675 -45.395 ;
        RECT -26.005 -47.085 -25.675 -46.755 ;
        RECT -26.005 -48.445 -25.675 -48.115 ;
        RECT -26.005 -49.805 -25.675 -49.475 ;
        RECT -26.005 -51.165 -25.675 -50.835 ;
        RECT -26.005 -52.525 -25.675 -52.195 ;
        RECT -26.005 -53.885 -25.675 -53.555 ;
        RECT -26.005 -55.245 -25.675 -54.915 ;
        RECT -26.005 -56.605 -25.675 -56.275 ;
        RECT -26.005 -57.965 -25.675 -57.635 ;
        RECT -26.005 -59.325 -25.675 -58.995 ;
        RECT -26.005 -60.685 -25.675 -60.355 ;
        RECT -26.005 -62.045 -25.675 -61.715 ;
        RECT -26.005 -63.405 -25.675 -63.075 ;
        RECT -26.005 -64.765 -25.675 -64.435 ;
        RECT -26.005 -66.125 -25.675 -65.795 ;
        RECT -26.005 -67.485 -25.675 -67.155 ;
        RECT -26.005 -68.845 -25.675 -68.515 ;
        RECT -26.005 -70.205 -25.675 -69.875 ;
        RECT -26.005 -71.565 -25.675 -71.235 ;
        RECT -26.005 -72.925 -25.675 -72.595 ;
        RECT -26.005 -74.285 -25.675 -73.955 ;
        RECT -26.005 -75.645 -25.675 -75.315 ;
        RECT -26.005 -77.005 -25.675 -76.675 ;
        RECT -26.005 -78.365 -25.675 -78.035 ;
        RECT -26.005 -79.725 -25.675 -79.395 ;
        RECT -26.005 -81.085 -25.675 -80.755 ;
        RECT -26.005 -82.445 -25.675 -82.115 ;
        RECT -26.005 -83.805 -25.675 -83.475 ;
        RECT -26.005 -85.165 -25.675 -84.835 ;
        RECT -26.005 -86.525 -25.675 -86.195 ;
        RECT -26.005 -87.885 -25.675 -87.555 ;
        RECT -26.005 -89.245 -25.675 -88.915 ;
        RECT -26.005 -90.605 -25.675 -90.275 ;
        RECT -26.005 -91.965 -25.675 -91.635 ;
        RECT -26.005 -93.325 -25.675 -92.995 ;
        RECT -26.005 -94.685 -25.675 -94.355 ;
        RECT -26.005 -96.045 -25.675 -95.715 ;
        RECT -26.005 -97.405 -25.675 -97.075 ;
        RECT -26.005 -98.765 -25.675 -98.435 ;
        RECT -26.005 -100.125 -25.675 -99.795 ;
        RECT -26.005 -101.485 -25.675 -101.155 ;
        RECT -26.005 -102.845 -25.675 -102.515 ;
        RECT -26.005 -104.205 -25.675 -103.875 ;
        RECT -26.005 -109.645 -25.675 -109.315 ;
        RECT -26.005 -111.005 -25.675 -110.675 ;
        RECT -26.005 -113.725 -25.675 -113.395 ;
        RECT -26.005 -116.445 -25.675 -116.115 ;
        RECT -26.005 -117.805 -25.675 -117.475 ;
        RECT -26.005 -119.165 -25.675 -118.835 ;
        RECT -26.005 -121.885 -25.675 -121.555 ;
        RECT -26.005 -123.245 -25.675 -122.915 ;
        RECT -26.005 -125.965 -25.675 -125.635 ;
        RECT -26.005 -127.325 -25.675 -126.995 ;
        RECT -26.005 -131.405 -25.675 -131.075 ;
        RECT -26.005 -132.765 -25.675 -132.435 ;
        RECT -26.005 -134.125 -25.675 -133.795 ;
        RECT -26.005 -135.485 -25.675 -135.155 ;
        RECT -26.005 -136.845 -25.675 -136.515 ;
        RECT -26.005 -138.205 -25.675 -137.875 ;
        RECT -26.005 -139.565 -25.675 -139.235 ;
        RECT -26.005 -140.925 -25.675 -140.595 ;
        RECT -26.005 -143.755 -25.675 -143.425 ;
        RECT -26.005 -145.005 -25.675 -144.675 ;
        RECT -26.005 -146.365 -25.675 -146.035 ;
        RECT -26.005 -147.725 -25.675 -147.395 ;
        RECT -26.005 -149.085 -25.675 -148.755 ;
        RECT -26.005 -151.805 -25.675 -151.475 ;
        RECT -26.005 -153.165 -25.675 -152.835 ;
        RECT -26.005 -158.81 -25.675 -157.68 ;
        RECT -26 -158.925 -25.68 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.645 44.8 -24.315 45.93 ;
        RECT -24.645 39.955 -24.315 40.285 ;
        RECT -24.645 38.595 -24.315 38.925 ;
        RECT -24.645 37.235 -24.315 37.565 ;
        RECT -24.645 35.875 -24.315 36.205 ;
        RECT -24.645 34.515 -24.315 34.845 ;
        RECT -24.645 33.155 -24.315 33.485 ;
        RECT -24.645 31.795 -24.315 32.125 ;
        RECT -24.645 30.435 -24.315 30.765 ;
        RECT -24.645 29.075 -24.315 29.405 ;
        RECT -24.645 27.715 -24.315 28.045 ;
        RECT -24.645 26.355 -24.315 26.685 ;
        RECT -24.645 24.995 -24.315 25.325 ;
        RECT -24.645 23.635 -24.315 23.965 ;
        RECT -24.645 22.275 -24.315 22.605 ;
        RECT -24.645 20.915 -24.315 21.245 ;
        RECT -24.645 19.555 -24.315 19.885 ;
        RECT -24.645 18.195 -24.315 18.525 ;
        RECT -24.645 16.835 -24.315 17.165 ;
        RECT -24.645 15.475 -24.315 15.805 ;
        RECT -24.645 14.115 -24.315 14.445 ;
        RECT -24.645 12.755 -24.315 13.085 ;
        RECT -24.645 11.395 -24.315 11.725 ;
        RECT -24.645 10.035 -24.315 10.365 ;
        RECT -24.645 8.675 -24.315 9.005 ;
        RECT -24.645 7.315 -24.315 7.645 ;
        RECT -24.645 5.955 -24.315 6.285 ;
        RECT -24.645 4.595 -24.315 4.925 ;
        RECT -24.645 3.235 -24.315 3.565 ;
        RECT -24.645 1.875 -24.315 2.205 ;
        RECT -24.645 -2.205 -24.315 -1.875 ;
        RECT -24.645 -4.925 -24.315 -4.595 ;
        RECT -24.645 -6.285 -24.315 -5.955 ;
        RECT -24.645 -7.645 -24.315 -7.315 ;
        RECT -24.645 -10.365 -24.315 -10.035 ;
        RECT -24.645 -11.725 -24.315 -11.395 ;
        RECT -24.645 -13.085 -24.315 -12.755 ;
        RECT -24.645 -14.445 -24.315 -14.115 ;
        RECT -24.645 -15.805 -24.315 -15.475 ;
        RECT -24.645 -17.165 -24.315 -16.835 ;
        RECT -24.645 -18.525 -24.315 -18.195 ;
        RECT -24.645 -25.325 -24.315 -24.995 ;
        RECT -24.645 -26.685 -24.315 -26.355 ;
        RECT -24.645 -28.045 -24.315 -27.715 ;
        RECT -24.645 -29.405 -24.315 -29.075 ;
        RECT -24.645 -30.765 -24.315 -30.435 ;
        RECT -24.645 -32.125 -24.315 -31.795 ;
        RECT -24.645 -33.485 -24.315 -33.155 ;
        RECT -24.645 -34.845 -24.315 -34.515 ;
        RECT -24.645 -36.205 -24.315 -35.875 ;
        RECT -24.645 -37.565 -24.315 -37.235 ;
        RECT -24.645 -38.925 -24.315 -38.595 ;
        RECT -24.645 -40.285 -24.315 -39.955 ;
        RECT -24.645 -44.365 -24.315 -44.035 ;
        RECT -24.645 -45.725 -24.315 -45.395 ;
        RECT -24.645 -47.085 -24.315 -46.755 ;
        RECT -24.645 -48.445 -24.315 -48.115 ;
        RECT -24.645 -49.805 -24.315 -49.475 ;
        RECT -24.645 -51.165 -24.315 -50.835 ;
        RECT -24.645 -52.525 -24.315 -52.195 ;
        RECT -24.645 -53.885 -24.315 -53.555 ;
        RECT -24.645 -55.245 -24.315 -54.915 ;
        RECT -24.645 -56.605 -24.315 -56.275 ;
        RECT -24.645 -57.965 -24.315 -57.635 ;
        RECT -24.645 -59.325 -24.315 -58.995 ;
        RECT -24.645 -60.685 -24.315 -60.355 ;
        RECT -24.645 -62.045 -24.315 -61.715 ;
        RECT -24.645 -63.405 -24.315 -63.075 ;
        RECT -24.645 -64.765 -24.315 -64.435 ;
        RECT -24.645 -66.125 -24.315 -65.795 ;
        RECT -24.645 -67.485 -24.315 -67.155 ;
        RECT -24.645 -68.845 -24.315 -68.515 ;
        RECT -24.645 -70.205 -24.315 -69.875 ;
        RECT -24.645 -71.565 -24.315 -71.235 ;
        RECT -24.645 -72.925 -24.315 -72.595 ;
        RECT -24.645 -74.285 -24.315 -73.955 ;
        RECT -24.645 -75.645 -24.315 -75.315 ;
        RECT -24.645 -77.005 -24.315 -76.675 ;
        RECT -24.645 -78.365 -24.315 -78.035 ;
        RECT -24.645 -79.725 -24.315 -79.395 ;
        RECT -24.645 -81.085 -24.315 -80.755 ;
        RECT -24.645 -82.445 -24.315 -82.115 ;
        RECT -24.645 -83.805 -24.315 -83.475 ;
        RECT -24.645 -85.165 -24.315 -84.835 ;
        RECT -24.645 -86.525 -24.315 -86.195 ;
        RECT -24.645 -87.885 -24.315 -87.555 ;
        RECT -24.645 -89.245 -24.315 -88.915 ;
        RECT -24.645 -90.605 -24.315 -90.275 ;
        RECT -24.645 -91.965 -24.315 -91.635 ;
        RECT -24.645 -93.325 -24.315 -92.995 ;
        RECT -24.645 -94.685 -24.315 -94.355 ;
        RECT -24.645 -96.045 -24.315 -95.715 ;
        RECT -24.645 -97.405 -24.315 -97.075 ;
        RECT -24.645 -98.765 -24.315 -98.435 ;
        RECT -24.645 -100.125 -24.315 -99.795 ;
        RECT -24.645 -101.485 -24.315 -101.155 ;
        RECT -24.645 -102.845 -24.315 -102.515 ;
        RECT -24.645 -109.645 -24.315 -109.315 ;
        RECT -24.645 -111.005 -24.315 -110.675 ;
        RECT -24.645 -113.725 -24.315 -113.395 ;
        RECT -24.645 -116.445 -24.315 -116.115 ;
        RECT -24.645 -117.805 -24.315 -117.475 ;
        RECT -24.645 -121.885 -24.315 -121.555 ;
        RECT -24.645 -123.245 -24.315 -122.915 ;
        RECT -24.645 -125.965 -24.315 -125.635 ;
        RECT -24.645 -127.325 -24.315 -126.995 ;
        RECT -24.645 -132.765 -24.315 -132.435 ;
        RECT -24.645 -134.125 -24.315 -133.795 ;
        RECT -24.645 -135.485 -24.315 -135.155 ;
        RECT -24.645 -136.845 -24.315 -136.515 ;
        RECT -24.645 -138.205 -24.315 -137.875 ;
        RECT -24.645 -139.565 -24.315 -139.235 ;
        RECT -24.645 -140.925 -24.315 -140.595 ;
        RECT -24.645 -143.755 -24.315 -143.425 ;
        RECT -24.645 -145.005 -24.315 -144.675 ;
        RECT -24.645 -146.365 -24.315 -146.035 ;
        RECT -24.645 -147.725 -24.315 -147.395 ;
        RECT -24.645 -149.085 -24.315 -148.755 ;
        RECT -24.645 -151.805 -24.315 -151.475 ;
        RECT -24.645 -153.165 -24.315 -152.835 ;
        RECT -24.645 -158.81 -24.315 -157.68 ;
        RECT -24.64 -158.925 -24.32 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.285 44.8 -22.955 45.93 ;
        RECT -23.285 39.955 -22.955 40.285 ;
        RECT -23.285 38.595 -22.955 38.925 ;
        RECT -23.285 37.235 -22.955 37.565 ;
        RECT -23.285 35.875 -22.955 36.205 ;
        RECT -23.285 34.515 -22.955 34.845 ;
        RECT -23.285 33.155 -22.955 33.485 ;
        RECT -23.285 31.795 -22.955 32.125 ;
        RECT -23.285 30.435 -22.955 30.765 ;
        RECT -23.285 29.075 -22.955 29.405 ;
        RECT -23.285 27.715 -22.955 28.045 ;
        RECT -23.285 26.355 -22.955 26.685 ;
        RECT -23.285 24.995 -22.955 25.325 ;
        RECT -23.285 23.635 -22.955 23.965 ;
        RECT -23.285 22.275 -22.955 22.605 ;
        RECT -23.285 20.915 -22.955 21.245 ;
        RECT -23.285 19.555 -22.955 19.885 ;
        RECT -23.285 18.195 -22.955 18.525 ;
        RECT -23.285 16.835 -22.955 17.165 ;
        RECT -23.285 15.475 -22.955 15.805 ;
        RECT -23.285 14.115 -22.955 14.445 ;
        RECT -23.285 12.755 -22.955 13.085 ;
        RECT -23.285 11.395 -22.955 11.725 ;
        RECT -23.285 10.035 -22.955 10.365 ;
        RECT -23.285 8.675 -22.955 9.005 ;
        RECT -23.285 7.315 -22.955 7.645 ;
        RECT -23.285 5.955 -22.955 6.285 ;
        RECT -23.285 4.595 -22.955 4.925 ;
        RECT -23.285 3.235 -22.955 3.565 ;
        RECT -23.285 1.875 -22.955 2.205 ;
        RECT -23.285 -2.205 -22.955 -1.875 ;
        RECT -23.285 -4.925 -22.955 -4.595 ;
        RECT -23.285 -6.285 -22.955 -5.955 ;
        RECT -23.285 -7.645 -22.955 -7.315 ;
        RECT -23.285 -10.365 -22.955 -10.035 ;
        RECT -23.285 -11.725 -22.955 -11.395 ;
        RECT -23.285 -13.085 -22.955 -12.755 ;
        RECT -23.285 -14.445 -22.955 -14.115 ;
        RECT -23.285 -15.805 -22.955 -15.475 ;
        RECT -23.285 -17.165 -22.955 -16.835 ;
        RECT -23.285 -18.525 -22.955 -18.195 ;
        RECT -23.285 -25.325 -22.955 -24.995 ;
        RECT -23.285 -26.685 -22.955 -26.355 ;
        RECT -23.285 -28.045 -22.955 -27.715 ;
        RECT -23.285 -29.405 -22.955 -29.075 ;
        RECT -23.285 -30.765 -22.955 -30.435 ;
        RECT -23.285 -32.125 -22.955 -31.795 ;
        RECT -23.285 -33.485 -22.955 -33.155 ;
        RECT -23.285 -34.845 -22.955 -34.515 ;
        RECT -23.285 -36.205 -22.955 -35.875 ;
        RECT -23.285 -37.565 -22.955 -37.235 ;
        RECT -23.285 -38.925 -22.955 -38.595 ;
        RECT -23.285 -40.285 -22.955 -39.955 ;
        RECT -23.285 -44.365 -22.955 -44.035 ;
        RECT -23.285 -45.725 -22.955 -45.395 ;
        RECT -23.285 -47.085 -22.955 -46.755 ;
        RECT -23.285 -48.445 -22.955 -48.115 ;
        RECT -23.285 -49.805 -22.955 -49.475 ;
        RECT -23.285 -51.165 -22.955 -50.835 ;
        RECT -23.285 -52.525 -22.955 -52.195 ;
        RECT -23.285 -53.885 -22.955 -53.555 ;
        RECT -23.285 -55.245 -22.955 -54.915 ;
        RECT -23.285 -56.605 -22.955 -56.275 ;
        RECT -23.285 -57.965 -22.955 -57.635 ;
        RECT -23.285 -59.325 -22.955 -58.995 ;
        RECT -23.285 -60.685 -22.955 -60.355 ;
        RECT -23.285 -62.045 -22.955 -61.715 ;
        RECT -23.285 -63.405 -22.955 -63.075 ;
        RECT -23.285 -64.765 -22.955 -64.435 ;
        RECT -23.285 -66.125 -22.955 -65.795 ;
        RECT -23.285 -67.485 -22.955 -67.155 ;
        RECT -23.285 -68.845 -22.955 -68.515 ;
        RECT -23.285 -70.205 -22.955 -69.875 ;
        RECT -23.285 -71.565 -22.955 -71.235 ;
        RECT -23.285 -72.925 -22.955 -72.595 ;
        RECT -23.285 -74.285 -22.955 -73.955 ;
        RECT -23.285 -75.645 -22.955 -75.315 ;
        RECT -23.285 -77.005 -22.955 -76.675 ;
        RECT -23.285 -78.365 -22.955 -78.035 ;
        RECT -23.285 -79.725 -22.955 -79.395 ;
        RECT -23.285 -81.085 -22.955 -80.755 ;
        RECT -23.285 -82.445 -22.955 -82.115 ;
        RECT -23.285 -83.805 -22.955 -83.475 ;
        RECT -23.285 -85.165 -22.955 -84.835 ;
        RECT -23.285 -86.525 -22.955 -86.195 ;
        RECT -23.28 -87.2 -22.96 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.285 -151.805 -22.955 -151.475 ;
        RECT -23.285 -153.165 -22.955 -152.835 ;
        RECT -23.285 -158.81 -22.955 -157.68 ;
        RECT -23.28 -158.925 -22.96 -147.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 44.8 -21.595 45.93 ;
        RECT -21.925 39.955 -21.595 40.285 ;
        RECT -21.925 38.595 -21.595 38.925 ;
        RECT -21.925 37.235 -21.595 37.565 ;
        RECT -21.925 35.875 -21.595 36.205 ;
        RECT -21.925 34.515 -21.595 34.845 ;
        RECT -21.925 33.155 -21.595 33.485 ;
        RECT -21.925 31.795 -21.595 32.125 ;
        RECT -21.925 30.435 -21.595 30.765 ;
        RECT -21.925 29.075 -21.595 29.405 ;
        RECT -21.925 27.715 -21.595 28.045 ;
        RECT -21.925 26.355 -21.595 26.685 ;
        RECT -21.925 24.995 -21.595 25.325 ;
        RECT -21.925 23.635 -21.595 23.965 ;
        RECT -21.925 22.275 -21.595 22.605 ;
        RECT -21.925 20.915 -21.595 21.245 ;
        RECT -21.925 19.555 -21.595 19.885 ;
        RECT -21.925 18.195 -21.595 18.525 ;
        RECT -21.925 16.835 -21.595 17.165 ;
        RECT -21.925 15.475 -21.595 15.805 ;
        RECT -21.925 14.115 -21.595 14.445 ;
        RECT -21.925 12.755 -21.595 13.085 ;
        RECT -21.925 11.395 -21.595 11.725 ;
        RECT -21.925 10.035 -21.595 10.365 ;
        RECT -21.925 8.675 -21.595 9.005 ;
        RECT -21.925 7.315 -21.595 7.645 ;
        RECT -21.925 5.955 -21.595 6.285 ;
        RECT -21.925 4.595 -21.595 4.925 ;
        RECT -21.925 3.235 -21.595 3.565 ;
        RECT -21.925 1.875 -21.595 2.205 ;
        RECT -21.925 -2.205 -21.595 -1.875 ;
        RECT -21.925 -4.925 -21.595 -4.595 ;
        RECT -21.925 -6.285 -21.595 -5.955 ;
        RECT -21.925 -7.645 -21.595 -7.315 ;
        RECT -21.925 -10.365 -21.595 -10.035 ;
        RECT -21.925 -11.725 -21.595 -11.395 ;
        RECT -21.925 -13.085 -21.595 -12.755 ;
        RECT -21.925 -14.445 -21.595 -14.115 ;
        RECT -21.925 -15.805 -21.595 -15.475 ;
        RECT -21.925 -17.165 -21.595 -16.835 ;
        RECT -21.925 -18.525 -21.595 -18.195 ;
        RECT -21.925 -25.325 -21.595 -24.995 ;
        RECT -21.925 -26.685 -21.595 -26.355 ;
        RECT -21.925 -28.045 -21.595 -27.715 ;
        RECT -21.925 -29.405 -21.595 -29.075 ;
        RECT -21.925 -30.765 -21.595 -30.435 ;
        RECT -21.925 -32.125 -21.595 -31.795 ;
        RECT -21.925 -33.485 -21.595 -33.155 ;
        RECT -21.925 -34.845 -21.595 -34.515 ;
        RECT -21.925 -36.205 -21.595 -35.875 ;
        RECT -21.925 -37.565 -21.595 -37.235 ;
        RECT -21.925 -38.925 -21.595 -38.595 ;
        RECT -21.925 -40.285 -21.595 -39.955 ;
        RECT -21.925 -44.365 -21.595 -44.035 ;
        RECT -21.925 -45.725 -21.595 -45.395 ;
        RECT -21.925 -47.085 -21.595 -46.755 ;
        RECT -21.925 -48.445 -21.595 -48.115 ;
        RECT -21.925 -49.805 -21.595 -49.475 ;
        RECT -21.925 -51.165 -21.595 -50.835 ;
        RECT -21.925 -52.525 -21.595 -52.195 ;
        RECT -21.925 -53.885 -21.595 -53.555 ;
        RECT -21.925 -55.245 -21.595 -54.915 ;
        RECT -21.925 -56.605 -21.595 -56.275 ;
        RECT -21.925 -57.965 -21.595 -57.635 ;
        RECT -21.925 -59.325 -21.595 -58.995 ;
        RECT -21.925 -60.685 -21.595 -60.355 ;
        RECT -21.925 -62.045 -21.595 -61.715 ;
        RECT -21.925 -63.405 -21.595 -63.075 ;
        RECT -21.925 -64.765 -21.595 -64.435 ;
        RECT -21.925 -66.125 -21.595 -65.795 ;
        RECT -21.925 -67.485 -21.595 -67.155 ;
        RECT -21.925 -68.845 -21.595 -68.515 ;
        RECT -21.925 -70.205 -21.595 -69.875 ;
        RECT -21.925 -71.565 -21.595 -71.235 ;
        RECT -21.925 -72.925 -21.595 -72.595 ;
        RECT -21.925 -74.285 -21.595 -73.955 ;
        RECT -21.925 -75.645 -21.595 -75.315 ;
        RECT -21.925 -77.005 -21.595 -76.675 ;
        RECT -21.925 -78.365 -21.595 -78.035 ;
        RECT -21.925 -79.725 -21.595 -79.395 ;
        RECT -21.925 -81.085 -21.595 -80.755 ;
        RECT -21.925 -82.445 -21.595 -82.115 ;
        RECT -21.925 -83.805 -21.595 -83.475 ;
        RECT -21.925 -85.165 -21.595 -84.835 ;
        RECT -21.925 -86.525 -21.595 -86.195 ;
        RECT -21.925 -89.245 -21.595 -88.915 ;
        RECT -21.925 -90.605 -21.595 -90.275 ;
        RECT -21.925 -91.965 -21.595 -91.635 ;
        RECT -21.925 -93.325 -21.595 -92.995 ;
        RECT -21.925 -94.685 -21.595 -94.355 ;
        RECT -21.925 -96.045 -21.595 -95.715 ;
        RECT -21.925 -97.405 -21.595 -97.075 ;
        RECT -21.925 -98.765 -21.595 -98.435 ;
        RECT -21.925 -100.125 -21.595 -99.795 ;
        RECT -21.925 -101.485 -21.595 -101.155 ;
        RECT -21.925 -102.845 -21.595 -102.515 ;
        RECT -21.925 -109.645 -21.595 -109.315 ;
        RECT -21.925 -113.725 -21.595 -113.395 ;
        RECT -21.925 -116.445 -21.595 -116.115 ;
        RECT -21.925 -117.805 -21.595 -117.475 ;
        RECT -21.925 -121.885 -21.595 -121.555 ;
        RECT -21.925 -123.245 -21.595 -122.915 ;
        RECT -21.925 -125.965 -21.595 -125.635 ;
        RECT -21.925 -127.325 -21.595 -126.995 ;
        RECT -21.925 -132.765 -21.595 -132.435 ;
        RECT -21.925 -134.125 -21.595 -133.795 ;
        RECT -21.925 -135.485 -21.595 -135.155 ;
        RECT -21.925 -136.845 -21.595 -136.515 ;
        RECT -21.925 -138.205 -21.595 -137.875 ;
        RECT -21.925 -139.565 -21.595 -139.235 ;
        RECT -21.925 -140.925 -21.595 -140.595 ;
        RECT -21.925 -143.755 -21.595 -143.425 ;
        RECT -21.925 -145.005 -21.595 -144.675 ;
        RECT -21.925 -146.365 -21.595 -146.035 ;
        RECT -21.92 -147.04 -21.6 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 -101.485 -20.235 -101.155 ;
        RECT -20.565 -102.845 -20.235 -102.515 ;
        RECT -20.565 -109.645 -20.235 -109.315 ;
        RECT -20.565 -113.725 -20.235 -113.395 ;
        RECT -20.565 -116.445 -20.235 -116.115 ;
        RECT -20.565 -119.165 -20.235 -118.835 ;
        RECT -20.565 -121.885 -20.235 -121.555 ;
        RECT -20.565 -123.245 -20.235 -122.915 ;
        RECT -20.565 -125.965 -20.235 -125.635 ;
        RECT -20.565 -127.325 -20.235 -126.995 ;
        RECT -20.565 -132.765 -20.235 -132.435 ;
        RECT -20.565 -134.125 -20.235 -133.795 ;
        RECT -20.565 -135.485 -20.235 -135.155 ;
        RECT -20.565 -136.845 -20.235 -136.515 ;
        RECT -20.565 -138.205 -20.235 -137.875 ;
        RECT -20.565 -139.565 -20.235 -139.235 ;
        RECT -20.565 -140.925 -20.235 -140.595 ;
        RECT -20.56 -141.6 -20.24 46.045 ;
        RECT -20.565 44.8 -20.235 45.93 ;
        RECT -20.565 39.955 -20.235 40.285 ;
        RECT -20.565 38.595 -20.235 38.925 ;
        RECT -20.565 37.235 -20.235 37.565 ;
        RECT -20.565 35.875 -20.235 36.205 ;
        RECT -20.565 34.515 -20.235 34.845 ;
        RECT -20.565 33.155 -20.235 33.485 ;
        RECT -20.565 31.795 -20.235 32.125 ;
        RECT -20.565 30.435 -20.235 30.765 ;
        RECT -20.565 29.075 -20.235 29.405 ;
        RECT -20.565 27.715 -20.235 28.045 ;
        RECT -20.565 26.355 -20.235 26.685 ;
        RECT -20.565 24.995 -20.235 25.325 ;
        RECT -20.565 23.635 -20.235 23.965 ;
        RECT -20.565 22.275 -20.235 22.605 ;
        RECT -20.565 20.915 -20.235 21.245 ;
        RECT -20.565 19.555 -20.235 19.885 ;
        RECT -20.565 18.195 -20.235 18.525 ;
        RECT -20.565 16.835 -20.235 17.165 ;
        RECT -20.565 15.475 -20.235 15.805 ;
        RECT -20.565 14.115 -20.235 14.445 ;
        RECT -20.565 12.755 -20.235 13.085 ;
        RECT -20.565 11.395 -20.235 11.725 ;
        RECT -20.565 10.035 -20.235 10.365 ;
        RECT -20.565 8.675 -20.235 9.005 ;
        RECT -20.565 7.315 -20.235 7.645 ;
        RECT -20.565 5.955 -20.235 6.285 ;
        RECT -20.565 4.595 -20.235 4.925 ;
        RECT -20.565 3.235 -20.235 3.565 ;
        RECT -20.565 1.875 -20.235 2.205 ;
        RECT -20.565 -2.205 -20.235 -1.875 ;
        RECT -20.565 -4.925 -20.235 -4.595 ;
        RECT -20.565 -5.65 -20.235 -5.32 ;
        RECT -20.565 -7.645 -20.235 -7.315 ;
        RECT -20.565 -11.69 -20.235 -11.36 ;
        RECT -20.565 -13.085 -20.235 -12.755 ;
        RECT -20.565 -15.805 -20.235 -15.475 ;
        RECT -20.565 -25.325 -20.235 -24.995 ;
        RECT -20.565 -26.685 -20.235 -26.355 ;
        RECT -20.565 -27.67 -20.235 -27.34 ;
        RECT -20.565 -29.405 -20.235 -29.075 ;
        RECT -20.565 -30.765 -20.235 -30.435 ;
        RECT -20.565 -33.71 -20.235 -33.38 ;
        RECT -20.565 -34.845 -20.235 -34.515 ;
        RECT -20.565 -37.565 -20.235 -37.235 ;
        RECT -20.565 -44.365 -20.235 -44.035 ;
        RECT -20.565 -45.725 -20.235 -45.395 ;
        RECT -20.565 -47.085 -20.235 -46.755 ;
        RECT -20.565 -48.29 -20.235 -47.96 ;
        RECT -20.565 -49.805 -20.235 -49.475 ;
        RECT -20.565 -52.525 -20.235 -52.195 ;
        RECT -20.565 -53.885 -20.235 -53.555 ;
        RECT -20.565 -55.83 -20.235 -55.5 ;
        RECT -20.565 -56.605 -20.235 -56.275 ;
        RECT -20.565 -57.965 -20.235 -57.635 ;
        RECT -20.565 -59.325 -20.235 -58.995 ;
        RECT -20.565 -62.045 -20.235 -61.715 ;
        RECT -20.565 -64.765 -20.235 -64.435 ;
        RECT -20.565 -66.125 -20.235 -65.795 ;
        RECT -20.565 -67.485 -20.235 -67.155 ;
        RECT -20.565 -68.845 -20.235 -68.515 ;
        RECT -20.565 -70.47 -20.235 -70.14 ;
        RECT -20.565 -71.565 -20.235 -71.235 ;
        RECT -20.565 -72.925 -20.235 -72.595 ;
        RECT -20.565 -75.645 -20.235 -75.315 ;
        RECT -20.565 -77.005 -20.235 -76.675 ;
        RECT -20.565 -78.01 -20.235 -77.68 ;
        RECT -20.565 -79.725 -20.235 -79.395 ;
        RECT -20.565 -81.085 -20.235 -80.755 ;
        RECT -20.565 -83.805 -20.235 -83.475 ;
        RECT -20.565 -89.245 -20.235 -88.915 ;
        RECT -20.565 -90.605 -20.235 -90.275 ;
        RECT -20.565 -91.965 -20.235 -91.635 ;
        RECT -20.565 -93.325 -20.235 -92.995 ;
        RECT -20.565 -96.045 -20.235 -95.715 ;
        RECT -20.565 -98.765 -20.235 -98.435 ;
        RECT -20.565 -100.125 -20.235 -99.795 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.325 44.8 -41.995 45.93 ;
        RECT -42.325 39.955 -41.995 40.285 ;
        RECT -42.325 38.595 -41.995 38.925 ;
        RECT -42.325 37.235 -41.995 37.565 ;
        RECT -42.325 35.875 -41.995 36.205 ;
        RECT -42.325 34.515 -41.995 34.845 ;
        RECT -42.325 33.155 -41.995 33.485 ;
        RECT -42.325 31.795 -41.995 32.125 ;
        RECT -42.325 30.435 -41.995 30.765 ;
        RECT -42.325 29.075 -41.995 29.405 ;
        RECT -42.325 27.715 -41.995 28.045 ;
        RECT -42.325 26.355 -41.995 26.685 ;
        RECT -42.325 24.995 -41.995 25.325 ;
        RECT -42.325 22.66 -41.995 22.99 ;
        RECT -42.325 20.485 -41.995 20.815 ;
        RECT -42.325 19.635 -41.995 19.965 ;
        RECT -42.325 17.325 -41.995 17.655 ;
        RECT -42.325 16.475 -41.995 16.805 ;
        RECT -42.325 14.3 -41.995 14.63 ;
        RECT -42.325 11.395 -41.995 11.725 ;
        RECT -42.325 10.035 -41.995 10.365 ;
        RECT -42.325 8.675 -41.995 9.005 ;
        RECT -42.325 7.315 -41.995 7.645 ;
        RECT -42.325 5.955 -41.995 6.285 ;
        RECT -42.325 4.595 -41.995 4.925 ;
        RECT -42.325 3.235 -41.995 3.565 ;
        RECT -42.325 1.875 -41.995 2.205 ;
        RECT -42.325 0.515 -41.995 0.845 ;
        RECT -42.325 -0.845 -41.995 -0.515 ;
        RECT -42.325 -2.205 -41.995 -1.875 ;
        RECT -42.325 -4.925 -41.995 -4.595 ;
        RECT -42.325 -6.285 -41.995 -5.955 ;
        RECT -42.325 -7.645 -41.995 -7.315 ;
        RECT -42.325 -10.365 -41.995 -10.035 ;
        RECT -42.325 -11.725 -41.995 -11.395 ;
        RECT -42.325 -13.085 -41.995 -12.755 ;
        RECT -42.325 -14.445 -41.995 -14.115 ;
        RECT -42.325 -15.805 -41.995 -15.475 ;
        RECT -42.325 -17.165 -41.995 -16.835 ;
        RECT -42.325 -18.525 -41.995 -18.195 ;
        RECT -42.325 -21.245 -41.995 -20.915 ;
        RECT -42.325 -22.605 -41.995 -22.275 ;
        RECT -42.325 -23.965 -41.995 -23.635 ;
        RECT -42.325 -25.325 -41.995 -24.995 ;
        RECT -42.325 -26.685 -41.995 -26.355 ;
        RECT -42.325 -28.045 -41.995 -27.715 ;
        RECT -42.325 -29.405 -41.995 -29.075 ;
        RECT -42.325 -30.765 -41.995 -30.435 ;
        RECT -42.325 -32.125 -41.995 -31.795 ;
        RECT -42.325 -33.485 -41.995 -33.155 ;
        RECT -42.325 -34.845 -41.995 -34.515 ;
        RECT -42.325 -36.205 -41.995 -35.875 ;
        RECT -42.325 -37.565 -41.995 -37.235 ;
        RECT -42.325 -38.925 -41.995 -38.595 ;
        RECT -42.325 -40.285 -41.995 -39.955 ;
        RECT -42.325 -41.645 -41.995 -41.315 ;
        RECT -42.325 -43.005 -41.995 -42.675 ;
        RECT -42.325 -44.365 -41.995 -44.035 ;
        RECT -42.325 -45.725 -41.995 -45.395 ;
        RECT -42.325 -47.085 -41.995 -46.755 ;
        RECT -42.325 -48.445 -41.995 -48.115 ;
        RECT -42.325 -49.805 -41.995 -49.475 ;
        RECT -42.325 -51.165 -41.995 -50.835 ;
        RECT -42.325 -52.525 -41.995 -52.195 ;
        RECT -42.325 -53.885 -41.995 -53.555 ;
        RECT -42.325 -55.245 -41.995 -54.915 ;
        RECT -42.325 -56.605 -41.995 -56.275 ;
        RECT -42.325 -57.965 -41.995 -57.635 ;
        RECT -42.325 -59.325 -41.995 -58.995 ;
        RECT -42.325 -60.685 -41.995 -60.355 ;
        RECT -42.325 -62.045 -41.995 -61.715 ;
        RECT -42.325 -63.405 -41.995 -63.075 ;
        RECT -42.325 -64.765 -41.995 -64.435 ;
        RECT -42.325 -65.91 -41.995 -65.58 ;
        RECT -42.325 -67.485 -41.995 -67.155 ;
        RECT -42.325 -68.845 -41.995 -68.515 ;
        RECT -42.325 -70.205 -41.995 -69.875 ;
        RECT -42.325 -71.565 -41.995 -71.235 ;
        RECT -42.325 -72.925 -41.995 -72.595 ;
        RECT -42.325 -75.645 -41.995 -75.315 ;
        RECT -42.325 -76.45 -41.995 -76.12 ;
        RECT -42.325 -78.365 -41.995 -78.035 ;
        RECT -42.325 -79.725 -41.995 -79.395 ;
        RECT -42.325 -81.085 -41.995 -80.755 ;
        RECT -42.325 -83.805 -41.995 -83.475 ;
        RECT -42.325 -85.165 -41.995 -84.835 ;
        RECT -42.325 -87.885 -41.995 -87.555 ;
        RECT -42.32 -87.885 -42 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.325 -151.805 -41.995 -151.475 ;
        RECT -42.325 -153.165 -41.995 -152.835 ;
        RECT -42.325 -158.81 -41.995 -157.68 ;
        RECT -42.32 -158.925 -42 -149.44 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.965 44.8 -40.635 45.93 ;
        RECT -40.965 39.955 -40.635 40.285 ;
        RECT -40.965 38.595 -40.635 38.925 ;
        RECT -40.965 37.235 -40.635 37.565 ;
        RECT -40.965 35.875 -40.635 36.205 ;
        RECT -40.965 34.515 -40.635 34.845 ;
        RECT -40.965 33.155 -40.635 33.485 ;
        RECT -40.965 31.795 -40.635 32.125 ;
        RECT -40.965 30.435 -40.635 30.765 ;
        RECT -40.965 29.075 -40.635 29.405 ;
        RECT -40.965 27.715 -40.635 28.045 ;
        RECT -40.965 26.355 -40.635 26.685 ;
        RECT -40.965 24.995 -40.635 25.325 ;
        RECT -40.965 22.66 -40.635 22.99 ;
        RECT -40.965 20.485 -40.635 20.815 ;
        RECT -40.965 19.635 -40.635 19.965 ;
        RECT -40.965 17.325 -40.635 17.655 ;
        RECT -40.965 16.475 -40.635 16.805 ;
        RECT -40.965 14.3 -40.635 14.63 ;
        RECT -40.965 11.395 -40.635 11.725 ;
        RECT -40.965 10.035 -40.635 10.365 ;
        RECT -40.965 8.675 -40.635 9.005 ;
        RECT -40.965 7.315 -40.635 7.645 ;
        RECT -40.965 5.955 -40.635 6.285 ;
        RECT -40.965 4.595 -40.635 4.925 ;
        RECT -40.965 3.235 -40.635 3.565 ;
        RECT -40.965 1.875 -40.635 2.205 ;
        RECT -40.965 0.515 -40.635 0.845 ;
        RECT -40.965 -0.845 -40.635 -0.515 ;
        RECT -40.965 -2.205 -40.635 -1.875 ;
        RECT -40.965 -4.925 -40.635 -4.595 ;
        RECT -40.965 -6.285 -40.635 -5.955 ;
        RECT -40.965 -7.645 -40.635 -7.315 ;
        RECT -40.965 -10.365 -40.635 -10.035 ;
        RECT -40.965 -11.725 -40.635 -11.395 ;
        RECT -40.965 -13.085 -40.635 -12.755 ;
        RECT -40.965 -14.445 -40.635 -14.115 ;
        RECT -40.965 -15.805 -40.635 -15.475 ;
        RECT -40.965 -17.165 -40.635 -16.835 ;
        RECT -40.965 -18.525 -40.635 -18.195 ;
        RECT -40.965 -21.245 -40.635 -20.915 ;
        RECT -40.965 -22.605 -40.635 -22.275 ;
        RECT -40.965 -25.325 -40.635 -24.995 ;
        RECT -40.965 -26.685 -40.635 -26.355 ;
        RECT -40.965 -28.045 -40.635 -27.715 ;
        RECT -40.965 -29.405 -40.635 -29.075 ;
        RECT -40.965 -30.765 -40.635 -30.435 ;
        RECT -40.965 -32.125 -40.635 -31.795 ;
        RECT -40.965 -33.485 -40.635 -33.155 ;
        RECT -40.965 -34.845 -40.635 -34.515 ;
        RECT -40.965 -36.205 -40.635 -35.875 ;
        RECT -40.965 -37.565 -40.635 -37.235 ;
        RECT -40.965 -38.925 -40.635 -38.595 ;
        RECT -40.965 -40.285 -40.635 -39.955 ;
        RECT -40.965 -41.645 -40.635 -41.315 ;
        RECT -40.965 -43.005 -40.635 -42.675 ;
        RECT -40.965 -44.365 -40.635 -44.035 ;
        RECT -40.965 -45.725 -40.635 -45.395 ;
        RECT -40.965 -47.085 -40.635 -46.755 ;
        RECT -40.965 -48.445 -40.635 -48.115 ;
        RECT -40.965 -49.805 -40.635 -49.475 ;
        RECT -40.965 -51.165 -40.635 -50.835 ;
        RECT -40.965 -52.525 -40.635 -52.195 ;
        RECT -40.965 -53.885 -40.635 -53.555 ;
        RECT -40.965 -55.245 -40.635 -54.915 ;
        RECT -40.965 -56.605 -40.635 -56.275 ;
        RECT -40.965 -57.965 -40.635 -57.635 ;
        RECT -40.965 -59.325 -40.635 -58.995 ;
        RECT -40.965 -60.685 -40.635 -60.355 ;
        RECT -40.965 -62.045 -40.635 -61.715 ;
        RECT -40.965 -63.405 -40.635 -63.075 ;
        RECT -40.965 -64.765 -40.635 -64.435 ;
        RECT -40.965 -65.91 -40.635 -65.58 ;
        RECT -40.965 -67.485 -40.635 -67.155 ;
        RECT -40.965 -68.845 -40.635 -68.515 ;
        RECT -40.965 -70.205 -40.635 -69.875 ;
        RECT -40.965 -71.565 -40.635 -71.235 ;
        RECT -40.965 -72.925 -40.635 -72.595 ;
        RECT -40.965 -75.645 -40.635 -75.315 ;
        RECT -40.965 -76.45 -40.635 -76.12 ;
        RECT -40.965 -78.365 -40.635 -78.035 ;
        RECT -40.965 -79.725 -40.635 -79.395 ;
        RECT -40.965 -81.085 -40.635 -80.755 ;
        RECT -40.965 -83.805 -40.635 -83.475 ;
        RECT -40.965 -85.165 -40.635 -84.835 ;
        RECT -40.965 -87.885 -40.635 -87.555 ;
        RECT -40.965 -89.245 -40.635 -88.915 ;
        RECT -40.965 -90.605 -40.635 -90.275 ;
        RECT -40.965 -91.965 -40.635 -91.635 ;
        RECT -40.965 -93.325 -40.635 -92.995 ;
        RECT -40.965 -94.685 -40.635 -94.355 ;
        RECT -40.965 -96.045 -40.635 -95.715 ;
        RECT -40.965 -97.405 -40.635 -97.075 ;
        RECT -40.965 -98.765 -40.635 -98.435 ;
        RECT -40.965 -100.125 -40.635 -99.795 ;
        RECT -40.965 -101.485 -40.635 -101.155 ;
        RECT -40.965 -102.845 -40.635 -102.515 ;
        RECT -40.965 -104.205 -40.635 -103.875 ;
        RECT -40.965 -105.565 -40.635 -105.235 ;
        RECT -40.965 -106.925 -40.635 -106.595 ;
        RECT -40.965 -108.285 -40.635 -107.955 ;
        RECT -40.965 -109.645 -40.635 -109.315 ;
        RECT -40.965 -111.005 -40.635 -110.675 ;
        RECT -40.965 -112.365 -40.635 -112.035 ;
        RECT -40.965 -113.725 -40.635 -113.395 ;
        RECT -40.965 -115.085 -40.635 -114.755 ;
        RECT -40.965 -116.445 -40.635 -116.115 ;
        RECT -40.965 -117.805 -40.635 -117.475 ;
        RECT -40.965 -119.165 -40.635 -118.835 ;
        RECT -40.965 -120.525 -40.635 -120.195 ;
        RECT -40.965 -121.885 -40.635 -121.555 ;
        RECT -40.965 -123.245 -40.635 -122.915 ;
        RECT -40.965 -125.965 -40.635 -125.635 ;
        RECT -40.965 -127.325 -40.635 -126.995 ;
        RECT -40.965 -128.685 -40.635 -128.355 ;
        RECT -40.965 -130.045 -40.635 -129.715 ;
        RECT -40.965 -132.765 -40.635 -132.435 ;
        RECT -40.965 -134.125 -40.635 -133.795 ;
        RECT -40.965 -135.485 -40.635 -135.155 ;
        RECT -40.965 -136.845 -40.635 -136.515 ;
        RECT -40.965 -138.205 -40.635 -137.875 ;
        RECT -40.965 -139.565 -40.635 -139.235 ;
        RECT -40.965 -140.925 -40.635 -140.595 ;
        RECT -40.965 -143.755 -40.635 -143.425 ;
        RECT -40.965 -145.005 -40.635 -144.675 ;
        RECT -40.965 -146.365 -40.635 -146.035 ;
        RECT -40.965 -149.085 -40.635 -148.755 ;
        RECT -40.965 -151.805 -40.635 -151.475 ;
        RECT -40.965 -153.165 -40.635 -152.835 ;
        RECT -40.965 -158.81 -40.635 -157.68 ;
        RECT -40.96 -158.925 -40.64 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.605 44.8 -39.275 45.93 ;
        RECT -39.605 39.955 -39.275 40.285 ;
        RECT -39.605 38.595 -39.275 38.925 ;
        RECT -39.605 37.235 -39.275 37.565 ;
        RECT -39.605 35.875 -39.275 36.205 ;
        RECT -39.605 34.515 -39.275 34.845 ;
        RECT -39.605 33.155 -39.275 33.485 ;
        RECT -39.605 31.795 -39.275 32.125 ;
        RECT -39.605 30.435 -39.275 30.765 ;
        RECT -39.605 29.075 -39.275 29.405 ;
        RECT -39.605 27.715 -39.275 28.045 ;
        RECT -39.605 26.355 -39.275 26.685 ;
        RECT -39.605 24.995 -39.275 25.325 ;
        RECT -39.605 23.635 -39.275 23.965 ;
        RECT -39.605 22.275 -39.275 22.605 ;
        RECT -39.605 20.915 -39.275 21.245 ;
        RECT -39.605 19.555 -39.275 19.885 ;
        RECT -39.605 18.195 -39.275 18.525 ;
        RECT -39.605 16.835 -39.275 17.165 ;
        RECT -39.605 15.475 -39.275 15.805 ;
        RECT -39.605 14.115 -39.275 14.445 ;
        RECT -39.605 12.755 -39.275 13.085 ;
        RECT -39.605 11.395 -39.275 11.725 ;
        RECT -39.605 10.035 -39.275 10.365 ;
        RECT -39.605 8.675 -39.275 9.005 ;
        RECT -39.605 7.315 -39.275 7.645 ;
        RECT -39.605 5.955 -39.275 6.285 ;
        RECT -39.605 4.595 -39.275 4.925 ;
        RECT -39.605 3.235 -39.275 3.565 ;
        RECT -39.605 1.875 -39.275 2.205 ;
        RECT -39.605 0.515 -39.275 0.845 ;
        RECT -39.605 -2.205 -39.275 -1.875 ;
        RECT -39.605 -4.925 -39.275 -4.595 ;
        RECT -39.605 -6.285 -39.275 -5.955 ;
        RECT -39.605 -7.645 -39.275 -7.315 ;
        RECT -39.605 -10.365 -39.275 -10.035 ;
        RECT -39.605 -11.725 -39.275 -11.395 ;
        RECT -39.605 -13.085 -39.275 -12.755 ;
        RECT -39.605 -14.445 -39.275 -14.115 ;
        RECT -39.605 -15.805 -39.275 -15.475 ;
        RECT -39.605 -17.165 -39.275 -16.835 ;
        RECT -39.605 -18.525 -39.275 -18.195 ;
        RECT -39.605 -25.325 -39.275 -24.995 ;
        RECT -39.605 -26.685 -39.275 -26.355 ;
        RECT -39.605 -28.045 -39.275 -27.715 ;
        RECT -39.605 -29.405 -39.275 -29.075 ;
        RECT -39.605 -30.765 -39.275 -30.435 ;
        RECT -39.605 -32.125 -39.275 -31.795 ;
        RECT -39.605 -33.485 -39.275 -33.155 ;
        RECT -39.605 -34.845 -39.275 -34.515 ;
        RECT -39.605 -36.205 -39.275 -35.875 ;
        RECT -39.605 -37.565 -39.275 -37.235 ;
        RECT -39.605 -38.925 -39.275 -38.595 ;
        RECT -39.605 -40.285 -39.275 -39.955 ;
        RECT -39.605 -41.645 -39.275 -41.315 ;
        RECT -39.605 -43.005 -39.275 -42.675 ;
        RECT -39.605 -44.365 -39.275 -44.035 ;
        RECT -39.605 -45.725 -39.275 -45.395 ;
        RECT -39.605 -47.085 -39.275 -46.755 ;
        RECT -39.605 -48.445 -39.275 -48.115 ;
        RECT -39.605 -49.805 -39.275 -49.475 ;
        RECT -39.605 -51.165 -39.275 -50.835 ;
        RECT -39.605 -52.525 -39.275 -52.195 ;
        RECT -39.605 -53.885 -39.275 -53.555 ;
        RECT -39.605 -55.245 -39.275 -54.915 ;
        RECT -39.605 -56.605 -39.275 -56.275 ;
        RECT -39.605 -57.965 -39.275 -57.635 ;
        RECT -39.605 -59.325 -39.275 -58.995 ;
        RECT -39.605 -60.685 -39.275 -60.355 ;
        RECT -39.605 -62.045 -39.275 -61.715 ;
        RECT -39.605 -63.405 -39.275 -63.075 ;
        RECT -39.605 -64.765 -39.275 -64.435 ;
        RECT -39.605 -65.91 -39.275 -65.58 ;
        RECT -39.605 -67.485 -39.275 -67.155 ;
        RECT -39.605 -68.845 -39.275 -68.515 ;
        RECT -39.605 -70.205 -39.275 -69.875 ;
        RECT -39.605 -71.565 -39.275 -71.235 ;
        RECT -39.605 -72.925 -39.275 -72.595 ;
        RECT -39.605 -75.645 -39.275 -75.315 ;
        RECT -39.605 -76.45 -39.275 -76.12 ;
        RECT -39.605 -78.365 -39.275 -78.035 ;
        RECT -39.605 -79.725 -39.275 -79.395 ;
        RECT -39.605 -81.085 -39.275 -80.755 ;
        RECT -39.605 -83.805 -39.275 -83.475 ;
        RECT -39.605 -85.165 -39.275 -84.835 ;
        RECT -39.605 -89.245 -39.275 -88.915 ;
        RECT -39.605 -90.605 -39.275 -90.275 ;
        RECT -39.605 -91.965 -39.275 -91.635 ;
        RECT -39.605 -93.325 -39.275 -92.995 ;
        RECT -39.605 -94.685 -39.275 -94.355 ;
        RECT -39.605 -96.045 -39.275 -95.715 ;
        RECT -39.605 -97.405 -39.275 -97.075 ;
        RECT -39.605 -98.765 -39.275 -98.435 ;
        RECT -39.605 -100.125 -39.275 -99.795 ;
        RECT -39.605 -101.485 -39.275 -101.155 ;
        RECT -39.605 -102.845 -39.275 -102.515 ;
        RECT -39.605 -104.205 -39.275 -103.875 ;
        RECT -39.605 -105.565 -39.275 -105.235 ;
        RECT -39.605 -108.285 -39.275 -107.955 ;
        RECT -39.605 -109.645 -39.275 -109.315 ;
        RECT -39.605 -111.005 -39.275 -110.675 ;
        RECT -39.605 -112.365 -39.275 -112.035 ;
        RECT -39.605 -113.725 -39.275 -113.395 ;
        RECT -39.605 -115.085 -39.275 -114.755 ;
        RECT -39.605 -116.445 -39.275 -116.115 ;
        RECT -39.605 -117.805 -39.275 -117.475 ;
        RECT -39.605 -119.165 -39.275 -118.835 ;
        RECT -39.605 -120.525 -39.275 -120.195 ;
        RECT -39.605 -121.885 -39.275 -121.555 ;
        RECT -39.605 -123.245 -39.275 -122.915 ;
        RECT -39.605 -125.965 -39.275 -125.635 ;
        RECT -39.605 -127.325 -39.275 -126.995 ;
        RECT -39.605 -130.045 -39.275 -129.715 ;
        RECT -39.605 -132.765 -39.275 -132.435 ;
        RECT -39.605 -134.125 -39.275 -133.795 ;
        RECT -39.605 -135.485 -39.275 -135.155 ;
        RECT -39.605 -136.845 -39.275 -136.515 ;
        RECT -39.605 -138.205 -39.275 -137.875 ;
        RECT -39.605 -139.565 -39.275 -139.235 ;
        RECT -39.605 -140.925 -39.275 -140.595 ;
        RECT -39.605 -143.755 -39.275 -143.425 ;
        RECT -39.605 -145.005 -39.275 -144.675 ;
        RECT -39.605 -146.365 -39.275 -146.035 ;
        RECT -39.605 -149.085 -39.275 -148.755 ;
        RECT -39.605 -151.805 -39.275 -151.475 ;
        RECT -39.605 -153.165 -39.275 -152.835 ;
        RECT -39.605 -158.81 -39.275 -157.68 ;
        RECT -39.6 -158.925 -39.28 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.245 44.8 -37.915 45.93 ;
        RECT -38.245 39.955 -37.915 40.285 ;
        RECT -38.245 38.595 -37.915 38.925 ;
        RECT -38.245 37.235 -37.915 37.565 ;
        RECT -38.245 35.875 -37.915 36.205 ;
        RECT -38.245 34.515 -37.915 34.845 ;
        RECT -38.245 33.155 -37.915 33.485 ;
        RECT -38.245 31.795 -37.915 32.125 ;
        RECT -38.245 30.435 -37.915 30.765 ;
        RECT -38.245 29.075 -37.915 29.405 ;
        RECT -38.245 27.715 -37.915 28.045 ;
        RECT -38.245 26.355 -37.915 26.685 ;
        RECT -38.245 24.995 -37.915 25.325 ;
        RECT -38.245 23.635 -37.915 23.965 ;
        RECT -38.245 22.275 -37.915 22.605 ;
        RECT -38.245 20.915 -37.915 21.245 ;
        RECT -38.245 19.555 -37.915 19.885 ;
        RECT -38.245 18.195 -37.915 18.525 ;
        RECT -38.245 16.835 -37.915 17.165 ;
        RECT -38.245 15.475 -37.915 15.805 ;
        RECT -38.245 14.115 -37.915 14.445 ;
        RECT -38.245 12.755 -37.915 13.085 ;
        RECT -38.245 11.395 -37.915 11.725 ;
        RECT -38.245 10.035 -37.915 10.365 ;
        RECT -38.245 8.675 -37.915 9.005 ;
        RECT -38.245 7.315 -37.915 7.645 ;
        RECT -38.245 5.955 -37.915 6.285 ;
        RECT -38.245 4.595 -37.915 4.925 ;
        RECT -38.245 3.235 -37.915 3.565 ;
        RECT -38.245 1.875 -37.915 2.205 ;
        RECT -38.245 -2.205 -37.915 -1.875 ;
        RECT -38.245 -4.925 -37.915 -4.595 ;
        RECT -38.245 -6.285 -37.915 -5.955 ;
        RECT -38.245 -7.645 -37.915 -7.315 ;
        RECT -38.245 -10.365 -37.915 -10.035 ;
        RECT -38.245 -11.725 -37.915 -11.395 ;
        RECT -38.245 -13.085 -37.915 -12.755 ;
        RECT -38.245 -14.445 -37.915 -14.115 ;
        RECT -38.245 -15.805 -37.915 -15.475 ;
        RECT -38.245 -17.165 -37.915 -16.835 ;
        RECT -38.245 -18.525 -37.915 -18.195 ;
        RECT -38.245 -25.325 -37.915 -24.995 ;
        RECT -38.245 -26.685 -37.915 -26.355 ;
        RECT -38.245 -28.045 -37.915 -27.715 ;
        RECT -38.245 -29.405 -37.915 -29.075 ;
        RECT -38.245 -30.765 -37.915 -30.435 ;
        RECT -38.245 -32.125 -37.915 -31.795 ;
        RECT -38.245 -33.485 -37.915 -33.155 ;
        RECT -38.245 -34.845 -37.915 -34.515 ;
        RECT -38.245 -36.205 -37.915 -35.875 ;
        RECT -38.245 -37.565 -37.915 -37.235 ;
        RECT -38.245 -38.925 -37.915 -38.595 ;
        RECT -38.245 -40.285 -37.915 -39.955 ;
        RECT -38.245 -41.645 -37.915 -41.315 ;
        RECT -38.245 -43.005 -37.915 -42.675 ;
        RECT -38.245 -44.365 -37.915 -44.035 ;
        RECT -38.245 -45.725 -37.915 -45.395 ;
        RECT -38.245 -47.085 -37.915 -46.755 ;
        RECT -38.245 -48.445 -37.915 -48.115 ;
        RECT -38.245 -49.805 -37.915 -49.475 ;
        RECT -38.245 -51.165 -37.915 -50.835 ;
        RECT -38.245 -52.525 -37.915 -52.195 ;
        RECT -38.245 -53.885 -37.915 -53.555 ;
        RECT -38.245 -55.245 -37.915 -54.915 ;
        RECT -38.245 -56.605 -37.915 -56.275 ;
        RECT -38.245 -57.965 -37.915 -57.635 ;
        RECT -38.245 -59.325 -37.915 -58.995 ;
        RECT -38.245 -60.685 -37.915 -60.355 ;
        RECT -38.245 -62.045 -37.915 -61.715 ;
        RECT -38.245 -63.405 -37.915 -63.075 ;
        RECT -38.245 -64.765 -37.915 -64.435 ;
        RECT -38.245 -65.91 -37.915 -65.58 ;
        RECT -38.245 -67.485 -37.915 -67.155 ;
        RECT -38.245 -68.845 -37.915 -68.515 ;
        RECT -38.245 -70.205 -37.915 -69.875 ;
        RECT -38.245 -71.565 -37.915 -71.235 ;
        RECT -38.245 -72.925 -37.915 -72.595 ;
        RECT -38.245 -75.645 -37.915 -75.315 ;
        RECT -38.245 -76.45 -37.915 -76.12 ;
        RECT -38.245 -78.365 -37.915 -78.035 ;
        RECT -38.245 -79.725 -37.915 -79.395 ;
        RECT -38.245 -81.085 -37.915 -80.755 ;
        RECT -38.245 -83.805 -37.915 -83.475 ;
        RECT -38.245 -85.165 -37.915 -84.835 ;
        RECT -38.245 -87.885 -37.915 -87.555 ;
        RECT -38.245 -89.245 -37.915 -88.915 ;
        RECT -38.245 -90.605 -37.915 -90.275 ;
        RECT -38.245 -91.965 -37.915 -91.635 ;
        RECT -38.245 -93.325 -37.915 -92.995 ;
        RECT -38.245 -94.685 -37.915 -94.355 ;
        RECT -38.245 -96.045 -37.915 -95.715 ;
        RECT -38.245 -97.405 -37.915 -97.075 ;
        RECT -38.245 -98.765 -37.915 -98.435 ;
        RECT -38.245 -100.125 -37.915 -99.795 ;
        RECT -38.245 -101.485 -37.915 -101.155 ;
        RECT -38.245 -102.845 -37.915 -102.515 ;
        RECT -38.245 -104.205 -37.915 -103.875 ;
        RECT -38.245 -108.285 -37.915 -107.955 ;
        RECT -38.245 -109.645 -37.915 -109.315 ;
        RECT -38.245 -111.005 -37.915 -110.675 ;
        RECT -38.245 -112.365 -37.915 -112.035 ;
        RECT -38.245 -113.725 -37.915 -113.395 ;
        RECT -38.245 -115.085 -37.915 -114.755 ;
        RECT -38.245 -116.445 -37.915 -116.115 ;
        RECT -38.245 -117.805 -37.915 -117.475 ;
        RECT -38.245 -119.165 -37.915 -118.835 ;
        RECT -38.245 -120.525 -37.915 -120.195 ;
        RECT -38.245 -121.885 -37.915 -121.555 ;
        RECT -38.245 -123.245 -37.915 -122.915 ;
        RECT -38.245 -125.965 -37.915 -125.635 ;
        RECT -38.245 -127.325 -37.915 -126.995 ;
        RECT -38.245 -131.405 -37.915 -131.075 ;
        RECT -38.245 -132.765 -37.915 -132.435 ;
        RECT -38.245 -134.125 -37.915 -133.795 ;
        RECT -38.245 -135.485 -37.915 -135.155 ;
        RECT -38.245 -136.845 -37.915 -136.515 ;
        RECT -38.245 -138.205 -37.915 -137.875 ;
        RECT -38.245 -139.565 -37.915 -139.235 ;
        RECT -38.245 -140.925 -37.915 -140.595 ;
        RECT -38.245 -143.755 -37.915 -143.425 ;
        RECT -38.245 -145.005 -37.915 -144.675 ;
        RECT -38.245 -146.365 -37.915 -146.035 ;
        RECT -38.245 -147.725 -37.915 -147.395 ;
        RECT -38.245 -149.085 -37.915 -148.755 ;
        RECT -38.245 -151.805 -37.915 -151.475 ;
        RECT -38.245 -153.165 -37.915 -152.835 ;
        RECT -38.245 -158.81 -37.915 -157.68 ;
        RECT -38.24 -158.925 -37.92 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.885 44.8 -36.555 45.93 ;
        RECT -36.885 39.955 -36.555 40.285 ;
        RECT -36.885 38.595 -36.555 38.925 ;
        RECT -36.885 37.235 -36.555 37.565 ;
        RECT -36.885 35.875 -36.555 36.205 ;
        RECT -36.885 34.515 -36.555 34.845 ;
        RECT -36.885 33.155 -36.555 33.485 ;
        RECT -36.885 31.795 -36.555 32.125 ;
        RECT -36.885 30.435 -36.555 30.765 ;
        RECT -36.885 29.075 -36.555 29.405 ;
        RECT -36.885 27.715 -36.555 28.045 ;
        RECT -36.885 26.355 -36.555 26.685 ;
        RECT -36.885 24.995 -36.555 25.325 ;
        RECT -36.885 23.635 -36.555 23.965 ;
        RECT -36.885 22.275 -36.555 22.605 ;
        RECT -36.885 20.915 -36.555 21.245 ;
        RECT -36.885 19.555 -36.555 19.885 ;
        RECT -36.885 18.195 -36.555 18.525 ;
        RECT -36.885 16.835 -36.555 17.165 ;
        RECT -36.885 15.475 -36.555 15.805 ;
        RECT -36.885 14.115 -36.555 14.445 ;
        RECT -36.885 12.755 -36.555 13.085 ;
        RECT -36.885 11.395 -36.555 11.725 ;
        RECT -36.885 10.035 -36.555 10.365 ;
        RECT -36.885 8.675 -36.555 9.005 ;
        RECT -36.885 7.315 -36.555 7.645 ;
        RECT -36.885 5.955 -36.555 6.285 ;
        RECT -36.885 4.595 -36.555 4.925 ;
        RECT -36.885 3.235 -36.555 3.565 ;
        RECT -36.885 1.875 -36.555 2.205 ;
        RECT -36.885 -2.205 -36.555 -1.875 ;
        RECT -36.885 -4.925 -36.555 -4.595 ;
        RECT -36.885 -6.285 -36.555 -5.955 ;
        RECT -36.885 -7.645 -36.555 -7.315 ;
        RECT -36.885 -10.365 -36.555 -10.035 ;
        RECT -36.885 -11.725 -36.555 -11.395 ;
        RECT -36.885 -13.085 -36.555 -12.755 ;
        RECT -36.885 -14.445 -36.555 -14.115 ;
        RECT -36.885 -15.805 -36.555 -15.475 ;
        RECT -36.885 -17.165 -36.555 -16.835 ;
        RECT -36.885 -18.525 -36.555 -18.195 ;
        RECT -36.885 -25.325 -36.555 -24.995 ;
        RECT -36.885 -26.685 -36.555 -26.355 ;
        RECT -36.885 -28.045 -36.555 -27.715 ;
        RECT -36.885 -29.405 -36.555 -29.075 ;
        RECT -36.885 -30.765 -36.555 -30.435 ;
        RECT -36.885 -32.125 -36.555 -31.795 ;
        RECT -36.885 -33.485 -36.555 -33.155 ;
        RECT -36.885 -34.845 -36.555 -34.515 ;
        RECT -36.885 -36.205 -36.555 -35.875 ;
        RECT -36.885 -37.565 -36.555 -37.235 ;
        RECT -36.885 -38.925 -36.555 -38.595 ;
        RECT -36.885 -40.285 -36.555 -39.955 ;
        RECT -36.885 -41.645 -36.555 -41.315 ;
        RECT -36.885 -43.005 -36.555 -42.675 ;
        RECT -36.885 -44.365 -36.555 -44.035 ;
        RECT -36.885 -45.725 -36.555 -45.395 ;
        RECT -36.885 -47.085 -36.555 -46.755 ;
        RECT -36.885 -48.445 -36.555 -48.115 ;
        RECT -36.885 -49.805 -36.555 -49.475 ;
        RECT -36.885 -51.165 -36.555 -50.835 ;
        RECT -36.885 -52.525 -36.555 -52.195 ;
        RECT -36.885 -53.885 -36.555 -53.555 ;
        RECT -36.885 -55.245 -36.555 -54.915 ;
        RECT -36.885 -56.605 -36.555 -56.275 ;
        RECT -36.885 -57.965 -36.555 -57.635 ;
        RECT -36.885 -59.325 -36.555 -58.995 ;
        RECT -36.885 -60.685 -36.555 -60.355 ;
        RECT -36.885 -62.045 -36.555 -61.715 ;
        RECT -36.885 -63.405 -36.555 -63.075 ;
        RECT -36.885 -64.765 -36.555 -64.435 ;
        RECT -36.885 -65.91 -36.555 -65.58 ;
        RECT -36.885 -67.485 -36.555 -67.155 ;
        RECT -36.885 -68.845 -36.555 -68.515 ;
        RECT -36.885 -70.205 -36.555 -69.875 ;
        RECT -36.885 -71.565 -36.555 -71.235 ;
        RECT -36.885 -72.925 -36.555 -72.595 ;
        RECT -36.885 -75.645 -36.555 -75.315 ;
        RECT -36.885 -76.45 -36.555 -76.12 ;
        RECT -36.885 -78.365 -36.555 -78.035 ;
        RECT -36.885 -79.725 -36.555 -79.395 ;
        RECT -36.885 -81.085 -36.555 -80.755 ;
        RECT -36.885 -83.805 -36.555 -83.475 ;
        RECT -36.885 -85.165 -36.555 -84.835 ;
        RECT -36.885 -87.885 -36.555 -87.555 ;
        RECT -36.885 -89.245 -36.555 -88.915 ;
        RECT -36.885 -90.605 -36.555 -90.275 ;
        RECT -36.885 -91.965 -36.555 -91.635 ;
        RECT -36.885 -93.325 -36.555 -92.995 ;
        RECT -36.885 -94.685 -36.555 -94.355 ;
        RECT -36.885 -96.045 -36.555 -95.715 ;
        RECT -36.885 -97.405 -36.555 -97.075 ;
        RECT -36.885 -98.765 -36.555 -98.435 ;
        RECT -36.885 -100.125 -36.555 -99.795 ;
        RECT -36.885 -101.485 -36.555 -101.155 ;
        RECT -36.885 -102.845 -36.555 -102.515 ;
        RECT -36.885 -104.205 -36.555 -103.875 ;
        RECT -36.885 -108.285 -36.555 -107.955 ;
        RECT -36.885 -109.645 -36.555 -109.315 ;
        RECT -36.885 -111.005 -36.555 -110.675 ;
        RECT -36.885 -112.365 -36.555 -112.035 ;
        RECT -36.885 -113.725 -36.555 -113.395 ;
        RECT -36.885 -115.085 -36.555 -114.755 ;
        RECT -36.885 -116.445 -36.555 -116.115 ;
        RECT -36.885 -117.805 -36.555 -117.475 ;
        RECT -36.885 -119.165 -36.555 -118.835 ;
        RECT -36.885 -120.525 -36.555 -120.195 ;
        RECT -36.885 -121.885 -36.555 -121.555 ;
        RECT -36.885 -123.245 -36.555 -122.915 ;
        RECT -36.885 -125.965 -36.555 -125.635 ;
        RECT -36.885 -127.325 -36.555 -126.995 ;
        RECT -36.885 -131.405 -36.555 -131.075 ;
        RECT -36.885 -132.765 -36.555 -132.435 ;
        RECT -36.885 -134.125 -36.555 -133.795 ;
        RECT -36.885 -135.485 -36.555 -135.155 ;
        RECT -36.885 -136.845 -36.555 -136.515 ;
        RECT -36.885 -138.205 -36.555 -137.875 ;
        RECT -36.885 -139.565 -36.555 -139.235 ;
        RECT -36.885 -140.925 -36.555 -140.595 ;
        RECT -36.885 -143.755 -36.555 -143.425 ;
        RECT -36.885 -145.005 -36.555 -144.675 ;
        RECT -36.885 -146.365 -36.555 -146.035 ;
        RECT -36.885 -147.725 -36.555 -147.395 ;
        RECT -36.885 -149.085 -36.555 -148.755 ;
        RECT -36.885 -151.805 -36.555 -151.475 ;
        RECT -36.885 -153.165 -36.555 -152.835 ;
        RECT -36.885 -158.81 -36.555 -157.68 ;
        RECT -36.88 -158.925 -36.56 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.525 44.8 -35.195 45.93 ;
        RECT -35.525 39.955 -35.195 40.285 ;
        RECT -35.525 38.595 -35.195 38.925 ;
        RECT -35.525 37.235 -35.195 37.565 ;
        RECT -35.525 35.875 -35.195 36.205 ;
        RECT -35.525 34.515 -35.195 34.845 ;
        RECT -35.525 33.155 -35.195 33.485 ;
        RECT -35.525 31.795 -35.195 32.125 ;
        RECT -35.525 30.435 -35.195 30.765 ;
        RECT -35.525 29.075 -35.195 29.405 ;
        RECT -35.525 27.715 -35.195 28.045 ;
        RECT -35.525 26.355 -35.195 26.685 ;
        RECT -35.525 24.995 -35.195 25.325 ;
        RECT -35.525 23.635 -35.195 23.965 ;
        RECT -35.525 22.275 -35.195 22.605 ;
        RECT -35.525 20.915 -35.195 21.245 ;
        RECT -35.525 19.555 -35.195 19.885 ;
        RECT -35.525 18.195 -35.195 18.525 ;
        RECT -35.525 16.835 -35.195 17.165 ;
        RECT -35.525 15.475 -35.195 15.805 ;
        RECT -35.525 14.115 -35.195 14.445 ;
        RECT -35.525 12.755 -35.195 13.085 ;
        RECT -35.525 11.395 -35.195 11.725 ;
        RECT -35.525 10.035 -35.195 10.365 ;
        RECT -35.525 8.675 -35.195 9.005 ;
        RECT -35.525 7.315 -35.195 7.645 ;
        RECT -35.525 5.955 -35.195 6.285 ;
        RECT -35.525 4.595 -35.195 4.925 ;
        RECT -35.525 3.235 -35.195 3.565 ;
        RECT -35.525 1.875 -35.195 2.205 ;
        RECT -35.525 -2.205 -35.195 -1.875 ;
        RECT -35.525 -4.925 -35.195 -4.595 ;
        RECT -35.525 -6.285 -35.195 -5.955 ;
        RECT -35.525 -7.645 -35.195 -7.315 ;
        RECT -35.525 -10.365 -35.195 -10.035 ;
        RECT -35.525 -11.725 -35.195 -11.395 ;
        RECT -35.525 -13.085 -35.195 -12.755 ;
        RECT -35.525 -14.445 -35.195 -14.115 ;
        RECT -35.525 -15.805 -35.195 -15.475 ;
        RECT -35.525 -17.165 -35.195 -16.835 ;
        RECT -35.525 -18.525 -35.195 -18.195 ;
        RECT -35.525 -25.325 -35.195 -24.995 ;
        RECT -35.525 -26.685 -35.195 -26.355 ;
        RECT -35.525 -28.045 -35.195 -27.715 ;
        RECT -35.525 -29.405 -35.195 -29.075 ;
        RECT -35.525 -30.765 -35.195 -30.435 ;
        RECT -35.525 -32.125 -35.195 -31.795 ;
        RECT -35.525 -33.485 -35.195 -33.155 ;
        RECT -35.525 -34.845 -35.195 -34.515 ;
        RECT -35.525 -36.205 -35.195 -35.875 ;
        RECT -35.525 -37.565 -35.195 -37.235 ;
        RECT -35.525 -38.925 -35.195 -38.595 ;
        RECT -35.525 -40.285 -35.195 -39.955 ;
        RECT -35.525 -41.645 -35.195 -41.315 ;
        RECT -35.525 -43.005 -35.195 -42.675 ;
        RECT -35.525 -44.365 -35.195 -44.035 ;
        RECT -35.525 -45.725 -35.195 -45.395 ;
        RECT -35.525 -47.085 -35.195 -46.755 ;
        RECT -35.525 -48.445 -35.195 -48.115 ;
        RECT -35.525 -49.805 -35.195 -49.475 ;
        RECT -35.525 -51.165 -35.195 -50.835 ;
        RECT -35.525 -52.525 -35.195 -52.195 ;
        RECT -35.525 -53.885 -35.195 -53.555 ;
        RECT -35.525 -55.245 -35.195 -54.915 ;
        RECT -35.525 -56.605 -35.195 -56.275 ;
        RECT -35.525 -57.965 -35.195 -57.635 ;
        RECT -35.525 -59.325 -35.195 -58.995 ;
        RECT -35.525 -60.685 -35.195 -60.355 ;
        RECT -35.525 -62.045 -35.195 -61.715 ;
        RECT -35.525 -63.405 -35.195 -63.075 ;
        RECT -35.525 -64.765 -35.195 -64.435 ;
        RECT -35.525 -65.91 -35.195 -65.58 ;
        RECT -35.525 -67.485 -35.195 -67.155 ;
        RECT -35.525 -68.845 -35.195 -68.515 ;
        RECT -35.525 -70.205 -35.195 -69.875 ;
        RECT -35.525 -71.565 -35.195 -71.235 ;
        RECT -35.525 -72.925 -35.195 -72.595 ;
        RECT -35.525 -75.645 -35.195 -75.315 ;
        RECT -35.525 -76.45 -35.195 -76.12 ;
        RECT -35.525 -78.365 -35.195 -78.035 ;
        RECT -35.525 -79.725 -35.195 -79.395 ;
        RECT -35.525 -81.085 -35.195 -80.755 ;
        RECT -35.525 -83.805 -35.195 -83.475 ;
        RECT -35.525 -85.165 -35.195 -84.835 ;
        RECT -35.525 -87.885 -35.195 -87.555 ;
        RECT -35.525 -89.245 -35.195 -88.915 ;
        RECT -35.525 -90.605 -35.195 -90.275 ;
        RECT -35.525 -91.965 -35.195 -91.635 ;
        RECT -35.525 -93.325 -35.195 -92.995 ;
        RECT -35.525 -94.685 -35.195 -94.355 ;
        RECT -35.525 -96.045 -35.195 -95.715 ;
        RECT -35.525 -97.405 -35.195 -97.075 ;
        RECT -35.525 -100.125 -35.195 -99.795 ;
        RECT -35.525 -101.485 -35.195 -101.155 ;
        RECT -35.525 -102.845 -35.195 -102.515 ;
        RECT -35.525 -104.205 -35.195 -103.875 ;
        RECT -35.525 -108.285 -35.195 -107.955 ;
        RECT -35.525 -109.645 -35.195 -109.315 ;
        RECT -35.525 -111.005 -35.195 -110.675 ;
        RECT -35.525 -112.365 -35.195 -112.035 ;
        RECT -35.525 -113.725 -35.195 -113.395 ;
        RECT -35.525 -116.445 -35.195 -116.115 ;
        RECT -35.525 -117.805 -35.195 -117.475 ;
        RECT -35.525 -119.165 -35.195 -118.835 ;
        RECT -35.525 -120.525 -35.195 -120.195 ;
        RECT -35.525 -121.885 -35.195 -121.555 ;
        RECT -35.525 -123.245 -35.195 -122.915 ;
        RECT -35.525 -125.965 -35.195 -125.635 ;
        RECT -35.525 -127.325 -35.195 -126.995 ;
        RECT -35.525 -131.405 -35.195 -131.075 ;
        RECT -35.525 -132.765 -35.195 -132.435 ;
        RECT -35.525 -134.125 -35.195 -133.795 ;
        RECT -35.525 -135.485 -35.195 -135.155 ;
        RECT -35.525 -136.845 -35.195 -136.515 ;
        RECT -35.525 -138.205 -35.195 -137.875 ;
        RECT -35.525 -139.565 -35.195 -139.235 ;
        RECT -35.525 -140.925 -35.195 -140.595 ;
        RECT -35.525 -143.755 -35.195 -143.425 ;
        RECT -35.525 -145.005 -35.195 -144.675 ;
        RECT -35.525 -146.365 -35.195 -146.035 ;
        RECT -35.525 -151.805 -35.195 -151.475 ;
        RECT -35.525 -153.165 -35.195 -152.835 ;
        RECT -35.525 -158.81 -35.195 -157.68 ;
        RECT -35.52 -158.925 -35.2 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.165 44.8 -33.835 45.93 ;
        RECT -34.165 39.955 -33.835 40.285 ;
        RECT -34.165 38.595 -33.835 38.925 ;
        RECT -34.165 37.235 -33.835 37.565 ;
        RECT -34.165 35.875 -33.835 36.205 ;
        RECT -34.165 34.515 -33.835 34.845 ;
        RECT -34.165 33.155 -33.835 33.485 ;
        RECT -34.165 31.795 -33.835 32.125 ;
        RECT -34.165 30.435 -33.835 30.765 ;
        RECT -34.165 29.075 -33.835 29.405 ;
        RECT -34.165 27.715 -33.835 28.045 ;
        RECT -34.165 26.355 -33.835 26.685 ;
        RECT -34.165 24.995 -33.835 25.325 ;
        RECT -34.165 23.635 -33.835 23.965 ;
        RECT -34.165 22.275 -33.835 22.605 ;
        RECT -34.165 20.915 -33.835 21.245 ;
        RECT -34.165 19.555 -33.835 19.885 ;
        RECT -34.165 18.195 -33.835 18.525 ;
        RECT -34.165 16.835 -33.835 17.165 ;
        RECT -34.165 15.475 -33.835 15.805 ;
        RECT -34.165 14.115 -33.835 14.445 ;
        RECT -34.165 12.755 -33.835 13.085 ;
        RECT -34.165 11.395 -33.835 11.725 ;
        RECT -34.165 10.035 -33.835 10.365 ;
        RECT -34.165 8.675 -33.835 9.005 ;
        RECT -34.165 7.315 -33.835 7.645 ;
        RECT -34.165 5.955 -33.835 6.285 ;
        RECT -34.165 4.595 -33.835 4.925 ;
        RECT -34.165 3.235 -33.835 3.565 ;
        RECT -34.165 1.875 -33.835 2.205 ;
        RECT -34.165 -2.205 -33.835 -1.875 ;
        RECT -34.165 -4.925 -33.835 -4.595 ;
        RECT -34.165 -6.285 -33.835 -5.955 ;
        RECT -34.165 -7.645 -33.835 -7.315 ;
        RECT -34.165 -10.365 -33.835 -10.035 ;
        RECT -34.165 -11.725 -33.835 -11.395 ;
        RECT -34.165 -13.085 -33.835 -12.755 ;
        RECT -34.165 -14.445 -33.835 -14.115 ;
        RECT -34.165 -15.805 -33.835 -15.475 ;
        RECT -34.165 -17.165 -33.835 -16.835 ;
        RECT -34.165 -18.525 -33.835 -18.195 ;
        RECT -34.165 -25.325 -33.835 -24.995 ;
        RECT -34.165 -26.685 -33.835 -26.355 ;
        RECT -34.165 -28.045 -33.835 -27.715 ;
        RECT -34.165 -29.405 -33.835 -29.075 ;
        RECT -34.165 -30.765 -33.835 -30.435 ;
        RECT -34.165 -32.125 -33.835 -31.795 ;
        RECT -34.165 -33.485 -33.835 -33.155 ;
        RECT -34.165 -34.845 -33.835 -34.515 ;
        RECT -34.165 -36.205 -33.835 -35.875 ;
        RECT -34.165 -37.565 -33.835 -37.235 ;
        RECT -34.165 -38.925 -33.835 -38.595 ;
        RECT -34.165 -40.285 -33.835 -39.955 ;
        RECT -34.165 -43.005 -33.835 -42.675 ;
        RECT -34.165 -44.365 -33.835 -44.035 ;
        RECT -34.165 -45.725 -33.835 -45.395 ;
        RECT -34.165 -47.085 -33.835 -46.755 ;
        RECT -34.165 -48.445 -33.835 -48.115 ;
        RECT -34.165 -49.805 -33.835 -49.475 ;
        RECT -34.165 -51.165 -33.835 -50.835 ;
        RECT -34.165 -52.525 -33.835 -52.195 ;
        RECT -34.165 -53.885 -33.835 -53.555 ;
        RECT -34.165 -55.245 -33.835 -54.915 ;
        RECT -34.165 -56.605 -33.835 -56.275 ;
        RECT -34.165 -57.965 -33.835 -57.635 ;
        RECT -34.165 -59.325 -33.835 -58.995 ;
        RECT -34.165 -60.685 -33.835 -60.355 ;
        RECT -34.165 -62.045 -33.835 -61.715 ;
        RECT -34.165 -63.405 -33.835 -63.075 ;
        RECT -34.165 -64.765 -33.835 -64.435 ;
        RECT -34.165 -65.91 -33.835 -65.58 ;
        RECT -34.165 -67.485 -33.835 -67.155 ;
        RECT -34.165 -68.845 -33.835 -68.515 ;
        RECT -34.165 -70.205 -33.835 -69.875 ;
        RECT -34.165 -71.565 -33.835 -71.235 ;
        RECT -34.165 -72.925 -33.835 -72.595 ;
        RECT -34.165 -75.645 -33.835 -75.315 ;
        RECT -34.165 -76.45 -33.835 -76.12 ;
        RECT -34.165 -78.365 -33.835 -78.035 ;
        RECT -34.165 -79.725 -33.835 -79.395 ;
        RECT -34.165 -81.085 -33.835 -80.755 ;
        RECT -34.165 -83.805 -33.835 -83.475 ;
        RECT -34.165 -85.165 -33.835 -84.835 ;
        RECT -34.165 -87.885 -33.835 -87.555 ;
        RECT -34.165 -89.245 -33.835 -88.915 ;
        RECT -34.165 -90.605 -33.835 -90.275 ;
        RECT -34.165 -91.965 -33.835 -91.635 ;
        RECT -34.165 -93.325 -33.835 -92.995 ;
        RECT -34.165 -94.685 -33.835 -94.355 ;
        RECT -34.165 -96.045 -33.835 -95.715 ;
        RECT -34.165 -97.405 -33.835 -97.075 ;
        RECT -34.165 -100.125 -33.835 -99.795 ;
        RECT -34.165 -101.485 -33.835 -101.155 ;
        RECT -34.165 -102.845 -33.835 -102.515 ;
        RECT -34.165 -104.205 -33.835 -103.875 ;
        RECT -34.165 -108.285 -33.835 -107.955 ;
        RECT -34.165 -109.645 -33.835 -109.315 ;
        RECT -34.165 -111.005 -33.835 -110.675 ;
        RECT -34.165 -112.365 -33.835 -112.035 ;
        RECT -34.165 -113.725 -33.835 -113.395 ;
        RECT -34.165 -116.445 -33.835 -116.115 ;
        RECT -34.165 -117.805 -33.835 -117.475 ;
        RECT -34.165 -119.165 -33.835 -118.835 ;
        RECT -34.165 -120.525 -33.835 -120.195 ;
        RECT -34.165 -121.885 -33.835 -121.555 ;
        RECT -34.165 -123.245 -33.835 -122.915 ;
        RECT -34.165 -125.965 -33.835 -125.635 ;
        RECT -34.165 -127.325 -33.835 -126.995 ;
        RECT -34.165 -131.405 -33.835 -131.075 ;
        RECT -34.165 -132.765 -33.835 -132.435 ;
        RECT -34.165 -134.125 -33.835 -133.795 ;
        RECT -34.165 -135.485 -33.835 -135.155 ;
        RECT -34.165 -136.845 -33.835 -136.515 ;
        RECT -34.165 -138.205 -33.835 -137.875 ;
        RECT -34.165 -139.565 -33.835 -139.235 ;
        RECT -34.165 -140.925 -33.835 -140.595 ;
        RECT -34.165 -143.755 -33.835 -143.425 ;
        RECT -34.165 -145.005 -33.835 -144.675 ;
        RECT -34.165 -146.365 -33.835 -146.035 ;
        RECT -34.16 -147.04 -33.84 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.805 -65.91 -32.475 -65.58 ;
        RECT -32.805 -67.485 -32.475 -67.155 ;
        RECT -32.805 -68.845 -32.475 -68.515 ;
        RECT -32.805 -70.205 -32.475 -69.875 ;
        RECT -32.805 -71.565 -32.475 -71.235 ;
        RECT -32.805 -72.925 -32.475 -72.595 ;
        RECT -32.805 -75.645 -32.475 -75.315 ;
        RECT -32.805 -76.45 -32.475 -76.12 ;
        RECT -32.805 -78.365 -32.475 -78.035 ;
        RECT -32.805 -79.725 -32.475 -79.395 ;
        RECT -32.805 -81.085 -32.475 -80.755 ;
        RECT -32.805 -83.805 -32.475 -83.475 ;
        RECT -32.805 -85.165 -32.475 -84.835 ;
        RECT -32.805 -87.885 -32.475 -87.555 ;
        RECT -32.805 -89.245 -32.475 -88.915 ;
        RECT -32.805 -90.605 -32.475 -90.275 ;
        RECT -32.805 -91.965 -32.475 -91.635 ;
        RECT -32.805 -93.325 -32.475 -92.995 ;
        RECT -32.805 -94.685 -32.475 -94.355 ;
        RECT -32.805 -96.045 -32.475 -95.715 ;
        RECT -32.805 -97.405 -32.475 -97.075 ;
        RECT -32.805 -100.125 -32.475 -99.795 ;
        RECT -32.805 -101.485 -32.475 -101.155 ;
        RECT -32.805 -102.845 -32.475 -102.515 ;
        RECT -32.805 -104.205 -32.475 -103.875 ;
        RECT -32.805 -108.285 -32.475 -107.955 ;
        RECT -32.805 -109.645 -32.475 -109.315 ;
        RECT -32.805 -111.005 -32.475 -110.675 ;
        RECT -32.805 -113.725 -32.475 -113.395 ;
        RECT -32.805 -116.445 -32.475 -116.115 ;
        RECT -32.805 -117.805 -32.475 -117.475 ;
        RECT -32.805 -119.165 -32.475 -118.835 ;
        RECT -32.805 -120.525 -32.475 -120.195 ;
        RECT -32.805 -121.885 -32.475 -121.555 ;
        RECT -32.805 -123.245 -32.475 -122.915 ;
        RECT -32.805 -125.965 -32.475 -125.635 ;
        RECT -32.805 -127.325 -32.475 -126.995 ;
        RECT -32.805 -131.405 -32.475 -131.075 ;
        RECT -32.805 -132.765 -32.475 -132.435 ;
        RECT -32.805 -134.125 -32.475 -133.795 ;
        RECT -32.805 -135.485 -32.475 -135.155 ;
        RECT -32.805 -136.845 -32.475 -136.515 ;
        RECT -32.805 -138.205 -32.475 -137.875 ;
        RECT -32.805 -139.565 -32.475 -139.235 ;
        RECT -32.805 -140.925 -32.475 -140.595 ;
        RECT -32.8 -141.6 -32.48 46.045 ;
        RECT -32.805 44.8 -32.475 45.93 ;
        RECT -32.805 39.955 -32.475 40.285 ;
        RECT -32.805 38.595 -32.475 38.925 ;
        RECT -32.805 37.235 -32.475 37.565 ;
        RECT -32.805 35.875 -32.475 36.205 ;
        RECT -32.805 34.515 -32.475 34.845 ;
        RECT -32.805 33.155 -32.475 33.485 ;
        RECT -32.805 31.795 -32.475 32.125 ;
        RECT -32.805 30.435 -32.475 30.765 ;
        RECT -32.805 29.075 -32.475 29.405 ;
        RECT -32.805 27.715 -32.475 28.045 ;
        RECT -32.805 26.355 -32.475 26.685 ;
        RECT -32.805 24.995 -32.475 25.325 ;
        RECT -32.805 23.635 -32.475 23.965 ;
        RECT -32.805 22.275 -32.475 22.605 ;
        RECT -32.805 20.915 -32.475 21.245 ;
        RECT -32.805 19.555 -32.475 19.885 ;
        RECT -32.805 18.195 -32.475 18.525 ;
        RECT -32.805 16.835 -32.475 17.165 ;
        RECT -32.805 15.475 -32.475 15.805 ;
        RECT -32.805 14.115 -32.475 14.445 ;
        RECT -32.805 12.755 -32.475 13.085 ;
        RECT -32.805 11.395 -32.475 11.725 ;
        RECT -32.805 10.035 -32.475 10.365 ;
        RECT -32.805 8.675 -32.475 9.005 ;
        RECT -32.805 7.315 -32.475 7.645 ;
        RECT -32.805 5.955 -32.475 6.285 ;
        RECT -32.805 4.595 -32.475 4.925 ;
        RECT -32.805 3.235 -32.475 3.565 ;
        RECT -32.805 1.875 -32.475 2.205 ;
        RECT -32.805 -2.205 -32.475 -1.875 ;
        RECT -32.805 -4.925 -32.475 -4.595 ;
        RECT -32.805 -6.285 -32.475 -5.955 ;
        RECT -32.805 -7.645 -32.475 -7.315 ;
        RECT -32.805 -10.365 -32.475 -10.035 ;
        RECT -32.805 -11.725 -32.475 -11.395 ;
        RECT -32.805 -13.085 -32.475 -12.755 ;
        RECT -32.805 -14.445 -32.475 -14.115 ;
        RECT -32.805 -15.805 -32.475 -15.475 ;
        RECT -32.805 -17.165 -32.475 -16.835 ;
        RECT -32.805 -18.525 -32.475 -18.195 ;
        RECT -32.805 -25.325 -32.475 -24.995 ;
        RECT -32.805 -26.685 -32.475 -26.355 ;
        RECT -32.805 -28.045 -32.475 -27.715 ;
        RECT -32.805 -29.405 -32.475 -29.075 ;
        RECT -32.805 -30.765 -32.475 -30.435 ;
        RECT -32.805 -32.125 -32.475 -31.795 ;
        RECT -32.805 -33.485 -32.475 -33.155 ;
        RECT -32.805 -34.845 -32.475 -34.515 ;
        RECT -32.805 -36.205 -32.475 -35.875 ;
        RECT -32.805 -37.565 -32.475 -37.235 ;
        RECT -32.805 -38.925 -32.475 -38.595 ;
        RECT -32.805 -40.285 -32.475 -39.955 ;
        RECT -32.805 -43.005 -32.475 -42.675 ;
        RECT -32.805 -44.365 -32.475 -44.035 ;
        RECT -32.805 -45.725 -32.475 -45.395 ;
        RECT -32.805 -47.085 -32.475 -46.755 ;
        RECT -32.805 -48.445 -32.475 -48.115 ;
        RECT -32.805 -49.805 -32.475 -49.475 ;
        RECT -32.805 -51.165 -32.475 -50.835 ;
        RECT -32.805 -52.525 -32.475 -52.195 ;
        RECT -32.805 -53.885 -32.475 -53.555 ;
        RECT -32.805 -55.245 -32.475 -54.915 ;
        RECT -32.805 -56.605 -32.475 -56.275 ;
        RECT -32.805 -57.965 -32.475 -57.635 ;
        RECT -32.805 -59.325 -32.475 -58.995 ;
        RECT -32.805 -60.685 -32.475 -60.355 ;
        RECT -32.805 -62.045 -32.475 -61.715 ;
        RECT -32.805 -63.405 -32.475 -63.075 ;
        RECT -32.805 -64.765 -32.475 -64.435 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 44.8 -54.235 45.93 ;
        RECT -54.565 39.955 -54.235 40.285 ;
        RECT -54.565 38.595 -54.235 38.925 ;
        RECT -54.565 37.235 -54.235 37.565 ;
        RECT -54.565 35.875 -54.235 36.205 ;
        RECT -54.565 34.515 -54.235 34.845 ;
        RECT -54.565 33.155 -54.235 33.485 ;
        RECT -54.565 31.795 -54.235 32.125 ;
        RECT -54.565 30.435 -54.235 30.765 ;
        RECT -54.565 29.075 -54.235 29.405 ;
        RECT -54.565 27.715 -54.235 28.045 ;
        RECT -54.565 26.355 -54.235 26.685 ;
        RECT -54.565 24.995 -54.235 25.325 ;
        RECT -54.565 22.66 -54.235 22.99 ;
        RECT -54.565 20.485 -54.235 20.815 ;
        RECT -54.565 19.635 -54.235 19.965 ;
        RECT -54.565 17.325 -54.235 17.655 ;
        RECT -54.565 16.475 -54.235 16.805 ;
        RECT -54.565 14.3 -54.235 14.63 ;
        RECT -54.565 11.395 -54.235 11.725 ;
        RECT -54.565 10.035 -54.235 10.365 ;
        RECT -54.565 8.675 -54.235 9.005 ;
        RECT -54.565 7.315 -54.235 7.645 ;
        RECT -54.565 5.955 -54.235 6.285 ;
        RECT -54.565 4.595 -54.235 4.925 ;
        RECT -54.565 3.235 -54.235 3.565 ;
        RECT -54.565 1.875 -54.235 2.205 ;
        RECT -54.565 0.515 -54.235 0.845 ;
        RECT -54.565 -0.845 -54.235 -0.515 ;
        RECT -54.565 -2.205 -54.235 -1.875 ;
        RECT -54.565 -3.565 -54.235 -3.235 ;
        RECT -54.565 -4.925 -54.235 -4.595 ;
        RECT -54.565 -6.285 -54.235 -5.955 ;
        RECT -54.565 -7.645 -54.235 -7.315 ;
        RECT -54.565 -9.005 -54.235 -8.675 ;
        RECT -54.565 -10.365 -54.235 -10.035 ;
        RECT -54.565 -11.725 -54.235 -11.395 ;
        RECT -54.565 -13.085 -54.235 -12.755 ;
        RECT -54.565 -14.445 -54.235 -14.115 ;
        RECT -54.565 -15.805 -54.235 -15.475 ;
        RECT -54.565 -17.165 -54.235 -16.835 ;
        RECT -54.565 -18.525 -54.235 -18.195 ;
        RECT -54.565 -19.885 -54.235 -19.555 ;
        RECT -54.565 -21.245 -54.235 -20.915 ;
        RECT -54.565 -22.605 -54.235 -22.275 ;
        RECT -54.565 -23.965 -54.235 -23.635 ;
        RECT -54.565 -25.325 -54.235 -24.995 ;
        RECT -54.565 -26.685 -54.235 -26.355 ;
        RECT -54.565 -28.045 -54.235 -27.715 ;
        RECT -54.565 -29.405 -54.235 -29.075 ;
        RECT -54.565 -30.765 -54.235 -30.435 ;
        RECT -54.565 -32.125 -54.235 -31.795 ;
        RECT -54.565 -33.485 -54.235 -33.155 ;
        RECT -54.565 -34.845 -54.235 -34.515 ;
        RECT -54.565 -36.205 -54.235 -35.875 ;
        RECT -54.565 -37.565 -54.235 -37.235 ;
        RECT -54.565 -38.925 -54.235 -38.595 ;
        RECT -54.565 -40.285 -54.235 -39.955 ;
        RECT -54.565 -41.645 -54.235 -41.315 ;
        RECT -54.565 -43.005 -54.235 -42.675 ;
        RECT -54.565 -44.365 -54.235 -44.035 ;
        RECT -54.565 -45.725 -54.235 -45.395 ;
        RECT -54.565 -47.085 -54.235 -46.755 ;
        RECT -54.565 -48.445 -54.235 -48.115 ;
        RECT -54.565 -49.805 -54.235 -49.475 ;
        RECT -54.565 -51.165 -54.235 -50.835 ;
        RECT -54.565 -52.525 -54.235 -52.195 ;
        RECT -54.565 -53.885 -54.235 -53.555 ;
        RECT -54.565 -55.245 -54.235 -54.915 ;
        RECT -54.565 -56.605 -54.235 -56.275 ;
        RECT -54.565 -57.965 -54.235 -57.635 ;
        RECT -54.565 -59.325 -54.235 -58.995 ;
        RECT -54.565 -60.685 -54.235 -60.355 ;
        RECT -54.565 -62.045 -54.235 -61.715 ;
        RECT -54.565 -63.405 -54.235 -63.075 ;
        RECT -54.565 -64.765 -54.235 -64.435 ;
        RECT -54.565 -66.125 -54.235 -65.795 ;
        RECT -54.565 -67.485 -54.235 -67.155 ;
        RECT -54.565 -68.845 -54.235 -68.515 ;
        RECT -54.565 -70.205 -54.235 -69.875 ;
        RECT -54.565 -71.565 -54.235 -71.235 ;
        RECT -54.565 -72.925 -54.235 -72.595 ;
        RECT -54.565 -74.285 -54.235 -73.955 ;
        RECT -54.565 -75.645 -54.235 -75.315 ;
        RECT -54.565 -77.005 -54.235 -76.675 ;
        RECT -54.565 -78.365 -54.235 -78.035 ;
        RECT -54.565 -79.725 -54.235 -79.395 ;
        RECT -54.565 -81.085 -54.235 -80.755 ;
        RECT -54.565 -82.445 -54.235 -82.115 ;
        RECT -54.565 -83.805 -54.235 -83.475 ;
        RECT -54.565 -85.165 -54.235 -84.835 ;
        RECT -54.565 -86.525 -54.235 -86.195 ;
        RECT -54.565 -87.885 -54.235 -87.555 ;
        RECT -54.565 -89.245 -54.235 -88.915 ;
        RECT -54.565 -90.605 -54.235 -90.275 ;
        RECT -54.565 -91.965 -54.235 -91.635 ;
        RECT -54.565 -93.325 -54.235 -92.995 ;
        RECT -54.565 -94.685 -54.235 -94.355 ;
        RECT -54.565 -96.045 -54.235 -95.715 ;
        RECT -54.565 -97.405 -54.235 -97.075 ;
        RECT -54.565 -98.765 -54.235 -98.435 ;
        RECT -54.565 -100.125 -54.235 -99.795 ;
        RECT -54.565 -101.485 -54.235 -101.155 ;
        RECT -54.565 -102.845 -54.235 -102.515 ;
        RECT -54.565 -104.205 -54.235 -103.875 ;
        RECT -54.565 -105.565 -54.235 -105.235 ;
        RECT -54.565 -106.925 -54.235 -106.595 ;
        RECT -54.565 -108.285 -54.235 -107.955 ;
        RECT -54.565 -109.645 -54.235 -109.315 ;
        RECT -54.565 -111.005 -54.235 -110.675 ;
        RECT -54.565 -112.365 -54.235 -112.035 ;
        RECT -54.565 -113.725 -54.235 -113.395 ;
        RECT -54.565 -115.085 -54.235 -114.755 ;
        RECT -54.565 -116.445 -54.235 -116.115 ;
        RECT -54.565 -117.805 -54.235 -117.475 ;
        RECT -54.565 -119.165 -54.235 -118.835 ;
        RECT -54.565 -120.525 -54.235 -120.195 ;
        RECT -54.565 -121.885 -54.235 -121.555 ;
        RECT -54.565 -123.245 -54.235 -122.915 ;
        RECT -54.565 -124.605 -54.235 -124.275 ;
        RECT -54.565 -125.965 -54.235 -125.635 ;
        RECT -54.565 -127.325 -54.235 -126.995 ;
        RECT -54.565 -128.685 -54.235 -128.355 ;
        RECT -54.565 -130.045 -54.235 -129.715 ;
        RECT -54.565 -131.405 -54.235 -131.075 ;
        RECT -54.565 -132.765 -54.235 -132.435 ;
        RECT -54.565 -134.125 -54.235 -133.795 ;
        RECT -54.565 -135.485 -54.235 -135.155 ;
        RECT -54.565 -136.845 -54.235 -136.515 ;
        RECT -54.565 -138.205 -54.235 -137.875 ;
        RECT -54.565 -139.565 -54.235 -139.235 ;
        RECT -54.565 -140.925 -54.235 -140.595 ;
        RECT -54.565 -142.285 -54.235 -141.955 ;
        RECT -54.565 -143.645 -54.235 -143.315 ;
        RECT -54.565 -145.005 -54.235 -144.675 ;
        RECT -54.565 -146.365 -54.235 -146.035 ;
        RECT -54.565 -147.725 -54.235 -147.395 ;
        RECT -54.565 -149.085 -54.235 -148.755 ;
        RECT -54.565 -150.445 -54.235 -150.115 ;
        RECT -54.565 -151.805 -54.235 -151.475 ;
        RECT -54.565 -153.165 -54.235 -152.835 ;
        RECT -54.565 -158.81 -54.235 -157.68 ;
        RECT -54.56 -158.925 -54.24 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.205 44.8 -52.875 45.93 ;
        RECT -53.205 39.955 -52.875 40.285 ;
        RECT -53.205 38.595 -52.875 38.925 ;
        RECT -53.205 37.235 -52.875 37.565 ;
        RECT -53.205 35.875 -52.875 36.205 ;
        RECT -53.205 34.515 -52.875 34.845 ;
        RECT -53.205 33.155 -52.875 33.485 ;
        RECT -53.205 31.795 -52.875 32.125 ;
        RECT -53.205 30.435 -52.875 30.765 ;
        RECT -53.205 29.075 -52.875 29.405 ;
        RECT -53.205 27.715 -52.875 28.045 ;
        RECT -53.205 26.355 -52.875 26.685 ;
        RECT -53.205 24.995 -52.875 25.325 ;
        RECT -53.205 22.66 -52.875 22.99 ;
        RECT -53.205 20.485 -52.875 20.815 ;
        RECT -53.205 19.635 -52.875 19.965 ;
        RECT -53.205 17.325 -52.875 17.655 ;
        RECT -53.205 16.475 -52.875 16.805 ;
        RECT -53.205 14.3 -52.875 14.63 ;
        RECT -53.205 11.395 -52.875 11.725 ;
        RECT -53.205 10.035 -52.875 10.365 ;
        RECT -53.205 8.675 -52.875 9.005 ;
        RECT -53.205 7.315 -52.875 7.645 ;
        RECT -53.205 5.955 -52.875 6.285 ;
        RECT -53.205 4.595 -52.875 4.925 ;
        RECT -53.205 3.235 -52.875 3.565 ;
        RECT -53.205 1.875 -52.875 2.205 ;
        RECT -53.205 0.515 -52.875 0.845 ;
        RECT -53.205 -0.845 -52.875 -0.515 ;
        RECT -53.205 -2.205 -52.875 -1.875 ;
        RECT -53.205 -3.565 -52.875 -3.235 ;
        RECT -53.205 -4.925 -52.875 -4.595 ;
        RECT -53.205 -6.285 -52.875 -5.955 ;
        RECT -53.205 -7.645 -52.875 -7.315 ;
        RECT -53.205 -9.005 -52.875 -8.675 ;
        RECT -53.205 -10.365 -52.875 -10.035 ;
        RECT -53.205 -11.725 -52.875 -11.395 ;
        RECT -53.205 -13.085 -52.875 -12.755 ;
        RECT -53.205 -14.445 -52.875 -14.115 ;
        RECT -53.205 -15.805 -52.875 -15.475 ;
        RECT -53.205 -17.165 -52.875 -16.835 ;
        RECT -53.205 -18.525 -52.875 -18.195 ;
        RECT -53.205 -19.885 -52.875 -19.555 ;
        RECT -53.205 -21.245 -52.875 -20.915 ;
        RECT -53.205 -22.605 -52.875 -22.275 ;
        RECT -53.205 -23.965 -52.875 -23.635 ;
        RECT -53.205 -25.325 -52.875 -24.995 ;
        RECT -53.205 -26.685 -52.875 -26.355 ;
        RECT -53.205 -28.045 -52.875 -27.715 ;
        RECT -53.205 -29.405 -52.875 -29.075 ;
        RECT -53.205 -30.765 -52.875 -30.435 ;
        RECT -53.205 -32.125 -52.875 -31.795 ;
        RECT -53.205 -33.485 -52.875 -33.155 ;
        RECT -53.205 -34.845 -52.875 -34.515 ;
        RECT -53.205 -36.205 -52.875 -35.875 ;
        RECT -53.205 -37.565 -52.875 -37.235 ;
        RECT -53.205 -38.925 -52.875 -38.595 ;
        RECT -53.205 -40.285 -52.875 -39.955 ;
        RECT -53.205 -41.645 -52.875 -41.315 ;
        RECT -53.205 -43.005 -52.875 -42.675 ;
        RECT -53.205 -44.365 -52.875 -44.035 ;
        RECT -53.205 -45.725 -52.875 -45.395 ;
        RECT -53.205 -47.085 -52.875 -46.755 ;
        RECT -53.205 -48.445 -52.875 -48.115 ;
        RECT -53.205 -49.805 -52.875 -49.475 ;
        RECT -53.205 -51.165 -52.875 -50.835 ;
        RECT -53.205 -52.525 -52.875 -52.195 ;
        RECT -53.205 -53.885 -52.875 -53.555 ;
        RECT -53.205 -55.245 -52.875 -54.915 ;
        RECT -53.205 -56.605 -52.875 -56.275 ;
        RECT -53.205 -57.965 -52.875 -57.635 ;
        RECT -53.205 -59.325 -52.875 -58.995 ;
        RECT -53.205 -60.685 -52.875 -60.355 ;
        RECT -53.205 -62.045 -52.875 -61.715 ;
        RECT -53.205 -63.405 -52.875 -63.075 ;
        RECT -53.205 -64.765 -52.875 -64.435 ;
        RECT -53.205 -66.125 -52.875 -65.795 ;
        RECT -53.205 -67.485 -52.875 -67.155 ;
        RECT -53.205 -68.845 -52.875 -68.515 ;
        RECT -53.205 -70.205 -52.875 -69.875 ;
        RECT -53.205 -71.565 -52.875 -71.235 ;
        RECT -53.205 -72.925 -52.875 -72.595 ;
        RECT -53.205 -74.285 -52.875 -73.955 ;
        RECT -53.205 -75.645 -52.875 -75.315 ;
        RECT -53.205 -77.005 -52.875 -76.675 ;
        RECT -53.205 -78.365 -52.875 -78.035 ;
        RECT -53.205 -79.725 -52.875 -79.395 ;
        RECT -53.205 -81.085 -52.875 -80.755 ;
        RECT -53.205 -82.445 -52.875 -82.115 ;
        RECT -53.205 -83.805 -52.875 -83.475 ;
        RECT -53.205 -85.165 -52.875 -84.835 ;
        RECT -53.205 -86.525 -52.875 -86.195 ;
        RECT -53.205 -87.885 -52.875 -87.555 ;
        RECT -53.205 -89.245 -52.875 -88.915 ;
        RECT -53.205 -90.605 -52.875 -90.275 ;
        RECT -53.205 -91.965 -52.875 -91.635 ;
        RECT -53.205 -93.325 -52.875 -92.995 ;
        RECT -53.205 -94.685 -52.875 -94.355 ;
        RECT -53.205 -96.045 -52.875 -95.715 ;
        RECT -53.205 -97.405 -52.875 -97.075 ;
        RECT -53.205 -98.765 -52.875 -98.435 ;
        RECT -53.205 -100.125 -52.875 -99.795 ;
        RECT -53.205 -101.485 -52.875 -101.155 ;
        RECT -53.205 -102.845 -52.875 -102.515 ;
        RECT -53.205 -104.205 -52.875 -103.875 ;
        RECT -53.205 -105.565 -52.875 -105.235 ;
        RECT -53.205 -106.925 -52.875 -106.595 ;
        RECT -53.205 -108.285 -52.875 -107.955 ;
        RECT -53.205 -109.645 -52.875 -109.315 ;
        RECT -53.205 -111.005 -52.875 -110.675 ;
        RECT -53.205 -112.365 -52.875 -112.035 ;
        RECT -53.205 -113.725 -52.875 -113.395 ;
        RECT -53.205 -115.085 -52.875 -114.755 ;
        RECT -53.205 -116.445 -52.875 -116.115 ;
        RECT -53.205 -117.805 -52.875 -117.475 ;
        RECT -53.205 -119.165 -52.875 -118.835 ;
        RECT -53.205 -120.525 -52.875 -120.195 ;
        RECT -53.205 -121.885 -52.875 -121.555 ;
        RECT -53.205 -123.245 -52.875 -122.915 ;
        RECT -53.205 -124.605 -52.875 -124.275 ;
        RECT -53.205 -125.965 -52.875 -125.635 ;
        RECT -53.205 -127.325 -52.875 -126.995 ;
        RECT -53.205 -128.685 -52.875 -128.355 ;
        RECT -53.205 -130.045 -52.875 -129.715 ;
        RECT -53.205 -131.405 -52.875 -131.075 ;
        RECT -53.205 -132.765 -52.875 -132.435 ;
        RECT -53.205 -134.125 -52.875 -133.795 ;
        RECT -53.205 -135.485 -52.875 -135.155 ;
        RECT -53.205 -136.845 -52.875 -136.515 ;
        RECT -53.205 -138.205 -52.875 -137.875 ;
        RECT -53.205 -139.565 -52.875 -139.235 ;
        RECT -53.205 -140.925 -52.875 -140.595 ;
        RECT -53.205 -142.285 -52.875 -141.955 ;
        RECT -53.205 -143.755 -52.875 -143.425 ;
        RECT -53.205 -145.005 -52.875 -144.675 ;
        RECT -53.205 -146.365 -52.875 -146.035 ;
        RECT -53.205 -149.085 -52.875 -148.755 ;
        RECT -53.205 -151.805 -52.875 -151.475 ;
        RECT -53.205 -153.165 -52.875 -152.835 ;
        RECT -53.205 -158.81 -52.875 -157.68 ;
        RECT -53.2 -158.925 -52.88 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.845 44.8 -51.515 45.93 ;
        RECT -51.845 39.955 -51.515 40.285 ;
        RECT -51.845 38.595 -51.515 38.925 ;
        RECT -51.845 37.235 -51.515 37.565 ;
        RECT -51.845 35.875 -51.515 36.205 ;
        RECT -51.845 34.515 -51.515 34.845 ;
        RECT -51.845 33.155 -51.515 33.485 ;
        RECT -51.845 31.795 -51.515 32.125 ;
        RECT -51.845 30.435 -51.515 30.765 ;
        RECT -51.845 29.075 -51.515 29.405 ;
        RECT -51.845 27.715 -51.515 28.045 ;
        RECT -51.845 26.355 -51.515 26.685 ;
        RECT -51.845 24.995 -51.515 25.325 ;
        RECT -51.845 22.66 -51.515 22.99 ;
        RECT -51.845 20.485 -51.515 20.815 ;
        RECT -51.845 19.635 -51.515 19.965 ;
        RECT -51.845 17.325 -51.515 17.655 ;
        RECT -51.845 16.475 -51.515 16.805 ;
        RECT -51.845 14.3 -51.515 14.63 ;
        RECT -51.845 11.395 -51.515 11.725 ;
        RECT -51.845 10.035 -51.515 10.365 ;
        RECT -51.845 8.675 -51.515 9.005 ;
        RECT -51.845 7.315 -51.515 7.645 ;
        RECT -51.845 5.955 -51.515 6.285 ;
        RECT -51.845 4.595 -51.515 4.925 ;
        RECT -51.845 3.235 -51.515 3.565 ;
        RECT -51.84 2.56 -51.52 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.845 -10.365 -51.515 -10.035 ;
        RECT -51.845 -11.725 -51.515 -11.395 ;
        RECT -51.845 -13.085 -51.515 -12.755 ;
        RECT -51.845 -14.445 -51.515 -14.115 ;
        RECT -51.845 -15.805 -51.515 -15.475 ;
        RECT -51.845 -17.165 -51.515 -16.835 ;
        RECT -51.845 -18.525 -51.515 -18.195 ;
        RECT -51.845 -19.885 -51.515 -19.555 ;
        RECT -51.845 -21.245 -51.515 -20.915 ;
        RECT -51.845 -22.605 -51.515 -22.275 ;
        RECT -51.845 -23.965 -51.515 -23.635 ;
        RECT -51.845 -25.325 -51.515 -24.995 ;
        RECT -51.845 -26.685 -51.515 -26.355 ;
        RECT -51.845 -28.045 -51.515 -27.715 ;
        RECT -51.845 -29.405 -51.515 -29.075 ;
        RECT -51.845 -30.765 -51.515 -30.435 ;
        RECT -51.845 -32.125 -51.515 -31.795 ;
        RECT -51.845 -33.485 -51.515 -33.155 ;
        RECT -51.845 -34.845 -51.515 -34.515 ;
        RECT -51.845 -36.205 -51.515 -35.875 ;
        RECT -51.845 -37.565 -51.515 -37.235 ;
        RECT -51.845 -38.925 -51.515 -38.595 ;
        RECT -51.845 -40.285 -51.515 -39.955 ;
        RECT -51.845 -41.645 -51.515 -41.315 ;
        RECT -51.845 -43.005 -51.515 -42.675 ;
        RECT -51.845 -44.365 -51.515 -44.035 ;
        RECT -51.845 -45.725 -51.515 -45.395 ;
        RECT -51.845 -47.085 -51.515 -46.755 ;
        RECT -51.845 -48.445 -51.515 -48.115 ;
        RECT -51.845 -49.805 -51.515 -49.475 ;
        RECT -51.845 -51.165 -51.515 -50.835 ;
        RECT -51.845 -52.525 -51.515 -52.195 ;
        RECT -51.845 -53.885 -51.515 -53.555 ;
        RECT -51.845 -55.245 -51.515 -54.915 ;
        RECT -51.845 -56.605 -51.515 -56.275 ;
        RECT -51.845 -57.965 -51.515 -57.635 ;
        RECT -51.845 -59.325 -51.515 -58.995 ;
        RECT -51.845 -60.685 -51.515 -60.355 ;
        RECT -51.845 -62.045 -51.515 -61.715 ;
        RECT -51.845 -63.405 -51.515 -63.075 ;
        RECT -51.845 -64.765 -51.515 -64.435 ;
        RECT -51.845 -66.125 -51.515 -65.795 ;
        RECT -51.845 -67.485 -51.515 -67.155 ;
        RECT -51.845 -68.845 -51.515 -68.515 ;
        RECT -51.845 -70.205 -51.515 -69.875 ;
        RECT -51.845 -71.565 -51.515 -71.235 ;
        RECT -51.845 -72.925 -51.515 -72.595 ;
        RECT -51.845 -74.285 -51.515 -73.955 ;
        RECT -51.845 -75.645 -51.515 -75.315 ;
        RECT -51.845 -77.005 -51.515 -76.675 ;
        RECT -51.845 -78.365 -51.515 -78.035 ;
        RECT -51.845 -79.725 -51.515 -79.395 ;
        RECT -51.845 -81.085 -51.515 -80.755 ;
        RECT -51.845 -82.445 -51.515 -82.115 ;
        RECT -51.845 -83.805 -51.515 -83.475 ;
        RECT -51.845 -85.165 -51.515 -84.835 ;
        RECT -51.845 -86.525 -51.515 -86.195 ;
        RECT -51.845 -87.885 -51.515 -87.555 ;
        RECT -51.845 -89.245 -51.515 -88.915 ;
        RECT -51.845 -90.605 -51.515 -90.275 ;
        RECT -51.845 -91.965 -51.515 -91.635 ;
        RECT -51.845 -93.325 -51.515 -92.995 ;
        RECT -51.845 -94.685 -51.515 -94.355 ;
        RECT -51.845 -96.045 -51.515 -95.715 ;
        RECT -51.845 -97.405 -51.515 -97.075 ;
        RECT -51.845 -98.765 -51.515 -98.435 ;
        RECT -51.845 -100.125 -51.515 -99.795 ;
        RECT -51.845 -101.485 -51.515 -101.155 ;
        RECT -51.845 -102.845 -51.515 -102.515 ;
        RECT -51.845 -104.205 -51.515 -103.875 ;
        RECT -51.845 -105.565 -51.515 -105.235 ;
        RECT -51.845 -106.925 -51.515 -106.595 ;
        RECT -51.845 -108.285 -51.515 -107.955 ;
        RECT -51.845 -109.645 -51.515 -109.315 ;
        RECT -51.845 -111.005 -51.515 -110.675 ;
        RECT -51.845 -112.365 -51.515 -112.035 ;
        RECT -51.845 -113.725 -51.515 -113.395 ;
        RECT -51.845 -115.085 -51.515 -114.755 ;
        RECT -51.845 -116.445 -51.515 -116.115 ;
        RECT -51.845 -117.805 -51.515 -117.475 ;
        RECT -51.845 -119.165 -51.515 -118.835 ;
        RECT -51.845 -120.525 -51.515 -120.195 ;
        RECT -51.845 -121.885 -51.515 -121.555 ;
        RECT -51.845 -123.245 -51.515 -122.915 ;
        RECT -51.845 -124.605 -51.515 -124.275 ;
        RECT -51.845 -125.965 -51.515 -125.635 ;
        RECT -51.845 -127.325 -51.515 -126.995 ;
        RECT -51.845 -128.685 -51.515 -128.355 ;
        RECT -51.845 -130.045 -51.515 -129.715 ;
        RECT -51.845 -131.405 -51.515 -131.075 ;
        RECT -51.845 -132.765 -51.515 -132.435 ;
        RECT -51.845 -134.125 -51.515 -133.795 ;
        RECT -51.845 -135.485 -51.515 -135.155 ;
        RECT -51.845 -136.845 -51.515 -136.515 ;
        RECT -51.845 -138.205 -51.515 -137.875 ;
        RECT -51.845 -139.565 -51.515 -139.235 ;
        RECT -51.845 -140.925 -51.515 -140.595 ;
        RECT -51.845 -142.285 -51.515 -141.955 ;
        RECT -51.845 -143.755 -51.515 -143.425 ;
        RECT -51.845 -145.005 -51.515 -144.675 ;
        RECT -51.845 -146.365 -51.515 -146.035 ;
        RECT -51.845 -149.085 -51.515 -148.755 ;
        RECT -51.845 -151.805 -51.515 -151.475 ;
        RECT -51.845 -153.165 -51.515 -152.835 ;
        RECT -51.845 -158.81 -51.515 -157.68 ;
        RECT -51.84 -158.925 -51.52 -9.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.485 44.8 -50.155 45.93 ;
        RECT -50.485 39.955 -50.155 40.285 ;
        RECT -50.485 38.595 -50.155 38.925 ;
        RECT -50.485 37.235 -50.155 37.565 ;
        RECT -50.485 35.875 -50.155 36.205 ;
        RECT -50.485 34.515 -50.155 34.845 ;
        RECT -50.485 33.155 -50.155 33.485 ;
        RECT -50.485 31.795 -50.155 32.125 ;
        RECT -50.485 30.435 -50.155 30.765 ;
        RECT -50.485 29.075 -50.155 29.405 ;
        RECT -50.485 27.715 -50.155 28.045 ;
        RECT -50.485 26.355 -50.155 26.685 ;
        RECT -50.485 24.995 -50.155 25.325 ;
        RECT -50.48 24.32 -50.16 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.485 11.395 -50.155 11.725 ;
        RECT -50.485 10.035 -50.155 10.365 ;
        RECT -50.485 8.675 -50.155 9.005 ;
        RECT -50.485 7.315 -50.155 7.645 ;
        RECT -50.485 4.595 -50.155 4.925 ;
        RECT -50.485 3.235 -50.155 3.565 ;
        RECT -50.485 -0.845 -50.155 -0.515 ;
        RECT -50.485 -2.205 -50.155 -1.875 ;
        RECT -50.485 -3.565 -50.155 -3.235 ;
        RECT -50.485 -4.925 -50.155 -4.595 ;
        RECT -50.485 -6.285 -50.155 -5.955 ;
        RECT -50.485 -7.645 -50.155 -7.315 ;
        RECT -50.485 -10.365 -50.155 -10.035 ;
        RECT -50.485 -11.725 -50.155 -11.395 ;
        RECT -50.485 -13.085 -50.155 -12.755 ;
        RECT -50.485 -14.445 -50.155 -14.115 ;
        RECT -50.485 -15.805 -50.155 -15.475 ;
        RECT -50.485 -17.165 -50.155 -16.835 ;
        RECT -50.485 -18.525 -50.155 -18.195 ;
        RECT -50.485 -19.885 -50.155 -19.555 ;
        RECT -50.485 -21.245 -50.155 -20.915 ;
        RECT -50.485 -22.605 -50.155 -22.275 ;
        RECT -50.485 -23.965 -50.155 -23.635 ;
        RECT -50.485 -25.325 -50.155 -24.995 ;
        RECT -50.485 -26.685 -50.155 -26.355 ;
        RECT -50.485 -28.045 -50.155 -27.715 ;
        RECT -50.485 -29.405 -50.155 -29.075 ;
        RECT -50.485 -30.765 -50.155 -30.435 ;
        RECT -50.485 -32.125 -50.155 -31.795 ;
        RECT -50.485 -33.485 -50.155 -33.155 ;
        RECT -50.485 -34.845 -50.155 -34.515 ;
        RECT -50.485 -36.205 -50.155 -35.875 ;
        RECT -50.485 -37.565 -50.155 -37.235 ;
        RECT -50.485 -38.925 -50.155 -38.595 ;
        RECT -50.485 -40.285 -50.155 -39.955 ;
        RECT -50.485 -41.645 -50.155 -41.315 ;
        RECT -50.485 -43.005 -50.155 -42.675 ;
        RECT -50.485 -44.365 -50.155 -44.035 ;
        RECT -50.485 -45.725 -50.155 -45.395 ;
        RECT -50.485 -47.085 -50.155 -46.755 ;
        RECT -50.485 -48.445 -50.155 -48.115 ;
        RECT -50.485 -49.805 -50.155 -49.475 ;
        RECT -50.485 -51.165 -50.155 -50.835 ;
        RECT -50.485 -52.525 -50.155 -52.195 ;
        RECT -50.485 -53.885 -50.155 -53.555 ;
        RECT -50.485 -55.245 -50.155 -54.915 ;
        RECT -50.485 -56.605 -50.155 -56.275 ;
        RECT -50.485 -57.965 -50.155 -57.635 ;
        RECT -50.485 -59.325 -50.155 -58.995 ;
        RECT -50.485 -60.685 -50.155 -60.355 ;
        RECT -50.485 -62.045 -50.155 -61.715 ;
        RECT -50.485 -63.405 -50.155 -63.075 ;
        RECT -50.485 -64.765 -50.155 -64.435 ;
        RECT -50.485 -66.125 -50.155 -65.795 ;
        RECT -50.485 -67.485 -50.155 -67.155 ;
        RECT -50.485 -68.845 -50.155 -68.515 ;
        RECT -50.485 -70.205 -50.155 -69.875 ;
        RECT -50.485 -71.565 -50.155 -71.235 ;
        RECT -50.485 -72.925 -50.155 -72.595 ;
        RECT -50.485 -74.285 -50.155 -73.955 ;
        RECT -50.485 -75.645 -50.155 -75.315 ;
        RECT -50.485 -77.005 -50.155 -76.675 ;
        RECT -50.485 -78.365 -50.155 -78.035 ;
        RECT -50.485 -79.725 -50.155 -79.395 ;
        RECT -50.485 -81.085 -50.155 -80.755 ;
        RECT -50.485 -82.445 -50.155 -82.115 ;
        RECT -50.485 -83.805 -50.155 -83.475 ;
        RECT -50.485 -85.165 -50.155 -84.835 ;
        RECT -50.485 -86.525 -50.155 -86.195 ;
        RECT -50.485 -87.885 -50.155 -87.555 ;
        RECT -50.485 -89.245 -50.155 -88.915 ;
        RECT -50.485 -90.605 -50.155 -90.275 ;
        RECT -50.485 -91.965 -50.155 -91.635 ;
        RECT -50.485 -93.325 -50.155 -92.995 ;
        RECT -50.485 -94.685 -50.155 -94.355 ;
        RECT -50.485 -96.045 -50.155 -95.715 ;
        RECT -50.485 -97.405 -50.155 -97.075 ;
        RECT -50.485 -98.765 -50.155 -98.435 ;
        RECT -50.485 -100.125 -50.155 -99.795 ;
        RECT -50.485 -101.485 -50.155 -101.155 ;
        RECT -50.485 -102.845 -50.155 -102.515 ;
        RECT -50.485 -104.205 -50.155 -103.875 ;
        RECT -50.485 -105.565 -50.155 -105.235 ;
        RECT -50.485 -106.925 -50.155 -106.595 ;
        RECT -50.485 -108.285 -50.155 -107.955 ;
        RECT -50.485 -109.645 -50.155 -109.315 ;
        RECT -50.485 -111.005 -50.155 -110.675 ;
        RECT -50.485 -112.365 -50.155 -112.035 ;
        RECT -50.485 -113.725 -50.155 -113.395 ;
        RECT -50.485 -115.085 -50.155 -114.755 ;
        RECT -50.485 -116.445 -50.155 -116.115 ;
        RECT -50.485 -117.805 -50.155 -117.475 ;
        RECT -50.485 -119.165 -50.155 -118.835 ;
        RECT -50.485 -120.525 -50.155 -120.195 ;
        RECT -50.485 -121.885 -50.155 -121.555 ;
        RECT -50.485 -123.245 -50.155 -122.915 ;
        RECT -50.485 -124.605 -50.155 -124.275 ;
        RECT -50.485 -125.965 -50.155 -125.635 ;
        RECT -50.485 -127.325 -50.155 -126.995 ;
        RECT -50.485 -128.685 -50.155 -128.355 ;
        RECT -50.485 -130.045 -50.155 -129.715 ;
        RECT -50.485 -131.405 -50.155 -131.075 ;
        RECT -50.485 -132.765 -50.155 -132.435 ;
        RECT -50.485 -134.125 -50.155 -133.795 ;
        RECT -50.485 -135.485 -50.155 -135.155 ;
        RECT -50.485 -136.845 -50.155 -136.515 ;
        RECT -50.485 -138.205 -50.155 -137.875 ;
        RECT -50.485 -139.565 -50.155 -139.235 ;
        RECT -50.485 -140.925 -50.155 -140.595 ;
        RECT -50.485 -142.285 -50.155 -141.955 ;
        RECT -50.485 -143.755 -50.155 -143.425 ;
        RECT -50.485 -145.005 -50.155 -144.675 ;
        RECT -50.485 -146.365 -50.155 -146.035 ;
        RECT -50.485 -147.725 -50.155 -147.395 ;
        RECT -50.485 -149.085 -50.155 -148.755 ;
        RECT -50.485 -151.805 -50.155 -151.475 ;
        RECT -50.485 -153.165 -50.155 -152.835 ;
        RECT -50.485 -158.81 -50.155 -157.68 ;
        RECT -50.48 -158.925 -50.16 12.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.125 44.8 -48.795 45.93 ;
        RECT -49.125 39.955 -48.795 40.285 ;
        RECT -49.125 38.595 -48.795 38.925 ;
        RECT -49.125 37.235 -48.795 37.565 ;
        RECT -49.125 35.875 -48.795 36.205 ;
        RECT -49.125 34.515 -48.795 34.845 ;
        RECT -49.125 33.155 -48.795 33.485 ;
        RECT -49.125 31.795 -48.795 32.125 ;
        RECT -49.125 30.435 -48.795 30.765 ;
        RECT -49.125 29.075 -48.795 29.405 ;
        RECT -49.125 27.715 -48.795 28.045 ;
        RECT -49.125 26.355 -48.795 26.685 ;
        RECT -49.125 24.995 -48.795 25.325 ;
        RECT -49.12 24.32 -48.8 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.125 11.395 -48.795 11.725 ;
        RECT -49.125 10.035 -48.795 10.365 ;
        RECT -49.125 8.675 -48.795 9.005 ;
        RECT -49.125 7.315 -48.795 7.645 ;
        RECT -49.125 4.595 -48.795 4.925 ;
        RECT -49.125 3.235 -48.795 3.565 ;
        RECT -49.125 -0.845 -48.795 -0.515 ;
        RECT -49.125 -2.205 -48.795 -1.875 ;
        RECT -49.125 -3.565 -48.795 -3.235 ;
        RECT -49.125 -4.925 -48.795 -4.595 ;
        RECT -49.125 -6.285 -48.795 -5.955 ;
        RECT -49.125 -7.645 -48.795 -7.315 ;
        RECT -49.125 -10.365 -48.795 -10.035 ;
        RECT -49.125 -11.725 -48.795 -11.395 ;
        RECT -49.125 -13.085 -48.795 -12.755 ;
        RECT -49.125 -14.445 -48.795 -14.115 ;
        RECT -49.125 -15.805 -48.795 -15.475 ;
        RECT -49.125 -17.165 -48.795 -16.835 ;
        RECT -49.125 -18.525 -48.795 -18.195 ;
        RECT -49.125 -19.885 -48.795 -19.555 ;
        RECT -49.125 -21.245 -48.795 -20.915 ;
        RECT -49.125 -22.605 -48.795 -22.275 ;
        RECT -49.125 -23.965 -48.795 -23.635 ;
        RECT -49.125 -25.325 -48.795 -24.995 ;
        RECT -49.125 -26.685 -48.795 -26.355 ;
        RECT -49.125 -28.045 -48.795 -27.715 ;
        RECT -49.125 -29.405 -48.795 -29.075 ;
        RECT -49.125 -30.765 -48.795 -30.435 ;
        RECT -49.125 -32.125 -48.795 -31.795 ;
        RECT -49.125 -33.485 -48.795 -33.155 ;
        RECT -49.125 -34.845 -48.795 -34.515 ;
        RECT -49.125 -36.205 -48.795 -35.875 ;
        RECT -49.125 -37.565 -48.795 -37.235 ;
        RECT -49.125 -38.925 -48.795 -38.595 ;
        RECT -49.125 -40.285 -48.795 -39.955 ;
        RECT -49.125 -41.645 -48.795 -41.315 ;
        RECT -49.125 -43.005 -48.795 -42.675 ;
        RECT -49.125 -44.365 -48.795 -44.035 ;
        RECT -49.125 -45.725 -48.795 -45.395 ;
        RECT -49.125 -47.085 -48.795 -46.755 ;
        RECT -49.125 -48.445 -48.795 -48.115 ;
        RECT -49.125 -49.805 -48.795 -49.475 ;
        RECT -49.125 -51.165 -48.795 -50.835 ;
        RECT -49.125 -52.525 -48.795 -52.195 ;
        RECT -49.125 -53.885 -48.795 -53.555 ;
        RECT -49.125 -55.245 -48.795 -54.915 ;
        RECT -49.125 -56.605 -48.795 -56.275 ;
        RECT -49.125 -57.965 -48.795 -57.635 ;
        RECT -49.125 -59.325 -48.795 -58.995 ;
        RECT -49.125 -60.685 -48.795 -60.355 ;
        RECT -49.125 -62.045 -48.795 -61.715 ;
        RECT -49.125 -63.405 -48.795 -63.075 ;
        RECT -49.125 -64.765 -48.795 -64.435 ;
        RECT -49.125 -66.125 -48.795 -65.795 ;
        RECT -49.125 -67.485 -48.795 -67.155 ;
        RECT -49.125 -68.845 -48.795 -68.515 ;
        RECT -49.125 -70.205 -48.795 -69.875 ;
        RECT -49.125 -71.565 -48.795 -71.235 ;
        RECT -49.125 -72.925 -48.795 -72.595 ;
        RECT -49.125 -74.285 -48.795 -73.955 ;
        RECT -49.125 -75.645 -48.795 -75.315 ;
        RECT -49.125 -77.005 -48.795 -76.675 ;
        RECT -49.125 -78.365 -48.795 -78.035 ;
        RECT -49.125 -79.725 -48.795 -79.395 ;
        RECT -49.125 -81.085 -48.795 -80.755 ;
        RECT -49.125 -82.445 -48.795 -82.115 ;
        RECT -49.125 -83.805 -48.795 -83.475 ;
        RECT -49.125 -85.165 -48.795 -84.835 ;
        RECT -49.125 -86.525 -48.795 -86.195 ;
        RECT -49.125 -87.885 -48.795 -87.555 ;
        RECT -49.125 -89.245 -48.795 -88.915 ;
        RECT -49.125 -90.605 -48.795 -90.275 ;
        RECT -49.125 -91.965 -48.795 -91.635 ;
        RECT -49.125 -93.325 -48.795 -92.995 ;
        RECT -49.125 -94.685 -48.795 -94.355 ;
        RECT -49.125 -96.045 -48.795 -95.715 ;
        RECT -49.125 -97.405 -48.795 -97.075 ;
        RECT -49.125 -98.765 -48.795 -98.435 ;
        RECT -49.125 -100.125 -48.795 -99.795 ;
        RECT -49.125 -101.485 -48.795 -101.155 ;
        RECT -49.125 -102.845 -48.795 -102.515 ;
        RECT -49.125 -104.205 -48.795 -103.875 ;
        RECT -49.125 -105.565 -48.795 -105.235 ;
        RECT -49.125 -106.925 -48.795 -106.595 ;
        RECT -49.125 -108.285 -48.795 -107.955 ;
        RECT -49.125 -109.645 -48.795 -109.315 ;
        RECT -49.125 -111.005 -48.795 -110.675 ;
        RECT -49.125 -112.365 -48.795 -112.035 ;
        RECT -49.125 -113.725 -48.795 -113.395 ;
        RECT -49.125 -115.085 -48.795 -114.755 ;
        RECT -49.125 -116.445 -48.795 -116.115 ;
        RECT -49.125 -117.805 -48.795 -117.475 ;
        RECT -49.125 -119.165 -48.795 -118.835 ;
        RECT -49.125 -120.525 -48.795 -120.195 ;
        RECT -49.125 -121.885 -48.795 -121.555 ;
        RECT -49.125 -123.245 -48.795 -122.915 ;
        RECT -49.125 -124.605 -48.795 -124.275 ;
        RECT -49.125 -125.965 -48.795 -125.635 ;
        RECT -49.125 -127.325 -48.795 -126.995 ;
        RECT -49.125 -128.685 -48.795 -128.355 ;
        RECT -49.125 -130.045 -48.795 -129.715 ;
        RECT -49.125 -131.405 -48.795 -131.075 ;
        RECT -49.125 -132.765 -48.795 -132.435 ;
        RECT -49.125 -134.125 -48.795 -133.795 ;
        RECT -49.125 -135.485 -48.795 -135.155 ;
        RECT -49.125 -136.845 -48.795 -136.515 ;
        RECT -49.125 -138.205 -48.795 -137.875 ;
        RECT -49.125 -139.565 -48.795 -139.235 ;
        RECT -49.125 -140.925 -48.795 -140.595 ;
        RECT -49.12 -141.6 -48.8 12.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.125 -147.725 -48.795 -147.395 ;
        RECT -49.125 -149.085 -48.795 -148.755 ;
        RECT -49.125 -151.805 -48.795 -151.475 ;
        RECT -49.125 -153.165 -48.795 -152.835 ;
        RECT -49.125 -158.81 -48.795 -157.68 ;
        RECT -49.12 -158.925 -48.8 -147.395 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.765 44.8 -47.435 45.93 ;
        RECT -47.765 39.955 -47.435 40.285 ;
        RECT -47.765 38.595 -47.435 38.925 ;
        RECT -47.765 37.235 -47.435 37.565 ;
        RECT -47.765 35.875 -47.435 36.205 ;
        RECT -47.765 34.515 -47.435 34.845 ;
        RECT -47.765 33.155 -47.435 33.485 ;
        RECT -47.765 31.795 -47.435 32.125 ;
        RECT -47.765 30.435 -47.435 30.765 ;
        RECT -47.765 29.075 -47.435 29.405 ;
        RECT -47.765 27.715 -47.435 28.045 ;
        RECT -47.765 26.355 -47.435 26.685 ;
        RECT -47.765 24.995 -47.435 25.325 ;
        RECT -47.76 24.32 -47.44 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.765 11.395 -47.435 11.725 ;
        RECT -47.765 10.035 -47.435 10.365 ;
        RECT -47.765 8.675 -47.435 9.005 ;
        RECT -47.765 7.315 -47.435 7.645 ;
        RECT -47.765 4.595 -47.435 4.925 ;
        RECT -47.765 3.235 -47.435 3.565 ;
        RECT -47.765 -0.845 -47.435 -0.515 ;
        RECT -47.765 -2.205 -47.435 -1.875 ;
        RECT -47.765 -3.565 -47.435 -3.235 ;
        RECT -47.765 -4.925 -47.435 -4.595 ;
        RECT -47.765 -6.285 -47.435 -5.955 ;
        RECT -47.765 -7.645 -47.435 -7.315 ;
        RECT -47.765 -10.365 -47.435 -10.035 ;
        RECT -47.765 -11.725 -47.435 -11.395 ;
        RECT -47.765 -13.085 -47.435 -12.755 ;
        RECT -47.765 -14.445 -47.435 -14.115 ;
        RECT -47.765 -15.805 -47.435 -15.475 ;
        RECT -47.765 -17.165 -47.435 -16.835 ;
        RECT -47.765 -18.525 -47.435 -18.195 ;
        RECT -47.765 -19.885 -47.435 -19.555 ;
        RECT -47.765 -21.245 -47.435 -20.915 ;
        RECT -47.765 -22.605 -47.435 -22.275 ;
        RECT -47.765 -23.965 -47.435 -23.635 ;
        RECT -47.765 -25.325 -47.435 -24.995 ;
        RECT -47.765 -26.685 -47.435 -26.355 ;
        RECT -47.765 -28.045 -47.435 -27.715 ;
        RECT -47.765 -29.405 -47.435 -29.075 ;
        RECT -47.765 -30.765 -47.435 -30.435 ;
        RECT -47.765 -32.125 -47.435 -31.795 ;
        RECT -47.765 -33.485 -47.435 -33.155 ;
        RECT -47.765 -34.845 -47.435 -34.515 ;
        RECT -47.765 -36.205 -47.435 -35.875 ;
        RECT -47.765 -37.565 -47.435 -37.235 ;
        RECT -47.765 -38.925 -47.435 -38.595 ;
        RECT -47.765 -40.285 -47.435 -39.955 ;
        RECT -47.765 -41.645 -47.435 -41.315 ;
        RECT -47.765 -43.005 -47.435 -42.675 ;
        RECT -47.765 -44.365 -47.435 -44.035 ;
        RECT -47.765 -45.725 -47.435 -45.395 ;
        RECT -47.765 -47.085 -47.435 -46.755 ;
        RECT -47.765 -48.445 -47.435 -48.115 ;
        RECT -47.765 -49.805 -47.435 -49.475 ;
        RECT -47.765 -51.165 -47.435 -50.835 ;
        RECT -47.765 -52.525 -47.435 -52.195 ;
        RECT -47.765 -53.885 -47.435 -53.555 ;
        RECT -47.765 -55.245 -47.435 -54.915 ;
        RECT -47.765 -56.605 -47.435 -56.275 ;
        RECT -47.765 -57.965 -47.435 -57.635 ;
        RECT -47.765 -59.325 -47.435 -58.995 ;
        RECT -47.765 -60.685 -47.435 -60.355 ;
        RECT -47.765 -62.045 -47.435 -61.715 ;
        RECT -47.765 -63.405 -47.435 -63.075 ;
        RECT -47.765 -64.765 -47.435 -64.435 ;
        RECT -47.765 -66.125 -47.435 -65.795 ;
        RECT -47.765 -67.485 -47.435 -67.155 ;
        RECT -47.765 -68.845 -47.435 -68.515 ;
        RECT -47.765 -70.205 -47.435 -69.875 ;
        RECT -47.765 -71.565 -47.435 -71.235 ;
        RECT -47.765 -72.925 -47.435 -72.595 ;
        RECT -47.765 -74.285 -47.435 -73.955 ;
        RECT -47.765 -75.645 -47.435 -75.315 ;
        RECT -47.765 -77.005 -47.435 -76.675 ;
        RECT -47.765 -78.365 -47.435 -78.035 ;
        RECT -47.765 -79.725 -47.435 -79.395 ;
        RECT -47.765 -81.085 -47.435 -80.755 ;
        RECT -47.765 -82.445 -47.435 -82.115 ;
        RECT -47.765 -83.805 -47.435 -83.475 ;
        RECT -47.765 -85.165 -47.435 -84.835 ;
        RECT -47.76 -86.52 -47.44 12.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.765 -96.045 -47.435 -95.715 ;
        RECT -47.765 -97.405 -47.435 -97.075 ;
        RECT -47.765 -98.765 -47.435 -98.435 ;
        RECT -47.765 -100.125 -47.435 -99.795 ;
        RECT -47.765 -101.485 -47.435 -101.155 ;
        RECT -47.765 -102.845 -47.435 -102.515 ;
        RECT -47.765 -104.205 -47.435 -103.875 ;
        RECT -47.765 -105.565 -47.435 -105.235 ;
        RECT -47.765 -106.925 -47.435 -106.595 ;
        RECT -47.765 -108.285 -47.435 -107.955 ;
        RECT -47.765 -109.645 -47.435 -109.315 ;
        RECT -47.765 -111.005 -47.435 -110.675 ;
        RECT -47.765 -112.365 -47.435 -112.035 ;
        RECT -47.765 -113.725 -47.435 -113.395 ;
        RECT -47.765 -115.085 -47.435 -114.755 ;
        RECT -47.765 -116.445 -47.435 -116.115 ;
        RECT -47.765 -117.805 -47.435 -117.475 ;
        RECT -47.765 -119.165 -47.435 -118.835 ;
        RECT -47.765 -120.525 -47.435 -120.195 ;
        RECT -47.765 -121.885 -47.435 -121.555 ;
        RECT -47.765 -123.245 -47.435 -122.915 ;
        RECT -47.765 -124.605 -47.435 -124.275 ;
        RECT -47.765 -125.965 -47.435 -125.635 ;
        RECT -47.765 -127.325 -47.435 -126.995 ;
        RECT -47.765 -128.685 -47.435 -128.355 ;
        RECT -47.765 -130.045 -47.435 -129.715 ;
        RECT -47.765 -131.405 -47.435 -131.075 ;
        RECT -47.765 -132.765 -47.435 -132.435 ;
        RECT -47.765 -134.125 -47.435 -133.795 ;
        RECT -47.765 -135.485 -47.435 -135.155 ;
        RECT -47.765 -136.845 -47.435 -136.515 ;
        RECT -47.765 -138.205 -47.435 -137.875 ;
        RECT -47.765 -139.565 -47.435 -139.235 ;
        RECT -47.765 -140.925 -47.435 -140.595 ;
        RECT -47.765 -145.005 -47.435 -144.675 ;
        RECT -47.765 -146.365 -47.435 -146.035 ;
        RECT -47.765 -151.805 -47.435 -151.475 ;
        RECT -47.765 -153.165 -47.435 -152.835 ;
        RECT -47.765 -158.81 -47.435 -157.68 ;
        RECT -47.76 -158.925 -47.44 -95.715 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.405 44.8 -46.075 45.93 ;
        RECT -46.405 39.955 -46.075 40.285 ;
        RECT -46.405 38.595 -46.075 38.925 ;
        RECT -46.405 37.235 -46.075 37.565 ;
        RECT -46.405 35.875 -46.075 36.205 ;
        RECT -46.405 34.515 -46.075 34.845 ;
        RECT -46.405 33.155 -46.075 33.485 ;
        RECT -46.405 31.795 -46.075 32.125 ;
        RECT -46.405 30.435 -46.075 30.765 ;
        RECT -46.405 29.075 -46.075 29.405 ;
        RECT -46.405 27.715 -46.075 28.045 ;
        RECT -46.405 26.355 -46.075 26.685 ;
        RECT -46.405 24.995 -46.075 25.325 ;
        RECT -46.4 24.32 -46.08 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.405 11.395 -46.075 11.725 ;
        RECT -46.405 10.035 -46.075 10.365 ;
        RECT -46.405 8.675 -46.075 9.005 ;
        RECT -46.405 7.315 -46.075 7.645 ;
        RECT -46.405 4.595 -46.075 4.925 ;
        RECT -46.405 3.235 -46.075 3.565 ;
        RECT -46.405 -0.845 -46.075 -0.515 ;
        RECT -46.405 -2.205 -46.075 -1.875 ;
        RECT -46.405 -3.565 -46.075 -3.235 ;
        RECT -46.405 -4.925 -46.075 -4.595 ;
        RECT -46.405 -6.285 -46.075 -5.955 ;
        RECT -46.405 -7.645 -46.075 -7.315 ;
        RECT -46.405 -10.365 -46.075 -10.035 ;
        RECT -46.405 -11.725 -46.075 -11.395 ;
        RECT -46.405 -13.085 -46.075 -12.755 ;
        RECT -46.405 -14.445 -46.075 -14.115 ;
        RECT -46.405 -15.805 -46.075 -15.475 ;
        RECT -46.405 -17.165 -46.075 -16.835 ;
        RECT -46.405 -18.525 -46.075 -18.195 ;
        RECT -46.405 -19.885 -46.075 -19.555 ;
        RECT -46.405 -21.245 -46.075 -20.915 ;
        RECT -46.405 -22.605 -46.075 -22.275 ;
        RECT -46.405 -23.965 -46.075 -23.635 ;
        RECT -46.405 -25.325 -46.075 -24.995 ;
        RECT -46.405 -26.685 -46.075 -26.355 ;
        RECT -46.405 -28.045 -46.075 -27.715 ;
        RECT -46.405 -29.405 -46.075 -29.075 ;
        RECT -46.405 -30.765 -46.075 -30.435 ;
        RECT -46.405 -32.125 -46.075 -31.795 ;
        RECT -46.405 -33.485 -46.075 -33.155 ;
        RECT -46.405 -34.845 -46.075 -34.515 ;
        RECT -46.405 -36.205 -46.075 -35.875 ;
        RECT -46.405 -37.565 -46.075 -37.235 ;
        RECT -46.405 -38.925 -46.075 -38.595 ;
        RECT -46.405 -40.285 -46.075 -39.955 ;
        RECT -46.405 -41.645 -46.075 -41.315 ;
        RECT -46.405 -43.005 -46.075 -42.675 ;
        RECT -46.405 -44.365 -46.075 -44.035 ;
        RECT -46.405 -45.725 -46.075 -45.395 ;
        RECT -46.405 -47.085 -46.075 -46.755 ;
        RECT -46.405 -48.445 -46.075 -48.115 ;
        RECT -46.405 -49.805 -46.075 -49.475 ;
        RECT -46.405 -51.165 -46.075 -50.835 ;
        RECT -46.405 -52.525 -46.075 -52.195 ;
        RECT -46.405 -53.885 -46.075 -53.555 ;
        RECT -46.405 -55.245 -46.075 -54.915 ;
        RECT -46.405 -56.605 -46.075 -56.275 ;
        RECT -46.405 -57.965 -46.075 -57.635 ;
        RECT -46.405 -59.325 -46.075 -58.995 ;
        RECT -46.405 -60.685 -46.075 -60.355 ;
        RECT -46.405 -62.045 -46.075 -61.715 ;
        RECT -46.405 -63.405 -46.075 -63.075 ;
        RECT -46.405 -64.765 -46.075 -64.435 ;
        RECT -46.405 -65.91 -46.075 -65.58 ;
        RECT -46.405 -67.485 -46.075 -67.155 ;
        RECT -46.405 -68.845 -46.075 -68.515 ;
        RECT -46.405 -70.205 -46.075 -69.875 ;
        RECT -46.405 -71.565 -46.075 -71.235 ;
        RECT -46.405 -72.925 -46.075 -72.595 ;
        RECT -46.405 -75.645 -46.075 -75.315 ;
        RECT -46.405 -76.45 -46.075 -76.12 ;
        RECT -46.405 -78.365 -46.075 -78.035 ;
        RECT -46.405 -79.725 -46.075 -79.395 ;
        RECT -46.405 -81.085 -46.075 -80.755 ;
        RECT -46.405 -83.805 -46.075 -83.475 ;
        RECT -46.405 -85.165 -46.075 -84.835 ;
        RECT -46.4 -87.2 -46.08 12.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.045 44.8 -44.715 45.93 ;
        RECT -45.045 39.955 -44.715 40.285 ;
        RECT -45.045 38.595 -44.715 38.925 ;
        RECT -45.045 37.235 -44.715 37.565 ;
        RECT -45.045 35.875 -44.715 36.205 ;
        RECT -45.045 34.515 -44.715 34.845 ;
        RECT -45.045 33.155 -44.715 33.485 ;
        RECT -45.045 31.795 -44.715 32.125 ;
        RECT -45.045 30.435 -44.715 30.765 ;
        RECT -45.045 29.075 -44.715 29.405 ;
        RECT -45.045 27.715 -44.715 28.045 ;
        RECT -45.045 26.355 -44.715 26.685 ;
        RECT -45.045 24.995 -44.715 25.325 ;
        RECT -45.045 22.66 -44.715 22.99 ;
        RECT -45.045 20.485 -44.715 20.815 ;
        RECT -45.045 19.635 -44.715 19.965 ;
        RECT -45.04 19.56 -44.72 46.045 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.045 -94.685 -44.715 -94.355 ;
        RECT -45.045 -96.045 -44.715 -95.715 ;
        RECT -45.045 -97.405 -44.715 -97.075 ;
        RECT -45.045 -98.765 -44.715 -98.435 ;
        RECT -45.045 -100.125 -44.715 -99.795 ;
        RECT -45.045 -101.485 -44.715 -101.155 ;
        RECT -45.045 -102.845 -44.715 -102.515 ;
        RECT -45.045 -104.205 -44.715 -103.875 ;
        RECT -45.045 -105.565 -44.715 -105.235 ;
        RECT -45.045 -106.925 -44.715 -106.595 ;
        RECT -45.045 -108.285 -44.715 -107.955 ;
        RECT -45.045 -109.645 -44.715 -109.315 ;
        RECT -45.045 -111.005 -44.715 -110.675 ;
        RECT -45.045 -112.365 -44.715 -112.035 ;
        RECT -45.045 -113.725 -44.715 -113.395 ;
        RECT -45.045 -115.085 -44.715 -114.755 ;
        RECT -45.045 -116.445 -44.715 -116.115 ;
        RECT -45.045 -117.805 -44.715 -117.475 ;
        RECT -45.045 -119.165 -44.715 -118.835 ;
        RECT -45.045 -120.525 -44.715 -120.195 ;
        RECT -45.045 -121.885 -44.715 -121.555 ;
        RECT -45.045 -123.245 -44.715 -122.915 ;
        RECT -45.045 -124.605 -44.715 -124.275 ;
        RECT -45.045 -125.965 -44.715 -125.635 ;
        RECT -45.045 -127.325 -44.715 -126.995 ;
        RECT -45.045 -128.685 -44.715 -128.355 ;
        RECT -45.045 -130.045 -44.715 -129.715 ;
        RECT -45.045 -131.405 -44.715 -131.075 ;
        RECT -45.045 -132.765 -44.715 -132.435 ;
        RECT -45.045 -134.125 -44.715 -133.795 ;
        RECT -45.045 -135.485 -44.715 -135.155 ;
        RECT -45.045 -136.845 -44.715 -136.515 ;
        RECT -45.045 -138.205 -44.715 -137.875 ;
        RECT -45.045 -139.565 -44.715 -139.235 ;
        RECT -45.045 -140.925 -44.715 -140.595 ;
        RECT -45.045 -143.755 -44.715 -143.425 ;
        RECT -45.045 -145.005 -44.715 -144.675 ;
        RECT -45.045 -146.365 -44.715 -146.035 ;
        RECT -45.045 -149.085 -44.715 -148.755 ;
        RECT -45.045 -151.805 -44.715 -151.475 ;
        RECT -45.045 -153.165 -44.715 -152.835 ;
        RECT -45.045 -158.81 -44.715 -157.68 ;
        RECT -45.04 -158.925 -44.72 -94.355 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.685 -109.645 -43.355 -109.315 ;
        RECT -43.685 -111.005 -43.355 -110.675 ;
        RECT -43.685 -112.365 -43.355 -112.035 ;
        RECT -43.685 -113.725 -43.355 -113.395 ;
        RECT -43.685 -115.085 -43.355 -114.755 ;
        RECT -43.685 -116.445 -43.355 -116.115 ;
        RECT -43.685 -117.805 -43.355 -117.475 ;
        RECT -43.685 -119.165 -43.355 -118.835 ;
        RECT -43.685 -120.525 -43.355 -120.195 ;
        RECT -43.685 -121.885 -43.355 -121.555 ;
        RECT -43.685 -123.245 -43.355 -122.915 ;
        RECT -43.685 -124.605 -43.355 -124.275 ;
        RECT -43.685 -125.965 -43.355 -125.635 ;
        RECT -43.685 -127.325 -43.355 -126.995 ;
        RECT -43.685 -128.685 -43.355 -128.355 ;
        RECT -43.685 -130.045 -43.355 -129.715 ;
        RECT -43.685 -131.405 -43.355 -131.075 ;
        RECT -43.685 -132.765 -43.355 -132.435 ;
        RECT -43.685 -134.125 -43.355 -133.795 ;
        RECT -43.685 -135.485 -43.355 -135.155 ;
        RECT -43.685 -136.845 -43.355 -136.515 ;
        RECT -43.685 -138.205 -43.355 -137.875 ;
        RECT -43.685 -139.565 -43.355 -139.235 ;
        RECT -43.685 -140.925 -43.355 -140.595 ;
        RECT -43.685 -143.755 -43.355 -143.425 ;
        RECT -43.685 -145.005 -43.355 -144.675 ;
        RECT -43.685 -146.365 -43.355 -146.035 ;
        RECT -43.685 -147.725 -43.355 -147.395 ;
        RECT -43.685 -149.085 -43.355 -148.755 ;
        RECT -43.685 -151.805 -43.355 -151.475 ;
        RECT -43.685 -153.165 -43.355 -152.835 ;
        RECT -43.685 -158.81 -43.355 -157.68 ;
        RECT -43.68 -158.925 -43.36 46.045 ;
        RECT -43.685 44.8 -43.355 45.93 ;
        RECT -43.685 39.955 -43.355 40.285 ;
        RECT -43.685 38.595 -43.355 38.925 ;
        RECT -43.685 37.235 -43.355 37.565 ;
        RECT -43.685 35.875 -43.355 36.205 ;
        RECT -43.685 34.515 -43.355 34.845 ;
        RECT -43.685 33.155 -43.355 33.485 ;
        RECT -43.685 31.795 -43.355 32.125 ;
        RECT -43.685 30.435 -43.355 30.765 ;
        RECT -43.685 29.075 -43.355 29.405 ;
        RECT -43.685 27.715 -43.355 28.045 ;
        RECT -43.685 26.355 -43.355 26.685 ;
        RECT -43.685 24.995 -43.355 25.325 ;
        RECT -43.685 22.66 -43.355 22.99 ;
        RECT -43.685 20.485 -43.355 20.815 ;
        RECT -43.685 19.635 -43.355 19.965 ;
        RECT -43.685 17.325 -43.355 17.655 ;
        RECT -43.685 16.475 -43.355 16.805 ;
        RECT -43.685 14.3 -43.355 14.63 ;
        RECT -43.685 11.395 -43.355 11.725 ;
        RECT -43.685 10.035 -43.355 10.365 ;
        RECT -43.685 8.675 -43.355 9.005 ;
        RECT -43.685 7.315 -43.355 7.645 ;
        RECT -43.685 5.955 -43.355 6.285 ;
        RECT -43.685 4.595 -43.355 4.925 ;
        RECT -43.685 3.235 -43.355 3.565 ;
        RECT -43.685 1.875 -43.355 2.205 ;
        RECT -43.685 0.515 -43.355 0.845 ;
        RECT -43.685 -0.845 -43.355 -0.515 ;
        RECT -43.685 -2.205 -43.355 -1.875 ;
        RECT -43.685 -3.565 -43.355 -3.235 ;
        RECT -43.685 -4.925 -43.355 -4.595 ;
        RECT -43.685 -6.285 -43.355 -5.955 ;
        RECT -43.685 -7.645 -43.355 -7.315 ;
        RECT -43.685 -10.365 -43.355 -10.035 ;
        RECT -43.685 -11.725 -43.355 -11.395 ;
        RECT -43.685 -13.085 -43.355 -12.755 ;
        RECT -43.685 -14.445 -43.355 -14.115 ;
        RECT -43.685 -15.805 -43.355 -15.475 ;
        RECT -43.685 -17.165 -43.355 -16.835 ;
        RECT -43.685 -18.525 -43.355 -18.195 ;
        RECT -43.685 -21.245 -43.355 -20.915 ;
        RECT -43.685 -22.605 -43.355 -22.275 ;
        RECT -43.685 -23.965 -43.355 -23.635 ;
        RECT -43.685 -25.325 -43.355 -24.995 ;
        RECT -43.685 -26.685 -43.355 -26.355 ;
        RECT -43.685 -28.045 -43.355 -27.715 ;
        RECT -43.685 -29.405 -43.355 -29.075 ;
        RECT -43.685 -30.765 -43.355 -30.435 ;
        RECT -43.685 -32.125 -43.355 -31.795 ;
        RECT -43.685 -33.485 -43.355 -33.155 ;
        RECT -43.685 -34.845 -43.355 -34.515 ;
        RECT -43.685 -36.205 -43.355 -35.875 ;
        RECT -43.685 -37.565 -43.355 -37.235 ;
        RECT -43.685 -38.925 -43.355 -38.595 ;
        RECT -43.685 -40.285 -43.355 -39.955 ;
        RECT -43.685 -41.645 -43.355 -41.315 ;
        RECT -43.685 -43.005 -43.355 -42.675 ;
        RECT -43.685 -44.365 -43.355 -44.035 ;
        RECT -43.685 -45.725 -43.355 -45.395 ;
        RECT -43.685 -47.085 -43.355 -46.755 ;
        RECT -43.685 -48.445 -43.355 -48.115 ;
        RECT -43.685 -49.805 -43.355 -49.475 ;
        RECT -43.685 -51.165 -43.355 -50.835 ;
        RECT -43.685 -52.525 -43.355 -52.195 ;
        RECT -43.685 -53.885 -43.355 -53.555 ;
        RECT -43.685 -55.245 -43.355 -54.915 ;
        RECT -43.685 -56.605 -43.355 -56.275 ;
        RECT -43.685 -57.965 -43.355 -57.635 ;
        RECT -43.685 -59.325 -43.355 -58.995 ;
        RECT -43.685 -60.685 -43.355 -60.355 ;
        RECT -43.685 -62.045 -43.355 -61.715 ;
        RECT -43.685 -63.405 -43.355 -63.075 ;
        RECT -43.685 -64.765 -43.355 -64.435 ;
        RECT -43.685 -65.91 -43.355 -65.58 ;
        RECT -43.685 -67.485 -43.355 -67.155 ;
        RECT -43.685 -68.845 -43.355 -68.515 ;
        RECT -43.685 -70.205 -43.355 -69.875 ;
        RECT -43.685 -71.565 -43.355 -71.235 ;
        RECT -43.685 -72.925 -43.355 -72.595 ;
        RECT -43.685 -75.645 -43.355 -75.315 ;
        RECT -43.685 -76.45 -43.355 -76.12 ;
        RECT -43.685 -78.365 -43.355 -78.035 ;
        RECT -43.685 -79.725 -43.355 -79.395 ;
        RECT -43.685 -81.085 -43.355 -80.755 ;
        RECT -43.685 -83.805 -43.355 -83.475 ;
        RECT -43.685 -85.165 -43.355 -84.835 ;
        RECT -43.685 -87.885 -43.355 -87.555 ;
        RECT -43.685 -89.245 -43.355 -88.915 ;
        RECT -43.685 -90.605 -43.355 -90.275 ;
        RECT -43.685 -91.965 -43.355 -91.635 ;
        RECT -43.685 -93.325 -43.355 -92.995 ;
        RECT -43.685 -94.685 -43.355 -94.355 ;
        RECT -43.685 -96.045 -43.355 -95.715 ;
        RECT -43.685 -97.405 -43.355 -97.075 ;
        RECT -43.685 -98.765 -43.355 -98.435 ;
        RECT -43.685 -100.125 -43.355 -99.795 ;
        RECT -43.685 -101.485 -43.355 -101.155 ;
        RECT -43.685 -102.845 -43.355 -102.515 ;
        RECT -43.685 -104.205 -43.355 -103.875 ;
        RECT -43.685 -105.565 -43.355 -105.235 ;
        RECT -43.685 -106.925 -43.355 -106.595 ;
        RECT -43.685 -108.285 -43.355 -107.955 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.925 5.955 -55.595 6.285 ;
        RECT -55.925 4.595 -55.595 4.925 ;
        RECT -55.925 3.235 -55.595 3.565 ;
        RECT -55.925 1.875 -55.595 2.205 ;
        RECT -55.925 0.515 -55.595 0.845 ;
        RECT -55.925 -0.845 -55.595 -0.515 ;
        RECT -55.925 -2.205 -55.595 -1.875 ;
        RECT -55.925 -3.565 -55.595 -3.235 ;
        RECT -55.925 -4.925 -55.595 -4.595 ;
        RECT -55.925 -6.285 -55.595 -5.955 ;
        RECT -55.925 -7.645 -55.595 -7.315 ;
        RECT -55.925 -9.005 -55.595 -8.675 ;
        RECT -55.925 -10.365 -55.595 -10.035 ;
        RECT -55.925 -11.725 -55.595 -11.395 ;
        RECT -55.925 -13.085 -55.595 -12.755 ;
        RECT -55.925 -14.445 -55.595 -14.115 ;
        RECT -55.925 -15.805 -55.595 -15.475 ;
        RECT -55.925 -17.165 -55.595 -16.835 ;
        RECT -55.925 -18.525 -55.595 -18.195 ;
        RECT -55.925 -19.885 -55.595 -19.555 ;
        RECT -55.925 -21.245 -55.595 -20.915 ;
        RECT -55.925 -22.605 -55.595 -22.275 ;
        RECT -55.925 -23.965 -55.595 -23.635 ;
        RECT -55.925 -25.325 -55.595 -24.995 ;
        RECT -55.925 -26.685 -55.595 -26.355 ;
        RECT -55.925 -28.045 -55.595 -27.715 ;
        RECT -55.925 -29.405 -55.595 -29.075 ;
        RECT -55.925 -30.765 -55.595 -30.435 ;
        RECT -55.925 -32.125 -55.595 -31.795 ;
        RECT -55.925 -33.485 -55.595 -33.155 ;
        RECT -55.925 -34.845 -55.595 -34.515 ;
        RECT -55.925 -36.205 -55.595 -35.875 ;
        RECT -55.925 -37.565 -55.595 -37.235 ;
        RECT -55.925 -38.925 -55.595 -38.595 ;
        RECT -55.925 -40.285 -55.595 -39.955 ;
        RECT -55.925 -41.645 -55.595 -41.315 ;
        RECT -55.925 -43.005 -55.595 -42.675 ;
        RECT -55.925 -44.365 -55.595 -44.035 ;
        RECT -55.925 -45.725 -55.595 -45.395 ;
        RECT -55.925 -47.085 -55.595 -46.755 ;
        RECT -55.925 -48.445 -55.595 -48.115 ;
        RECT -55.925 -49.805 -55.595 -49.475 ;
        RECT -55.925 -51.165 -55.595 -50.835 ;
        RECT -55.925 -52.525 -55.595 -52.195 ;
        RECT -55.925 -53.885 -55.595 -53.555 ;
        RECT -55.925 -55.245 -55.595 -54.915 ;
        RECT -55.925 -56.605 -55.595 -56.275 ;
        RECT -55.925 -57.965 -55.595 -57.635 ;
        RECT -55.925 -59.325 -55.595 -58.995 ;
        RECT -55.925 -60.685 -55.595 -60.355 ;
        RECT -55.925 -62.045 -55.595 -61.715 ;
        RECT -55.925 -63.405 -55.595 -63.075 ;
        RECT -55.925 -64.765 -55.595 -64.435 ;
        RECT -55.925 -66.125 -55.595 -65.795 ;
        RECT -55.925 -67.485 -55.595 -67.155 ;
        RECT -55.925 -68.845 -55.595 -68.515 ;
        RECT -55.925 -70.205 -55.595 -69.875 ;
        RECT -55.925 -71.565 -55.595 -71.235 ;
        RECT -55.925 -72.925 -55.595 -72.595 ;
        RECT -55.925 -74.285 -55.595 -73.955 ;
        RECT -55.925 -75.645 -55.595 -75.315 ;
        RECT -55.925 -77.005 -55.595 -76.675 ;
        RECT -55.925 -78.365 -55.595 -78.035 ;
        RECT -55.925 -79.725 -55.595 -79.395 ;
        RECT -55.925 -81.085 -55.595 -80.755 ;
        RECT -55.925 -82.445 -55.595 -82.115 ;
        RECT -55.925 -83.805 -55.595 -83.475 ;
        RECT -55.925 -85.165 -55.595 -84.835 ;
        RECT -55.925 -86.525 -55.595 -86.195 ;
        RECT -55.925 -87.885 -55.595 -87.555 ;
        RECT -55.925 -89.245 -55.595 -88.915 ;
        RECT -55.925 -90.605 -55.595 -90.275 ;
        RECT -55.925 -91.965 -55.595 -91.635 ;
        RECT -55.925 -93.325 -55.595 -92.995 ;
        RECT -55.925 -94.685 -55.595 -94.355 ;
        RECT -55.925 -96.045 -55.595 -95.715 ;
        RECT -55.925 -97.405 -55.595 -97.075 ;
        RECT -55.925 -98.765 -55.595 -98.435 ;
        RECT -55.925 -100.125 -55.595 -99.795 ;
        RECT -55.925 -101.485 -55.595 -101.155 ;
        RECT -55.925 -102.845 -55.595 -102.515 ;
        RECT -55.925 -104.205 -55.595 -103.875 ;
        RECT -55.925 -105.565 -55.595 -105.235 ;
        RECT -55.925 -106.925 -55.595 -106.595 ;
        RECT -55.925 -108.285 -55.595 -107.955 ;
        RECT -55.925 -109.645 -55.595 -109.315 ;
        RECT -55.925 -111.005 -55.595 -110.675 ;
        RECT -55.925 -112.365 -55.595 -112.035 ;
        RECT -55.925 -113.725 -55.595 -113.395 ;
        RECT -55.925 -115.085 -55.595 -114.755 ;
        RECT -55.925 -116.445 -55.595 -116.115 ;
        RECT -55.925 -117.805 -55.595 -117.475 ;
        RECT -55.925 -119.165 -55.595 -118.835 ;
        RECT -55.925 -120.525 -55.595 -120.195 ;
        RECT -55.925 -121.885 -55.595 -121.555 ;
        RECT -55.925 -123.245 -55.595 -122.915 ;
        RECT -55.925 -124.605 -55.595 -124.275 ;
        RECT -55.925 -125.965 -55.595 -125.635 ;
        RECT -55.925 -127.325 -55.595 -126.995 ;
        RECT -55.925 -128.685 -55.595 -128.355 ;
        RECT -55.925 -130.045 -55.595 -129.715 ;
        RECT -55.925 -131.405 -55.595 -131.075 ;
        RECT -55.925 -132.765 -55.595 -132.435 ;
        RECT -55.925 -134.125 -55.595 -133.795 ;
        RECT -55.925 -135.485 -55.595 -135.155 ;
        RECT -55.925 -136.845 -55.595 -136.515 ;
        RECT -55.925 -138.205 -55.595 -137.875 ;
        RECT -55.925 -139.565 -55.595 -139.235 ;
        RECT -55.925 -140.925 -55.595 -140.595 ;
        RECT -55.925 -142.285 -55.595 -141.955 ;
        RECT -55.925 -143.645 -55.595 -143.315 ;
        RECT -55.925 -145.005 -55.595 -144.675 ;
        RECT -55.925 -146.365 -55.595 -146.035 ;
        RECT -55.925 -147.725 -55.595 -147.395 ;
        RECT -55.925 -149.085 -55.595 -148.755 ;
        RECT -55.925 -150.445 -55.595 -150.115 ;
        RECT -55.925 -151.805 -55.595 -151.475 ;
        RECT -55.925 -153.165 -55.595 -152.835 ;
        RECT -55.925 -158.81 -55.595 -157.68 ;
        RECT -55.92 -158.925 -55.6 46.045 ;
        RECT -55.925 44.8 -55.595 45.93 ;
        RECT -55.925 39.955 -55.595 40.285 ;
        RECT -55.925 38.595 -55.595 38.925 ;
        RECT -55.925 37.235 -55.595 37.565 ;
        RECT -55.925 35.875 -55.595 36.205 ;
        RECT -55.925 34.515 -55.595 34.845 ;
        RECT -55.925 33.155 -55.595 33.485 ;
        RECT -55.925 31.795 -55.595 32.125 ;
        RECT -55.925 30.435 -55.595 30.765 ;
        RECT -55.925 29.075 -55.595 29.405 ;
        RECT -55.925 27.715 -55.595 28.045 ;
        RECT -55.925 26.355 -55.595 26.685 ;
        RECT -55.925 24.995 -55.595 25.325 ;
        RECT -55.925 22.66 -55.595 22.99 ;
        RECT -55.925 20.485 -55.595 20.815 ;
        RECT -55.925 19.635 -55.595 19.965 ;
        RECT -55.925 17.325 -55.595 17.655 ;
        RECT -55.925 16.475 -55.595 16.805 ;
        RECT -55.925 14.3 -55.595 14.63 ;
        RECT -55.925 11.395 -55.595 11.725 ;
        RECT -55.925 10.035 -55.595 10.365 ;
        RECT -55.925 8.675 -55.595 9.005 ;
        RECT -55.925 7.315 -55.595 7.645 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 15.51 -94.075 15.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 42.08 17.165 43.21 ;
        RECT 16.835 40.635 17.165 40.965 ;
        RECT 16.835 39.275 17.165 39.605 ;
        RECT 16.835 37.915 17.165 38.245 ;
        RECT 16.84 37.915 17.16 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 -1.525 17.165 -1.195 ;
        RECT 16.835 -2.885 17.165 -2.555 ;
        RECT 16.84 -3.56 17.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 42.08 18.525 43.21 ;
        RECT 18.195 40.635 18.525 40.965 ;
        RECT 18.195 39.275 18.525 39.605 ;
        RECT 18.195 37.915 18.525 38.245 ;
        RECT 18.2 37.915 18.52 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 -1.525 18.525 -1.195 ;
        RECT 18.195 -2.885 18.525 -2.555 ;
        RECT 18.2 -3.56 18.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 42.08 19.885 43.21 ;
        RECT 19.555 40.635 19.885 40.965 ;
        RECT 19.555 39.275 19.885 39.605 ;
        RECT 19.555 37.915 19.885 38.245 ;
        RECT 19.56 37.915 19.88 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 -1.525 19.885 -1.195 ;
        RECT 19.555 -2.885 19.885 -2.555 ;
        RECT 19.56 -3.56 19.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 -91.285 19.885 -90.955 ;
        RECT 19.555 -92.645 19.885 -92.315 ;
        RECT 19.555 -94.005 19.885 -93.675 ;
        RECT 19.555 -95.365 19.885 -95.035 ;
        RECT 19.555 -96.725 19.885 -96.395 ;
        RECT 19.555 -98.085 19.885 -97.755 ;
        RECT 19.555 -99.445 19.885 -99.115 ;
        RECT 19.555 -100.805 19.885 -100.475 ;
        RECT 19.555 -102.165 19.885 -101.835 ;
        RECT 19.555 -103.525 19.885 -103.195 ;
        RECT 19.555 -104.885 19.885 -104.555 ;
        RECT 19.555 -106.245 19.885 -105.915 ;
        RECT 19.555 -107.605 19.885 -107.275 ;
        RECT 19.555 -108.965 19.885 -108.635 ;
        RECT 19.555 -110.325 19.885 -109.995 ;
        RECT 19.555 -111.685 19.885 -111.355 ;
        RECT 19.555 -113.045 19.885 -112.715 ;
        RECT 19.555 -114.405 19.885 -114.075 ;
        RECT 19.555 -115.765 19.885 -115.435 ;
        RECT 19.555 -117.125 19.885 -116.795 ;
        RECT 19.555 -118.485 19.885 -118.155 ;
        RECT 19.555 -119.845 19.885 -119.515 ;
        RECT 19.555 -121.205 19.885 -120.875 ;
        RECT 19.555 -122.565 19.885 -122.235 ;
        RECT 19.555 -123.925 19.885 -123.595 ;
        RECT 19.555 -125.285 19.885 -124.955 ;
        RECT 19.555 -126.645 19.885 -126.315 ;
        RECT 19.555 -128.005 19.885 -127.675 ;
        RECT 19.555 -129.365 19.885 -129.035 ;
        RECT 19.555 -130.725 19.885 -130.395 ;
        RECT 19.555 -132.085 19.885 -131.755 ;
        RECT 19.555 -133.445 19.885 -133.115 ;
        RECT 19.555 -134.805 19.885 -134.475 ;
        RECT 19.555 -136.165 19.885 -135.835 ;
        RECT 19.555 -137.525 19.885 -137.195 ;
        RECT 19.555 -138.885 19.885 -138.555 ;
        RECT 19.555 -140.245 19.885 -139.915 ;
        RECT 19.555 -141.605 19.885 -141.275 ;
        RECT 19.555 -142.965 19.885 -142.635 ;
        RECT 19.555 -144.325 19.885 -143.995 ;
        RECT 19.555 -145.685 19.885 -145.355 ;
        RECT 19.555 -147.045 19.885 -146.715 ;
        RECT 19.555 -148.405 19.885 -148.075 ;
        RECT 19.555 -149.765 19.885 -149.435 ;
        RECT 19.555 -151.125 19.885 -150.795 ;
        RECT 19.555 -152.485 19.885 -152.155 ;
        RECT 19.555 -153.845 19.885 -153.515 ;
        RECT 19.555 -156.09 19.885 -154.96 ;
        RECT 19.56 -156.205 19.88 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 42.08 21.245 43.21 ;
        RECT 20.915 40.635 21.245 40.965 ;
        RECT 20.915 39.275 21.245 39.605 ;
        RECT 20.915 37.915 21.245 38.245 ;
        RECT 20.92 37.915 21.24 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 -95.365 21.245 -95.035 ;
        RECT 20.915 -96.725 21.245 -96.395 ;
        RECT 20.915 -98.085 21.245 -97.755 ;
        RECT 20.915 -99.445 21.245 -99.115 ;
        RECT 20.915 -100.805 21.245 -100.475 ;
        RECT 20.915 -102.165 21.245 -101.835 ;
        RECT 20.915 -103.525 21.245 -103.195 ;
        RECT 20.915 -104.885 21.245 -104.555 ;
        RECT 20.915 -106.245 21.245 -105.915 ;
        RECT 20.915 -107.605 21.245 -107.275 ;
        RECT 20.915 -108.965 21.245 -108.635 ;
        RECT 20.915 -110.325 21.245 -109.995 ;
        RECT 20.915 -111.685 21.245 -111.355 ;
        RECT 20.915 -113.045 21.245 -112.715 ;
        RECT 20.915 -114.405 21.245 -114.075 ;
        RECT 20.915 -115.765 21.245 -115.435 ;
        RECT 20.915 -117.125 21.245 -116.795 ;
        RECT 20.915 -118.485 21.245 -118.155 ;
        RECT 20.915 -119.845 21.245 -119.515 ;
        RECT 20.915 -121.205 21.245 -120.875 ;
        RECT 20.915 -122.565 21.245 -122.235 ;
        RECT 20.915 -123.925 21.245 -123.595 ;
        RECT 20.915 -125.285 21.245 -124.955 ;
        RECT 20.915 -126.645 21.245 -126.315 ;
        RECT 20.915 -128.005 21.245 -127.675 ;
        RECT 20.915 -129.365 21.245 -129.035 ;
        RECT 20.915 -130.725 21.245 -130.395 ;
        RECT 20.915 -132.085 21.245 -131.755 ;
        RECT 20.915 -133.445 21.245 -133.115 ;
        RECT 20.915 -134.805 21.245 -134.475 ;
        RECT 20.915 -136.165 21.245 -135.835 ;
        RECT 20.915 -137.525 21.245 -137.195 ;
        RECT 20.915 -138.885 21.245 -138.555 ;
        RECT 20.915 -140.245 21.245 -139.915 ;
        RECT 20.915 -141.605 21.245 -141.275 ;
        RECT 20.915 -142.965 21.245 -142.635 ;
        RECT 20.915 -144.325 21.245 -143.995 ;
        RECT 20.915 -145.685 21.245 -145.355 ;
        RECT 20.915 -147.045 21.245 -146.715 ;
        RECT 20.915 -148.405 21.245 -148.075 ;
        RECT 20.915 -149.765 21.245 -149.435 ;
        RECT 20.915 -151.125 21.245 -150.795 ;
        RECT 20.915 -152.485 21.245 -152.155 ;
        RECT 20.915 -153.845 21.245 -153.515 ;
        RECT 20.915 -156.09 21.245 -154.96 ;
        RECT 20.92 -156.205 21.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.61 -94.075 21.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 42.08 22.605 43.21 ;
        RECT 22.275 40.635 22.605 40.965 ;
        RECT 22.275 39.275 22.605 39.605 ;
        RECT 22.275 37.915 22.605 38.245 ;
        RECT 22.28 37.915 22.6 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 42.08 23.965 43.21 ;
        RECT 23.635 40.635 23.965 40.965 ;
        RECT 23.635 39.275 23.965 39.605 ;
        RECT 23.635 37.915 23.965 38.245 ;
        RECT 23.64 37.915 23.96 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 -1.525 23.965 -1.195 ;
        RECT 23.635 -2.885 23.965 -2.555 ;
        RECT 23.64 -3.56 23.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 42.08 25.325 43.21 ;
        RECT 24.995 40.635 25.325 40.965 ;
        RECT 24.995 39.275 25.325 39.605 ;
        RECT 24.995 37.915 25.325 38.245 ;
        RECT 25 37.915 25.32 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 -1.525 25.325 -1.195 ;
        RECT 24.995 -2.885 25.325 -2.555 ;
        RECT 25 -3.56 25.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 -91.285 25.325 -90.955 ;
        RECT 24.995 -92.645 25.325 -92.315 ;
        RECT 24.995 -94.005 25.325 -93.675 ;
        RECT 24.995 -95.365 25.325 -95.035 ;
        RECT 24.995 -96.725 25.325 -96.395 ;
        RECT 24.995 -98.085 25.325 -97.755 ;
        RECT 24.995 -99.445 25.325 -99.115 ;
        RECT 24.995 -100.805 25.325 -100.475 ;
        RECT 24.995 -102.165 25.325 -101.835 ;
        RECT 24.995 -103.525 25.325 -103.195 ;
        RECT 24.995 -104.885 25.325 -104.555 ;
        RECT 24.995 -106.245 25.325 -105.915 ;
        RECT 24.995 -107.605 25.325 -107.275 ;
        RECT 24.995 -108.965 25.325 -108.635 ;
        RECT 24.995 -110.325 25.325 -109.995 ;
        RECT 24.995 -111.685 25.325 -111.355 ;
        RECT 24.995 -113.045 25.325 -112.715 ;
        RECT 24.995 -114.405 25.325 -114.075 ;
        RECT 24.995 -115.765 25.325 -115.435 ;
        RECT 24.995 -117.125 25.325 -116.795 ;
        RECT 24.995 -118.485 25.325 -118.155 ;
        RECT 24.995 -119.845 25.325 -119.515 ;
        RECT 24.995 -121.205 25.325 -120.875 ;
        RECT 24.995 -122.565 25.325 -122.235 ;
        RECT 24.995 -123.925 25.325 -123.595 ;
        RECT 24.995 -125.285 25.325 -124.955 ;
        RECT 24.995 -126.645 25.325 -126.315 ;
        RECT 24.995 -128.005 25.325 -127.675 ;
        RECT 24.995 -129.365 25.325 -129.035 ;
        RECT 24.995 -130.725 25.325 -130.395 ;
        RECT 24.995 -132.085 25.325 -131.755 ;
        RECT 24.995 -133.445 25.325 -133.115 ;
        RECT 24.995 -134.805 25.325 -134.475 ;
        RECT 24.995 -136.165 25.325 -135.835 ;
        RECT 24.995 -137.525 25.325 -137.195 ;
        RECT 24.995 -138.885 25.325 -138.555 ;
        RECT 24.995 -140.245 25.325 -139.915 ;
        RECT 24.995 -141.605 25.325 -141.275 ;
        RECT 24.995 -142.965 25.325 -142.635 ;
        RECT 24.995 -144.325 25.325 -143.995 ;
        RECT 24.995 -145.685 25.325 -145.355 ;
        RECT 24.995 -147.045 25.325 -146.715 ;
        RECT 24.995 -148.405 25.325 -148.075 ;
        RECT 24.995 -149.765 25.325 -149.435 ;
        RECT 24.995 -151.125 25.325 -150.795 ;
        RECT 24.995 -152.485 25.325 -152.155 ;
        RECT 24.995 -153.845 25.325 -153.515 ;
        RECT 24.995 -156.09 25.325 -154.96 ;
        RECT 25 -156.205 25.32 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 42.08 26.685 43.21 ;
        RECT 26.355 40.635 26.685 40.965 ;
        RECT 26.355 39.275 26.685 39.605 ;
        RECT 26.355 37.915 26.685 38.245 ;
        RECT 26.36 37.915 26.68 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 -1.525 26.685 -1.195 ;
        RECT 26.355 -2.885 26.685 -2.555 ;
        RECT 26.36 -3.56 26.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 -91.285 26.685 -90.955 ;
        RECT 26.355 -92.645 26.685 -92.315 ;
        RECT 26.355 -94.005 26.685 -93.675 ;
        RECT 26.355 -95.365 26.685 -95.035 ;
        RECT 26.355 -96.725 26.685 -96.395 ;
        RECT 26.355 -98.085 26.685 -97.755 ;
        RECT 26.355 -99.445 26.685 -99.115 ;
        RECT 26.355 -100.805 26.685 -100.475 ;
        RECT 26.355 -102.165 26.685 -101.835 ;
        RECT 26.355 -103.525 26.685 -103.195 ;
        RECT 26.355 -104.885 26.685 -104.555 ;
        RECT 26.355 -106.245 26.685 -105.915 ;
        RECT 26.355 -107.605 26.685 -107.275 ;
        RECT 26.355 -108.965 26.685 -108.635 ;
        RECT 26.355 -110.325 26.685 -109.995 ;
        RECT 26.355 -111.685 26.685 -111.355 ;
        RECT 26.355 -113.045 26.685 -112.715 ;
        RECT 26.355 -114.405 26.685 -114.075 ;
        RECT 26.355 -115.765 26.685 -115.435 ;
        RECT 26.355 -117.125 26.685 -116.795 ;
        RECT 26.355 -118.485 26.685 -118.155 ;
        RECT 26.355 -119.845 26.685 -119.515 ;
        RECT 26.355 -121.205 26.685 -120.875 ;
        RECT 26.355 -122.565 26.685 -122.235 ;
        RECT 26.355 -123.925 26.685 -123.595 ;
        RECT 26.355 -125.285 26.685 -124.955 ;
        RECT 26.355 -126.645 26.685 -126.315 ;
        RECT 26.355 -128.005 26.685 -127.675 ;
        RECT 26.355 -129.365 26.685 -129.035 ;
        RECT 26.355 -130.725 26.685 -130.395 ;
        RECT 26.355 -132.085 26.685 -131.755 ;
        RECT 26.355 -133.445 26.685 -133.115 ;
        RECT 26.355 -134.805 26.685 -134.475 ;
        RECT 26.355 -136.165 26.685 -135.835 ;
        RECT 26.355 -137.525 26.685 -137.195 ;
        RECT 26.355 -138.885 26.685 -138.555 ;
        RECT 26.355 -140.245 26.685 -139.915 ;
        RECT 26.355 -141.605 26.685 -141.275 ;
        RECT 26.355 -142.965 26.685 -142.635 ;
        RECT 26.355 -144.325 26.685 -143.995 ;
        RECT 26.355 -145.685 26.685 -145.355 ;
        RECT 26.355 -147.045 26.685 -146.715 ;
        RECT 26.355 -148.405 26.685 -148.075 ;
        RECT 26.355 -149.765 26.685 -149.435 ;
        RECT 26.355 -151.125 26.685 -150.795 ;
        RECT 26.355 -152.485 26.685 -152.155 ;
        RECT 26.355 -153.845 26.685 -153.515 ;
        RECT 26.355 -156.09 26.685 -154.96 ;
        RECT 26.36 -156.205 26.68 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.06 -94.075 27.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 42.08 28.045 43.21 ;
        RECT 27.715 40.635 28.045 40.965 ;
        RECT 27.715 39.275 28.045 39.605 ;
        RECT 27.715 37.915 28.045 38.245 ;
        RECT 27.72 37.915 28.04 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 -95.365 28.045 -95.035 ;
        RECT 27.715 -96.725 28.045 -96.395 ;
        RECT 27.715 -98.085 28.045 -97.755 ;
        RECT 27.715 -99.445 28.045 -99.115 ;
        RECT 27.715 -100.805 28.045 -100.475 ;
        RECT 27.715 -102.165 28.045 -101.835 ;
        RECT 27.715 -103.525 28.045 -103.195 ;
        RECT 27.715 -104.885 28.045 -104.555 ;
        RECT 27.715 -106.245 28.045 -105.915 ;
        RECT 27.715 -107.605 28.045 -107.275 ;
        RECT 27.715 -108.965 28.045 -108.635 ;
        RECT 27.715 -110.325 28.045 -109.995 ;
        RECT 27.715 -111.685 28.045 -111.355 ;
        RECT 27.715 -113.045 28.045 -112.715 ;
        RECT 27.715 -114.405 28.045 -114.075 ;
        RECT 27.715 -115.765 28.045 -115.435 ;
        RECT 27.715 -117.125 28.045 -116.795 ;
        RECT 27.715 -118.485 28.045 -118.155 ;
        RECT 27.715 -119.845 28.045 -119.515 ;
        RECT 27.715 -121.205 28.045 -120.875 ;
        RECT 27.715 -122.565 28.045 -122.235 ;
        RECT 27.715 -123.925 28.045 -123.595 ;
        RECT 27.715 -125.285 28.045 -124.955 ;
        RECT 27.715 -126.645 28.045 -126.315 ;
        RECT 27.715 -128.005 28.045 -127.675 ;
        RECT 27.715 -129.365 28.045 -129.035 ;
        RECT 27.715 -130.725 28.045 -130.395 ;
        RECT 27.715 -132.085 28.045 -131.755 ;
        RECT 27.715 -133.445 28.045 -133.115 ;
        RECT 27.715 -134.805 28.045 -134.475 ;
        RECT 27.715 -136.165 28.045 -135.835 ;
        RECT 27.715 -137.525 28.045 -137.195 ;
        RECT 27.715 -138.885 28.045 -138.555 ;
        RECT 27.715 -140.245 28.045 -139.915 ;
        RECT 27.715 -141.605 28.045 -141.275 ;
        RECT 27.715 -142.965 28.045 -142.635 ;
        RECT 27.715 -144.325 28.045 -143.995 ;
        RECT 27.715 -145.685 28.045 -145.355 ;
        RECT 27.715 -147.045 28.045 -146.715 ;
        RECT 27.715 -148.405 28.045 -148.075 ;
        RECT 27.715 -149.765 28.045 -149.435 ;
        RECT 27.715 -151.125 28.045 -150.795 ;
        RECT 27.715 -152.485 28.045 -152.155 ;
        RECT 27.715 -153.845 28.045 -153.515 ;
        RECT 27.715 -156.09 28.045 -154.96 ;
        RECT 27.72 -156.205 28.04 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 42.08 29.405 43.21 ;
        RECT 29.075 40.635 29.405 40.965 ;
        RECT 29.075 39.275 29.405 39.605 ;
        RECT 29.075 37.915 29.405 38.245 ;
        RECT 29.08 37.915 29.4 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 -1.525 29.405 -1.195 ;
        RECT 29.075 -2.885 29.405 -2.555 ;
        RECT 29.08 -3.56 29.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 -91.285 29.405 -90.955 ;
        RECT 29.075 -92.645 29.405 -92.315 ;
        RECT 29.075 -94.005 29.405 -93.675 ;
        RECT 29.075 -95.365 29.405 -95.035 ;
        RECT 29.075 -96.725 29.405 -96.395 ;
        RECT 29.075 -98.085 29.405 -97.755 ;
        RECT 29.075 -99.445 29.405 -99.115 ;
        RECT 29.075 -100.805 29.405 -100.475 ;
        RECT 29.075 -102.165 29.405 -101.835 ;
        RECT 29.075 -103.525 29.405 -103.195 ;
        RECT 29.075 -104.885 29.405 -104.555 ;
        RECT 29.075 -106.245 29.405 -105.915 ;
        RECT 29.075 -107.605 29.405 -107.275 ;
        RECT 29.075 -108.965 29.405 -108.635 ;
        RECT 29.075 -110.325 29.405 -109.995 ;
        RECT 29.075 -111.685 29.405 -111.355 ;
        RECT 29.075 -113.045 29.405 -112.715 ;
        RECT 29.075 -114.405 29.405 -114.075 ;
        RECT 29.075 -115.765 29.405 -115.435 ;
        RECT 29.075 -117.125 29.405 -116.795 ;
        RECT 29.075 -118.485 29.405 -118.155 ;
        RECT 29.075 -119.845 29.405 -119.515 ;
        RECT 29.075 -121.205 29.405 -120.875 ;
        RECT 29.075 -122.565 29.405 -122.235 ;
        RECT 29.075 -123.925 29.405 -123.595 ;
        RECT 29.075 -125.285 29.405 -124.955 ;
        RECT 29.075 -126.645 29.405 -126.315 ;
        RECT 29.075 -128.005 29.405 -127.675 ;
        RECT 29.075 -129.365 29.405 -129.035 ;
        RECT 29.075 -130.725 29.405 -130.395 ;
        RECT 29.075 -132.085 29.405 -131.755 ;
        RECT 29.075 -133.445 29.405 -133.115 ;
        RECT 29.075 -134.805 29.405 -134.475 ;
        RECT 29.075 -136.165 29.405 -135.835 ;
        RECT 29.075 -137.525 29.405 -137.195 ;
        RECT 29.075 -138.885 29.405 -138.555 ;
        RECT 29.075 -140.245 29.405 -139.915 ;
        RECT 29.075 -141.605 29.405 -141.275 ;
        RECT 29.075 -142.965 29.405 -142.635 ;
        RECT 29.075 -144.325 29.405 -143.995 ;
        RECT 29.075 -145.685 29.405 -145.355 ;
        RECT 29.075 -147.045 29.405 -146.715 ;
        RECT 29.075 -148.405 29.405 -148.075 ;
        RECT 29.075 -149.765 29.405 -149.435 ;
        RECT 29.075 -151.125 29.405 -150.795 ;
        RECT 29.075 -152.485 29.405 -152.155 ;
        RECT 29.075 -153.845 29.405 -153.515 ;
        RECT 29.075 -156.09 29.405 -154.96 ;
        RECT 29.08 -156.205 29.4 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 42.08 30.765 43.21 ;
        RECT 30.435 40.635 30.765 40.965 ;
        RECT 30.435 39.275 30.765 39.605 ;
        RECT 30.435 37.915 30.765 38.245 ;
        RECT 30.44 37.915 30.76 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 -1.525 30.765 -1.195 ;
        RECT 30.435 -2.885 30.765 -2.555 ;
        RECT 30.44 -3.56 30.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 -91.285 30.765 -90.955 ;
        RECT 30.435 -92.645 30.765 -92.315 ;
        RECT 30.435 -94.005 30.765 -93.675 ;
        RECT 30.435 -95.365 30.765 -95.035 ;
        RECT 30.435 -96.725 30.765 -96.395 ;
        RECT 30.435 -98.085 30.765 -97.755 ;
        RECT 30.435 -99.445 30.765 -99.115 ;
        RECT 30.435 -100.805 30.765 -100.475 ;
        RECT 30.435 -102.165 30.765 -101.835 ;
        RECT 30.435 -103.525 30.765 -103.195 ;
        RECT 30.435 -104.885 30.765 -104.555 ;
        RECT 30.435 -106.245 30.765 -105.915 ;
        RECT 30.435 -107.605 30.765 -107.275 ;
        RECT 30.435 -108.965 30.765 -108.635 ;
        RECT 30.435 -110.325 30.765 -109.995 ;
        RECT 30.435 -111.685 30.765 -111.355 ;
        RECT 30.435 -113.045 30.765 -112.715 ;
        RECT 30.435 -114.405 30.765 -114.075 ;
        RECT 30.435 -115.765 30.765 -115.435 ;
        RECT 30.435 -117.125 30.765 -116.795 ;
        RECT 30.435 -118.485 30.765 -118.155 ;
        RECT 30.435 -119.845 30.765 -119.515 ;
        RECT 30.435 -121.205 30.765 -120.875 ;
        RECT 30.435 -122.565 30.765 -122.235 ;
        RECT 30.435 -123.925 30.765 -123.595 ;
        RECT 30.435 -125.285 30.765 -124.955 ;
        RECT 30.435 -126.645 30.765 -126.315 ;
        RECT 30.435 -128.005 30.765 -127.675 ;
        RECT 30.435 -129.365 30.765 -129.035 ;
        RECT 30.435 -130.725 30.765 -130.395 ;
        RECT 30.435 -132.085 30.765 -131.755 ;
        RECT 30.435 -133.445 30.765 -133.115 ;
        RECT 30.435 -134.805 30.765 -134.475 ;
        RECT 30.435 -136.165 30.765 -135.835 ;
        RECT 30.435 -137.525 30.765 -137.195 ;
        RECT 30.435 -138.885 30.765 -138.555 ;
        RECT 30.435 -140.245 30.765 -139.915 ;
        RECT 30.435 -141.605 30.765 -141.275 ;
        RECT 30.435 -142.965 30.765 -142.635 ;
        RECT 30.435 -144.325 30.765 -143.995 ;
        RECT 30.435 -145.685 30.765 -145.355 ;
        RECT 30.435 -147.045 30.765 -146.715 ;
        RECT 30.435 -148.405 30.765 -148.075 ;
        RECT 30.435 -149.765 30.765 -149.435 ;
        RECT 30.435 -151.125 30.765 -150.795 ;
        RECT 30.435 -152.485 30.765 -152.155 ;
        RECT 30.435 -153.845 30.765 -153.515 ;
        RECT 30.435 -156.09 30.765 -154.96 ;
        RECT 30.44 -156.205 30.76 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 42.08 32.125 43.21 ;
        RECT 31.795 40.635 32.125 40.965 ;
        RECT 31.795 39.275 32.125 39.605 ;
        RECT 31.795 37.915 32.125 38.245 ;
        RECT 31.795 36.895 32.125 37.225 ;
        RECT 31.795 34.845 32.125 35.175 ;
        RECT 31.795 32.915 32.125 33.245 ;
        RECT 31.795 31.075 32.125 31.405 ;
        RECT 31.795 29.585 32.125 29.915 ;
        RECT 31.795 27.915 32.125 28.245 ;
        RECT 31.795 26.425 32.125 26.755 ;
        RECT 31.795 24.755 32.125 25.085 ;
        RECT 31.795 23.265 32.125 23.595 ;
        RECT 31.795 21.595 32.125 21.925 ;
        RECT 31.795 20.105 32.125 20.435 ;
        RECT 31.795 18.695 32.125 19.025 ;
        RECT 31.795 16.855 32.125 17.185 ;
        RECT 31.795 15.365 32.125 15.695 ;
        RECT 31.795 13.695 32.125 14.025 ;
        RECT 31.795 12.205 32.125 12.535 ;
        RECT 31.795 10.535 32.125 10.865 ;
        RECT 31.795 9.045 32.125 9.375 ;
        RECT 31.795 7.375 32.125 7.705 ;
        RECT 31.795 5.885 32.125 6.215 ;
        RECT 31.795 4.475 32.125 4.805 ;
        RECT 31.795 2.115 32.125 2.445 ;
        RECT 31.795 0.06 32.125 0.39 ;
        RECT 31.795 -1.525 32.125 -1.195 ;
        RECT 31.795 -2.885 32.125 -2.555 ;
        RECT 31.795 -4.245 32.125 -3.915 ;
        RECT 31.795 -5.605 32.125 -5.275 ;
        RECT 31.795 -6.965 32.125 -6.635 ;
        RECT 31.795 -8.325 32.125 -7.995 ;
        RECT 31.795 -9.685 32.125 -9.355 ;
        RECT 31.795 -11.045 32.125 -10.715 ;
        RECT 31.795 -12.405 32.125 -12.075 ;
        RECT 31.795 -13.765 32.125 -13.435 ;
        RECT 31.795 -15.125 32.125 -14.795 ;
        RECT 31.795 -16.485 32.125 -16.155 ;
        RECT 31.795 -17.845 32.125 -17.515 ;
        RECT 31.795 -19.205 32.125 -18.875 ;
        RECT 31.795 -20.565 32.125 -20.235 ;
        RECT 31.795 -21.925 32.125 -21.595 ;
        RECT 31.795 -23.285 32.125 -22.955 ;
        RECT 31.795 -24.645 32.125 -24.315 ;
        RECT 31.795 -26.005 32.125 -25.675 ;
        RECT 31.795 -27.365 32.125 -27.035 ;
        RECT 31.795 -28.725 32.125 -28.395 ;
        RECT 31.795 -30.085 32.125 -29.755 ;
        RECT 31.795 -31.445 32.125 -31.115 ;
        RECT 31.795 -32.805 32.125 -32.475 ;
        RECT 31.795 -34.165 32.125 -33.835 ;
        RECT 31.795 -35.525 32.125 -35.195 ;
        RECT 31.795 -36.885 32.125 -36.555 ;
        RECT 31.795 -38.245 32.125 -37.915 ;
        RECT 31.795 -39.605 32.125 -39.275 ;
        RECT 31.795 -40.965 32.125 -40.635 ;
        RECT 31.795 -42.325 32.125 -41.995 ;
        RECT 31.795 -43.685 32.125 -43.355 ;
        RECT 31.795 -45.045 32.125 -44.715 ;
        RECT 31.795 -46.405 32.125 -46.075 ;
        RECT 31.795 -47.765 32.125 -47.435 ;
        RECT 31.795 -49.125 32.125 -48.795 ;
        RECT 31.795 -50.485 32.125 -50.155 ;
        RECT 31.795 -51.845 32.125 -51.515 ;
        RECT 31.795 -53.205 32.125 -52.875 ;
        RECT 31.795 -54.565 32.125 -54.235 ;
        RECT 31.795 -55.925 32.125 -55.595 ;
        RECT 31.795 -57.285 32.125 -56.955 ;
        RECT 31.795 -58.645 32.125 -58.315 ;
        RECT 31.795 -60.005 32.125 -59.675 ;
        RECT 31.795 -61.365 32.125 -61.035 ;
        RECT 31.795 -62.725 32.125 -62.395 ;
        RECT 31.795 -64.085 32.125 -63.755 ;
        RECT 31.795 -65.445 32.125 -65.115 ;
        RECT 31.795 -66.805 32.125 -66.475 ;
        RECT 31.795 -68.165 32.125 -67.835 ;
        RECT 31.795 -69.525 32.125 -69.195 ;
        RECT 31.795 -70.885 32.125 -70.555 ;
        RECT 31.795 -72.245 32.125 -71.915 ;
        RECT 31.795 -73.605 32.125 -73.275 ;
        RECT 31.795 -74.965 32.125 -74.635 ;
        RECT 31.795 -76.325 32.125 -75.995 ;
        RECT 31.795 -77.685 32.125 -77.355 ;
        RECT 31.795 -79.045 32.125 -78.715 ;
        RECT 31.795 -80.405 32.125 -80.075 ;
        RECT 31.795 -81.765 32.125 -81.435 ;
        RECT 31.795 -83.125 32.125 -82.795 ;
        RECT 31.795 -84.485 32.125 -84.155 ;
        RECT 31.795 -85.845 32.125 -85.515 ;
        RECT 31.795 -87.205 32.125 -86.875 ;
        RECT 31.795 -88.565 32.125 -88.235 ;
        RECT 31.795 -89.925 32.125 -89.595 ;
        RECT 31.795 -91.285 32.125 -90.955 ;
        RECT 31.795 -92.645 32.125 -92.315 ;
        RECT 31.795 -94.005 32.125 -93.675 ;
        RECT 31.795 -95.365 32.125 -95.035 ;
        RECT 31.795 -96.725 32.125 -96.395 ;
        RECT 31.795 -98.085 32.125 -97.755 ;
        RECT 31.795 -99.445 32.125 -99.115 ;
        RECT 31.795 -100.805 32.125 -100.475 ;
        RECT 31.795 -102.165 32.125 -101.835 ;
        RECT 31.795 -103.525 32.125 -103.195 ;
        RECT 31.795 -104.885 32.125 -104.555 ;
        RECT 31.795 -106.245 32.125 -105.915 ;
        RECT 31.795 -107.605 32.125 -107.275 ;
        RECT 31.795 -108.965 32.125 -108.635 ;
        RECT 31.795 -110.325 32.125 -109.995 ;
        RECT 31.795 -111.685 32.125 -111.355 ;
        RECT 31.795 -113.045 32.125 -112.715 ;
        RECT 31.795 -114.405 32.125 -114.075 ;
        RECT 31.795 -115.765 32.125 -115.435 ;
        RECT 31.795 -117.125 32.125 -116.795 ;
        RECT 31.795 -118.485 32.125 -118.155 ;
        RECT 31.795 -119.845 32.125 -119.515 ;
        RECT 31.795 -121.205 32.125 -120.875 ;
        RECT 31.795 -122.565 32.125 -122.235 ;
        RECT 31.795 -123.925 32.125 -123.595 ;
        RECT 31.795 -125.285 32.125 -124.955 ;
        RECT 31.795 -126.645 32.125 -126.315 ;
        RECT 31.795 -128.005 32.125 -127.675 ;
        RECT 31.795 -129.365 32.125 -129.035 ;
        RECT 31.795 -130.725 32.125 -130.395 ;
        RECT 31.795 -132.085 32.125 -131.755 ;
        RECT 31.795 -133.445 32.125 -133.115 ;
        RECT 31.795 -134.805 32.125 -134.475 ;
        RECT 31.795 -136.165 32.125 -135.835 ;
        RECT 31.795 -137.525 32.125 -137.195 ;
        RECT 31.795 -138.885 32.125 -138.555 ;
        RECT 31.795 -140.245 32.125 -139.915 ;
        RECT 31.795 -141.605 32.125 -141.275 ;
        RECT 31.795 -142.965 32.125 -142.635 ;
        RECT 31.795 -144.325 32.125 -143.995 ;
        RECT 31.795 -145.685 32.125 -145.355 ;
        RECT 31.795 -147.045 32.125 -146.715 ;
        RECT 31.795 -148.405 32.125 -148.075 ;
        RECT 31.795 -149.765 32.125 -149.435 ;
        RECT 31.795 -151.125 32.125 -150.795 ;
        RECT 31.795 -152.485 32.125 -152.155 ;
        RECT 31.795 -153.845 32.125 -153.515 ;
        RECT 31.795 -156.09 32.125 -154.96 ;
        RECT 31.8 -156.205 32.12 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 42.08 33.485 43.21 ;
        RECT 33.155 40.635 33.485 40.965 ;
        RECT 33.155 39.275 33.485 39.605 ;
        RECT 33.155 37.915 33.485 38.245 ;
        RECT 33.155 36.895 33.485 37.225 ;
        RECT 33.155 34.845 33.485 35.175 ;
        RECT 33.155 32.915 33.485 33.245 ;
        RECT 33.155 31.075 33.485 31.405 ;
        RECT 33.155 29.585 33.485 29.915 ;
        RECT 33.155 27.915 33.485 28.245 ;
        RECT 33.155 26.425 33.485 26.755 ;
        RECT 33.155 24.755 33.485 25.085 ;
        RECT 33.155 23.265 33.485 23.595 ;
        RECT 33.155 21.595 33.485 21.925 ;
        RECT 33.155 20.105 33.485 20.435 ;
        RECT 33.155 18.695 33.485 19.025 ;
        RECT 33.155 16.855 33.485 17.185 ;
        RECT 33.155 15.365 33.485 15.695 ;
        RECT 33.155 13.695 33.485 14.025 ;
        RECT 33.155 12.205 33.485 12.535 ;
        RECT 33.155 10.535 33.485 10.865 ;
        RECT 33.155 9.045 33.485 9.375 ;
        RECT 33.155 7.375 33.485 7.705 ;
        RECT 33.155 5.885 33.485 6.215 ;
        RECT 33.155 4.475 33.485 4.805 ;
        RECT 33.155 2.115 33.485 2.445 ;
        RECT 33.155 0.06 33.485 0.39 ;
        RECT 33.155 -1.525 33.485 -1.195 ;
        RECT 33.155 -2.885 33.485 -2.555 ;
        RECT 33.155 -4.245 33.485 -3.915 ;
        RECT 33.155 -5.605 33.485 -5.275 ;
        RECT 33.155 -6.965 33.485 -6.635 ;
        RECT 33.155 -8.325 33.485 -7.995 ;
        RECT 33.155 -9.685 33.485 -9.355 ;
        RECT 33.155 -11.045 33.485 -10.715 ;
        RECT 33.155 -12.405 33.485 -12.075 ;
        RECT 33.155 -13.765 33.485 -13.435 ;
        RECT 33.155 -15.125 33.485 -14.795 ;
        RECT 33.155 -16.485 33.485 -16.155 ;
        RECT 33.155 -17.845 33.485 -17.515 ;
        RECT 33.155 -19.205 33.485 -18.875 ;
        RECT 33.155 -20.565 33.485 -20.235 ;
        RECT 33.155 -21.925 33.485 -21.595 ;
        RECT 33.155 -23.285 33.485 -22.955 ;
        RECT 33.155 -24.645 33.485 -24.315 ;
        RECT 33.155 -26.005 33.485 -25.675 ;
        RECT 33.155 -27.365 33.485 -27.035 ;
        RECT 33.155 -28.725 33.485 -28.395 ;
        RECT 33.155 -30.085 33.485 -29.755 ;
        RECT 33.155 -31.445 33.485 -31.115 ;
        RECT 33.155 -32.805 33.485 -32.475 ;
        RECT 33.155 -34.165 33.485 -33.835 ;
        RECT 33.155 -35.525 33.485 -35.195 ;
        RECT 33.155 -36.885 33.485 -36.555 ;
        RECT 33.155 -38.245 33.485 -37.915 ;
        RECT 33.155 -39.605 33.485 -39.275 ;
        RECT 33.155 -40.965 33.485 -40.635 ;
        RECT 33.155 -42.325 33.485 -41.995 ;
        RECT 33.155 -43.685 33.485 -43.355 ;
        RECT 33.155 -45.045 33.485 -44.715 ;
        RECT 33.155 -46.405 33.485 -46.075 ;
        RECT 33.155 -47.765 33.485 -47.435 ;
        RECT 33.155 -49.125 33.485 -48.795 ;
        RECT 33.155 -50.485 33.485 -50.155 ;
        RECT 33.155 -51.845 33.485 -51.515 ;
        RECT 33.155 -53.205 33.485 -52.875 ;
        RECT 33.155 -54.565 33.485 -54.235 ;
        RECT 33.155 -55.925 33.485 -55.595 ;
        RECT 33.155 -57.285 33.485 -56.955 ;
        RECT 33.155 -58.645 33.485 -58.315 ;
        RECT 33.155 -60.005 33.485 -59.675 ;
        RECT 33.155 -61.365 33.485 -61.035 ;
        RECT 33.155 -62.725 33.485 -62.395 ;
        RECT 33.155 -64.085 33.485 -63.755 ;
        RECT 33.155 -65.445 33.485 -65.115 ;
        RECT 33.155 -66.805 33.485 -66.475 ;
        RECT 33.155 -68.165 33.485 -67.835 ;
        RECT 33.155 -69.525 33.485 -69.195 ;
        RECT 33.155 -70.885 33.485 -70.555 ;
        RECT 33.155 -72.245 33.485 -71.915 ;
        RECT 33.155 -73.605 33.485 -73.275 ;
        RECT 33.155 -74.965 33.485 -74.635 ;
        RECT 33.155 -76.325 33.485 -75.995 ;
        RECT 33.155 -77.685 33.485 -77.355 ;
        RECT 33.155 -79.045 33.485 -78.715 ;
        RECT 33.155 -80.405 33.485 -80.075 ;
        RECT 33.155 -81.765 33.485 -81.435 ;
        RECT 33.155 -83.125 33.485 -82.795 ;
        RECT 33.155 -84.485 33.485 -84.155 ;
        RECT 33.155 -85.845 33.485 -85.515 ;
        RECT 33.155 -87.205 33.485 -86.875 ;
        RECT 33.155 -88.565 33.485 -88.235 ;
        RECT 33.155 -89.925 33.485 -89.595 ;
        RECT 33.155 -91.285 33.485 -90.955 ;
        RECT 33.155 -92.645 33.485 -92.315 ;
        RECT 33.155 -94.005 33.485 -93.675 ;
        RECT 33.155 -95.365 33.485 -95.035 ;
        RECT 33.155 -96.725 33.485 -96.395 ;
        RECT 33.155 -98.085 33.485 -97.755 ;
        RECT 33.155 -99.445 33.485 -99.115 ;
        RECT 33.155 -100.805 33.485 -100.475 ;
        RECT 33.155 -102.165 33.485 -101.835 ;
        RECT 33.155 -103.525 33.485 -103.195 ;
        RECT 33.155 -104.885 33.485 -104.555 ;
        RECT 33.155 -106.245 33.485 -105.915 ;
        RECT 33.155 -107.605 33.485 -107.275 ;
        RECT 33.155 -108.965 33.485 -108.635 ;
        RECT 33.155 -110.325 33.485 -109.995 ;
        RECT 33.155 -111.685 33.485 -111.355 ;
        RECT 33.155 -113.045 33.485 -112.715 ;
        RECT 33.155 -114.405 33.485 -114.075 ;
        RECT 33.155 -115.765 33.485 -115.435 ;
        RECT 33.155 -117.125 33.485 -116.795 ;
        RECT 33.155 -118.485 33.485 -118.155 ;
        RECT 33.155 -119.845 33.485 -119.515 ;
        RECT 33.155 -121.205 33.485 -120.875 ;
        RECT 33.155 -122.565 33.485 -122.235 ;
        RECT 33.155 -123.925 33.485 -123.595 ;
        RECT 33.155 -125.285 33.485 -124.955 ;
        RECT 33.155 -126.645 33.485 -126.315 ;
        RECT 33.155 -128.005 33.485 -127.675 ;
        RECT 33.155 -129.365 33.485 -129.035 ;
        RECT 33.155 -130.725 33.485 -130.395 ;
        RECT 33.155 -132.085 33.485 -131.755 ;
        RECT 33.155 -133.445 33.485 -133.115 ;
        RECT 33.155 -134.805 33.485 -134.475 ;
        RECT 33.155 -136.165 33.485 -135.835 ;
        RECT 33.155 -137.525 33.485 -137.195 ;
        RECT 33.155 -138.885 33.485 -138.555 ;
        RECT 33.155 -140.245 33.485 -139.915 ;
        RECT 33.155 -141.605 33.485 -141.275 ;
        RECT 33.155 -142.965 33.485 -142.635 ;
        RECT 33.155 -144.325 33.485 -143.995 ;
        RECT 33.155 -145.685 33.485 -145.355 ;
        RECT 33.155 -147.045 33.485 -146.715 ;
        RECT 33.155 -148.405 33.485 -148.075 ;
        RECT 33.155 -149.765 33.485 -149.435 ;
        RECT 33.155 -151.125 33.485 -150.795 ;
        RECT 33.155 -152.485 33.485 -152.155 ;
        RECT 33.155 -153.845 33.485 -153.515 ;
        RECT 33.155 -156.09 33.485 -154.96 ;
        RECT 33.16 -156.205 33.48 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 42.08 34.845 43.21 ;
        RECT 34.515 40.635 34.845 40.965 ;
        RECT 34.515 39.275 34.845 39.605 ;
        RECT 34.515 37.915 34.845 38.245 ;
        RECT 34.515 36.895 34.845 37.225 ;
        RECT 34.515 34.845 34.845 35.175 ;
        RECT 34.515 32.915 34.845 33.245 ;
        RECT 34.515 31.075 34.845 31.405 ;
        RECT 34.515 29.585 34.845 29.915 ;
        RECT 34.515 27.915 34.845 28.245 ;
        RECT 34.515 26.425 34.845 26.755 ;
        RECT 34.515 24.755 34.845 25.085 ;
        RECT 34.515 23.265 34.845 23.595 ;
        RECT 34.515 21.595 34.845 21.925 ;
        RECT 34.515 20.105 34.845 20.435 ;
        RECT 34.515 18.695 34.845 19.025 ;
        RECT 34.515 16.855 34.845 17.185 ;
        RECT 34.515 15.365 34.845 15.695 ;
        RECT 34.515 13.695 34.845 14.025 ;
        RECT 34.515 12.205 34.845 12.535 ;
        RECT 34.515 10.535 34.845 10.865 ;
        RECT 34.515 9.045 34.845 9.375 ;
        RECT 34.515 7.375 34.845 7.705 ;
        RECT 34.515 5.885 34.845 6.215 ;
        RECT 34.515 4.475 34.845 4.805 ;
        RECT 34.515 2.115 34.845 2.445 ;
        RECT 34.515 0.06 34.845 0.39 ;
        RECT 34.515 -1.525 34.845 -1.195 ;
        RECT 34.515 -2.885 34.845 -2.555 ;
        RECT 34.515 -4.245 34.845 -3.915 ;
        RECT 34.515 -5.605 34.845 -5.275 ;
        RECT 34.515 -6.965 34.845 -6.635 ;
        RECT 34.515 -8.325 34.845 -7.995 ;
        RECT 34.515 -9.685 34.845 -9.355 ;
        RECT 34.515 -11.045 34.845 -10.715 ;
        RECT 34.515 -12.405 34.845 -12.075 ;
        RECT 34.515 -13.765 34.845 -13.435 ;
        RECT 34.515 -15.125 34.845 -14.795 ;
        RECT 34.515 -16.485 34.845 -16.155 ;
        RECT 34.515 -17.845 34.845 -17.515 ;
        RECT 34.515 -19.205 34.845 -18.875 ;
        RECT 34.515 -20.565 34.845 -20.235 ;
        RECT 34.515 -21.925 34.845 -21.595 ;
        RECT 34.515 -23.285 34.845 -22.955 ;
        RECT 34.515 -24.645 34.845 -24.315 ;
        RECT 34.515 -26.005 34.845 -25.675 ;
        RECT 34.515 -27.365 34.845 -27.035 ;
        RECT 34.515 -28.725 34.845 -28.395 ;
        RECT 34.515 -30.085 34.845 -29.755 ;
        RECT 34.515 -31.445 34.845 -31.115 ;
        RECT 34.515 -32.805 34.845 -32.475 ;
        RECT 34.515 -34.165 34.845 -33.835 ;
        RECT 34.515 -35.525 34.845 -35.195 ;
        RECT 34.515 -36.885 34.845 -36.555 ;
        RECT 34.515 -38.245 34.845 -37.915 ;
        RECT 34.515 -39.605 34.845 -39.275 ;
        RECT 34.515 -40.965 34.845 -40.635 ;
        RECT 34.515 -42.325 34.845 -41.995 ;
        RECT 34.515 -43.685 34.845 -43.355 ;
        RECT 34.515 -45.045 34.845 -44.715 ;
        RECT 34.515 -46.405 34.845 -46.075 ;
        RECT 34.515 -47.765 34.845 -47.435 ;
        RECT 34.515 -49.125 34.845 -48.795 ;
        RECT 34.515 -50.485 34.845 -50.155 ;
        RECT 34.515 -51.845 34.845 -51.515 ;
        RECT 34.515 -53.205 34.845 -52.875 ;
        RECT 34.515 -54.565 34.845 -54.235 ;
        RECT 34.515 -55.925 34.845 -55.595 ;
        RECT 34.515 -57.285 34.845 -56.955 ;
        RECT 34.515 -58.645 34.845 -58.315 ;
        RECT 34.515 -60.005 34.845 -59.675 ;
        RECT 34.515 -61.365 34.845 -61.035 ;
        RECT 34.515 -62.725 34.845 -62.395 ;
        RECT 34.515 -64.085 34.845 -63.755 ;
        RECT 34.515 -65.445 34.845 -65.115 ;
        RECT 34.515 -66.805 34.845 -66.475 ;
        RECT 34.515 -68.165 34.845 -67.835 ;
        RECT 34.515 -69.525 34.845 -69.195 ;
        RECT 34.515 -70.885 34.845 -70.555 ;
        RECT 34.515 -72.245 34.845 -71.915 ;
        RECT 34.515 -73.605 34.845 -73.275 ;
        RECT 34.515 -74.965 34.845 -74.635 ;
        RECT 34.515 -76.325 34.845 -75.995 ;
        RECT 34.515 -77.685 34.845 -77.355 ;
        RECT 34.515 -79.045 34.845 -78.715 ;
        RECT 34.515 -80.405 34.845 -80.075 ;
        RECT 34.515 -81.765 34.845 -81.435 ;
        RECT 34.515 -83.125 34.845 -82.795 ;
        RECT 34.515 -84.485 34.845 -84.155 ;
        RECT 34.515 -85.845 34.845 -85.515 ;
        RECT 34.515 -87.205 34.845 -86.875 ;
        RECT 34.515 -88.565 34.845 -88.235 ;
        RECT 34.515 -89.925 34.845 -89.595 ;
        RECT 34.515 -91.285 34.845 -90.955 ;
        RECT 34.515 -92.645 34.845 -92.315 ;
        RECT 34.515 -94.005 34.845 -93.675 ;
        RECT 34.515 -95.365 34.845 -95.035 ;
        RECT 34.515 -96.725 34.845 -96.395 ;
        RECT 34.515 -98.085 34.845 -97.755 ;
        RECT 34.515 -99.445 34.845 -99.115 ;
        RECT 34.515 -100.805 34.845 -100.475 ;
        RECT 34.515 -102.165 34.845 -101.835 ;
        RECT 34.515 -103.525 34.845 -103.195 ;
        RECT 34.515 -104.885 34.845 -104.555 ;
        RECT 34.515 -106.245 34.845 -105.915 ;
        RECT 34.515 -107.605 34.845 -107.275 ;
        RECT 34.515 -108.965 34.845 -108.635 ;
        RECT 34.515 -110.325 34.845 -109.995 ;
        RECT 34.515 -111.685 34.845 -111.355 ;
        RECT 34.515 -113.045 34.845 -112.715 ;
        RECT 34.515 -114.405 34.845 -114.075 ;
        RECT 34.515 -115.765 34.845 -115.435 ;
        RECT 34.515 -117.125 34.845 -116.795 ;
        RECT 34.515 -118.485 34.845 -118.155 ;
        RECT 34.515 -119.845 34.845 -119.515 ;
        RECT 34.515 -121.205 34.845 -120.875 ;
        RECT 34.515 -122.565 34.845 -122.235 ;
        RECT 34.515 -123.925 34.845 -123.595 ;
        RECT 34.515 -125.285 34.845 -124.955 ;
        RECT 34.515 -126.645 34.845 -126.315 ;
        RECT 34.515 -128.005 34.845 -127.675 ;
        RECT 34.515 -129.365 34.845 -129.035 ;
        RECT 34.515 -130.725 34.845 -130.395 ;
        RECT 34.515 -132.085 34.845 -131.755 ;
        RECT 34.515 -133.445 34.845 -133.115 ;
        RECT 34.515 -134.805 34.845 -134.475 ;
        RECT 34.515 -136.165 34.845 -135.835 ;
        RECT 34.515 -137.525 34.845 -137.195 ;
        RECT 34.515 -138.885 34.845 -138.555 ;
        RECT 34.515 -140.245 34.845 -139.915 ;
        RECT 34.515 -141.605 34.845 -141.275 ;
        RECT 34.515 -142.965 34.845 -142.635 ;
        RECT 34.515 -144.325 34.845 -143.995 ;
        RECT 34.515 -145.685 34.845 -145.355 ;
        RECT 34.515 -147.045 34.845 -146.715 ;
        RECT 34.515 -148.405 34.845 -148.075 ;
        RECT 34.515 -149.765 34.845 -149.435 ;
        RECT 34.515 -151.125 34.845 -150.795 ;
        RECT 34.515 -152.485 34.845 -152.155 ;
        RECT 34.515 -153.845 34.845 -153.515 ;
        RECT 34.515 -156.09 34.845 -154.96 ;
        RECT 34.52 -156.205 34.84 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 42.08 36.205 43.21 ;
        RECT 35.875 40.635 36.205 40.965 ;
        RECT 35.875 39.275 36.205 39.605 ;
        RECT 35.875 37.915 36.205 38.245 ;
        RECT 35.875 36.895 36.205 37.225 ;
        RECT 35.875 34.845 36.205 35.175 ;
        RECT 35.875 32.915 36.205 33.245 ;
        RECT 35.875 31.075 36.205 31.405 ;
        RECT 35.875 29.585 36.205 29.915 ;
        RECT 35.875 27.915 36.205 28.245 ;
        RECT 35.875 26.425 36.205 26.755 ;
        RECT 35.875 24.755 36.205 25.085 ;
        RECT 35.875 23.265 36.205 23.595 ;
        RECT 35.875 21.595 36.205 21.925 ;
        RECT 35.875 20.105 36.205 20.435 ;
        RECT 35.875 18.695 36.205 19.025 ;
        RECT 35.875 16.855 36.205 17.185 ;
        RECT 35.875 15.365 36.205 15.695 ;
        RECT 35.875 13.695 36.205 14.025 ;
        RECT 35.875 12.205 36.205 12.535 ;
        RECT 35.875 10.535 36.205 10.865 ;
        RECT 35.875 9.045 36.205 9.375 ;
        RECT 35.875 7.375 36.205 7.705 ;
        RECT 35.875 5.885 36.205 6.215 ;
        RECT 35.875 4.475 36.205 4.805 ;
        RECT 35.875 2.115 36.205 2.445 ;
        RECT 35.875 0.06 36.205 0.39 ;
        RECT 35.875 -1.525 36.205 -1.195 ;
        RECT 35.875 -2.885 36.205 -2.555 ;
        RECT 35.875 -4.245 36.205 -3.915 ;
        RECT 35.875 -5.605 36.205 -5.275 ;
        RECT 35.875 -6.965 36.205 -6.635 ;
        RECT 35.875 -8.325 36.205 -7.995 ;
        RECT 35.875 -9.685 36.205 -9.355 ;
        RECT 35.875 -11.045 36.205 -10.715 ;
        RECT 35.875 -12.405 36.205 -12.075 ;
        RECT 35.875 -13.765 36.205 -13.435 ;
        RECT 35.875 -15.125 36.205 -14.795 ;
        RECT 35.875 -16.485 36.205 -16.155 ;
        RECT 35.875 -17.845 36.205 -17.515 ;
        RECT 35.875 -19.205 36.205 -18.875 ;
        RECT 35.875 -20.565 36.205 -20.235 ;
        RECT 35.875 -21.925 36.205 -21.595 ;
        RECT 35.875 -23.285 36.205 -22.955 ;
        RECT 35.875 -24.645 36.205 -24.315 ;
        RECT 35.875 -26.005 36.205 -25.675 ;
        RECT 35.875 -27.365 36.205 -27.035 ;
        RECT 35.875 -28.725 36.205 -28.395 ;
        RECT 35.875 -30.085 36.205 -29.755 ;
        RECT 35.875 -31.445 36.205 -31.115 ;
        RECT 35.875 -32.805 36.205 -32.475 ;
        RECT 35.875 -34.165 36.205 -33.835 ;
        RECT 35.875 -35.525 36.205 -35.195 ;
        RECT 35.875 -36.885 36.205 -36.555 ;
        RECT 35.875 -38.245 36.205 -37.915 ;
        RECT 35.875 -39.605 36.205 -39.275 ;
        RECT 35.875 -40.965 36.205 -40.635 ;
        RECT 35.875 -42.325 36.205 -41.995 ;
        RECT 35.875 -43.685 36.205 -43.355 ;
        RECT 35.875 -45.045 36.205 -44.715 ;
        RECT 35.875 -46.405 36.205 -46.075 ;
        RECT 35.875 -47.765 36.205 -47.435 ;
        RECT 35.875 -49.125 36.205 -48.795 ;
        RECT 35.875 -50.485 36.205 -50.155 ;
        RECT 35.875 -51.845 36.205 -51.515 ;
        RECT 35.875 -53.205 36.205 -52.875 ;
        RECT 35.875 -54.565 36.205 -54.235 ;
        RECT 35.875 -55.925 36.205 -55.595 ;
        RECT 35.875 -57.285 36.205 -56.955 ;
        RECT 35.875 -58.645 36.205 -58.315 ;
        RECT 35.875 -60.005 36.205 -59.675 ;
        RECT 35.875 -61.365 36.205 -61.035 ;
        RECT 35.875 -62.725 36.205 -62.395 ;
        RECT 35.875 -64.085 36.205 -63.755 ;
        RECT 35.875 -65.445 36.205 -65.115 ;
        RECT 35.875 -66.805 36.205 -66.475 ;
        RECT 35.875 -68.165 36.205 -67.835 ;
        RECT 35.875 -69.525 36.205 -69.195 ;
        RECT 35.875 -70.885 36.205 -70.555 ;
        RECT 35.875 -72.245 36.205 -71.915 ;
        RECT 35.875 -73.605 36.205 -73.275 ;
        RECT 35.875 -74.965 36.205 -74.635 ;
        RECT 35.875 -76.325 36.205 -75.995 ;
        RECT 35.875 -77.685 36.205 -77.355 ;
        RECT 35.875 -79.045 36.205 -78.715 ;
        RECT 35.875 -80.405 36.205 -80.075 ;
        RECT 35.875 -81.765 36.205 -81.435 ;
        RECT 35.875 -83.125 36.205 -82.795 ;
        RECT 35.875 -84.485 36.205 -84.155 ;
        RECT 35.875 -85.845 36.205 -85.515 ;
        RECT 35.875 -87.205 36.205 -86.875 ;
        RECT 35.875 -88.565 36.205 -88.235 ;
        RECT 35.875 -89.925 36.205 -89.595 ;
        RECT 35.875 -91.285 36.205 -90.955 ;
        RECT 35.875 -92.645 36.205 -92.315 ;
        RECT 35.875 -94.005 36.205 -93.675 ;
        RECT 35.875 -95.365 36.205 -95.035 ;
        RECT 35.875 -96.725 36.205 -96.395 ;
        RECT 35.875 -98.085 36.205 -97.755 ;
        RECT 35.875 -99.445 36.205 -99.115 ;
        RECT 35.875 -100.805 36.205 -100.475 ;
        RECT 35.875 -102.165 36.205 -101.835 ;
        RECT 35.875 -103.525 36.205 -103.195 ;
        RECT 35.875 -104.885 36.205 -104.555 ;
        RECT 35.875 -106.245 36.205 -105.915 ;
        RECT 35.875 -107.605 36.205 -107.275 ;
        RECT 35.875 -108.965 36.205 -108.635 ;
        RECT 35.875 -110.325 36.205 -109.995 ;
        RECT 35.875 -111.685 36.205 -111.355 ;
        RECT 35.875 -113.045 36.205 -112.715 ;
        RECT 35.875 -114.405 36.205 -114.075 ;
        RECT 35.875 -115.765 36.205 -115.435 ;
        RECT 35.875 -117.125 36.205 -116.795 ;
        RECT 35.875 -118.485 36.205 -118.155 ;
        RECT 35.875 -119.845 36.205 -119.515 ;
        RECT 35.875 -121.205 36.205 -120.875 ;
        RECT 35.875 -122.565 36.205 -122.235 ;
        RECT 35.875 -123.925 36.205 -123.595 ;
        RECT 35.875 -125.285 36.205 -124.955 ;
        RECT 35.875 -126.645 36.205 -126.315 ;
        RECT 35.875 -128.005 36.205 -127.675 ;
        RECT 35.875 -129.365 36.205 -129.035 ;
        RECT 35.875 -130.725 36.205 -130.395 ;
        RECT 35.875 -132.085 36.205 -131.755 ;
        RECT 35.875 -133.445 36.205 -133.115 ;
        RECT 35.875 -134.805 36.205 -134.475 ;
        RECT 35.875 -136.165 36.205 -135.835 ;
        RECT 35.875 -137.525 36.205 -137.195 ;
        RECT 35.875 -138.885 36.205 -138.555 ;
        RECT 35.875 -140.245 36.205 -139.915 ;
        RECT 35.875 -141.605 36.205 -141.275 ;
        RECT 35.875 -142.965 36.205 -142.635 ;
        RECT 35.875 -144.325 36.205 -143.995 ;
        RECT 35.875 -145.685 36.205 -145.355 ;
        RECT 35.875 -147.045 36.205 -146.715 ;
        RECT 35.875 -148.405 36.205 -148.075 ;
        RECT 35.875 -149.765 36.205 -149.435 ;
        RECT 35.875 -151.125 36.205 -150.795 ;
        RECT 35.875 -152.485 36.205 -152.155 ;
        RECT 35.875 -153.845 36.205 -153.515 ;
        RECT 35.875 -156.09 36.205 -154.96 ;
        RECT 35.88 -156.205 36.2 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.925 42.08 -4.595 43.21 ;
        RECT -4.925 40.635 -4.595 40.965 ;
        RECT -4.925 39.275 -4.595 39.605 ;
        RECT -4.925 37.915 -4.595 38.245 ;
        RECT -4.925 36.895 -4.595 37.225 ;
        RECT -4.925 34.845 -4.595 35.175 ;
        RECT -4.925 32.915 -4.595 33.245 ;
        RECT -4.925 31.075 -4.595 31.405 ;
        RECT -4.925 29.585 -4.595 29.915 ;
        RECT -4.925 27.915 -4.595 28.245 ;
        RECT -4.925 26.425 -4.595 26.755 ;
        RECT -4.925 24.755 -4.595 25.085 ;
        RECT -4.925 23.265 -4.595 23.595 ;
        RECT -4.925 21.595 -4.595 21.925 ;
        RECT -4.925 20.105 -4.595 20.435 ;
        RECT -4.925 18.695 -4.595 19.025 ;
        RECT -4.925 16.855 -4.595 17.185 ;
        RECT -4.925 15.365 -4.595 15.695 ;
        RECT -4.925 13.695 -4.595 14.025 ;
        RECT -4.925 12.205 -4.595 12.535 ;
        RECT -4.925 10.535 -4.595 10.865 ;
        RECT -4.925 9.045 -4.595 9.375 ;
        RECT -4.925 7.375 -4.595 7.705 ;
        RECT -4.925 5.885 -4.595 6.215 ;
        RECT -4.925 4.475 -4.595 4.805 ;
        RECT -4.925 2.115 -4.595 2.445 ;
        RECT -4.925 0.06 -4.595 0.39 ;
        RECT -4.925 -1.525 -4.595 -1.195 ;
        RECT -4.925 -2.885 -4.595 -2.555 ;
        RECT -4.925 -4.245 -4.595 -3.915 ;
        RECT -4.925 -5.605 -4.595 -5.275 ;
        RECT -4.925 -6.965 -4.595 -6.635 ;
        RECT -4.925 -8.325 -4.595 -7.995 ;
        RECT -4.925 -9.685 -4.595 -9.355 ;
        RECT -4.925 -12.405 -4.595 -12.075 ;
        RECT -4.925 -13.765 -4.595 -13.435 ;
        RECT -4.925 -15.125 -4.595 -14.795 ;
        RECT -4.925 -16.485 -4.595 -16.155 ;
        RECT -4.925 -17.845 -4.595 -17.515 ;
        RECT -4.925 -21.925 -4.595 -21.595 ;
        RECT -4.925 -23.285 -4.595 -22.955 ;
        RECT -4.925 -24.645 -4.595 -24.315 ;
        RECT -4.925 -26.005 -4.595 -25.675 ;
        RECT -4.925 -27.365 -4.595 -27.035 ;
        RECT -4.925 -28.725 -4.595 -28.395 ;
        RECT -4.925 -30.085 -4.595 -29.755 ;
        RECT -4.925 -31.445 -4.595 -31.115 ;
        RECT -4.925 -34.165 -4.595 -33.835 ;
        RECT -4.925 -35.525 -4.595 -35.195 ;
        RECT -4.925 -36.885 -4.595 -36.555 ;
        RECT -4.925 -38.245 -4.595 -37.915 ;
        RECT -4.925 -40.965 -4.595 -40.635 ;
        RECT -4.925 -42.325 -4.595 -41.995 ;
        RECT -4.925 -43.685 -4.595 -43.355 ;
        RECT -4.925 -46.405 -4.595 -46.075 ;
        RECT -4.925 -47.765 -4.595 -47.435 ;
        RECT -4.925 -49.125 -4.595 -48.795 ;
        RECT -4.925 -50.485 -4.595 -50.155 ;
        RECT -4.925 -51.845 -4.595 -51.515 ;
        RECT -4.925 -53.205 -4.595 -52.875 ;
        RECT -4.925 -54.565 -4.595 -54.235 ;
        RECT -4.925 -55.925 -4.595 -55.595 ;
        RECT -4.925 -57.285 -4.595 -56.955 ;
        RECT -4.925 -58.645 -4.595 -58.315 ;
        RECT -4.925 -60.005 -4.595 -59.675 ;
        RECT -4.925 -61.365 -4.595 -61.035 ;
        RECT -4.925 -62.725 -4.595 -62.395 ;
        RECT -4.925 -64.085 -4.595 -63.755 ;
        RECT -4.925 -65.445 -4.595 -65.115 ;
        RECT -4.925 -66.805 -4.595 -66.475 ;
        RECT -4.925 -68.165 -4.595 -67.835 ;
        RECT -4.925 -69.525 -4.595 -69.195 ;
        RECT -4.925 -70.885 -4.595 -70.555 ;
        RECT -4.925 -72.245 -4.595 -71.915 ;
        RECT -4.925 -73.605 -4.595 -73.275 ;
        RECT -4.925 -74.965 -4.595 -74.635 ;
        RECT -4.925 -76.325 -4.595 -75.995 ;
        RECT -4.925 -77.685 -4.595 -77.355 ;
        RECT -4.925 -79.045 -4.595 -78.715 ;
        RECT -4.925 -80.405 -4.595 -80.075 ;
        RECT -4.925 -81.765 -4.595 -81.435 ;
        RECT -4.925 -83.125 -4.595 -82.795 ;
        RECT -4.925 -84.485 -4.595 -84.155 ;
        RECT -4.925 -85.845 -4.595 -85.515 ;
        RECT -4.925 -87.205 -4.595 -86.875 ;
        RECT -4.925 -88.565 -4.595 -88.235 ;
        RECT -4.925 -89.925 -4.595 -89.595 ;
        RECT -4.925 -91.285 -4.595 -90.955 ;
        RECT -4.925 -92.645 -4.595 -92.315 ;
        RECT -4.925 -94.005 -4.595 -93.675 ;
        RECT -4.925 -95.365 -4.595 -95.035 ;
        RECT -4.925 -96.725 -4.595 -96.395 ;
        RECT -4.925 -98.085 -4.595 -97.755 ;
        RECT -4.925 -99.445 -4.595 -99.115 ;
        RECT -4.925 -100.805 -4.595 -100.475 ;
        RECT -4.925 -102.165 -4.595 -101.835 ;
        RECT -4.925 -103.525 -4.595 -103.195 ;
        RECT -4.925 -104.885 -4.595 -104.555 ;
        RECT -4.925 -106.245 -4.595 -105.915 ;
        RECT -4.925 -107.605 -4.595 -107.275 ;
        RECT -4.925 -108.965 -4.595 -108.635 ;
        RECT -4.925 -110.325 -4.595 -109.995 ;
        RECT -4.925 -111.685 -4.595 -111.355 ;
        RECT -4.925 -113.045 -4.595 -112.715 ;
        RECT -4.925 -114.405 -4.595 -114.075 ;
        RECT -4.925 -115.765 -4.595 -115.435 ;
        RECT -4.925 -117.125 -4.595 -116.795 ;
        RECT -4.925 -118.485 -4.595 -118.155 ;
        RECT -4.925 -119.845 -4.595 -119.515 ;
        RECT -4.925 -121.205 -4.595 -120.875 ;
        RECT -4.925 -122.565 -4.595 -122.235 ;
        RECT -4.925 -123.925 -4.595 -123.595 ;
        RECT -4.925 -125.285 -4.595 -124.955 ;
        RECT -4.925 -126.645 -4.595 -126.315 ;
        RECT -4.925 -128.005 -4.595 -127.675 ;
        RECT -4.925 -129.365 -4.595 -129.035 ;
        RECT -4.925 -130.725 -4.595 -130.395 ;
        RECT -4.925 -132.085 -4.595 -131.755 ;
        RECT -4.925 -133.445 -4.595 -133.115 ;
        RECT -4.925 -134.805 -4.595 -134.475 ;
        RECT -4.925 -136.165 -4.595 -135.835 ;
        RECT -4.925 -137.525 -4.595 -137.195 ;
        RECT -4.925 -138.885 -4.595 -138.555 ;
        RECT -4.925 -140.245 -4.595 -139.915 ;
        RECT -4.925 -141.605 -4.595 -141.275 ;
        RECT -4.925 -142.965 -4.595 -142.635 ;
        RECT -4.925 -144.325 -4.595 -143.995 ;
        RECT -4.925 -145.685 -4.595 -145.355 ;
        RECT -4.925 -147.045 -4.595 -146.715 ;
        RECT -4.925 -148.405 -4.595 -148.075 ;
        RECT -4.925 -149.765 -4.595 -149.435 ;
        RECT -4.925 -151.125 -4.595 -150.795 ;
        RECT -4.925 -152.485 -4.595 -152.155 ;
        RECT -4.925 -153.845 -4.595 -153.515 ;
        RECT -4.925 -156.09 -4.595 -154.96 ;
        RECT -4.92 -156.205 -4.6 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.565 42.08 -3.235 43.21 ;
        RECT -3.565 40.635 -3.235 40.965 ;
        RECT -3.565 39.275 -3.235 39.605 ;
        RECT -3.565 37.915 -3.235 38.245 ;
        RECT -3.565 36.895 -3.235 37.225 ;
        RECT -3.565 34.845 -3.235 35.175 ;
        RECT -3.565 32.915 -3.235 33.245 ;
        RECT -3.565 31.075 -3.235 31.405 ;
        RECT -3.565 29.585 -3.235 29.915 ;
        RECT -3.565 27.915 -3.235 28.245 ;
        RECT -3.565 26.425 -3.235 26.755 ;
        RECT -3.565 24.755 -3.235 25.085 ;
        RECT -3.565 23.265 -3.235 23.595 ;
        RECT -3.565 21.595 -3.235 21.925 ;
        RECT -3.565 20.105 -3.235 20.435 ;
        RECT -3.565 18.695 -3.235 19.025 ;
        RECT -3.565 16.855 -3.235 17.185 ;
        RECT -3.565 15.365 -3.235 15.695 ;
        RECT -3.565 13.695 -3.235 14.025 ;
        RECT -3.565 12.205 -3.235 12.535 ;
        RECT -3.565 10.535 -3.235 10.865 ;
        RECT -3.565 9.045 -3.235 9.375 ;
        RECT -3.565 7.375 -3.235 7.705 ;
        RECT -3.565 5.885 -3.235 6.215 ;
        RECT -3.565 4.475 -3.235 4.805 ;
        RECT -3.565 2.115 -3.235 2.445 ;
        RECT -3.565 0.06 -3.235 0.39 ;
        RECT -3.565 -1.525 -3.235 -1.195 ;
        RECT -3.565 -2.885 -3.235 -2.555 ;
        RECT -3.565 -4.245 -3.235 -3.915 ;
        RECT -3.565 -5.605 -3.235 -5.275 ;
        RECT -3.565 -6.965 -3.235 -6.635 ;
        RECT -3.565 -8.325 -3.235 -7.995 ;
        RECT -3.565 -9.685 -3.235 -9.355 ;
        RECT -3.565 -12.405 -3.235 -12.075 ;
        RECT -3.565 -13.765 -3.235 -13.435 ;
        RECT -3.565 -15.125 -3.235 -14.795 ;
        RECT -3.565 -16.485 -3.235 -16.155 ;
        RECT -3.565 -17.845 -3.235 -17.515 ;
        RECT -3.565 -21.925 -3.235 -21.595 ;
        RECT -3.565 -23.285 -3.235 -22.955 ;
        RECT -3.565 -24.645 -3.235 -24.315 ;
        RECT -3.565 -26.005 -3.235 -25.675 ;
        RECT -3.565 -27.365 -3.235 -27.035 ;
        RECT -3.565 -28.725 -3.235 -28.395 ;
        RECT -3.565 -30.085 -3.235 -29.755 ;
        RECT -3.565 -31.445 -3.235 -31.115 ;
        RECT -3.565 -34.165 -3.235 -33.835 ;
        RECT -3.565 -35.525 -3.235 -35.195 ;
        RECT -3.565 -36.885 -3.235 -36.555 ;
        RECT -3.565 -38.245 -3.235 -37.915 ;
        RECT -3.565 -40.965 -3.235 -40.635 ;
        RECT -3.565 -42.325 -3.235 -41.995 ;
        RECT -3.565 -43.685 -3.235 -43.355 ;
        RECT -3.565 -46.405 -3.235 -46.075 ;
        RECT -3.565 -47.765 -3.235 -47.435 ;
        RECT -3.565 -49.125 -3.235 -48.795 ;
        RECT -3.565 -50.485 -3.235 -50.155 ;
        RECT -3.565 -51.845 -3.235 -51.515 ;
        RECT -3.565 -53.205 -3.235 -52.875 ;
        RECT -3.565 -54.565 -3.235 -54.235 ;
        RECT -3.565 -55.925 -3.235 -55.595 ;
        RECT -3.565 -57.285 -3.235 -56.955 ;
        RECT -3.565 -58.645 -3.235 -58.315 ;
        RECT -3.565 -60.005 -3.235 -59.675 ;
        RECT -3.565 -61.365 -3.235 -61.035 ;
        RECT -3.565 -62.725 -3.235 -62.395 ;
        RECT -3.565 -64.085 -3.235 -63.755 ;
        RECT -3.565 -65.445 -3.235 -65.115 ;
        RECT -3.565 -66.805 -3.235 -66.475 ;
        RECT -3.565 -68.165 -3.235 -67.835 ;
        RECT -3.565 -69.525 -3.235 -69.195 ;
        RECT -3.565 -70.885 -3.235 -70.555 ;
        RECT -3.565 -72.245 -3.235 -71.915 ;
        RECT -3.565 -73.605 -3.235 -73.275 ;
        RECT -3.565 -74.965 -3.235 -74.635 ;
        RECT -3.565 -76.325 -3.235 -75.995 ;
        RECT -3.565 -77.685 -3.235 -77.355 ;
        RECT -3.565 -79.045 -3.235 -78.715 ;
        RECT -3.565 -80.405 -3.235 -80.075 ;
        RECT -3.565 -81.765 -3.235 -81.435 ;
        RECT -3.565 -83.125 -3.235 -82.795 ;
        RECT -3.565 -84.485 -3.235 -84.155 ;
        RECT -3.565 -85.845 -3.235 -85.515 ;
        RECT -3.565 -87.205 -3.235 -86.875 ;
        RECT -3.565 -88.565 -3.235 -88.235 ;
        RECT -3.565 -89.925 -3.235 -89.595 ;
        RECT -3.565 -91.285 -3.235 -90.955 ;
        RECT -3.565 -92.645 -3.235 -92.315 ;
        RECT -3.565 -94.005 -3.235 -93.675 ;
        RECT -3.565 -95.365 -3.235 -95.035 ;
        RECT -3.565 -96.725 -3.235 -96.395 ;
        RECT -3.565 -98.085 -3.235 -97.755 ;
        RECT -3.565 -99.445 -3.235 -99.115 ;
        RECT -3.565 -100.805 -3.235 -100.475 ;
        RECT -3.565 -102.165 -3.235 -101.835 ;
        RECT -3.565 -103.525 -3.235 -103.195 ;
        RECT -3.565 -104.885 -3.235 -104.555 ;
        RECT -3.565 -106.245 -3.235 -105.915 ;
        RECT -3.565 -107.605 -3.235 -107.275 ;
        RECT -3.565 -108.965 -3.235 -108.635 ;
        RECT -3.565 -110.325 -3.235 -109.995 ;
        RECT -3.565 -111.685 -3.235 -111.355 ;
        RECT -3.565 -113.045 -3.235 -112.715 ;
        RECT -3.565 -114.405 -3.235 -114.075 ;
        RECT -3.565 -115.765 -3.235 -115.435 ;
        RECT -3.565 -117.125 -3.235 -116.795 ;
        RECT -3.565 -118.485 -3.235 -118.155 ;
        RECT -3.565 -119.845 -3.235 -119.515 ;
        RECT -3.565 -121.205 -3.235 -120.875 ;
        RECT -3.565 -122.565 -3.235 -122.235 ;
        RECT -3.565 -123.925 -3.235 -123.595 ;
        RECT -3.565 -125.285 -3.235 -124.955 ;
        RECT -3.565 -126.645 -3.235 -126.315 ;
        RECT -3.565 -128.005 -3.235 -127.675 ;
        RECT -3.565 -129.365 -3.235 -129.035 ;
        RECT -3.565 -130.725 -3.235 -130.395 ;
        RECT -3.565 -132.085 -3.235 -131.755 ;
        RECT -3.565 -133.445 -3.235 -133.115 ;
        RECT -3.565 -134.805 -3.235 -134.475 ;
        RECT -3.565 -136.165 -3.235 -135.835 ;
        RECT -3.565 -137.525 -3.235 -137.195 ;
        RECT -3.565 -138.885 -3.235 -138.555 ;
        RECT -3.565 -140.245 -3.235 -139.915 ;
        RECT -3.565 -141.605 -3.235 -141.275 ;
        RECT -3.565 -142.965 -3.235 -142.635 ;
        RECT -3.565 -144.325 -3.235 -143.995 ;
        RECT -3.565 -145.685 -3.235 -145.355 ;
        RECT -3.565 -147.045 -3.235 -146.715 ;
        RECT -3.565 -148.405 -3.235 -148.075 ;
        RECT -3.565 -149.765 -3.235 -149.435 ;
        RECT -3.565 -151.125 -3.235 -150.795 ;
        RECT -3.565 -152.485 -3.235 -152.155 ;
        RECT -3.565 -153.845 -3.235 -153.515 ;
        RECT -3.565 -156.09 -3.235 -154.96 ;
        RECT -3.56 -156.205 -3.24 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.205 42.08 -1.875 43.21 ;
        RECT -2.205 40.635 -1.875 40.965 ;
        RECT -2.205 39.275 -1.875 39.605 ;
        RECT -2.205 37.915 -1.875 38.245 ;
        RECT -2.205 36.895 -1.875 37.225 ;
        RECT -2.205 34.845 -1.875 35.175 ;
        RECT -2.205 32.915 -1.875 33.245 ;
        RECT -2.205 31.075 -1.875 31.405 ;
        RECT -2.205 29.585 -1.875 29.915 ;
        RECT -2.205 27.915 -1.875 28.245 ;
        RECT -2.205 26.425 -1.875 26.755 ;
        RECT -2.205 24.755 -1.875 25.085 ;
        RECT -2.205 23.265 -1.875 23.595 ;
        RECT -2.205 21.595 -1.875 21.925 ;
        RECT -2.205 20.105 -1.875 20.435 ;
        RECT -2.205 18.695 -1.875 19.025 ;
        RECT -2.205 16.855 -1.875 17.185 ;
        RECT -2.205 15.365 -1.875 15.695 ;
        RECT -2.205 13.695 -1.875 14.025 ;
        RECT -2.205 12.205 -1.875 12.535 ;
        RECT -2.205 10.535 -1.875 10.865 ;
        RECT -2.205 9.045 -1.875 9.375 ;
        RECT -2.205 7.375 -1.875 7.705 ;
        RECT -2.205 5.885 -1.875 6.215 ;
        RECT -2.205 4.475 -1.875 4.805 ;
        RECT -2.205 2.115 -1.875 2.445 ;
        RECT -2.205 0.06 -1.875 0.39 ;
        RECT -2.205 -1.525 -1.875 -1.195 ;
        RECT -2.205 -2.885 -1.875 -2.555 ;
        RECT -2.205 -4.245 -1.875 -3.915 ;
        RECT -2.205 -5.605 -1.875 -5.275 ;
        RECT -2.205 -6.965 -1.875 -6.635 ;
        RECT -2.205 -8.325 -1.875 -7.995 ;
        RECT -2.205 -9.685 -1.875 -9.355 ;
        RECT -2.205 -12.405 -1.875 -12.075 ;
        RECT -2.205 -13.765 -1.875 -13.435 ;
        RECT -2.205 -15.125 -1.875 -14.795 ;
        RECT -2.205 -16.485 -1.875 -16.155 ;
        RECT -2.205 -17.845 -1.875 -17.515 ;
        RECT -2.205 -21.925 -1.875 -21.595 ;
        RECT -2.205 -23.285 -1.875 -22.955 ;
        RECT -2.205 -24.645 -1.875 -24.315 ;
        RECT -2.205 -26.005 -1.875 -25.675 ;
        RECT -2.205 -27.365 -1.875 -27.035 ;
        RECT -2.205 -28.725 -1.875 -28.395 ;
        RECT -2.205 -30.085 -1.875 -29.755 ;
        RECT -2.205 -31.445 -1.875 -31.115 ;
        RECT -2.205 -34.165 -1.875 -33.835 ;
        RECT -2.205 -35.525 -1.875 -35.195 ;
        RECT -2.205 -36.885 -1.875 -36.555 ;
        RECT -2.205 -38.245 -1.875 -37.915 ;
        RECT -2.205 -40.965 -1.875 -40.635 ;
        RECT -2.205 -42.325 -1.875 -41.995 ;
        RECT -2.205 -43.685 -1.875 -43.355 ;
        RECT -2.205 -46.405 -1.875 -46.075 ;
        RECT -2.205 -47.765 -1.875 -47.435 ;
        RECT -2.205 -49.125 -1.875 -48.795 ;
        RECT -2.205 -50.485 -1.875 -50.155 ;
        RECT -2.205 -51.845 -1.875 -51.515 ;
        RECT -2.205 -53.205 -1.875 -52.875 ;
        RECT -2.205 -54.565 -1.875 -54.235 ;
        RECT -2.205 -55.925 -1.875 -55.595 ;
        RECT -2.205 -57.285 -1.875 -56.955 ;
        RECT -2.205 -58.645 -1.875 -58.315 ;
        RECT -2.205 -60.005 -1.875 -59.675 ;
        RECT -2.205 -61.365 -1.875 -61.035 ;
        RECT -2.205 -62.725 -1.875 -62.395 ;
        RECT -2.205 -64.085 -1.875 -63.755 ;
        RECT -2.205 -65.445 -1.875 -65.115 ;
        RECT -2.205 -66.805 -1.875 -66.475 ;
        RECT -2.205 -68.165 -1.875 -67.835 ;
        RECT -2.205 -69.525 -1.875 -69.195 ;
        RECT -2.205 -70.885 -1.875 -70.555 ;
        RECT -2.205 -72.245 -1.875 -71.915 ;
        RECT -2.205 -73.605 -1.875 -73.275 ;
        RECT -2.205 -74.965 -1.875 -74.635 ;
        RECT -2.205 -76.325 -1.875 -75.995 ;
        RECT -2.205 -77.685 -1.875 -77.355 ;
        RECT -2.205 -79.045 -1.875 -78.715 ;
        RECT -2.205 -80.405 -1.875 -80.075 ;
        RECT -2.205 -81.765 -1.875 -81.435 ;
        RECT -2.205 -83.125 -1.875 -82.795 ;
        RECT -2.205 -84.485 -1.875 -84.155 ;
        RECT -2.205 -85.845 -1.875 -85.515 ;
        RECT -2.205 -87.205 -1.875 -86.875 ;
        RECT -2.205 -88.565 -1.875 -88.235 ;
        RECT -2.205 -89.925 -1.875 -89.595 ;
        RECT -2.205 -91.285 -1.875 -90.955 ;
        RECT -2.205 -92.645 -1.875 -92.315 ;
        RECT -2.205 -94.005 -1.875 -93.675 ;
        RECT -2.205 -95.365 -1.875 -95.035 ;
        RECT -2.205 -96.725 -1.875 -96.395 ;
        RECT -2.205 -98.085 -1.875 -97.755 ;
        RECT -2.205 -99.445 -1.875 -99.115 ;
        RECT -2.205 -100.805 -1.875 -100.475 ;
        RECT -2.205 -102.165 -1.875 -101.835 ;
        RECT -2.205 -103.525 -1.875 -103.195 ;
        RECT -2.205 -104.885 -1.875 -104.555 ;
        RECT -2.205 -106.245 -1.875 -105.915 ;
        RECT -2.205 -107.605 -1.875 -107.275 ;
        RECT -2.205 -108.965 -1.875 -108.635 ;
        RECT -2.205 -110.325 -1.875 -109.995 ;
        RECT -2.205 -111.685 -1.875 -111.355 ;
        RECT -2.205 -113.045 -1.875 -112.715 ;
        RECT -2.205 -114.405 -1.875 -114.075 ;
        RECT -2.205 -115.765 -1.875 -115.435 ;
        RECT -2.205 -117.125 -1.875 -116.795 ;
        RECT -2.205 -118.485 -1.875 -118.155 ;
        RECT -2.205 -119.845 -1.875 -119.515 ;
        RECT -2.205 -121.205 -1.875 -120.875 ;
        RECT -2.205 -122.565 -1.875 -122.235 ;
        RECT -2.205 -123.925 -1.875 -123.595 ;
        RECT -2.205 -125.285 -1.875 -124.955 ;
        RECT -2.205 -126.645 -1.875 -126.315 ;
        RECT -2.205 -128.005 -1.875 -127.675 ;
        RECT -2.205 -129.365 -1.875 -129.035 ;
        RECT -2.205 -130.725 -1.875 -130.395 ;
        RECT -2.205 -132.085 -1.875 -131.755 ;
        RECT -2.205 -133.445 -1.875 -133.115 ;
        RECT -2.205 -134.805 -1.875 -134.475 ;
        RECT -2.205 -136.165 -1.875 -135.835 ;
        RECT -2.205 -137.525 -1.875 -137.195 ;
        RECT -2.205 -138.885 -1.875 -138.555 ;
        RECT -2.205 -140.245 -1.875 -139.915 ;
        RECT -2.205 -141.605 -1.875 -141.275 ;
        RECT -2.205 -142.965 -1.875 -142.635 ;
        RECT -2.205 -144.325 -1.875 -143.995 ;
        RECT -2.205 -145.685 -1.875 -145.355 ;
        RECT -2.205 -147.045 -1.875 -146.715 ;
        RECT -2.205 -148.405 -1.875 -148.075 ;
        RECT -2.205 -149.765 -1.875 -149.435 ;
        RECT -2.205 -151.125 -1.875 -150.795 ;
        RECT -2.205 -152.485 -1.875 -152.155 ;
        RECT -2.205 -153.845 -1.875 -153.515 ;
        RECT -2.205 -156.09 -1.875 -154.96 ;
        RECT -2.2 -156.205 -1.88 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.845 42.08 -0.515 43.21 ;
        RECT -0.845 40.635 -0.515 40.965 ;
        RECT -0.845 39.275 -0.515 39.605 ;
        RECT -0.845 37.915 -0.515 38.245 ;
        RECT -0.845 36.895 -0.515 37.225 ;
        RECT -0.845 34.845 -0.515 35.175 ;
        RECT -0.845 32.915 -0.515 33.245 ;
        RECT -0.845 31.075 -0.515 31.405 ;
        RECT -0.845 29.585 -0.515 29.915 ;
        RECT -0.845 27.915 -0.515 28.245 ;
        RECT -0.845 26.425 -0.515 26.755 ;
        RECT -0.845 24.755 -0.515 25.085 ;
        RECT -0.845 23.265 -0.515 23.595 ;
        RECT -0.845 21.595 -0.515 21.925 ;
        RECT -0.845 20.105 -0.515 20.435 ;
        RECT -0.845 18.695 -0.515 19.025 ;
        RECT -0.845 16.855 -0.515 17.185 ;
        RECT -0.845 15.365 -0.515 15.695 ;
        RECT -0.845 13.695 -0.515 14.025 ;
        RECT -0.845 12.205 -0.515 12.535 ;
        RECT -0.845 10.535 -0.515 10.865 ;
        RECT -0.845 9.045 -0.515 9.375 ;
        RECT -0.845 7.375 -0.515 7.705 ;
        RECT -0.845 5.885 -0.515 6.215 ;
        RECT -0.845 4.475 -0.515 4.805 ;
        RECT -0.845 2.115 -0.515 2.445 ;
        RECT -0.845 0.06 -0.515 0.39 ;
        RECT -0.845 -1.525 -0.515 -1.195 ;
        RECT -0.845 -2.885 -0.515 -2.555 ;
        RECT -0.845 -4.245 -0.515 -3.915 ;
        RECT -0.845 -5.605 -0.515 -5.275 ;
        RECT -0.845 -6.965 -0.515 -6.635 ;
        RECT -0.845 -8.325 -0.515 -7.995 ;
        RECT -0.845 -9.685 -0.515 -9.355 ;
        RECT -0.845 -12.405 -0.515 -12.075 ;
        RECT -0.845 -13.765 -0.515 -13.435 ;
        RECT -0.845 -15.125 -0.515 -14.795 ;
        RECT -0.845 -16.485 -0.515 -16.155 ;
        RECT -0.845 -17.845 -0.515 -17.515 ;
        RECT -0.845 -21.925 -0.515 -21.595 ;
        RECT -0.845 -23.285 -0.515 -22.955 ;
        RECT -0.845 -24.645 -0.515 -24.315 ;
        RECT -0.845 -26.005 -0.515 -25.675 ;
        RECT -0.845 -27.365 -0.515 -27.035 ;
        RECT -0.845 -28.725 -0.515 -28.395 ;
        RECT -0.845 -30.085 -0.515 -29.755 ;
        RECT -0.845 -31.445 -0.515 -31.115 ;
        RECT -0.845 -34.165 -0.515 -33.835 ;
        RECT -0.845 -35.525 -0.515 -35.195 ;
        RECT -0.845 -36.885 -0.515 -36.555 ;
        RECT -0.845 -38.245 -0.515 -37.915 ;
        RECT -0.845 -40.965 -0.515 -40.635 ;
        RECT -0.845 -42.325 -0.515 -41.995 ;
        RECT -0.845 -43.685 -0.515 -43.355 ;
        RECT -0.845 -46.405 -0.515 -46.075 ;
        RECT -0.845 -47.765 -0.515 -47.435 ;
        RECT -0.845 -49.125 -0.515 -48.795 ;
        RECT -0.845 -50.485 -0.515 -50.155 ;
        RECT -0.845 -51.845 -0.515 -51.515 ;
        RECT -0.845 -53.205 -0.515 -52.875 ;
        RECT -0.845 -54.565 -0.515 -54.235 ;
        RECT -0.845 -55.925 -0.515 -55.595 ;
        RECT -0.845 -57.285 -0.515 -56.955 ;
        RECT -0.845 -58.645 -0.515 -58.315 ;
        RECT -0.845 -60.005 -0.515 -59.675 ;
        RECT -0.845 -61.365 -0.515 -61.035 ;
        RECT -0.845 -62.725 -0.515 -62.395 ;
        RECT -0.845 -64.085 -0.515 -63.755 ;
        RECT -0.845 -65.445 -0.515 -65.115 ;
        RECT -0.845 -66.805 -0.515 -66.475 ;
        RECT -0.845 -68.165 -0.515 -67.835 ;
        RECT -0.845 -69.525 -0.515 -69.195 ;
        RECT -0.845 -70.885 -0.515 -70.555 ;
        RECT -0.845 -72.245 -0.515 -71.915 ;
        RECT -0.845 -73.605 -0.515 -73.275 ;
        RECT -0.845 -74.965 -0.515 -74.635 ;
        RECT -0.845 -76.325 -0.515 -75.995 ;
        RECT -0.845 -77.685 -0.515 -77.355 ;
        RECT -0.845 -79.045 -0.515 -78.715 ;
        RECT -0.845 -80.405 -0.515 -80.075 ;
        RECT -0.845 -81.765 -0.515 -81.435 ;
        RECT -0.845 -83.125 -0.515 -82.795 ;
        RECT -0.845 -84.485 -0.515 -84.155 ;
        RECT -0.845 -85.845 -0.515 -85.515 ;
        RECT -0.845 -87.205 -0.515 -86.875 ;
        RECT -0.845 -88.565 -0.515 -88.235 ;
        RECT -0.845 -89.925 -0.515 -89.595 ;
        RECT -0.845 -91.285 -0.515 -90.955 ;
        RECT -0.845 -92.645 -0.515 -92.315 ;
        RECT -0.845 -94.005 -0.515 -93.675 ;
        RECT -0.845 -95.365 -0.515 -95.035 ;
        RECT -0.845 -96.725 -0.515 -96.395 ;
        RECT -0.845 -98.085 -0.515 -97.755 ;
        RECT -0.845 -99.445 -0.515 -99.115 ;
        RECT -0.845 -100.805 -0.515 -100.475 ;
        RECT -0.845 -102.165 -0.515 -101.835 ;
        RECT -0.845 -103.525 -0.515 -103.195 ;
        RECT -0.845 -104.885 -0.515 -104.555 ;
        RECT -0.845 -106.245 -0.515 -105.915 ;
        RECT -0.845 -107.605 -0.515 -107.275 ;
        RECT -0.845 -108.965 -0.515 -108.635 ;
        RECT -0.845 -110.325 -0.515 -109.995 ;
        RECT -0.845 -111.685 -0.515 -111.355 ;
        RECT -0.845 -113.045 -0.515 -112.715 ;
        RECT -0.845 -114.405 -0.515 -114.075 ;
        RECT -0.845 -115.765 -0.515 -115.435 ;
        RECT -0.845 -117.125 -0.515 -116.795 ;
        RECT -0.845 -118.485 -0.515 -118.155 ;
        RECT -0.845 -119.845 -0.515 -119.515 ;
        RECT -0.845 -121.205 -0.515 -120.875 ;
        RECT -0.845 -122.565 -0.515 -122.235 ;
        RECT -0.845 -123.925 -0.515 -123.595 ;
        RECT -0.845 -125.285 -0.515 -124.955 ;
        RECT -0.845 -126.645 -0.515 -126.315 ;
        RECT -0.845 -128.005 -0.515 -127.675 ;
        RECT -0.845 -129.365 -0.515 -129.035 ;
        RECT -0.845 -130.725 -0.515 -130.395 ;
        RECT -0.845 -132.085 -0.515 -131.755 ;
        RECT -0.845 -133.445 -0.515 -133.115 ;
        RECT -0.845 -134.805 -0.515 -134.475 ;
        RECT -0.845 -136.165 -0.515 -135.835 ;
        RECT -0.845 -137.525 -0.515 -137.195 ;
        RECT -0.845 -138.885 -0.515 -138.555 ;
        RECT -0.845 -140.245 -0.515 -139.915 ;
        RECT -0.845 -141.605 -0.515 -141.275 ;
        RECT -0.845 -142.965 -0.515 -142.635 ;
        RECT -0.845 -144.325 -0.515 -143.995 ;
        RECT -0.845 -145.685 -0.515 -145.355 ;
        RECT -0.845 -147.045 -0.515 -146.715 ;
        RECT -0.845 -148.405 -0.515 -148.075 ;
        RECT -0.845 -149.765 -0.515 -149.435 ;
        RECT -0.845 -151.125 -0.515 -150.795 ;
        RECT -0.845 -152.485 -0.515 -152.155 ;
        RECT -0.845 -153.845 -0.515 -153.515 ;
        RECT -0.845 -156.09 -0.515 -154.96 ;
        RECT -0.84 -156.205 -0.52 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 42.08 0.845 43.21 ;
        RECT 0.515 40.635 0.845 40.965 ;
        RECT 0.515 39.275 0.845 39.605 ;
        RECT 0.515 37.915 0.845 38.245 ;
        RECT 0.52 37.915 0.84 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 -1.525 0.845 -1.195 ;
        RECT 0.515 -2.885 0.845 -2.555 ;
        RECT 0.52 -3.56 0.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 -91.285 0.845 -90.955 ;
        RECT 0.515 -92.645 0.845 -92.315 ;
        RECT 0.515 -94.005 0.845 -93.675 ;
        RECT 0.515 -95.365 0.845 -95.035 ;
        RECT 0.515 -96.725 0.845 -96.395 ;
        RECT 0.515 -98.085 0.845 -97.755 ;
        RECT 0.515 -99.445 0.845 -99.115 ;
        RECT 0.515 -100.805 0.845 -100.475 ;
        RECT 0.515 -102.165 0.845 -101.835 ;
        RECT 0.515 -103.525 0.845 -103.195 ;
        RECT 0.515 -104.885 0.845 -104.555 ;
        RECT 0.515 -106.245 0.845 -105.915 ;
        RECT 0.515 -107.605 0.845 -107.275 ;
        RECT 0.515 -108.965 0.845 -108.635 ;
        RECT 0.515 -110.325 0.845 -109.995 ;
        RECT 0.515 -111.685 0.845 -111.355 ;
        RECT 0.515 -113.045 0.845 -112.715 ;
        RECT 0.515 -114.405 0.845 -114.075 ;
        RECT 0.515 -115.765 0.845 -115.435 ;
        RECT 0.515 -117.125 0.845 -116.795 ;
        RECT 0.515 -118.485 0.845 -118.155 ;
        RECT 0.515 -119.845 0.845 -119.515 ;
        RECT 0.515 -121.205 0.845 -120.875 ;
        RECT 0.515 -122.565 0.845 -122.235 ;
        RECT 0.515 -123.925 0.845 -123.595 ;
        RECT 0.515 -125.285 0.845 -124.955 ;
        RECT 0.515 -126.645 0.845 -126.315 ;
        RECT 0.515 -128.005 0.845 -127.675 ;
        RECT 0.515 -129.365 0.845 -129.035 ;
        RECT 0.515 -130.725 0.845 -130.395 ;
        RECT 0.515 -132.085 0.845 -131.755 ;
        RECT 0.515 -133.445 0.845 -133.115 ;
        RECT 0.515 -134.805 0.845 -134.475 ;
        RECT 0.515 -136.165 0.845 -135.835 ;
        RECT 0.515 -137.525 0.845 -137.195 ;
        RECT 0.515 -138.885 0.845 -138.555 ;
        RECT 0.515 -140.245 0.845 -139.915 ;
        RECT 0.515 -141.605 0.845 -141.275 ;
        RECT 0.515 -142.965 0.845 -142.635 ;
        RECT 0.515 -144.325 0.845 -143.995 ;
        RECT 0.515 -145.685 0.845 -145.355 ;
        RECT 0.515 -147.045 0.845 -146.715 ;
        RECT 0.515 -148.405 0.845 -148.075 ;
        RECT 0.515 -149.765 0.845 -149.435 ;
        RECT 0.515 -151.125 0.845 -150.795 ;
        RECT 0.515 -152.485 0.845 -152.155 ;
        RECT 0.515 -153.845 0.845 -153.515 ;
        RECT 0.515 -156.09 0.845 -154.96 ;
        RECT 0.52 -156.205 0.84 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 42.08 2.205 43.21 ;
        RECT 1.875 40.635 2.205 40.965 ;
        RECT 1.875 39.275 2.205 39.605 ;
        RECT 1.875 37.915 2.205 38.245 ;
        RECT 1.88 37.915 2.2 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 -1.525 2.205 -1.195 ;
        RECT 1.875 -2.885 2.205 -2.555 ;
        RECT 1.88 -3.56 2.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 -91.285 2.205 -90.955 ;
        RECT 1.875 -92.645 2.205 -92.315 ;
        RECT 1.875 -94.005 2.205 -93.675 ;
        RECT 1.875 -95.365 2.205 -95.035 ;
        RECT 1.875 -96.725 2.205 -96.395 ;
        RECT 1.875 -98.085 2.205 -97.755 ;
        RECT 1.875 -99.445 2.205 -99.115 ;
        RECT 1.875 -100.805 2.205 -100.475 ;
        RECT 1.875 -102.165 2.205 -101.835 ;
        RECT 1.875 -103.525 2.205 -103.195 ;
        RECT 1.875 -104.885 2.205 -104.555 ;
        RECT 1.875 -106.245 2.205 -105.915 ;
        RECT 1.875 -107.605 2.205 -107.275 ;
        RECT 1.875 -108.965 2.205 -108.635 ;
        RECT 1.875 -110.325 2.205 -109.995 ;
        RECT 1.875 -111.685 2.205 -111.355 ;
        RECT 1.875 -113.045 2.205 -112.715 ;
        RECT 1.875 -114.405 2.205 -114.075 ;
        RECT 1.875 -115.765 2.205 -115.435 ;
        RECT 1.875 -117.125 2.205 -116.795 ;
        RECT 1.875 -118.485 2.205 -118.155 ;
        RECT 1.875 -119.845 2.205 -119.515 ;
        RECT 1.875 -121.205 2.205 -120.875 ;
        RECT 1.875 -122.565 2.205 -122.235 ;
        RECT 1.875 -123.925 2.205 -123.595 ;
        RECT 1.875 -125.285 2.205 -124.955 ;
        RECT 1.875 -126.645 2.205 -126.315 ;
        RECT 1.875 -128.005 2.205 -127.675 ;
        RECT 1.875 -129.365 2.205 -129.035 ;
        RECT 1.875 -130.725 2.205 -130.395 ;
        RECT 1.875 -132.085 2.205 -131.755 ;
        RECT 1.875 -133.445 2.205 -133.115 ;
        RECT 1.875 -134.805 2.205 -134.475 ;
        RECT 1.875 -136.165 2.205 -135.835 ;
        RECT 1.875 -137.525 2.205 -137.195 ;
        RECT 1.875 -138.885 2.205 -138.555 ;
        RECT 1.875 -140.245 2.205 -139.915 ;
        RECT 1.875 -141.605 2.205 -141.275 ;
        RECT 1.875 -142.965 2.205 -142.635 ;
        RECT 1.875 -144.325 2.205 -143.995 ;
        RECT 1.875 -145.685 2.205 -145.355 ;
        RECT 1.875 -147.045 2.205 -146.715 ;
        RECT 1.875 -148.405 2.205 -148.075 ;
        RECT 1.875 -149.765 2.205 -149.435 ;
        RECT 1.875 -151.125 2.205 -150.795 ;
        RECT 1.875 -152.485 2.205 -152.155 ;
        RECT 1.875 -153.845 2.205 -153.515 ;
        RECT 1.875 -156.09 2.205 -154.96 ;
        RECT 1.88 -156.205 2.2 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 42.08 3.565 43.21 ;
        RECT 3.235 40.635 3.565 40.965 ;
        RECT 3.235 39.275 3.565 39.605 ;
        RECT 3.235 37.915 3.565 38.245 ;
        RECT 3.24 37.915 3.56 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 -95.365 3.565 -95.035 ;
        RECT 3.235 -96.725 3.565 -96.395 ;
        RECT 3.235 -98.085 3.565 -97.755 ;
        RECT 3.235 -99.445 3.565 -99.115 ;
        RECT 3.235 -100.805 3.565 -100.475 ;
        RECT 3.235 -102.165 3.565 -101.835 ;
        RECT 3.235 -103.525 3.565 -103.195 ;
        RECT 3.235 -104.885 3.565 -104.555 ;
        RECT 3.235 -106.245 3.565 -105.915 ;
        RECT 3.235 -107.605 3.565 -107.275 ;
        RECT 3.235 -108.965 3.565 -108.635 ;
        RECT 3.235 -110.325 3.565 -109.995 ;
        RECT 3.235 -111.685 3.565 -111.355 ;
        RECT 3.235 -113.045 3.565 -112.715 ;
        RECT 3.235 -114.405 3.565 -114.075 ;
        RECT 3.235 -115.765 3.565 -115.435 ;
        RECT 3.235 -117.125 3.565 -116.795 ;
        RECT 3.235 -118.485 3.565 -118.155 ;
        RECT 3.235 -119.845 3.565 -119.515 ;
        RECT 3.235 -121.205 3.565 -120.875 ;
        RECT 3.235 -122.565 3.565 -122.235 ;
        RECT 3.235 -123.925 3.565 -123.595 ;
        RECT 3.235 -125.285 3.565 -124.955 ;
        RECT 3.235 -126.645 3.565 -126.315 ;
        RECT 3.235 -128.005 3.565 -127.675 ;
        RECT 3.235 -129.365 3.565 -129.035 ;
        RECT 3.235 -130.725 3.565 -130.395 ;
        RECT 3.235 -132.085 3.565 -131.755 ;
        RECT 3.235 -133.445 3.565 -133.115 ;
        RECT 3.235 -134.805 3.565 -134.475 ;
        RECT 3.235 -136.165 3.565 -135.835 ;
        RECT 3.235 -137.525 3.565 -137.195 ;
        RECT 3.235 -138.885 3.565 -138.555 ;
        RECT 3.235 -140.245 3.565 -139.915 ;
        RECT 3.235 -141.605 3.565 -141.275 ;
        RECT 3.235 -142.965 3.565 -142.635 ;
        RECT 3.235 -144.325 3.565 -143.995 ;
        RECT 3.235 -145.685 3.565 -145.355 ;
        RECT 3.235 -147.045 3.565 -146.715 ;
        RECT 3.235 -148.405 3.565 -148.075 ;
        RECT 3.235 -149.765 3.565 -149.435 ;
        RECT 3.235 -151.125 3.565 -150.795 ;
        RECT 3.235 -152.485 3.565 -152.155 ;
        RECT 3.235 -153.845 3.565 -153.515 ;
        RECT 3.235 -156.09 3.565 -154.96 ;
        RECT 3.24 -156.205 3.56 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.31 -94.075 3.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 42.08 4.925 43.21 ;
        RECT 4.595 40.635 4.925 40.965 ;
        RECT 4.595 39.275 4.925 39.605 ;
        RECT 4.595 37.915 4.925 38.245 ;
        RECT 4.6 37.915 4.92 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 -1.525 4.925 -1.195 ;
        RECT 4.595 -2.885 4.925 -2.555 ;
        RECT 4.6 -3.56 4.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 42.08 6.285 43.21 ;
        RECT 5.955 40.635 6.285 40.965 ;
        RECT 5.955 39.275 6.285 39.605 ;
        RECT 5.955 37.915 6.285 38.245 ;
        RECT 5.96 37.915 6.28 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 -1.525 6.285 -1.195 ;
        RECT 5.955 -2.885 6.285 -2.555 ;
        RECT 5.96 -3.56 6.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 42.08 7.645 43.21 ;
        RECT 7.315 40.635 7.645 40.965 ;
        RECT 7.315 39.275 7.645 39.605 ;
        RECT 7.315 37.915 7.645 38.245 ;
        RECT 7.32 37.915 7.64 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 -1.525 7.645 -1.195 ;
        RECT 7.315 -2.885 7.645 -2.555 ;
        RECT 7.32 -3.56 7.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 -91.285 7.645 -90.955 ;
        RECT 7.315 -92.645 7.645 -92.315 ;
        RECT 7.315 -94.005 7.645 -93.675 ;
        RECT 7.315 -95.365 7.645 -95.035 ;
        RECT 7.315 -96.725 7.645 -96.395 ;
        RECT 7.315 -98.085 7.645 -97.755 ;
        RECT 7.315 -99.445 7.645 -99.115 ;
        RECT 7.315 -100.805 7.645 -100.475 ;
        RECT 7.315 -102.165 7.645 -101.835 ;
        RECT 7.315 -103.525 7.645 -103.195 ;
        RECT 7.315 -104.885 7.645 -104.555 ;
        RECT 7.315 -106.245 7.645 -105.915 ;
        RECT 7.315 -107.605 7.645 -107.275 ;
        RECT 7.315 -108.965 7.645 -108.635 ;
        RECT 7.315 -110.325 7.645 -109.995 ;
        RECT 7.315 -111.685 7.645 -111.355 ;
        RECT 7.315 -113.045 7.645 -112.715 ;
        RECT 7.315 -114.405 7.645 -114.075 ;
        RECT 7.315 -115.765 7.645 -115.435 ;
        RECT 7.315 -117.125 7.645 -116.795 ;
        RECT 7.315 -118.485 7.645 -118.155 ;
        RECT 7.315 -119.845 7.645 -119.515 ;
        RECT 7.315 -121.205 7.645 -120.875 ;
        RECT 7.315 -122.565 7.645 -122.235 ;
        RECT 7.315 -123.925 7.645 -123.595 ;
        RECT 7.315 -125.285 7.645 -124.955 ;
        RECT 7.315 -126.645 7.645 -126.315 ;
        RECT 7.315 -128.005 7.645 -127.675 ;
        RECT 7.315 -129.365 7.645 -129.035 ;
        RECT 7.315 -130.725 7.645 -130.395 ;
        RECT 7.315 -132.085 7.645 -131.755 ;
        RECT 7.315 -133.445 7.645 -133.115 ;
        RECT 7.315 -134.805 7.645 -134.475 ;
        RECT 7.315 -136.165 7.645 -135.835 ;
        RECT 7.315 -137.525 7.645 -137.195 ;
        RECT 7.315 -138.885 7.645 -138.555 ;
        RECT 7.315 -140.245 7.645 -139.915 ;
        RECT 7.315 -141.605 7.645 -141.275 ;
        RECT 7.315 -142.965 7.645 -142.635 ;
        RECT 7.315 -144.325 7.645 -143.995 ;
        RECT 7.315 -145.685 7.645 -145.355 ;
        RECT 7.315 -147.045 7.645 -146.715 ;
        RECT 7.315 -148.405 7.645 -148.075 ;
        RECT 7.315 -149.765 7.645 -149.435 ;
        RECT 7.315 -151.125 7.645 -150.795 ;
        RECT 7.315 -152.485 7.645 -152.155 ;
        RECT 7.315 -153.845 7.645 -153.515 ;
        RECT 7.315 -156.09 7.645 -154.96 ;
        RECT 7.32 -156.205 7.64 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 42.08 9.005 43.21 ;
        RECT 8.675 40.635 9.005 40.965 ;
        RECT 8.675 39.275 9.005 39.605 ;
        RECT 8.675 37.915 9.005 38.245 ;
        RECT 8.68 37.915 9 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 -95.365 9.005 -95.035 ;
        RECT 8.675 -96.725 9.005 -96.395 ;
        RECT 8.675 -98.085 9.005 -97.755 ;
        RECT 8.675 -99.445 9.005 -99.115 ;
        RECT 8.675 -100.805 9.005 -100.475 ;
        RECT 8.675 -102.165 9.005 -101.835 ;
        RECT 8.675 -103.525 9.005 -103.195 ;
        RECT 8.675 -104.885 9.005 -104.555 ;
        RECT 8.675 -106.245 9.005 -105.915 ;
        RECT 8.675 -107.605 9.005 -107.275 ;
        RECT 8.675 -108.965 9.005 -108.635 ;
        RECT 8.675 -110.325 9.005 -109.995 ;
        RECT 8.675 -111.685 9.005 -111.355 ;
        RECT 8.675 -113.045 9.005 -112.715 ;
        RECT 8.675 -114.405 9.005 -114.075 ;
        RECT 8.675 -115.765 9.005 -115.435 ;
        RECT 8.675 -117.125 9.005 -116.795 ;
        RECT 8.675 -118.485 9.005 -118.155 ;
        RECT 8.675 -119.845 9.005 -119.515 ;
        RECT 8.675 -121.205 9.005 -120.875 ;
        RECT 8.675 -122.565 9.005 -122.235 ;
        RECT 8.675 -123.925 9.005 -123.595 ;
        RECT 8.675 -125.285 9.005 -124.955 ;
        RECT 8.675 -126.645 9.005 -126.315 ;
        RECT 8.675 -128.005 9.005 -127.675 ;
        RECT 8.675 -129.365 9.005 -129.035 ;
        RECT 8.675 -130.725 9.005 -130.395 ;
        RECT 8.675 -132.085 9.005 -131.755 ;
        RECT 8.675 -133.445 9.005 -133.115 ;
        RECT 8.675 -134.805 9.005 -134.475 ;
        RECT 8.675 -136.165 9.005 -135.835 ;
        RECT 8.675 -137.525 9.005 -137.195 ;
        RECT 8.675 -138.885 9.005 -138.555 ;
        RECT 8.675 -140.245 9.005 -139.915 ;
        RECT 8.675 -141.605 9.005 -141.275 ;
        RECT 8.675 -142.965 9.005 -142.635 ;
        RECT 8.675 -144.325 9.005 -143.995 ;
        RECT 8.675 -145.685 9.005 -145.355 ;
        RECT 8.675 -147.045 9.005 -146.715 ;
        RECT 8.675 -148.405 9.005 -148.075 ;
        RECT 8.675 -149.765 9.005 -149.435 ;
        RECT 8.675 -151.125 9.005 -150.795 ;
        RECT 8.675 -152.485 9.005 -152.155 ;
        RECT 8.675 -153.845 9.005 -153.515 ;
        RECT 8.675 -156.09 9.005 -154.96 ;
        RECT 8.68 -156.205 9 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.41 -94.075 9.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 42.08 10.365 43.21 ;
        RECT 10.035 40.635 10.365 40.965 ;
        RECT 10.035 39.275 10.365 39.605 ;
        RECT 10.035 37.915 10.365 38.245 ;
        RECT 10.04 37.915 10.36 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 42.08 11.725 43.21 ;
        RECT 11.395 40.635 11.725 40.965 ;
        RECT 11.395 39.275 11.725 39.605 ;
        RECT 11.395 37.915 11.725 38.245 ;
        RECT 11.4 37.915 11.72 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 -1.525 11.725 -1.195 ;
        RECT 11.395 -2.885 11.725 -2.555 ;
        RECT 11.4 -3.56 11.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 42.08 13.085 43.21 ;
        RECT 12.755 40.635 13.085 40.965 ;
        RECT 12.755 39.275 13.085 39.605 ;
        RECT 12.755 37.915 13.085 38.245 ;
        RECT 12.76 37.915 13.08 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 -1.525 13.085 -1.195 ;
        RECT 12.755 -2.885 13.085 -2.555 ;
        RECT 12.76 -3.56 13.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 -91.285 13.085 -90.955 ;
        RECT 12.755 -92.645 13.085 -92.315 ;
        RECT 12.755 -94.005 13.085 -93.675 ;
        RECT 12.755 -95.365 13.085 -95.035 ;
        RECT 12.755 -96.725 13.085 -96.395 ;
        RECT 12.755 -98.085 13.085 -97.755 ;
        RECT 12.755 -99.445 13.085 -99.115 ;
        RECT 12.755 -100.805 13.085 -100.475 ;
        RECT 12.755 -102.165 13.085 -101.835 ;
        RECT 12.755 -103.525 13.085 -103.195 ;
        RECT 12.755 -104.885 13.085 -104.555 ;
        RECT 12.755 -106.245 13.085 -105.915 ;
        RECT 12.755 -107.605 13.085 -107.275 ;
        RECT 12.755 -108.965 13.085 -108.635 ;
        RECT 12.755 -110.325 13.085 -109.995 ;
        RECT 12.755 -111.685 13.085 -111.355 ;
        RECT 12.755 -113.045 13.085 -112.715 ;
        RECT 12.755 -114.405 13.085 -114.075 ;
        RECT 12.755 -115.765 13.085 -115.435 ;
        RECT 12.755 -117.125 13.085 -116.795 ;
        RECT 12.755 -118.485 13.085 -118.155 ;
        RECT 12.755 -119.845 13.085 -119.515 ;
        RECT 12.755 -121.205 13.085 -120.875 ;
        RECT 12.755 -122.565 13.085 -122.235 ;
        RECT 12.755 -123.925 13.085 -123.595 ;
        RECT 12.755 -125.285 13.085 -124.955 ;
        RECT 12.755 -126.645 13.085 -126.315 ;
        RECT 12.755 -128.005 13.085 -127.675 ;
        RECT 12.755 -129.365 13.085 -129.035 ;
        RECT 12.755 -130.725 13.085 -130.395 ;
        RECT 12.755 -132.085 13.085 -131.755 ;
        RECT 12.755 -133.445 13.085 -133.115 ;
        RECT 12.755 -134.805 13.085 -134.475 ;
        RECT 12.755 -136.165 13.085 -135.835 ;
        RECT 12.755 -137.525 13.085 -137.195 ;
        RECT 12.755 -138.885 13.085 -138.555 ;
        RECT 12.755 -140.245 13.085 -139.915 ;
        RECT 12.755 -141.605 13.085 -141.275 ;
        RECT 12.755 -142.965 13.085 -142.635 ;
        RECT 12.755 -144.325 13.085 -143.995 ;
        RECT 12.755 -145.685 13.085 -145.355 ;
        RECT 12.755 -147.045 13.085 -146.715 ;
        RECT 12.755 -148.405 13.085 -148.075 ;
        RECT 12.755 -149.765 13.085 -149.435 ;
        RECT 12.755 -151.125 13.085 -150.795 ;
        RECT 12.755 -152.485 13.085 -152.155 ;
        RECT 12.755 -153.845 13.085 -153.515 ;
        RECT 12.755 -156.09 13.085 -154.96 ;
        RECT 12.76 -156.205 13.08 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 42.08 14.445 43.21 ;
        RECT 14.115 40.635 14.445 40.965 ;
        RECT 14.115 39.275 14.445 39.605 ;
        RECT 14.115 37.915 14.445 38.245 ;
        RECT 14.12 37.915 14.44 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 -1.525 14.445 -1.195 ;
        RECT 14.115 -2.885 14.445 -2.555 ;
        RECT 14.12 -3.56 14.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 -91.285 14.445 -90.955 ;
        RECT 14.115 -92.645 14.445 -92.315 ;
        RECT 14.115 -94.005 14.445 -93.675 ;
        RECT 14.115 -95.365 14.445 -95.035 ;
        RECT 14.115 -96.725 14.445 -96.395 ;
        RECT 14.115 -98.085 14.445 -97.755 ;
        RECT 14.115 -99.445 14.445 -99.115 ;
        RECT 14.115 -100.805 14.445 -100.475 ;
        RECT 14.115 -102.165 14.445 -101.835 ;
        RECT 14.115 -103.525 14.445 -103.195 ;
        RECT 14.115 -104.885 14.445 -104.555 ;
        RECT 14.115 -106.245 14.445 -105.915 ;
        RECT 14.115 -107.605 14.445 -107.275 ;
        RECT 14.115 -108.965 14.445 -108.635 ;
        RECT 14.115 -110.325 14.445 -109.995 ;
        RECT 14.115 -111.685 14.445 -111.355 ;
        RECT 14.115 -113.045 14.445 -112.715 ;
        RECT 14.115 -114.405 14.445 -114.075 ;
        RECT 14.115 -115.765 14.445 -115.435 ;
        RECT 14.115 -117.125 14.445 -116.795 ;
        RECT 14.115 -118.485 14.445 -118.155 ;
        RECT 14.115 -119.845 14.445 -119.515 ;
        RECT 14.115 -121.205 14.445 -120.875 ;
        RECT 14.115 -122.565 14.445 -122.235 ;
        RECT 14.115 -123.925 14.445 -123.595 ;
        RECT 14.115 -125.285 14.445 -124.955 ;
        RECT 14.115 -126.645 14.445 -126.315 ;
        RECT 14.115 -128.005 14.445 -127.675 ;
        RECT 14.115 -129.365 14.445 -129.035 ;
        RECT 14.115 -130.725 14.445 -130.395 ;
        RECT 14.115 -132.085 14.445 -131.755 ;
        RECT 14.115 -133.445 14.445 -133.115 ;
        RECT 14.115 -134.805 14.445 -134.475 ;
        RECT 14.115 -136.165 14.445 -135.835 ;
        RECT 14.115 -137.525 14.445 -137.195 ;
        RECT 14.115 -138.885 14.445 -138.555 ;
        RECT 14.115 -140.245 14.445 -139.915 ;
        RECT 14.115 -141.605 14.445 -141.275 ;
        RECT 14.115 -142.965 14.445 -142.635 ;
        RECT 14.115 -144.325 14.445 -143.995 ;
        RECT 14.115 -145.685 14.445 -145.355 ;
        RECT 14.115 -147.045 14.445 -146.715 ;
        RECT 14.115 -148.405 14.445 -148.075 ;
        RECT 14.115 -149.765 14.445 -149.435 ;
        RECT 14.115 -151.125 14.445 -150.795 ;
        RECT 14.115 -152.485 14.445 -152.155 ;
        RECT 14.115 -153.845 14.445 -153.515 ;
        RECT 14.115 -156.09 14.445 -154.96 ;
        RECT 14.12 -156.205 14.44 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 42.08 15.805 43.21 ;
        RECT 15.475 40.635 15.805 40.965 ;
        RECT 15.475 39.275 15.805 39.605 ;
        RECT 15.475 37.915 15.805 38.245 ;
        RECT 15.48 37.915 15.8 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 -113.045 15.805 -112.715 ;
        RECT 15.475 -114.405 15.805 -114.075 ;
        RECT 15.475 -115.765 15.805 -115.435 ;
        RECT 15.475 -117.125 15.805 -116.795 ;
        RECT 15.475 -118.485 15.805 -118.155 ;
        RECT 15.475 -119.845 15.805 -119.515 ;
        RECT 15.475 -121.205 15.805 -120.875 ;
        RECT 15.475 -122.565 15.805 -122.235 ;
        RECT 15.475 -123.925 15.805 -123.595 ;
        RECT 15.475 -125.285 15.805 -124.955 ;
        RECT 15.475 -126.645 15.805 -126.315 ;
        RECT 15.475 -128.005 15.805 -127.675 ;
        RECT 15.475 -129.365 15.805 -129.035 ;
        RECT 15.475 -130.725 15.805 -130.395 ;
        RECT 15.475 -132.085 15.805 -131.755 ;
        RECT 15.475 -133.445 15.805 -133.115 ;
        RECT 15.475 -134.805 15.805 -134.475 ;
        RECT 15.475 -136.165 15.805 -135.835 ;
        RECT 15.475 -137.525 15.805 -137.195 ;
        RECT 15.475 -138.885 15.805 -138.555 ;
        RECT 15.475 -140.245 15.805 -139.915 ;
        RECT 15.475 -141.605 15.805 -141.275 ;
        RECT 15.475 -142.965 15.805 -142.635 ;
        RECT 15.475 -144.325 15.805 -143.995 ;
        RECT 15.475 -145.685 15.805 -145.355 ;
        RECT 15.475 -147.045 15.805 -146.715 ;
        RECT 15.475 -148.405 15.805 -148.075 ;
        RECT 15.475 -149.765 15.805 -149.435 ;
        RECT 15.475 -151.125 15.805 -150.795 ;
        RECT 15.475 -152.485 15.805 -152.155 ;
        RECT 15.475 -153.845 15.805 -153.515 ;
        RECT 15.475 -156.09 15.805 -154.96 ;
        RECT 15.48 -156.205 15.8 -95.035 ;
        RECT 15.475 -95.365 15.805 -95.035 ;
        RECT 15.475 -96.725 15.805 -96.395 ;
        RECT 15.475 -98.085 15.805 -97.755 ;
        RECT 15.475 -99.445 15.805 -99.115 ;
        RECT 15.475 -100.805 15.805 -100.475 ;
        RECT 15.475 -102.165 15.805 -101.835 ;
        RECT 15.475 -103.525 15.805 -103.195 ;
        RECT 15.475 -104.885 15.805 -104.555 ;
        RECT 15.475 -106.245 15.805 -105.915 ;
        RECT 15.475 -107.605 15.805 -107.275 ;
        RECT 15.475 -108.965 15.805 -108.635 ;
        RECT 15.475 -110.325 15.805 -109.995 ;
        RECT 15.475 -111.685 15.805 -111.355 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 42.08 -18.195 43.21 ;
        RECT -18.525 40.635 -18.195 40.965 ;
        RECT -18.525 39.275 -18.195 39.605 ;
        RECT -18.525 37.915 -18.195 38.245 ;
        RECT -18.525 36.555 -18.195 36.885 ;
        RECT -18.525 35.195 -18.195 35.525 ;
        RECT -18.525 33.835 -18.195 34.165 ;
        RECT -18.525 32.475 -18.195 32.805 ;
        RECT -18.525 31.115 -18.195 31.445 ;
        RECT -18.525 29.755 -18.195 30.085 ;
        RECT -18.525 28.395 -18.195 28.725 ;
        RECT -18.525 27.035 -18.195 27.365 ;
        RECT -18.525 25.675 -18.195 26.005 ;
        RECT -18.525 24.315 -18.195 24.645 ;
        RECT -18.525 22.955 -18.195 23.285 ;
        RECT -18.525 21.595 -18.195 21.925 ;
        RECT -18.525 20.235 -18.195 20.565 ;
        RECT -18.525 18.875 -18.195 19.205 ;
        RECT -18.525 17.515 -18.195 17.845 ;
        RECT -18.525 16.155 -18.195 16.485 ;
        RECT -18.525 14.795 -18.195 15.125 ;
        RECT -18.525 13.435 -18.195 13.765 ;
        RECT -18.525 12.075 -18.195 12.405 ;
        RECT -18.525 10.715 -18.195 11.045 ;
        RECT -18.525 9.355 -18.195 9.685 ;
        RECT -18.525 7.995 -18.195 8.325 ;
        RECT -18.525 6.635 -18.195 6.965 ;
        RECT -18.525 5.275 -18.195 5.605 ;
        RECT -18.525 3.915 -18.195 4.245 ;
        RECT -18.525 2.555 -18.195 2.885 ;
        RECT -18.525 -1.525 -18.195 -1.195 ;
        RECT -18.525 -2.885 -18.195 -2.555 ;
        RECT -18.525 -4.245 -18.195 -3.915 ;
        RECT -18.525 -6.965 -18.195 -6.635 ;
        RECT -18.525 -8.325 -18.195 -7.995 ;
        RECT -18.525 -9.87 -18.195 -9.54 ;
        RECT -18.525 -12.405 -18.195 -12.075 ;
        RECT -18.525 -13.765 -18.195 -13.435 ;
        RECT -18.525 -14.71 -18.195 -14.38 ;
        RECT -18.525 -16.485 -18.195 -16.155 ;
        RECT -18.525 -24.645 -18.195 -24.315 ;
        RECT -18.525 -26.005 -18.195 -25.675 ;
        RECT -18.525 -28.725 -18.195 -28.395 ;
        RECT -18.525 -30.085 -18.195 -29.755 ;
        RECT -18.525 -31.89 -18.195 -31.56 ;
        RECT -18.525 -35.525 -18.195 -35.195 ;
        RECT -18.525 -36.73 -18.195 -36.4 ;
        RECT -18.525 -38.245 -18.195 -37.915 ;
        RECT -18.525 -45.045 -18.195 -44.715 ;
        RECT -18.525 -46.405 -18.195 -46.075 ;
        RECT -18.525 -49.125 -18.195 -48.795 ;
        RECT -18.525 -50.485 -18.195 -50.155 ;
        RECT -18.525 -51.81 -18.195 -51.48 ;
        RECT -18.525 -53.205 -18.195 -52.875 ;
        RECT -18.525 -54.565 -18.195 -54.235 ;
        RECT -18.525 -57.285 -18.195 -56.955 ;
        RECT -18.525 -58.645 -18.195 -58.315 ;
        RECT -18.525 -60.35 -18.195 -60.02 ;
        RECT -18.525 -61.365 -18.195 -61.035 ;
        RECT -18.525 -64.085 -18.195 -63.755 ;
        RECT -18.525 -65.445 -18.195 -65.115 ;
        RECT -18.525 -66.805 -18.195 -66.475 ;
        RECT -18.525 -68.165 -18.195 -67.835 ;
        RECT -18.525 -69.525 -18.195 -69.195 ;
        RECT -18.525 -72.245 -18.195 -71.915 ;
        RECT -18.525 -73.99 -18.195 -73.66 ;
        RECT -18.525 -74.965 -18.195 -74.635 ;
        RECT -18.525 -76.325 -18.195 -75.995 ;
        RECT -18.525 -79.045 -18.195 -78.715 ;
        RECT -18.525 -80.405 -18.195 -80.075 ;
        RECT -18.525 -81.765 -18.195 -81.435 ;
        RECT -18.525 -82.53 -18.195 -82.2 ;
        RECT -18.525 -84.485 -18.195 -84.155 ;
        RECT -18.52 -87.88 -18.2 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 -149.765 -18.195 -149.435 ;
        RECT -18.525 -150.825 -18.195 -150.495 ;
        RECT -18.525 -152.485 -18.195 -152.155 ;
        RECT -18.525 -153.845 -18.195 -153.515 ;
        RECT -18.525 -156.09 -18.195 -154.96 ;
        RECT -18.52 -156.205 -18.2 -149.435 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 42.08 -16.835 43.21 ;
        RECT -17.165 40.635 -16.835 40.965 ;
        RECT -17.165 39.275 -16.835 39.605 ;
        RECT -17.165 37.915 -16.835 38.245 ;
        RECT -17.165 36.555 -16.835 36.885 ;
        RECT -17.165 35.195 -16.835 35.525 ;
        RECT -17.165 33.835 -16.835 34.165 ;
        RECT -17.165 32.475 -16.835 32.805 ;
        RECT -17.165 31.115 -16.835 31.445 ;
        RECT -17.165 29.755 -16.835 30.085 ;
        RECT -17.165 28.395 -16.835 28.725 ;
        RECT -17.165 27.035 -16.835 27.365 ;
        RECT -17.165 25.675 -16.835 26.005 ;
        RECT -17.165 24.315 -16.835 24.645 ;
        RECT -17.165 22.955 -16.835 23.285 ;
        RECT -17.165 21.595 -16.835 21.925 ;
        RECT -17.165 20.235 -16.835 20.565 ;
        RECT -17.165 18.875 -16.835 19.205 ;
        RECT -17.165 17.515 -16.835 17.845 ;
        RECT -17.165 16.155 -16.835 16.485 ;
        RECT -17.165 14.795 -16.835 15.125 ;
        RECT -17.165 13.435 -16.835 13.765 ;
        RECT -17.165 12.075 -16.835 12.405 ;
        RECT -17.165 10.715 -16.835 11.045 ;
        RECT -17.165 9.355 -16.835 9.685 ;
        RECT -17.165 7.995 -16.835 8.325 ;
        RECT -17.165 6.635 -16.835 6.965 ;
        RECT -17.165 5.275 -16.835 5.605 ;
        RECT -17.165 3.915 -16.835 4.245 ;
        RECT -17.165 2.555 -16.835 2.885 ;
        RECT -17.165 1.195 -16.835 1.525 ;
        RECT -17.165 -1.525 -16.835 -1.195 ;
        RECT -17.165 -2.885 -16.835 -2.555 ;
        RECT -17.165 -4.245 -16.835 -3.915 ;
        RECT -17.165 -6.965 -16.835 -6.635 ;
        RECT -17.165 -8.325 -16.835 -7.995 ;
        RECT -17.165 -9.87 -16.835 -9.54 ;
        RECT -17.165 -12.405 -16.835 -12.075 ;
        RECT -17.165 -13.765 -16.835 -13.435 ;
        RECT -17.165 -14.71 -16.835 -14.38 ;
        RECT -17.165 -16.485 -16.835 -16.155 ;
        RECT -17.165 -23.285 -16.835 -22.955 ;
        RECT -17.165 -24.645 -16.835 -24.315 ;
        RECT -17.165 -26.005 -16.835 -25.675 ;
        RECT -17.165 -28.725 -16.835 -28.395 ;
        RECT -17.165 -30.085 -16.835 -29.755 ;
        RECT -17.165 -31.89 -16.835 -31.56 ;
        RECT -17.165 -35.525 -16.835 -35.195 ;
        RECT -17.165 -36.73 -16.835 -36.4 ;
        RECT -17.165 -38.245 -16.835 -37.915 ;
        RECT -17.165 -46.405 -16.835 -46.075 ;
        RECT -17.165 -49.125 -16.835 -48.795 ;
        RECT -17.165 -50.485 -16.835 -50.155 ;
        RECT -17.165 -51.81 -16.835 -51.48 ;
        RECT -17.165 -53.205 -16.835 -52.875 ;
        RECT -17.165 -54.565 -16.835 -54.235 ;
        RECT -17.165 -57.285 -16.835 -56.955 ;
        RECT -17.165 -58.645 -16.835 -58.315 ;
        RECT -17.165 -60.35 -16.835 -60.02 ;
        RECT -17.165 -61.365 -16.835 -61.035 ;
        RECT -17.165 -64.085 -16.835 -63.755 ;
        RECT -17.165 -65.445 -16.835 -65.115 ;
        RECT -17.165 -66.805 -16.835 -66.475 ;
        RECT -17.165 -68.165 -16.835 -67.835 ;
        RECT -17.165 -69.525 -16.835 -69.195 ;
        RECT -17.165 -72.245 -16.835 -71.915 ;
        RECT -17.165 -73.99 -16.835 -73.66 ;
        RECT -17.165 -74.965 -16.835 -74.635 ;
        RECT -17.165 -79.045 -16.835 -78.715 ;
        RECT -17.165 -80.405 -16.835 -80.075 ;
        RECT -17.165 -81.765 -16.835 -81.435 ;
        RECT -17.165 -82.53 -16.835 -82.2 ;
        RECT -17.165 -84.485 -16.835 -84.155 ;
        RECT -17.16 -88.56 -16.84 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 -149.765 -16.835 -149.435 ;
        RECT -17.165 -150.825 -16.835 -150.495 ;
        RECT -17.165 -152.485 -16.835 -152.155 ;
        RECT -17.165 -153.845 -16.835 -153.515 ;
        RECT -17.165 -156.09 -16.835 -154.96 ;
        RECT -17.16 -156.205 -16.84 -147.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 42.08 -15.475 43.21 ;
        RECT -15.805 40.635 -15.475 40.965 ;
        RECT -15.805 39.275 -15.475 39.605 ;
        RECT -15.805 37.915 -15.475 38.245 ;
        RECT -15.805 36.555 -15.475 36.885 ;
        RECT -15.805 35.195 -15.475 35.525 ;
        RECT -15.805 33.835 -15.475 34.165 ;
        RECT -15.805 32.475 -15.475 32.805 ;
        RECT -15.805 31.115 -15.475 31.445 ;
        RECT -15.805 29.755 -15.475 30.085 ;
        RECT -15.805 28.395 -15.475 28.725 ;
        RECT -15.805 27.035 -15.475 27.365 ;
        RECT -15.805 25.675 -15.475 26.005 ;
        RECT -15.805 24.315 -15.475 24.645 ;
        RECT -15.805 22.955 -15.475 23.285 ;
        RECT -15.805 21.595 -15.475 21.925 ;
        RECT -15.805 20.235 -15.475 20.565 ;
        RECT -15.805 18.875 -15.475 19.205 ;
        RECT -15.805 17.515 -15.475 17.845 ;
        RECT -15.805 16.155 -15.475 16.485 ;
        RECT -15.805 14.795 -15.475 15.125 ;
        RECT -15.805 13.435 -15.475 13.765 ;
        RECT -15.805 12.075 -15.475 12.405 ;
        RECT -15.805 10.715 -15.475 11.045 ;
        RECT -15.805 9.355 -15.475 9.685 ;
        RECT -15.805 7.995 -15.475 8.325 ;
        RECT -15.805 6.635 -15.475 6.965 ;
        RECT -15.805 5.275 -15.475 5.605 ;
        RECT -15.805 3.915 -15.475 4.245 ;
        RECT -15.805 2.555 -15.475 2.885 ;
        RECT -15.805 1.195 -15.475 1.525 ;
        RECT -15.805 -1.525 -15.475 -1.195 ;
        RECT -15.805 -2.885 -15.475 -2.555 ;
        RECT -15.805 -4.245 -15.475 -3.915 ;
        RECT -15.805 -6.965 -15.475 -6.635 ;
        RECT -15.805 -8.325 -15.475 -7.995 ;
        RECT -15.805 -9.87 -15.475 -9.54 ;
        RECT -15.805 -12.405 -15.475 -12.075 ;
        RECT -15.805 -13.765 -15.475 -13.435 ;
        RECT -15.805 -14.71 -15.475 -14.38 ;
        RECT -15.805 -16.485 -15.475 -16.155 ;
        RECT -15.8 -17.16 -15.48 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 -21.925 -15.475 -21.595 ;
        RECT -15.805 -23.285 -15.475 -22.955 ;
        RECT -15.805 -24.645 -15.475 -24.315 ;
        RECT -15.805 -26.005 -15.475 -25.675 ;
        RECT -15.805 -28.725 -15.475 -28.395 ;
        RECT -15.805 -30.085 -15.475 -29.755 ;
        RECT -15.805 -31.89 -15.475 -31.56 ;
        RECT -15.805 -35.525 -15.475 -35.195 ;
        RECT -15.805 -36.73 -15.475 -36.4 ;
        RECT -15.805 -38.245 -15.475 -37.915 ;
        RECT -15.8 -39.6 -15.48 -21.595 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 -43.685 -15.475 -43.355 ;
        RECT -15.805 -46.405 -15.475 -46.075 ;
        RECT -15.805 -49.125 -15.475 -48.795 ;
        RECT -15.805 -50.485 -15.475 -50.155 ;
        RECT -15.805 -51.81 -15.475 -51.48 ;
        RECT -15.805 -53.205 -15.475 -52.875 ;
        RECT -15.805 -54.565 -15.475 -54.235 ;
        RECT -15.805 -57.285 -15.475 -56.955 ;
        RECT -15.805 -58.645 -15.475 -58.315 ;
        RECT -15.805 -60.35 -15.475 -60.02 ;
        RECT -15.805 -61.365 -15.475 -61.035 ;
        RECT -15.805 -64.085 -15.475 -63.755 ;
        RECT -15.805 -65.445 -15.475 -65.115 ;
        RECT -15.805 -66.805 -15.475 -66.475 ;
        RECT -15.805 -68.165 -15.475 -67.835 ;
        RECT -15.805 -69.525 -15.475 -69.195 ;
        RECT -15.805 -72.245 -15.475 -71.915 ;
        RECT -15.805 -73.99 -15.475 -73.66 ;
        RECT -15.805 -74.965 -15.475 -74.635 ;
        RECT -15.805 -79.045 -15.475 -78.715 ;
        RECT -15.805 -80.405 -15.475 -80.075 ;
        RECT -15.805 -81.765 -15.475 -81.435 ;
        RECT -15.805 -82.53 -15.475 -82.2 ;
        RECT -15.805 -84.485 -15.475 -84.155 ;
        RECT -15.8 -85.16 -15.48 -43.355 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 -89.925 -15.475 -89.595 ;
        RECT -15.805 -91.285 -15.475 -90.955 ;
        RECT -15.805 -92.645 -15.475 -92.315 ;
        RECT -15.805 -96.725 -15.475 -96.395 ;
        RECT -15.805 -100.805 -15.475 -100.475 ;
        RECT -15.805 -102.165 -15.475 -101.835 ;
        RECT -15.805 -111.685 -15.475 -111.355 ;
        RECT -15.805 -115.765 -15.475 -115.435 ;
        RECT -15.805 -125.285 -15.475 -124.955 ;
        RECT -15.805 -132.085 -15.475 -131.755 ;
        RECT -15.805 -133.445 -15.475 -133.115 ;
        RECT -15.805 -134.805 -15.475 -134.475 ;
        RECT -15.805 -136.165 -15.475 -135.835 ;
        RECT -15.805 -137.525 -15.475 -137.195 ;
        RECT -15.805 -138.885 -15.475 -138.555 ;
        RECT -15.805 -140.245 -15.475 -139.915 ;
        RECT -15.805 -141.605 -15.475 -141.275 ;
        RECT -15.805 -142.965 -15.475 -142.635 ;
        RECT -15.805 -145.685 -15.475 -145.355 ;
        RECT -15.805 -147.045 -15.475 -146.715 ;
        RECT -15.8 -147.045 -15.48 -89.595 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 42.08 -14.115 43.21 ;
        RECT -14.445 40.635 -14.115 40.965 ;
        RECT -14.445 39.275 -14.115 39.605 ;
        RECT -14.445 37.915 -14.115 38.245 ;
        RECT -14.445 36.555 -14.115 36.885 ;
        RECT -14.445 35.195 -14.115 35.525 ;
        RECT -14.445 33.835 -14.115 34.165 ;
        RECT -14.445 32.475 -14.115 32.805 ;
        RECT -14.445 31.115 -14.115 31.445 ;
        RECT -14.445 29.755 -14.115 30.085 ;
        RECT -14.445 28.395 -14.115 28.725 ;
        RECT -14.445 27.035 -14.115 27.365 ;
        RECT -14.445 25.675 -14.115 26.005 ;
        RECT -14.445 24.315 -14.115 24.645 ;
        RECT -14.445 22.955 -14.115 23.285 ;
        RECT -14.445 21.595 -14.115 21.925 ;
        RECT -14.445 20.235 -14.115 20.565 ;
        RECT -14.445 18.875 -14.115 19.205 ;
        RECT -14.445 17.515 -14.115 17.845 ;
        RECT -14.445 16.155 -14.115 16.485 ;
        RECT -14.445 14.795 -14.115 15.125 ;
        RECT -14.445 13.435 -14.115 13.765 ;
        RECT -14.445 12.075 -14.115 12.405 ;
        RECT -14.445 10.715 -14.115 11.045 ;
        RECT -14.445 9.355 -14.115 9.685 ;
        RECT -14.445 7.995 -14.115 8.325 ;
        RECT -14.445 6.635 -14.115 6.965 ;
        RECT -14.445 5.275 -14.115 5.605 ;
        RECT -14.445 3.915 -14.115 4.245 ;
        RECT -14.445 2.555 -14.115 2.885 ;
        RECT -14.445 1.195 -14.115 1.525 ;
        RECT -14.445 -1.525 -14.115 -1.195 ;
        RECT -14.445 -2.885 -14.115 -2.555 ;
        RECT -14.445 -4.245 -14.115 -3.915 ;
        RECT -14.445 -6.965 -14.115 -6.635 ;
        RECT -14.445 -8.325 -14.115 -7.995 ;
        RECT -14.445 -9.87 -14.115 -9.54 ;
        RECT -14.445 -12.405 -14.115 -12.075 ;
        RECT -14.445 -13.765 -14.115 -13.435 ;
        RECT -14.445 -14.71 -14.115 -14.38 ;
        RECT -14.445 -16.485 -14.115 -16.155 ;
        RECT -14.44 -16.485 -14.12 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 -21.925 -14.115 -21.595 ;
        RECT -14.445 -23.285 -14.115 -22.955 ;
        RECT -14.445 -24.645 -14.115 -24.315 ;
        RECT -14.445 -26.005 -14.115 -25.675 ;
        RECT -14.445 -28.725 -14.115 -28.395 ;
        RECT -14.445 -30.085 -14.115 -29.755 ;
        RECT -14.445 -31.89 -14.115 -31.56 ;
        RECT -14.445 -35.525 -14.115 -35.195 ;
        RECT -14.445 -36.73 -14.115 -36.4 ;
        RECT -14.445 -38.245 -14.115 -37.915 ;
        RECT -14.44 -38.245 -14.12 -20.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 -42.325 -14.115 -41.995 ;
        RECT -14.445 -43.685 -14.115 -43.355 ;
        RECT -14.445 -46.405 -14.115 -46.075 ;
        RECT -14.445 -49.125 -14.115 -48.795 ;
        RECT -14.445 -50.485 -14.115 -50.155 ;
        RECT -14.445 -51.81 -14.115 -51.48 ;
        RECT -14.445 -53.205 -14.115 -52.875 ;
        RECT -14.445 -54.565 -14.115 -54.235 ;
        RECT -14.445 -57.285 -14.115 -56.955 ;
        RECT -14.445 -58.645 -14.115 -58.315 ;
        RECT -14.445 -60.35 -14.115 -60.02 ;
        RECT -14.445 -61.365 -14.115 -61.035 ;
        RECT -14.445 -64.085 -14.115 -63.755 ;
        RECT -14.445 -65.445 -14.115 -65.115 ;
        RECT -14.445 -66.805 -14.115 -66.475 ;
        RECT -14.445 -68.165 -14.115 -67.835 ;
        RECT -14.445 -69.525 -14.115 -69.195 ;
        RECT -14.445 -72.245 -14.115 -71.915 ;
        RECT -14.445 -73.99 -14.115 -73.66 ;
        RECT -14.445 -74.965 -14.115 -74.635 ;
        RECT -14.445 -79.045 -14.115 -78.715 ;
        RECT -14.445 -80.405 -14.115 -80.075 ;
        RECT -14.445 -81.765 -14.115 -81.435 ;
        RECT -14.445 -82.53 -14.115 -82.2 ;
        RECT -14.445 -84.485 -14.115 -84.155 ;
        RECT -14.44 -84.485 -14.12 -41.995 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 -88.565 -14.115 -88.235 ;
        RECT -14.445 -89.925 -14.115 -89.595 ;
        RECT -14.445 -91.285 -14.115 -90.955 ;
        RECT -14.445 -92.645 -14.115 -92.315 ;
        RECT -14.445 -95.365 -14.115 -95.035 ;
        RECT -14.445 -96.725 -14.115 -96.395 ;
        RECT -14.445 -100.805 -14.115 -100.475 ;
        RECT -14.445 -106.245 -14.115 -105.915 ;
        RECT -14.445 -108.965 -14.115 -108.635 ;
        RECT -14.445 -111.685 -14.115 -111.355 ;
        RECT -14.445 -115.765 -14.115 -115.435 ;
        RECT -14.445 -117.125 -14.115 -116.795 ;
        RECT -14.445 -121.205 -14.115 -120.875 ;
        RECT -14.445 -122.565 -14.115 -122.235 ;
        RECT -14.445 -125.285 -14.115 -124.955 ;
        RECT -14.445 -129.365 -14.115 -129.035 ;
        RECT -14.445 -132.085 -14.115 -131.755 ;
        RECT -14.445 -133.445 -14.115 -133.115 ;
        RECT -14.445 -134.805 -14.115 -134.475 ;
        RECT -14.445 -136.165 -14.115 -135.835 ;
        RECT -14.445 -137.525 -14.115 -137.195 ;
        RECT -14.445 -138.885 -14.115 -138.555 ;
        RECT -14.445 -140.245 -14.115 -139.915 ;
        RECT -14.445 -141.605 -14.115 -141.275 ;
        RECT -14.44 -141.605 -14.12 -88.235 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 -148.405 -14.115 -148.075 ;
        RECT -14.445 -149.765 -14.115 -149.435 ;
        RECT -14.445 -150.825 -14.115 -150.495 ;
        RECT -14.445 -152.485 -14.115 -152.155 ;
        RECT -14.445 -153.845 -14.115 -153.515 ;
        RECT -14.445 -156.09 -14.115 -154.96 ;
        RECT -14.44 -156.205 -14.12 -147.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.085 42.08 -12.755 43.21 ;
        RECT -13.085 40.635 -12.755 40.965 ;
        RECT -13.085 39.275 -12.755 39.605 ;
        RECT -13.085 37.915 -12.755 38.245 ;
        RECT -13.085 36.555 -12.755 36.885 ;
        RECT -13.085 35.195 -12.755 35.525 ;
        RECT -13.085 33.835 -12.755 34.165 ;
        RECT -13.085 32.475 -12.755 32.805 ;
        RECT -13.085 31.115 -12.755 31.445 ;
        RECT -13.085 29.755 -12.755 30.085 ;
        RECT -13.085 28.395 -12.755 28.725 ;
        RECT -13.085 27.035 -12.755 27.365 ;
        RECT -13.085 25.675 -12.755 26.005 ;
        RECT -13.085 24.315 -12.755 24.645 ;
        RECT -13.085 22.955 -12.755 23.285 ;
        RECT -13.085 21.595 -12.755 21.925 ;
        RECT -13.085 20.235 -12.755 20.565 ;
        RECT -13.085 18.875 -12.755 19.205 ;
        RECT -13.085 17.515 -12.755 17.845 ;
        RECT -13.085 16.155 -12.755 16.485 ;
        RECT -13.085 14.795 -12.755 15.125 ;
        RECT -13.085 13.435 -12.755 13.765 ;
        RECT -13.085 12.075 -12.755 12.405 ;
        RECT -13.085 10.715 -12.755 11.045 ;
        RECT -13.085 9.355 -12.755 9.685 ;
        RECT -13.085 7.995 -12.755 8.325 ;
        RECT -13.085 6.635 -12.755 6.965 ;
        RECT -13.085 5.275 -12.755 5.605 ;
        RECT -13.085 3.915 -12.755 4.245 ;
        RECT -13.085 2.555 -12.755 2.885 ;
        RECT -13.085 1.195 -12.755 1.525 ;
        RECT -13.085 -0.165 -12.755 0.165 ;
        RECT -13.085 -1.525 -12.755 -1.195 ;
        RECT -13.085 -2.885 -12.755 -2.555 ;
        RECT -13.085 -4.245 -12.755 -3.915 ;
        RECT -13.085 -6.965 -12.755 -6.635 ;
        RECT -13.085 -8.325 -12.755 -7.995 ;
        RECT -13.085 -9.87 -12.755 -9.54 ;
        RECT -13.085 -12.405 -12.755 -12.075 ;
        RECT -13.085 -13.765 -12.755 -13.435 ;
        RECT -13.085 -14.71 -12.755 -14.38 ;
        RECT -13.085 -16.485 -12.755 -16.155 ;
        RECT -13.08 -19.2 -12.76 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.085 -84.485 -12.755 -84.155 ;
        RECT -13.085 -88.565 -12.755 -88.235 ;
        RECT -13.085 -89.925 -12.755 -89.595 ;
        RECT -13.085 -91.285 -12.755 -90.955 ;
        RECT -13.085 -92.645 -12.755 -92.315 ;
        RECT -13.085 -94.005 -12.755 -93.675 ;
        RECT -13.085 -95.365 -12.755 -95.035 ;
        RECT -13.085 -100.805 -12.755 -100.475 ;
        RECT -13.085 -106.245 -12.755 -105.915 ;
        RECT -13.085 -108.965 -12.755 -108.635 ;
        RECT -13.085 -111.685 -12.755 -111.355 ;
        RECT -13.085 -114.405 -12.755 -114.075 ;
        RECT -13.085 -115.765 -12.755 -115.435 ;
        RECT -13.085 -117.125 -12.755 -116.795 ;
        RECT -13.085 -121.205 -12.755 -120.875 ;
        RECT -13.085 -122.565 -12.755 -122.235 ;
        RECT -13.085 -123.925 -12.755 -123.595 ;
        RECT -13.085 -125.285 -12.755 -124.955 ;
        RECT -13.085 -128.005 -12.755 -127.675 ;
        RECT -13.085 -129.365 -12.755 -129.035 ;
        RECT -13.085 -130.725 -12.755 -130.395 ;
        RECT -13.085 -132.085 -12.755 -131.755 ;
        RECT -13.085 -134.805 -12.755 -134.475 ;
        RECT -13.085 -136.165 -12.755 -135.835 ;
        RECT -13.085 -137.525 -12.755 -137.195 ;
        RECT -13.085 -138.885 -12.755 -138.555 ;
        RECT -13.085 -140.245 -12.755 -139.915 ;
        RECT -13.085 -141.605 -12.755 -141.275 ;
        RECT -13.085 -145.685 -12.755 -145.355 ;
        RECT -13.085 -147.045 -12.755 -146.715 ;
        RECT -13.085 -148.405 -12.755 -148.075 ;
        RECT -13.085 -149.765 -12.755 -149.435 ;
        RECT -13.085 -150.825 -12.755 -150.495 ;
        RECT -13.085 -152.485 -12.755 -152.155 ;
        RECT -13.085 -153.845 -12.755 -153.515 ;
        RECT -13.085 -156.09 -12.755 -154.96 ;
        RECT -13.08 -156.205 -12.76 -84.155 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.725 42.08 -11.395 43.21 ;
        RECT -11.725 40.635 -11.395 40.965 ;
        RECT -11.725 39.275 -11.395 39.605 ;
        RECT -11.725 37.915 -11.395 38.245 ;
        RECT -11.725 36.555 -11.395 36.885 ;
        RECT -11.725 35.195 -11.395 35.525 ;
        RECT -11.725 33.835 -11.395 34.165 ;
        RECT -11.725 32.475 -11.395 32.805 ;
        RECT -11.725 31.115 -11.395 31.445 ;
        RECT -11.725 29.755 -11.395 30.085 ;
        RECT -11.725 28.395 -11.395 28.725 ;
        RECT -11.725 27.035 -11.395 27.365 ;
        RECT -11.725 25.675 -11.395 26.005 ;
        RECT -11.725 24.315 -11.395 24.645 ;
        RECT -11.725 22.955 -11.395 23.285 ;
        RECT -11.725 21.595 -11.395 21.925 ;
        RECT -11.725 20.235 -11.395 20.565 ;
        RECT -11.725 18.875 -11.395 19.205 ;
        RECT -11.725 17.515 -11.395 17.845 ;
        RECT -11.725 16.155 -11.395 16.485 ;
        RECT -11.725 14.795 -11.395 15.125 ;
        RECT -11.725 13.435 -11.395 13.765 ;
        RECT -11.725 12.075 -11.395 12.405 ;
        RECT -11.725 10.715 -11.395 11.045 ;
        RECT -11.725 9.355 -11.395 9.685 ;
        RECT -11.725 7.995 -11.395 8.325 ;
        RECT -11.725 6.635 -11.395 6.965 ;
        RECT -11.725 5.275 -11.395 5.605 ;
        RECT -11.725 3.915 -11.395 4.245 ;
        RECT -11.725 2.555 -11.395 2.885 ;
        RECT -11.725 1.195 -11.395 1.525 ;
        RECT -11.725 -0.165 -11.395 0.165 ;
        RECT -11.725 -1.525 -11.395 -1.195 ;
        RECT -11.725 -2.885 -11.395 -2.555 ;
        RECT -11.725 -4.245 -11.395 -3.915 ;
        RECT -11.725 -6.965 -11.395 -6.635 ;
        RECT -11.725 -8.325 -11.395 -7.995 ;
        RECT -11.725 -9.87 -11.395 -9.54 ;
        RECT -11.725 -12.405 -11.395 -12.075 ;
        RECT -11.725 -13.765 -11.395 -13.435 ;
        RECT -11.725 -14.71 -11.395 -14.38 ;
        RECT -11.725 -16.485 -11.395 -16.155 ;
        RECT -11.725 -21.925 -11.395 -21.595 ;
        RECT -11.725 -23.285 -11.395 -22.955 ;
        RECT -11.725 -24.645 -11.395 -24.315 ;
        RECT -11.725 -26.005 -11.395 -25.675 ;
        RECT -11.725 -28.725 -11.395 -28.395 ;
        RECT -11.725 -30.085 -11.395 -29.755 ;
        RECT -11.725 -31.89 -11.395 -31.56 ;
        RECT -11.725 -35.525 -11.395 -35.195 ;
        RECT -11.725 -36.73 -11.395 -36.4 ;
        RECT -11.725 -38.245 -11.395 -37.915 ;
        RECT -11.725 -42.325 -11.395 -41.995 ;
        RECT -11.725 -43.685 -11.395 -43.355 ;
        RECT -11.725 -46.405 -11.395 -46.075 ;
        RECT -11.725 -49.125 -11.395 -48.795 ;
        RECT -11.725 -50.485 -11.395 -50.155 ;
        RECT -11.725 -51.81 -11.395 -51.48 ;
        RECT -11.725 -53.205 -11.395 -52.875 ;
        RECT -11.725 -54.565 -11.395 -54.235 ;
        RECT -11.725 -57.285 -11.395 -56.955 ;
        RECT -11.725 -58.645 -11.395 -58.315 ;
        RECT -11.725 -60.35 -11.395 -60.02 ;
        RECT -11.725 -61.365 -11.395 -61.035 ;
        RECT -11.725 -64.085 -11.395 -63.755 ;
        RECT -11.725 -65.445 -11.395 -65.115 ;
        RECT -11.725 -66.805 -11.395 -66.475 ;
        RECT -11.725 -68.165 -11.395 -67.835 ;
        RECT -11.725 -69.525 -11.395 -69.195 ;
        RECT -11.725 -72.245 -11.395 -71.915 ;
        RECT -11.725 -73.99 -11.395 -73.66 ;
        RECT -11.725 -74.965 -11.395 -74.635 ;
        RECT -11.725 -79.045 -11.395 -78.715 ;
        RECT -11.725 -80.405 -11.395 -80.075 ;
        RECT -11.725 -82.53 -11.395 -82.2 ;
        RECT -11.725 -84.485 -11.395 -84.155 ;
        RECT -11.725 -88.565 -11.395 -88.235 ;
        RECT -11.725 -89.925 -11.395 -89.595 ;
        RECT -11.725 -91.285 -11.395 -90.955 ;
        RECT -11.725 -92.645 -11.395 -92.315 ;
        RECT -11.725 -94.005 -11.395 -93.675 ;
        RECT -11.725 -95.365 -11.395 -95.035 ;
        RECT -11.725 -100.805 -11.395 -100.475 ;
        RECT -11.725 -102.165 -11.395 -101.835 ;
        RECT -11.725 -104.885 -11.395 -104.555 ;
        RECT -11.725 -106.245 -11.395 -105.915 ;
        RECT -11.725 -108.965 -11.395 -108.635 ;
        RECT -11.725 -110.325 -11.395 -109.995 ;
        RECT -11.725 -111.685 -11.395 -111.355 ;
        RECT -11.725 -113.045 -11.395 -112.715 ;
        RECT -11.725 -114.405 -11.395 -114.075 ;
        RECT -11.725 -115.765 -11.395 -115.435 ;
        RECT -11.725 -117.125 -11.395 -116.795 ;
        RECT -11.725 -121.205 -11.395 -120.875 ;
        RECT -11.725 -122.565 -11.395 -122.235 ;
        RECT -11.725 -123.925 -11.395 -123.595 ;
        RECT -11.725 -125.285 -11.395 -124.955 ;
        RECT -11.725 -126.645 -11.395 -126.315 ;
        RECT -11.725 -128.005 -11.395 -127.675 ;
        RECT -11.725 -129.365 -11.395 -129.035 ;
        RECT -11.725 -130.725 -11.395 -130.395 ;
        RECT -11.725 -132.085 -11.395 -131.755 ;
        RECT -11.725 -134.805 -11.395 -134.475 ;
        RECT -11.725 -136.165 -11.395 -135.835 ;
        RECT -11.725 -137.525 -11.395 -137.195 ;
        RECT -11.725 -138.885 -11.395 -138.555 ;
        RECT -11.725 -140.245 -11.395 -139.915 ;
        RECT -11.725 -141.605 -11.395 -141.275 ;
        RECT -11.725 -145.685 -11.395 -145.355 ;
        RECT -11.725 -147.045 -11.395 -146.715 ;
        RECT -11.725 -149.765 -11.395 -149.435 ;
        RECT -11.725 -150.825 -11.395 -150.495 ;
        RECT -11.725 -152.485 -11.395 -152.155 ;
        RECT -11.725 -153.845 -11.395 -153.515 ;
        RECT -11.725 -156.09 -11.395 -154.96 ;
        RECT -11.72 -156.205 -11.4 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.365 42.08 -10.035 43.21 ;
        RECT -10.365 40.635 -10.035 40.965 ;
        RECT -10.365 39.275 -10.035 39.605 ;
        RECT -10.365 37.915 -10.035 38.245 ;
        RECT -10.365 36.555 -10.035 36.885 ;
        RECT -10.365 35.195 -10.035 35.525 ;
        RECT -10.365 33.835 -10.035 34.165 ;
        RECT -10.365 32.475 -10.035 32.805 ;
        RECT -10.365 28.395 -10.035 28.725 ;
        RECT -10.365 25.675 -10.035 26.005 ;
        RECT -10.365 18.875 -10.035 19.205 ;
        RECT -10.365 17.515 -10.035 17.845 ;
        RECT -10.365 14.795 -10.035 15.125 ;
        RECT -10.365 7.995 -10.035 8.325 ;
        RECT -10.365 5.275 -10.035 5.605 ;
        RECT -10.365 3.915 -10.035 4.245 ;
        RECT -10.365 2.555 -10.035 2.885 ;
        RECT -10.365 1.195 -10.035 1.525 ;
        RECT -10.365 -0.165 -10.035 0.165 ;
        RECT -10.365 -1.525 -10.035 -1.195 ;
        RECT -10.365 -2.885 -10.035 -2.555 ;
        RECT -10.365 -4.245 -10.035 -3.915 ;
        RECT -10.365 -6.965 -10.035 -6.635 ;
        RECT -10.365 -8.325 -10.035 -7.995 ;
        RECT -10.365 -12.405 -10.035 -12.075 ;
        RECT -10.365 -13.765 -10.035 -13.435 ;
        RECT -10.365 -16.485 -10.035 -16.155 ;
        RECT -10.365 -21.925 -10.035 -21.595 ;
        RECT -10.365 -23.285 -10.035 -22.955 ;
        RECT -10.365 -24.645 -10.035 -24.315 ;
        RECT -10.365 -26.005 -10.035 -25.675 ;
        RECT -10.365 -28.725 -10.035 -28.395 ;
        RECT -10.365 -30.085 -10.035 -29.755 ;
        RECT -10.365 -35.525 -10.035 -35.195 ;
        RECT -10.365 -38.245 -10.035 -37.915 ;
        RECT -10.365 -42.325 -10.035 -41.995 ;
        RECT -10.365 -43.685 -10.035 -43.355 ;
        RECT -10.365 -46.405 -10.035 -46.075 ;
        RECT -10.365 -49.125 -10.035 -48.795 ;
        RECT -10.365 -50.485 -10.035 -50.155 ;
        RECT -10.365 -53.205 -10.035 -52.875 ;
        RECT -10.365 -54.565 -10.035 -54.235 ;
        RECT -10.365 -57.285 -10.035 -56.955 ;
        RECT -10.365 -58.645 -10.035 -58.315 ;
        RECT -10.365 -61.365 -10.035 -61.035 ;
        RECT -10.365 -64.085 -10.035 -63.755 ;
        RECT -10.365 -65.445 -10.035 -65.115 ;
        RECT -10.365 -66.805 -10.035 -66.475 ;
        RECT -10.365 -68.165 -10.035 -67.835 ;
        RECT -10.365 -69.525 -10.035 -69.195 ;
        RECT -10.365 -72.245 -10.035 -71.915 ;
        RECT -10.365 -74.965 -10.035 -74.635 ;
        RECT -10.365 -79.045 -10.035 -78.715 ;
        RECT -10.365 -80.405 -10.035 -80.075 ;
        RECT -10.365 -84.485 -10.035 -84.155 ;
        RECT -10.365 -88.565 -10.035 -88.235 ;
        RECT -10.365 -89.925 -10.035 -89.595 ;
        RECT -10.365 -91.285 -10.035 -90.955 ;
        RECT -10.365 -92.645 -10.035 -92.315 ;
        RECT -10.365 -94.005 -10.035 -93.675 ;
        RECT -10.365 -95.365 -10.035 -95.035 ;
        RECT -10.365 -100.805 -10.035 -100.475 ;
        RECT -10.365 -102.165 -10.035 -101.835 ;
        RECT -10.365 -103.525 -10.035 -103.195 ;
        RECT -10.365 -104.885 -10.035 -104.555 ;
        RECT -10.365 -106.245 -10.035 -105.915 ;
        RECT -10.365 -108.965 -10.035 -108.635 ;
        RECT -10.365 -110.325 -10.035 -109.995 ;
        RECT -10.365 -111.685 -10.035 -111.355 ;
        RECT -10.365 -113.045 -10.035 -112.715 ;
        RECT -10.365 -114.405 -10.035 -114.075 ;
        RECT -10.365 -115.765 -10.035 -115.435 ;
        RECT -10.365 -117.125 -10.035 -116.795 ;
        RECT -10.365 -119.845 -10.035 -119.515 ;
        RECT -10.365 -121.205 -10.035 -120.875 ;
        RECT -10.365 -122.565 -10.035 -122.235 ;
        RECT -10.365 -123.925 -10.035 -123.595 ;
        RECT -10.365 -125.285 -10.035 -124.955 ;
        RECT -10.365 -126.645 -10.035 -126.315 ;
        RECT -10.365 -128.005 -10.035 -127.675 ;
        RECT -10.365 -129.365 -10.035 -129.035 ;
        RECT -10.365 -130.725 -10.035 -130.395 ;
        RECT -10.365 -132.085 -10.035 -131.755 ;
        RECT -10.365 -134.805 -10.035 -134.475 ;
        RECT -10.365 -136.165 -10.035 -135.835 ;
        RECT -10.365 -137.525 -10.035 -137.195 ;
        RECT -10.365 -138.885 -10.035 -138.555 ;
        RECT -10.365 -140.245 -10.035 -139.915 ;
        RECT -10.365 -141.605 -10.035 -141.275 ;
        RECT -10.365 -142.965 -10.035 -142.635 ;
        RECT -10.365 -145.685 -10.035 -145.355 ;
        RECT -10.365 -148.405 -10.035 -148.075 ;
        RECT -10.365 -149.765 -10.035 -149.435 ;
        RECT -10.365 -152.485 -10.035 -152.155 ;
        RECT -10.365 -153.845 -10.035 -153.515 ;
        RECT -10.365 -156.09 -10.035 -154.96 ;
        RECT -10.36 -156.205 -10.04 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.005 42.08 -8.675 43.21 ;
        RECT -9.005 40.635 -8.675 40.965 ;
        RECT -9.005 39.275 -8.675 39.605 ;
        RECT -9.005 37.915 -8.675 38.245 ;
        RECT -9.005 36.555 -8.675 36.885 ;
        RECT -9.005 35.195 -8.675 35.525 ;
        RECT -9.005 33.835 -8.675 34.165 ;
        RECT -9.005 32.475 -8.675 32.805 ;
        RECT -9.005 28.395 -8.675 28.725 ;
        RECT -9.005 25.675 -8.675 26.005 ;
        RECT -9.005 18.875 -8.675 19.205 ;
        RECT -9.005 17.515 -8.675 17.845 ;
        RECT -9.005 14.795 -8.675 15.125 ;
        RECT -9.005 7.995 -8.675 8.325 ;
        RECT -9.005 5.275 -8.675 5.605 ;
        RECT -9.005 3.915 -8.675 4.245 ;
        RECT -9.005 2.555 -8.675 2.885 ;
        RECT -9.005 1.195 -8.675 1.525 ;
        RECT -9.005 -0.165 -8.675 0.165 ;
        RECT -9.005 -1.525 -8.675 -1.195 ;
        RECT -9.005 -2.885 -8.675 -2.555 ;
        RECT -9.005 -4.245 -8.675 -3.915 ;
        RECT -9.005 -5.605 -8.675 -5.275 ;
        RECT -9.005 -6.965 -8.675 -6.635 ;
        RECT -9.005 -8.325 -8.675 -7.995 ;
        RECT -9 -8.325 -8.68 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.005 -98.085 -8.675 -97.755 ;
        RECT -9.005 -99.445 -8.675 -99.115 ;
        RECT -9.005 -100.805 -8.675 -100.475 ;
        RECT -9.005 -102.165 -8.675 -101.835 ;
        RECT -9.005 -103.525 -8.675 -103.195 ;
        RECT -9.005 -104.885 -8.675 -104.555 ;
        RECT -9.005 -106.245 -8.675 -105.915 ;
        RECT -9.005 -107.605 -8.675 -107.275 ;
        RECT -9.005 -108.965 -8.675 -108.635 ;
        RECT -9.005 -110.325 -8.675 -109.995 ;
        RECT -9.005 -111.685 -8.675 -111.355 ;
        RECT -9.005 -113.045 -8.675 -112.715 ;
        RECT -9.005 -114.405 -8.675 -114.075 ;
        RECT -9.005 -115.765 -8.675 -115.435 ;
        RECT -9.005 -117.125 -8.675 -116.795 ;
        RECT -9.005 -118.485 -8.675 -118.155 ;
        RECT -9.005 -119.845 -8.675 -119.515 ;
        RECT -9.005 -121.205 -8.675 -120.875 ;
        RECT -9.005 -122.565 -8.675 -122.235 ;
        RECT -9.005 -123.925 -8.675 -123.595 ;
        RECT -9.005 -125.285 -8.675 -124.955 ;
        RECT -9.005 -126.645 -8.675 -126.315 ;
        RECT -9.005 -128.005 -8.675 -127.675 ;
        RECT -9.005 -129.365 -8.675 -129.035 ;
        RECT -9.005 -130.725 -8.675 -130.395 ;
        RECT -9.005 -132.085 -8.675 -131.755 ;
        RECT -9.005 -133.445 -8.675 -133.115 ;
        RECT -9.005 -134.805 -8.675 -134.475 ;
        RECT -9.005 -136.165 -8.675 -135.835 ;
        RECT -9.005 -137.525 -8.675 -137.195 ;
        RECT -9.005 -138.885 -8.675 -138.555 ;
        RECT -9.005 -140.245 -8.675 -139.915 ;
        RECT -9.005 -141.605 -8.675 -141.275 ;
        RECT -9.005 -142.965 -8.675 -142.635 ;
        RECT -9.005 -144.325 -8.675 -143.995 ;
        RECT -9.005 -145.685 -8.675 -145.355 ;
        RECT -9.005 -147.045 -8.675 -146.715 ;
        RECT -9.005 -148.405 -8.675 -148.075 ;
        RECT -9.005 -149.765 -8.675 -149.435 ;
        RECT -9.005 -151.125 -8.675 -150.795 ;
        RECT -9.005 -152.485 -8.675 -152.155 ;
        RECT -9.005 -153.845 -8.675 -153.515 ;
        RECT -9.005 -156.09 -8.675 -154.96 ;
        RECT -9 -156.205 -8.68 -97.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.645 42.08 -7.315 43.21 ;
        RECT -7.645 40.635 -7.315 40.965 ;
        RECT -7.645 39.275 -7.315 39.605 ;
        RECT -7.645 37.915 -7.315 38.245 ;
        RECT -7.645 36.555 -7.315 36.885 ;
        RECT -7.645 35.195 -7.315 35.525 ;
        RECT -7.645 33.835 -7.315 34.165 ;
        RECT -7.645 32.475 -7.315 32.805 ;
        RECT -7.645 28.395 -7.315 28.725 ;
        RECT -7.645 25.675 -7.315 26.005 ;
        RECT -7.645 18.875 -7.315 19.205 ;
        RECT -7.645 17.515 -7.315 17.845 ;
        RECT -7.645 14.795 -7.315 15.125 ;
        RECT -7.645 7.995 -7.315 8.325 ;
        RECT -7.645 5.275 -7.315 5.605 ;
        RECT -7.645 3.915 -7.315 4.245 ;
        RECT -7.645 2.555 -7.315 2.885 ;
        RECT -7.645 1.195 -7.315 1.525 ;
        RECT -7.645 -0.165 -7.315 0.165 ;
        RECT -7.645 -1.525 -7.315 -1.195 ;
        RECT -7.645 -2.885 -7.315 -2.555 ;
        RECT -7.645 -4.245 -7.315 -3.915 ;
        RECT -7.645 -5.605 -7.315 -5.275 ;
        RECT -7.645 -6.965 -7.315 -6.635 ;
        RECT -7.645 -8.325 -7.315 -7.995 ;
        RECT -7.645 -9.685 -7.315 -9.355 ;
        RECT -7.645 -12.405 -7.315 -12.075 ;
        RECT -7.645 -13.765 -7.315 -13.435 ;
        RECT -7.645 -15.125 -7.315 -14.795 ;
        RECT -7.645 -16.485 -7.315 -16.155 ;
        RECT -7.645 -17.845 -7.315 -17.515 ;
        RECT -7.645 -21.925 -7.315 -21.595 ;
        RECT -7.645 -23.285 -7.315 -22.955 ;
        RECT -7.645 -24.645 -7.315 -24.315 ;
        RECT -7.645 -26.005 -7.315 -25.675 ;
        RECT -7.645 -27.365 -7.315 -27.035 ;
        RECT -7.645 -28.725 -7.315 -28.395 ;
        RECT -7.645 -30.085 -7.315 -29.755 ;
        RECT -7.645 -31.445 -7.315 -31.115 ;
        RECT -7.645 -34.165 -7.315 -33.835 ;
        RECT -7.645 -35.525 -7.315 -35.195 ;
        RECT -7.645 -36.885 -7.315 -36.555 ;
        RECT -7.645 -38.245 -7.315 -37.915 ;
        RECT -7.645 -40.965 -7.315 -40.635 ;
        RECT -7.645 -42.325 -7.315 -41.995 ;
        RECT -7.645 -43.685 -7.315 -43.355 ;
        RECT -7.645 -46.405 -7.315 -46.075 ;
        RECT -7.645 -47.765 -7.315 -47.435 ;
        RECT -7.645 -49.125 -7.315 -48.795 ;
        RECT -7.645 -50.485 -7.315 -50.155 ;
        RECT -7.645 -51.845 -7.315 -51.515 ;
        RECT -7.645 -53.205 -7.315 -52.875 ;
        RECT -7.645 -54.565 -7.315 -54.235 ;
        RECT -7.645 -55.925 -7.315 -55.595 ;
        RECT -7.645 -57.285 -7.315 -56.955 ;
        RECT -7.645 -58.645 -7.315 -58.315 ;
        RECT -7.645 -60.005 -7.315 -59.675 ;
        RECT -7.645 -61.365 -7.315 -61.035 ;
        RECT -7.645 -62.725 -7.315 -62.395 ;
        RECT -7.645 -64.085 -7.315 -63.755 ;
        RECT -7.645 -65.445 -7.315 -65.115 ;
        RECT -7.645 -66.805 -7.315 -66.475 ;
        RECT -7.645 -68.165 -7.315 -67.835 ;
        RECT -7.645 -69.525 -7.315 -69.195 ;
        RECT -7.645 -70.885 -7.315 -70.555 ;
        RECT -7.645 -72.245 -7.315 -71.915 ;
        RECT -7.645 -73.605 -7.315 -73.275 ;
        RECT -7.645 -74.965 -7.315 -74.635 ;
        RECT -7.645 -76.325 -7.315 -75.995 ;
        RECT -7.645 -77.685 -7.315 -77.355 ;
        RECT -7.645 -79.045 -7.315 -78.715 ;
        RECT -7.645 -80.405 -7.315 -80.075 ;
        RECT -7.645 -81.765 -7.315 -81.435 ;
        RECT -7.645 -83.125 -7.315 -82.795 ;
        RECT -7.645 -84.485 -7.315 -84.155 ;
        RECT -7.645 -85.845 -7.315 -85.515 ;
        RECT -7.645 -87.205 -7.315 -86.875 ;
        RECT -7.645 -88.565 -7.315 -88.235 ;
        RECT -7.645 -89.925 -7.315 -89.595 ;
        RECT -7.645 -91.285 -7.315 -90.955 ;
        RECT -7.645 -92.645 -7.315 -92.315 ;
        RECT -7.645 -94.005 -7.315 -93.675 ;
        RECT -7.645 -95.365 -7.315 -95.035 ;
        RECT -7.645 -96.725 -7.315 -96.395 ;
        RECT -7.645 -98.085 -7.315 -97.755 ;
        RECT -7.645 -99.445 -7.315 -99.115 ;
        RECT -7.645 -100.805 -7.315 -100.475 ;
        RECT -7.645 -102.165 -7.315 -101.835 ;
        RECT -7.645 -103.525 -7.315 -103.195 ;
        RECT -7.645 -104.885 -7.315 -104.555 ;
        RECT -7.645 -106.245 -7.315 -105.915 ;
        RECT -7.645 -107.605 -7.315 -107.275 ;
        RECT -7.645 -108.965 -7.315 -108.635 ;
        RECT -7.645 -110.325 -7.315 -109.995 ;
        RECT -7.645 -111.685 -7.315 -111.355 ;
        RECT -7.645 -113.045 -7.315 -112.715 ;
        RECT -7.645 -114.405 -7.315 -114.075 ;
        RECT -7.645 -115.765 -7.315 -115.435 ;
        RECT -7.645 -117.125 -7.315 -116.795 ;
        RECT -7.645 -118.485 -7.315 -118.155 ;
        RECT -7.645 -119.845 -7.315 -119.515 ;
        RECT -7.645 -121.205 -7.315 -120.875 ;
        RECT -7.645 -122.565 -7.315 -122.235 ;
        RECT -7.645 -123.925 -7.315 -123.595 ;
        RECT -7.645 -125.285 -7.315 -124.955 ;
        RECT -7.645 -126.645 -7.315 -126.315 ;
        RECT -7.645 -128.005 -7.315 -127.675 ;
        RECT -7.645 -129.365 -7.315 -129.035 ;
        RECT -7.645 -130.725 -7.315 -130.395 ;
        RECT -7.645 -132.085 -7.315 -131.755 ;
        RECT -7.645 -133.445 -7.315 -133.115 ;
        RECT -7.645 -134.805 -7.315 -134.475 ;
        RECT -7.645 -136.165 -7.315 -135.835 ;
        RECT -7.645 -137.525 -7.315 -137.195 ;
        RECT -7.645 -138.885 -7.315 -138.555 ;
        RECT -7.645 -140.245 -7.315 -139.915 ;
        RECT -7.645 -141.605 -7.315 -141.275 ;
        RECT -7.645 -142.965 -7.315 -142.635 ;
        RECT -7.645 -144.325 -7.315 -143.995 ;
        RECT -7.645 -145.685 -7.315 -145.355 ;
        RECT -7.645 -147.045 -7.315 -146.715 ;
        RECT -7.645 -148.405 -7.315 -148.075 ;
        RECT -7.645 -149.765 -7.315 -149.435 ;
        RECT -7.645 -151.125 -7.315 -150.795 ;
        RECT -7.645 -152.485 -7.315 -152.155 ;
        RECT -7.645 -153.845 -7.315 -153.515 ;
        RECT -7.645 -156.09 -7.315 -154.96 ;
        RECT -7.64 -156.205 -7.32 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.285 42.08 -5.955 43.21 ;
        RECT -6.285 40.635 -5.955 40.965 ;
        RECT -6.285 39.275 -5.955 39.605 ;
        RECT -6.285 37.915 -5.955 38.245 ;
        RECT -6.285 -1.525 -5.955 -1.195 ;
        RECT -6.285 -2.885 -5.955 -2.555 ;
        RECT -6.285 -4.245 -5.955 -3.915 ;
        RECT -6.285 -5.605 -5.955 -5.275 ;
        RECT -6.285 -6.965 -5.955 -6.635 ;
        RECT -6.285 -8.325 -5.955 -7.995 ;
        RECT -6.285 -9.685 -5.955 -9.355 ;
        RECT -6.285 -12.405 -5.955 -12.075 ;
        RECT -6.285 -13.765 -5.955 -13.435 ;
        RECT -6.285 -15.125 -5.955 -14.795 ;
        RECT -6.285 -16.485 -5.955 -16.155 ;
        RECT -6.285 -17.845 -5.955 -17.515 ;
        RECT -6.285 -21.925 -5.955 -21.595 ;
        RECT -6.285 -23.285 -5.955 -22.955 ;
        RECT -6.285 -24.645 -5.955 -24.315 ;
        RECT -6.285 -26.005 -5.955 -25.675 ;
        RECT -6.285 -27.365 -5.955 -27.035 ;
        RECT -6.285 -28.725 -5.955 -28.395 ;
        RECT -6.285 -30.085 -5.955 -29.755 ;
        RECT -6.285 -31.445 -5.955 -31.115 ;
        RECT -6.285 -34.165 -5.955 -33.835 ;
        RECT -6.285 -35.525 -5.955 -35.195 ;
        RECT -6.285 -36.885 -5.955 -36.555 ;
        RECT -6.285 -38.245 -5.955 -37.915 ;
        RECT -6.285 -40.965 -5.955 -40.635 ;
        RECT -6.285 -42.325 -5.955 -41.995 ;
        RECT -6.285 -43.685 -5.955 -43.355 ;
        RECT -6.285 -46.405 -5.955 -46.075 ;
        RECT -6.285 -47.765 -5.955 -47.435 ;
        RECT -6.285 -49.125 -5.955 -48.795 ;
        RECT -6.285 -50.485 -5.955 -50.155 ;
        RECT -6.285 -51.845 -5.955 -51.515 ;
        RECT -6.285 -53.205 -5.955 -52.875 ;
        RECT -6.285 -54.565 -5.955 -54.235 ;
        RECT -6.285 -55.925 -5.955 -55.595 ;
        RECT -6.285 -57.285 -5.955 -56.955 ;
        RECT -6.285 -58.645 -5.955 -58.315 ;
        RECT -6.285 -60.005 -5.955 -59.675 ;
        RECT -6.285 -61.365 -5.955 -61.035 ;
        RECT -6.285 -62.725 -5.955 -62.395 ;
        RECT -6.285 -64.085 -5.955 -63.755 ;
        RECT -6.285 -65.445 -5.955 -65.115 ;
        RECT -6.285 -66.805 -5.955 -66.475 ;
        RECT -6.285 -68.165 -5.955 -67.835 ;
        RECT -6.285 -69.525 -5.955 -69.195 ;
        RECT -6.285 -70.885 -5.955 -70.555 ;
        RECT -6.285 -72.245 -5.955 -71.915 ;
        RECT -6.285 -73.605 -5.955 -73.275 ;
        RECT -6.285 -74.965 -5.955 -74.635 ;
        RECT -6.285 -76.325 -5.955 -75.995 ;
        RECT -6.285 -77.685 -5.955 -77.355 ;
        RECT -6.285 -79.045 -5.955 -78.715 ;
        RECT -6.285 -80.405 -5.955 -80.075 ;
        RECT -6.285 -81.765 -5.955 -81.435 ;
        RECT -6.285 -83.125 -5.955 -82.795 ;
        RECT -6.285 -84.485 -5.955 -84.155 ;
        RECT -6.285 -85.845 -5.955 -85.515 ;
        RECT -6.285 -87.205 -5.955 -86.875 ;
        RECT -6.285 -88.565 -5.955 -88.235 ;
        RECT -6.285 -89.925 -5.955 -89.595 ;
        RECT -6.285 -91.285 -5.955 -90.955 ;
        RECT -6.285 -92.645 -5.955 -92.315 ;
        RECT -6.285 -94.005 -5.955 -93.675 ;
        RECT -6.285 -95.365 -5.955 -95.035 ;
        RECT -6.285 -96.725 -5.955 -96.395 ;
        RECT -6.285 -98.085 -5.955 -97.755 ;
        RECT -6.285 -99.445 -5.955 -99.115 ;
        RECT -6.285 -100.805 -5.955 -100.475 ;
        RECT -6.285 -102.165 -5.955 -101.835 ;
        RECT -6.285 -103.525 -5.955 -103.195 ;
        RECT -6.285 -104.885 -5.955 -104.555 ;
        RECT -6.285 -106.245 -5.955 -105.915 ;
        RECT -6.285 -107.605 -5.955 -107.275 ;
        RECT -6.285 -108.965 -5.955 -108.635 ;
        RECT -6.285 -110.325 -5.955 -109.995 ;
        RECT -6.285 -111.685 -5.955 -111.355 ;
        RECT -6.285 -113.045 -5.955 -112.715 ;
        RECT -6.285 -114.405 -5.955 -114.075 ;
        RECT -6.285 -115.765 -5.955 -115.435 ;
        RECT -6.285 -117.125 -5.955 -116.795 ;
        RECT -6.285 -118.485 -5.955 -118.155 ;
        RECT -6.285 -119.845 -5.955 -119.515 ;
        RECT -6.285 -121.205 -5.955 -120.875 ;
        RECT -6.285 -122.565 -5.955 -122.235 ;
        RECT -6.285 -123.925 -5.955 -123.595 ;
        RECT -6.285 -125.285 -5.955 -124.955 ;
        RECT -6.285 -126.645 -5.955 -126.315 ;
        RECT -6.285 -128.005 -5.955 -127.675 ;
        RECT -6.285 -129.365 -5.955 -129.035 ;
        RECT -6.285 -130.725 -5.955 -130.395 ;
        RECT -6.285 -132.085 -5.955 -131.755 ;
        RECT -6.285 -133.445 -5.955 -133.115 ;
        RECT -6.285 -134.805 -5.955 -134.475 ;
        RECT -6.285 -136.165 -5.955 -135.835 ;
        RECT -6.285 -137.525 -5.955 -137.195 ;
        RECT -6.285 -138.885 -5.955 -138.555 ;
        RECT -6.285 -140.245 -5.955 -139.915 ;
        RECT -6.285 -141.605 -5.955 -141.275 ;
        RECT -6.285 -142.965 -5.955 -142.635 ;
        RECT -6.285 -144.325 -5.955 -143.995 ;
        RECT -6.285 -145.685 -5.955 -145.355 ;
        RECT -6.285 -147.045 -5.955 -146.715 ;
        RECT -6.285 -148.405 -5.955 -148.075 ;
        RECT -6.285 -149.765 -5.955 -149.435 ;
        RECT -6.285 -151.125 -5.955 -150.795 ;
        RECT -6.285 -152.485 -5.955 -152.155 ;
        RECT -6.285 -153.845 -5.955 -153.515 ;
        RECT -6.285 -156.09 -5.955 -154.96 ;
        RECT -6.28 -156.205 -5.96 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.765 42.08 -30.435 43.21 ;
        RECT -30.765 40.635 -30.435 40.965 ;
        RECT -30.765 39.275 -30.435 39.605 ;
        RECT -30.765 37.915 -30.435 38.245 ;
        RECT -30.765 36.555 -30.435 36.885 ;
        RECT -30.765 35.195 -30.435 35.525 ;
        RECT -30.765 33.835 -30.435 34.165 ;
        RECT -30.765 32.475 -30.435 32.805 ;
        RECT -30.765 31.115 -30.435 31.445 ;
        RECT -30.765 29.755 -30.435 30.085 ;
        RECT -30.765 28.395 -30.435 28.725 ;
        RECT -30.765 27.035 -30.435 27.365 ;
        RECT -30.765 25.675 -30.435 26.005 ;
        RECT -30.765 24.315 -30.435 24.645 ;
        RECT -30.765 22.955 -30.435 23.285 ;
        RECT -30.765 21.595 -30.435 21.925 ;
        RECT -30.765 20.235 -30.435 20.565 ;
        RECT -30.765 18.875 -30.435 19.205 ;
        RECT -30.765 17.515 -30.435 17.845 ;
        RECT -30.765 16.155 -30.435 16.485 ;
        RECT -30.765 14.795 -30.435 15.125 ;
        RECT -30.765 13.435 -30.435 13.765 ;
        RECT -30.765 12.075 -30.435 12.405 ;
        RECT -30.765 10.715 -30.435 11.045 ;
        RECT -30.765 9.355 -30.435 9.685 ;
        RECT -30.765 7.995 -30.435 8.325 ;
        RECT -30.765 6.635 -30.435 6.965 ;
        RECT -30.765 5.275 -30.435 5.605 ;
        RECT -30.765 3.915 -30.435 4.245 ;
        RECT -30.765 2.555 -30.435 2.885 ;
        RECT -30.765 -1.525 -30.435 -1.195 ;
        RECT -30.765 -2.885 -30.435 -2.555 ;
        RECT -30.765 -4.245 -30.435 -3.915 ;
        RECT -30.765 -5.605 -30.435 -5.275 ;
        RECT -30.765 -6.965 -30.435 -6.635 ;
        RECT -30.765 -8.325 -30.435 -7.995 ;
        RECT -30.765 -9.685 -30.435 -9.355 ;
        RECT -30.765 -11.045 -30.435 -10.715 ;
        RECT -30.765 -12.405 -30.435 -12.075 ;
        RECT -30.765 -13.765 -30.435 -13.435 ;
        RECT -30.765 -15.125 -30.435 -14.795 ;
        RECT -30.765 -16.485 -30.435 -16.155 ;
        RECT -30.765 -17.845 -30.435 -17.515 ;
        RECT -30.765 -19.205 -30.435 -18.875 ;
        RECT -30.765 -24.645 -30.435 -24.315 ;
        RECT -30.765 -26.005 -30.435 -25.675 ;
        RECT -30.765 -27.365 -30.435 -27.035 ;
        RECT -30.765 -28.725 -30.435 -28.395 ;
        RECT -30.765 -30.085 -30.435 -29.755 ;
        RECT -30.765 -31.445 -30.435 -31.115 ;
        RECT -30.765 -32.805 -30.435 -32.475 ;
        RECT -30.765 -34.165 -30.435 -33.835 ;
        RECT -30.765 -35.525 -30.435 -35.195 ;
        RECT -30.765 -36.885 -30.435 -36.555 ;
        RECT -30.765 -38.245 -30.435 -37.915 ;
        RECT -30.765 -39.605 -30.435 -39.275 ;
        RECT -30.765 -40.965 -30.435 -40.635 ;
        RECT -30.765 -43.685 -30.435 -43.355 ;
        RECT -30.765 -45.045 -30.435 -44.715 ;
        RECT -30.765 -46.405 -30.435 -46.075 ;
        RECT -30.765 -47.765 -30.435 -47.435 ;
        RECT -30.765 -49.125 -30.435 -48.795 ;
        RECT -30.765 -50.485 -30.435 -50.155 ;
        RECT -30.765 -51.845 -30.435 -51.515 ;
        RECT -30.765 -53.205 -30.435 -52.875 ;
        RECT -30.765 -54.565 -30.435 -54.235 ;
        RECT -30.765 -55.925 -30.435 -55.595 ;
        RECT -30.765 -57.285 -30.435 -56.955 ;
        RECT -30.765 -58.645 -30.435 -58.315 ;
        RECT -30.765 -60.005 -30.435 -59.675 ;
        RECT -30.765 -61.365 -30.435 -61.035 ;
        RECT -30.765 -62.725 -30.435 -62.395 ;
        RECT -30.765 -64.085 -30.435 -63.755 ;
        RECT -30.765 -66.805 -30.435 -66.475 ;
        RECT -30.765 -68.165 -30.435 -67.835 ;
        RECT -30.765 -69.525 -30.435 -69.195 ;
        RECT -30.765 -70.885 -30.435 -70.555 ;
        RECT -30.765 -72.245 -30.435 -71.915 ;
        RECT -30.765 -73.83 -30.435 -73.5 ;
        RECT -30.765 -74.965 -30.435 -74.635 ;
        RECT -30.765 -77.685 -30.435 -77.355 ;
        RECT -30.765 -79.045 -30.435 -78.715 ;
        RECT -30.765 -80.405 -30.435 -80.075 ;
        RECT -30.765 -81.97 -30.435 -81.64 ;
        RECT -30.765 -83.125 -30.435 -82.795 ;
        RECT -30.765 -84.485 -30.435 -84.155 ;
        RECT -30.765 -85.845 -30.435 -85.515 ;
        RECT -30.765 -88.565 -30.435 -88.235 ;
        RECT -30.765 -89.925 -30.435 -89.595 ;
        RECT -30.765 -91.285 -30.435 -90.955 ;
        RECT -30.765 -92.645 -30.435 -92.315 ;
        RECT -30.765 -98.085 -30.435 -97.755 ;
        RECT -30.765 -99.445 -30.435 -99.115 ;
        RECT -30.765 -100.805 -30.435 -100.475 ;
        RECT -30.765 -102.165 -30.435 -101.835 ;
        RECT -30.765 -103.525 -30.435 -103.195 ;
        RECT -30.765 -104.885 -30.435 -104.555 ;
        RECT -30.765 -107.605 -30.435 -107.275 ;
        RECT -30.765 -108.965 -30.435 -108.635 ;
        RECT -30.765 -110.325 -30.435 -109.995 ;
        RECT -30.765 -111.685 -30.435 -111.355 ;
        RECT -30.765 -115.765 -30.435 -115.435 ;
        RECT -30.765 -117.125 -30.435 -116.795 ;
        RECT -30.765 -118.485 -30.435 -118.155 ;
        RECT -30.765 -119.845 -30.435 -119.515 ;
        RECT -30.765 -121.205 -30.435 -120.875 ;
        RECT -30.765 -122.565 -30.435 -122.235 ;
        RECT -30.765 -125.285 -30.435 -124.955 ;
        RECT -30.765 -126.645 -30.435 -126.315 ;
        RECT -30.765 -128.005 -30.435 -127.675 ;
        RECT -30.765 -132.085 -30.435 -131.755 ;
        RECT -30.765 -133.445 -30.435 -133.115 ;
        RECT -30.765 -134.805 -30.435 -134.475 ;
        RECT -30.765 -136.165 -30.435 -135.835 ;
        RECT -30.765 -137.525 -30.435 -137.195 ;
        RECT -30.765 -138.885 -30.435 -138.555 ;
        RECT -30.765 -140.245 -30.435 -139.915 ;
        RECT -30.765 -141.605 -30.435 -141.275 ;
        RECT -30.765 -142.965 -30.435 -142.635 ;
        RECT -30.765 -145.685 -30.435 -145.355 ;
        RECT -30.765 -147.045 -30.435 -146.715 ;
        RECT -30.765 -148.405 -30.435 -148.075 ;
        RECT -30.765 -149.765 -30.435 -149.435 ;
        RECT -30.765 -150.825 -30.435 -150.495 ;
        RECT -30.765 -152.485 -30.435 -152.155 ;
        RECT -30.765 -153.845 -30.435 -153.515 ;
        RECT -30.765 -156.09 -30.435 -154.96 ;
        RECT -30.76 -156.205 -30.44 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 42.08 -29.075 43.21 ;
        RECT -29.405 40.635 -29.075 40.965 ;
        RECT -29.405 39.275 -29.075 39.605 ;
        RECT -29.405 37.915 -29.075 38.245 ;
        RECT -29.405 36.555 -29.075 36.885 ;
        RECT -29.405 35.195 -29.075 35.525 ;
        RECT -29.405 33.835 -29.075 34.165 ;
        RECT -29.405 32.475 -29.075 32.805 ;
        RECT -29.405 31.115 -29.075 31.445 ;
        RECT -29.405 29.755 -29.075 30.085 ;
        RECT -29.405 28.395 -29.075 28.725 ;
        RECT -29.405 27.035 -29.075 27.365 ;
        RECT -29.405 25.675 -29.075 26.005 ;
        RECT -29.405 24.315 -29.075 24.645 ;
        RECT -29.405 22.955 -29.075 23.285 ;
        RECT -29.405 21.595 -29.075 21.925 ;
        RECT -29.405 20.235 -29.075 20.565 ;
        RECT -29.405 18.875 -29.075 19.205 ;
        RECT -29.405 17.515 -29.075 17.845 ;
        RECT -29.405 16.155 -29.075 16.485 ;
        RECT -29.405 14.795 -29.075 15.125 ;
        RECT -29.405 13.435 -29.075 13.765 ;
        RECT -29.405 12.075 -29.075 12.405 ;
        RECT -29.405 10.715 -29.075 11.045 ;
        RECT -29.405 9.355 -29.075 9.685 ;
        RECT -29.405 7.995 -29.075 8.325 ;
        RECT -29.405 6.635 -29.075 6.965 ;
        RECT -29.405 5.275 -29.075 5.605 ;
        RECT -29.405 3.915 -29.075 4.245 ;
        RECT -29.405 2.555 -29.075 2.885 ;
        RECT -29.405 -1.525 -29.075 -1.195 ;
        RECT -29.405 -2.885 -29.075 -2.555 ;
        RECT -29.405 -4.245 -29.075 -3.915 ;
        RECT -29.405 -5.605 -29.075 -5.275 ;
        RECT -29.405 -6.965 -29.075 -6.635 ;
        RECT -29.405 -8.325 -29.075 -7.995 ;
        RECT -29.405 -9.685 -29.075 -9.355 ;
        RECT -29.405 -11.045 -29.075 -10.715 ;
        RECT -29.405 -12.405 -29.075 -12.075 ;
        RECT -29.405 -13.765 -29.075 -13.435 ;
        RECT -29.405 -15.125 -29.075 -14.795 ;
        RECT -29.405 -16.485 -29.075 -16.155 ;
        RECT -29.405 -17.845 -29.075 -17.515 ;
        RECT -29.405 -19.205 -29.075 -18.875 ;
        RECT -29.405 -24.645 -29.075 -24.315 ;
        RECT -29.405 -26.005 -29.075 -25.675 ;
        RECT -29.405 -27.365 -29.075 -27.035 ;
        RECT -29.405 -28.725 -29.075 -28.395 ;
        RECT -29.405 -30.085 -29.075 -29.755 ;
        RECT -29.405 -31.445 -29.075 -31.115 ;
        RECT -29.405 -32.805 -29.075 -32.475 ;
        RECT -29.405 -34.165 -29.075 -33.835 ;
        RECT -29.405 -35.525 -29.075 -35.195 ;
        RECT -29.405 -36.885 -29.075 -36.555 ;
        RECT -29.405 -38.245 -29.075 -37.915 ;
        RECT -29.405 -39.605 -29.075 -39.275 ;
        RECT -29.405 -40.965 -29.075 -40.635 ;
        RECT -29.405 -45.045 -29.075 -44.715 ;
        RECT -29.405 -46.405 -29.075 -46.075 ;
        RECT -29.405 -47.765 -29.075 -47.435 ;
        RECT -29.405 -49.125 -29.075 -48.795 ;
        RECT -29.405 -50.485 -29.075 -50.155 ;
        RECT -29.405 -51.845 -29.075 -51.515 ;
        RECT -29.405 -53.205 -29.075 -52.875 ;
        RECT -29.405 -54.565 -29.075 -54.235 ;
        RECT -29.405 -55.925 -29.075 -55.595 ;
        RECT -29.405 -57.285 -29.075 -56.955 ;
        RECT -29.405 -58.645 -29.075 -58.315 ;
        RECT -29.405 -60.005 -29.075 -59.675 ;
        RECT -29.405 -61.365 -29.075 -61.035 ;
        RECT -29.405 -62.725 -29.075 -62.395 ;
        RECT -29.405 -64.085 -29.075 -63.755 ;
        RECT -29.405 -66.805 -29.075 -66.475 ;
        RECT -29.405 -68.165 -29.075 -67.835 ;
        RECT -29.405 -69.525 -29.075 -69.195 ;
        RECT -29.405 -70.885 -29.075 -70.555 ;
        RECT -29.405 -72.245 -29.075 -71.915 ;
        RECT -29.405 -73.83 -29.075 -73.5 ;
        RECT -29.405 -74.965 -29.075 -74.635 ;
        RECT -29.405 -77.685 -29.075 -77.355 ;
        RECT -29.405 -79.045 -29.075 -78.715 ;
        RECT -29.405 -80.405 -29.075 -80.075 ;
        RECT -29.405 -81.97 -29.075 -81.64 ;
        RECT -29.405 -83.125 -29.075 -82.795 ;
        RECT -29.405 -84.485 -29.075 -84.155 ;
        RECT -29.405 -85.845 -29.075 -85.515 ;
        RECT -29.4 -87.2 -29.08 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 -149.765 -29.075 -149.435 ;
        RECT -29.405 -150.825 -29.075 -150.495 ;
        RECT -29.405 -152.485 -29.075 -152.155 ;
        RECT -29.405 -153.845 -29.075 -153.515 ;
        RECT -29.405 -156.09 -29.075 -154.96 ;
        RECT -29.4 -156.205 -29.08 -147.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.045 42.08 -27.715 43.21 ;
        RECT -28.045 40.635 -27.715 40.965 ;
        RECT -28.045 39.275 -27.715 39.605 ;
        RECT -28.045 37.915 -27.715 38.245 ;
        RECT -28.045 36.555 -27.715 36.885 ;
        RECT -28.045 35.195 -27.715 35.525 ;
        RECT -28.045 33.835 -27.715 34.165 ;
        RECT -28.045 32.475 -27.715 32.805 ;
        RECT -28.045 31.115 -27.715 31.445 ;
        RECT -28.045 29.755 -27.715 30.085 ;
        RECT -28.045 28.395 -27.715 28.725 ;
        RECT -28.045 27.035 -27.715 27.365 ;
        RECT -28.045 25.675 -27.715 26.005 ;
        RECT -28.045 24.315 -27.715 24.645 ;
        RECT -28.045 22.955 -27.715 23.285 ;
        RECT -28.045 21.595 -27.715 21.925 ;
        RECT -28.045 20.235 -27.715 20.565 ;
        RECT -28.045 18.875 -27.715 19.205 ;
        RECT -28.045 17.515 -27.715 17.845 ;
        RECT -28.045 16.155 -27.715 16.485 ;
        RECT -28.045 14.795 -27.715 15.125 ;
        RECT -28.045 13.435 -27.715 13.765 ;
        RECT -28.045 12.075 -27.715 12.405 ;
        RECT -28.045 10.715 -27.715 11.045 ;
        RECT -28.045 9.355 -27.715 9.685 ;
        RECT -28.045 7.995 -27.715 8.325 ;
        RECT -28.045 6.635 -27.715 6.965 ;
        RECT -28.045 5.275 -27.715 5.605 ;
        RECT -28.045 3.915 -27.715 4.245 ;
        RECT -28.045 2.555 -27.715 2.885 ;
        RECT -28.045 -1.525 -27.715 -1.195 ;
        RECT -28.045 -2.885 -27.715 -2.555 ;
        RECT -28.045 -4.245 -27.715 -3.915 ;
        RECT -28.045 -5.605 -27.715 -5.275 ;
        RECT -28.045 -6.965 -27.715 -6.635 ;
        RECT -28.045 -8.325 -27.715 -7.995 ;
        RECT -28.045 -9.685 -27.715 -9.355 ;
        RECT -28.045 -11.045 -27.715 -10.715 ;
        RECT -28.045 -12.405 -27.715 -12.075 ;
        RECT -28.045 -13.765 -27.715 -13.435 ;
        RECT -28.045 -15.125 -27.715 -14.795 ;
        RECT -28.045 -16.485 -27.715 -16.155 ;
        RECT -28.045 -17.845 -27.715 -17.515 ;
        RECT -28.045 -19.205 -27.715 -18.875 ;
        RECT -28.045 -24.645 -27.715 -24.315 ;
        RECT -28.045 -26.005 -27.715 -25.675 ;
        RECT -28.045 -27.365 -27.715 -27.035 ;
        RECT -28.045 -28.725 -27.715 -28.395 ;
        RECT -28.045 -30.085 -27.715 -29.755 ;
        RECT -28.045 -31.445 -27.715 -31.115 ;
        RECT -28.045 -32.805 -27.715 -32.475 ;
        RECT -28.045 -34.165 -27.715 -33.835 ;
        RECT -28.045 -35.525 -27.715 -35.195 ;
        RECT -28.045 -36.885 -27.715 -36.555 ;
        RECT -28.045 -38.245 -27.715 -37.915 ;
        RECT -28.045 -39.605 -27.715 -39.275 ;
        RECT -28.045 -40.965 -27.715 -40.635 ;
        RECT -28.045 -45.045 -27.715 -44.715 ;
        RECT -28.045 -46.405 -27.715 -46.075 ;
        RECT -28.045 -47.765 -27.715 -47.435 ;
        RECT -28.045 -49.125 -27.715 -48.795 ;
        RECT -28.045 -50.485 -27.715 -50.155 ;
        RECT -28.045 -51.845 -27.715 -51.515 ;
        RECT -28.045 -53.205 -27.715 -52.875 ;
        RECT -28.045 -54.565 -27.715 -54.235 ;
        RECT -28.045 -55.925 -27.715 -55.595 ;
        RECT -28.045 -57.285 -27.715 -56.955 ;
        RECT -28.045 -58.645 -27.715 -58.315 ;
        RECT -28.045 -60.005 -27.715 -59.675 ;
        RECT -28.045 -61.365 -27.715 -61.035 ;
        RECT -28.045 -62.725 -27.715 -62.395 ;
        RECT -28.045 -64.085 -27.715 -63.755 ;
        RECT -28.045 -66.805 -27.715 -66.475 ;
        RECT -28.045 -68.165 -27.715 -67.835 ;
        RECT -28.045 -69.525 -27.715 -69.195 ;
        RECT -28.045 -70.885 -27.715 -70.555 ;
        RECT -28.045 -72.245 -27.715 -71.915 ;
        RECT -28.045 -73.83 -27.715 -73.5 ;
        RECT -28.045 -74.965 -27.715 -74.635 ;
        RECT -28.045 -77.685 -27.715 -77.355 ;
        RECT -28.045 -79.045 -27.715 -78.715 ;
        RECT -28.045 -80.405 -27.715 -80.075 ;
        RECT -28.045 -81.97 -27.715 -81.64 ;
        RECT -28.045 -83.125 -27.715 -82.795 ;
        RECT -28.045 -84.485 -27.715 -84.155 ;
        RECT -28.045 -85.845 -27.715 -85.515 ;
        RECT -28.045 -88.565 -27.715 -88.235 ;
        RECT -28.045 -89.925 -27.715 -89.595 ;
        RECT -28.045 -91.285 -27.715 -90.955 ;
        RECT -28.045 -92.645 -27.715 -92.315 ;
        RECT -28.045 -98.085 -27.715 -97.755 ;
        RECT -28.045 -100.805 -27.715 -100.475 ;
        RECT -28.045 -102.165 -27.715 -101.835 ;
        RECT -28.045 -103.525 -27.715 -103.195 ;
        RECT -28.045 -104.885 -27.715 -104.555 ;
        RECT -28.045 -107.605 -27.715 -107.275 ;
        RECT -28.045 -108.965 -27.715 -108.635 ;
        RECT -28.045 -110.325 -27.715 -109.995 ;
        RECT -28.045 -111.685 -27.715 -111.355 ;
        RECT -28.045 -115.765 -27.715 -115.435 ;
        RECT -28.045 -117.125 -27.715 -116.795 ;
        RECT -28.045 -118.485 -27.715 -118.155 ;
        RECT -28.045 -119.845 -27.715 -119.515 ;
        RECT -28.045 -121.205 -27.715 -120.875 ;
        RECT -28.045 -122.565 -27.715 -122.235 ;
        RECT -28.045 -126.645 -27.715 -126.315 ;
        RECT -28.045 -128.005 -27.715 -127.675 ;
        RECT -28.045 -132.085 -27.715 -131.755 ;
        RECT -28.045 -133.445 -27.715 -133.115 ;
        RECT -28.045 -134.805 -27.715 -134.475 ;
        RECT -28.045 -136.165 -27.715 -135.835 ;
        RECT -28.045 -137.525 -27.715 -137.195 ;
        RECT -28.045 -138.885 -27.715 -138.555 ;
        RECT -28.045 -140.245 -27.715 -139.915 ;
        RECT -28.045 -141.605 -27.715 -141.275 ;
        RECT -28.045 -142.965 -27.715 -142.635 ;
        RECT -28.045 -145.685 -27.715 -145.355 ;
        RECT -28.045 -147.045 -27.715 -146.715 ;
        RECT -28.04 -147.045 -27.72 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.685 42.08 -26.355 43.21 ;
        RECT -26.685 40.635 -26.355 40.965 ;
        RECT -26.685 39.275 -26.355 39.605 ;
        RECT -26.685 37.915 -26.355 38.245 ;
        RECT -26.685 36.555 -26.355 36.885 ;
        RECT -26.685 35.195 -26.355 35.525 ;
        RECT -26.685 33.835 -26.355 34.165 ;
        RECT -26.685 32.475 -26.355 32.805 ;
        RECT -26.685 31.115 -26.355 31.445 ;
        RECT -26.685 29.755 -26.355 30.085 ;
        RECT -26.685 28.395 -26.355 28.725 ;
        RECT -26.685 27.035 -26.355 27.365 ;
        RECT -26.685 25.675 -26.355 26.005 ;
        RECT -26.685 24.315 -26.355 24.645 ;
        RECT -26.685 22.955 -26.355 23.285 ;
        RECT -26.685 21.595 -26.355 21.925 ;
        RECT -26.685 20.235 -26.355 20.565 ;
        RECT -26.685 18.875 -26.355 19.205 ;
        RECT -26.685 17.515 -26.355 17.845 ;
        RECT -26.685 16.155 -26.355 16.485 ;
        RECT -26.685 14.795 -26.355 15.125 ;
        RECT -26.685 13.435 -26.355 13.765 ;
        RECT -26.685 12.075 -26.355 12.405 ;
        RECT -26.685 10.715 -26.355 11.045 ;
        RECT -26.685 9.355 -26.355 9.685 ;
        RECT -26.685 7.995 -26.355 8.325 ;
        RECT -26.685 6.635 -26.355 6.965 ;
        RECT -26.685 5.275 -26.355 5.605 ;
        RECT -26.685 3.915 -26.355 4.245 ;
        RECT -26.685 2.555 -26.355 2.885 ;
        RECT -26.685 -1.525 -26.355 -1.195 ;
        RECT -26.685 -2.885 -26.355 -2.555 ;
        RECT -26.685 -4.245 -26.355 -3.915 ;
        RECT -26.685 -5.605 -26.355 -5.275 ;
        RECT -26.685 -6.965 -26.355 -6.635 ;
        RECT -26.685 -8.325 -26.355 -7.995 ;
        RECT -26.685 -9.685 -26.355 -9.355 ;
        RECT -26.685 -11.045 -26.355 -10.715 ;
        RECT -26.685 -12.405 -26.355 -12.075 ;
        RECT -26.685 -13.765 -26.355 -13.435 ;
        RECT -26.685 -15.125 -26.355 -14.795 ;
        RECT -26.685 -16.485 -26.355 -16.155 ;
        RECT -26.685 -17.845 -26.355 -17.515 ;
        RECT -26.685 -19.205 -26.355 -18.875 ;
        RECT -26.685 -24.645 -26.355 -24.315 ;
        RECT -26.685 -26.005 -26.355 -25.675 ;
        RECT -26.685 -27.365 -26.355 -27.035 ;
        RECT -26.685 -28.725 -26.355 -28.395 ;
        RECT -26.685 -30.085 -26.355 -29.755 ;
        RECT -26.685 -31.445 -26.355 -31.115 ;
        RECT -26.685 -32.805 -26.355 -32.475 ;
        RECT -26.685 -34.165 -26.355 -33.835 ;
        RECT -26.685 -35.525 -26.355 -35.195 ;
        RECT -26.685 -36.885 -26.355 -36.555 ;
        RECT -26.685 -38.245 -26.355 -37.915 ;
        RECT -26.685 -39.605 -26.355 -39.275 ;
        RECT -26.685 -40.965 -26.355 -40.635 ;
        RECT -26.685 -45.045 -26.355 -44.715 ;
        RECT -26.685 -46.405 -26.355 -46.075 ;
        RECT -26.685 -47.765 -26.355 -47.435 ;
        RECT -26.685 -49.125 -26.355 -48.795 ;
        RECT -26.685 -50.485 -26.355 -50.155 ;
        RECT -26.685 -51.845 -26.355 -51.515 ;
        RECT -26.685 -53.205 -26.355 -52.875 ;
        RECT -26.685 -54.565 -26.355 -54.235 ;
        RECT -26.685 -55.925 -26.355 -55.595 ;
        RECT -26.685 -57.285 -26.355 -56.955 ;
        RECT -26.685 -58.645 -26.355 -58.315 ;
        RECT -26.685 -60.005 -26.355 -59.675 ;
        RECT -26.685 -61.365 -26.355 -61.035 ;
        RECT -26.685 -62.725 -26.355 -62.395 ;
        RECT -26.685 -64.085 -26.355 -63.755 ;
        RECT -26.685 -66.805 -26.355 -66.475 ;
        RECT -26.685 -68.165 -26.355 -67.835 ;
        RECT -26.685 -69.525 -26.355 -69.195 ;
        RECT -26.685 -70.885 -26.355 -70.555 ;
        RECT -26.685 -72.245 -26.355 -71.915 ;
        RECT -26.685 -74.965 -26.355 -74.635 ;
        RECT -26.685 -77.685 -26.355 -77.355 ;
        RECT -26.685 -79.045 -26.355 -78.715 ;
        RECT -26.685 -80.405 -26.355 -80.075 ;
        RECT -26.685 -83.125 -26.355 -82.795 ;
        RECT -26.685 -84.485 -26.355 -84.155 ;
        RECT -26.685 -85.845 -26.355 -85.515 ;
        RECT -26.685 -88.565 -26.355 -88.235 ;
        RECT -26.685 -89.925 -26.355 -89.595 ;
        RECT -26.685 -91.285 -26.355 -90.955 ;
        RECT -26.685 -92.645 -26.355 -92.315 ;
        RECT -26.685 -98.085 -26.355 -97.755 ;
        RECT -26.685 -100.805 -26.355 -100.475 ;
        RECT -26.685 -102.165 -26.355 -101.835 ;
        RECT -26.685 -103.525 -26.355 -103.195 ;
        RECT -26.685 -104.885 -26.355 -104.555 ;
        RECT -26.685 -110.325 -26.355 -109.995 ;
        RECT -26.685 -111.685 -26.355 -111.355 ;
        RECT -26.685 -115.765 -26.355 -115.435 ;
        RECT -26.685 -117.125 -26.355 -116.795 ;
        RECT -26.685 -118.485 -26.355 -118.155 ;
        RECT -26.685 -121.205 -26.355 -120.875 ;
        RECT -26.685 -122.565 -26.355 -122.235 ;
        RECT -26.685 -126.645 -26.355 -126.315 ;
        RECT -26.685 -128.005 -26.355 -127.675 ;
        RECT -26.685 -132.085 -26.355 -131.755 ;
        RECT -26.685 -133.445 -26.355 -133.115 ;
        RECT -26.685 -134.805 -26.355 -134.475 ;
        RECT -26.685 -136.165 -26.355 -135.835 ;
        RECT -26.685 -137.525 -26.355 -137.195 ;
        RECT -26.685 -138.885 -26.355 -138.555 ;
        RECT -26.685 -140.245 -26.355 -139.915 ;
        RECT -26.685 -141.605 -26.355 -141.275 ;
        RECT -26.68 -141.605 -26.36 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.685 -148.405 -26.355 -148.075 ;
        RECT -26.685 -149.765 -26.355 -149.435 ;
        RECT -26.685 -150.825 -26.355 -150.495 ;
        RECT -26.685 -152.485 -26.355 -152.155 ;
        RECT -26.685 -153.845 -26.355 -153.515 ;
        RECT -26.685 -156.09 -26.355 -154.96 ;
        RECT -26.68 -156.205 -26.36 -147.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.325 42.08 -24.995 43.21 ;
        RECT -25.325 40.635 -24.995 40.965 ;
        RECT -25.325 39.275 -24.995 39.605 ;
        RECT -25.325 37.915 -24.995 38.245 ;
        RECT -25.325 36.555 -24.995 36.885 ;
        RECT -25.325 35.195 -24.995 35.525 ;
        RECT -25.325 33.835 -24.995 34.165 ;
        RECT -25.325 32.475 -24.995 32.805 ;
        RECT -25.325 31.115 -24.995 31.445 ;
        RECT -25.325 29.755 -24.995 30.085 ;
        RECT -25.325 28.395 -24.995 28.725 ;
        RECT -25.325 27.035 -24.995 27.365 ;
        RECT -25.325 25.675 -24.995 26.005 ;
        RECT -25.325 24.315 -24.995 24.645 ;
        RECT -25.325 22.955 -24.995 23.285 ;
        RECT -25.325 21.595 -24.995 21.925 ;
        RECT -25.325 20.235 -24.995 20.565 ;
        RECT -25.325 18.875 -24.995 19.205 ;
        RECT -25.325 17.515 -24.995 17.845 ;
        RECT -25.325 16.155 -24.995 16.485 ;
        RECT -25.325 14.795 -24.995 15.125 ;
        RECT -25.325 13.435 -24.995 13.765 ;
        RECT -25.325 12.075 -24.995 12.405 ;
        RECT -25.325 10.715 -24.995 11.045 ;
        RECT -25.325 9.355 -24.995 9.685 ;
        RECT -25.325 7.995 -24.995 8.325 ;
        RECT -25.325 6.635 -24.995 6.965 ;
        RECT -25.325 5.275 -24.995 5.605 ;
        RECT -25.325 3.915 -24.995 4.245 ;
        RECT -25.325 2.555 -24.995 2.885 ;
        RECT -25.325 -1.525 -24.995 -1.195 ;
        RECT -25.325 -2.885 -24.995 -2.555 ;
        RECT -25.325 -4.245 -24.995 -3.915 ;
        RECT -25.325 -5.605 -24.995 -5.275 ;
        RECT -25.325 -6.965 -24.995 -6.635 ;
        RECT -25.325 -8.325 -24.995 -7.995 ;
        RECT -25.325 -9.685 -24.995 -9.355 ;
        RECT -25.325 -11.045 -24.995 -10.715 ;
        RECT -25.325 -12.405 -24.995 -12.075 ;
        RECT -25.325 -13.765 -24.995 -13.435 ;
        RECT -25.325 -15.125 -24.995 -14.795 ;
        RECT -25.325 -16.485 -24.995 -16.155 ;
        RECT -25.325 -17.845 -24.995 -17.515 ;
        RECT -25.325 -19.205 -24.995 -18.875 ;
        RECT -25.325 -24.645 -24.995 -24.315 ;
        RECT -25.325 -26.005 -24.995 -25.675 ;
        RECT -25.325 -27.365 -24.995 -27.035 ;
        RECT -25.325 -28.725 -24.995 -28.395 ;
        RECT -25.325 -30.085 -24.995 -29.755 ;
        RECT -25.325 -31.445 -24.995 -31.115 ;
        RECT -25.325 -32.805 -24.995 -32.475 ;
        RECT -25.325 -34.165 -24.995 -33.835 ;
        RECT -25.325 -35.525 -24.995 -35.195 ;
        RECT -25.325 -36.885 -24.995 -36.555 ;
        RECT -25.325 -38.245 -24.995 -37.915 ;
        RECT -25.325 -39.605 -24.995 -39.275 ;
        RECT -25.325 -40.965 -24.995 -40.635 ;
        RECT -25.325 -45.045 -24.995 -44.715 ;
        RECT -25.325 -46.405 -24.995 -46.075 ;
        RECT -25.325 -47.765 -24.995 -47.435 ;
        RECT -25.325 -49.125 -24.995 -48.795 ;
        RECT -25.325 -50.485 -24.995 -50.155 ;
        RECT -25.325 -51.845 -24.995 -51.515 ;
        RECT -25.325 -53.205 -24.995 -52.875 ;
        RECT -25.325 -54.565 -24.995 -54.235 ;
        RECT -25.325 -55.925 -24.995 -55.595 ;
        RECT -25.325 -57.285 -24.995 -56.955 ;
        RECT -25.325 -58.645 -24.995 -58.315 ;
        RECT -25.325 -60.005 -24.995 -59.675 ;
        RECT -25.325 -61.365 -24.995 -61.035 ;
        RECT -25.325 -62.725 -24.995 -62.395 ;
        RECT -25.325 -64.085 -24.995 -63.755 ;
        RECT -25.325 -65.445 -24.995 -65.115 ;
        RECT -25.325 -66.805 -24.995 -66.475 ;
        RECT -25.325 -68.165 -24.995 -67.835 ;
        RECT -25.325 -69.525 -24.995 -69.195 ;
        RECT -25.325 -70.885 -24.995 -70.555 ;
        RECT -25.325 -72.245 -24.995 -71.915 ;
        RECT -25.325 -73.605 -24.995 -73.275 ;
        RECT -25.325 -74.965 -24.995 -74.635 ;
        RECT -25.325 -76.325 -24.995 -75.995 ;
        RECT -25.325 -77.685 -24.995 -77.355 ;
        RECT -25.325 -79.045 -24.995 -78.715 ;
        RECT -25.325 -80.405 -24.995 -80.075 ;
        RECT -25.325 -81.765 -24.995 -81.435 ;
        RECT -25.325 -83.125 -24.995 -82.795 ;
        RECT -25.325 -84.485 -24.995 -84.155 ;
        RECT -25.325 -85.845 -24.995 -85.515 ;
        RECT -25.325 -87.205 -24.995 -86.875 ;
        RECT -25.325 -88.565 -24.995 -88.235 ;
        RECT -25.325 -89.925 -24.995 -89.595 ;
        RECT -25.325 -91.285 -24.995 -90.955 ;
        RECT -25.325 -92.645 -24.995 -92.315 ;
        RECT -25.325 -98.085 -24.995 -97.755 ;
        RECT -25.325 -99.445 -24.995 -99.115 ;
        RECT -25.325 -100.805 -24.995 -100.475 ;
        RECT -25.325 -102.165 -24.995 -101.835 ;
        RECT -25.325 -103.525 -24.995 -103.195 ;
        RECT -25.325 -104.885 -24.995 -104.555 ;
        RECT -25.325 -110.325 -24.995 -109.995 ;
        RECT -25.325 -111.685 -24.995 -111.355 ;
        RECT -25.325 -115.765 -24.995 -115.435 ;
        RECT -25.325 -117.125 -24.995 -116.795 ;
        RECT -25.325 -118.485 -24.995 -118.155 ;
        RECT -25.325 -121.205 -24.995 -120.875 ;
        RECT -25.325 -122.565 -24.995 -122.235 ;
        RECT -25.325 -126.645 -24.995 -126.315 ;
        RECT -25.325 -128.005 -24.995 -127.675 ;
        RECT -25.325 -132.085 -24.995 -131.755 ;
        RECT -25.325 -133.445 -24.995 -133.115 ;
        RECT -25.325 -134.805 -24.995 -134.475 ;
        RECT -25.325 -136.165 -24.995 -135.835 ;
        RECT -25.325 -137.525 -24.995 -137.195 ;
        RECT -25.325 -138.885 -24.995 -138.555 ;
        RECT -25.325 -140.245 -24.995 -139.915 ;
        RECT -25.325 -141.605 -24.995 -141.275 ;
        RECT -25.325 -142.965 -24.995 -142.635 ;
        RECT -25.325 -145.685 -24.995 -145.355 ;
        RECT -25.325 -147.045 -24.995 -146.715 ;
        RECT -25.325 -148.405 -24.995 -148.075 ;
        RECT -25.325 -149.765 -24.995 -149.435 ;
        RECT -25.325 -150.825 -24.995 -150.495 ;
        RECT -25.325 -152.485 -24.995 -152.155 ;
        RECT -25.325 -153.845 -24.995 -153.515 ;
        RECT -25.325 -156.09 -24.995 -154.96 ;
        RECT -25.32 -156.205 -25 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.965 42.08 -23.635 43.21 ;
        RECT -23.965 40.635 -23.635 40.965 ;
        RECT -23.965 39.275 -23.635 39.605 ;
        RECT -23.965 37.915 -23.635 38.245 ;
        RECT -23.965 36.555 -23.635 36.885 ;
        RECT -23.965 35.195 -23.635 35.525 ;
        RECT -23.965 33.835 -23.635 34.165 ;
        RECT -23.965 32.475 -23.635 32.805 ;
        RECT -23.965 31.115 -23.635 31.445 ;
        RECT -23.965 29.755 -23.635 30.085 ;
        RECT -23.965 28.395 -23.635 28.725 ;
        RECT -23.965 27.035 -23.635 27.365 ;
        RECT -23.965 25.675 -23.635 26.005 ;
        RECT -23.965 24.315 -23.635 24.645 ;
        RECT -23.965 22.955 -23.635 23.285 ;
        RECT -23.965 21.595 -23.635 21.925 ;
        RECT -23.965 20.235 -23.635 20.565 ;
        RECT -23.965 18.875 -23.635 19.205 ;
        RECT -23.965 17.515 -23.635 17.845 ;
        RECT -23.965 16.155 -23.635 16.485 ;
        RECT -23.965 14.795 -23.635 15.125 ;
        RECT -23.965 13.435 -23.635 13.765 ;
        RECT -23.965 12.075 -23.635 12.405 ;
        RECT -23.965 10.715 -23.635 11.045 ;
        RECT -23.965 9.355 -23.635 9.685 ;
        RECT -23.965 7.995 -23.635 8.325 ;
        RECT -23.965 6.635 -23.635 6.965 ;
        RECT -23.965 5.275 -23.635 5.605 ;
        RECT -23.965 3.915 -23.635 4.245 ;
        RECT -23.965 2.555 -23.635 2.885 ;
        RECT -23.965 -1.525 -23.635 -1.195 ;
        RECT -23.965 -2.885 -23.635 -2.555 ;
        RECT -23.965 -4.245 -23.635 -3.915 ;
        RECT -23.965 -5.605 -23.635 -5.275 ;
        RECT -23.965 -6.965 -23.635 -6.635 ;
        RECT -23.965 -8.325 -23.635 -7.995 ;
        RECT -23.965 -9.685 -23.635 -9.355 ;
        RECT -23.965 -11.045 -23.635 -10.715 ;
        RECT -23.965 -12.405 -23.635 -12.075 ;
        RECT -23.965 -13.765 -23.635 -13.435 ;
        RECT -23.965 -15.125 -23.635 -14.795 ;
        RECT -23.965 -16.485 -23.635 -16.155 ;
        RECT -23.965 -17.845 -23.635 -17.515 ;
        RECT -23.965 -19.205 -23.635 -18.875 ;
        RECT -23.965 -24.645 -23.635 -24.315 ;
        RECT -23.965 -26.005 -23.635 -25.675 ;
        RECT -23.965 -27.365 -23.635 -27.035 ;
        RECT -23.965 -28.725 -23.635 -28.395 ;
        RECT -23.965 -30.085 -23.635 -29.755 ;
        RECT -23.965 -31.445 -23.635 -31.115 ;
        RECT -23.965 -32.805 -23.635 -32.475 ;
        RECT -23.965 -34.165 -23.635 -33.835 ;
        RECT -23.965 -35.525 -23.635 -35.195 ;
        RECT -23.965 -36.885 -23.635 -36.555 ;
        RECT -23.965 -38.245 -23.635 -37.915 ;
        RECT -23.965 -39.605 -23.635 -39.275 ;
        RECT -23.965 -40.965 -23.635 -40.635 ;
        RECT -23.965 -45.045 -23.635 -44.715 ;
        RECT -23.965 -46.405 -23.635 -46.075 ;
        RECT -23.965 -47.765 -23.635 -47.435 ;
        RECT -23.965 -49.125 -23.635 -48.795 ;
        RECT -23.965 -50.485 -23.635 -50.155 ;
        RECT -23.965 -51.845 -23.635 -51.515 ;
        RECT -23.965 -53.205 -23.635 -52.875 ;
        RECT -23.965 -54.565 -23.635 -54.235 ;
        RECT -23.965 -55.925 -23.635 -55.595 ;
        RECT -23.965 -57.285 -23.635 -56.955 ;
        RECT -23.965 -58.645 -23.635 -58.315 ;
        RECT -23.965 -60.005 -23.635 -59.675 ;
        RECT -23.965 -61.365 -23.635 -61.035 ;
        RECT -23.965 -62.725 -23.635 -62.395 ;
        RECT -23.965 -64.085 -23.635 -63.755 ;
        RECT -23.965 -65.445 -23.635 -65.115 ;
        RECT -23.965 -66.805 -23.635 -66.475 ;
        RECT -23.965 -68.165 -23.635 -67.835 ;
        RECT -23.965 -69.525 -23.635 -69.195 ;
        RECT -23.965 -70.885 -23.635 -70.555 ;
        RECT -23.965 -72.245 -23.635 -71.915 ;
        RECT -23.965 -73.605 -23.635 -73.275 ;
        RECT -23.965 -74.965 -23.635 -74.635 ;
        RECT -23.965 -76.325 -23.635 -75.995 ;
        RECT -23.965 -77.685 -23.635 -77.355 ;
        RECT -23.965 -79.045 -23.635 -78.715 ;
        RECT -23.965 -80.405 -23.635 -80.075 ;
        RECT -23.965 -81.765 -23.635 -81.435 ;
        RECT -23.965 -83.125 -23.635 -82.795 ;
        RECT -23.965 -84.485 -23.635 -84.155 ;
        RECT -23.965 -85.845 -23.635 -85.515 ;
        RECT -23.965 -87.205 -23.635 -86.875 ;
        RECT -23.965 -88.565 -23.635 -88.235 ;
        RECT -23.965 -89.925 -23.635 -89.595 ;
        RECT -23.965 -91.285 -23.635 -90.955 ;
        RECT -23.965 -92.645 -23.635 -92.315 ;
        RECT -23.965 -98.085 -23.635 -97.755 ;
        RECT -23.965 -99.445 -23.635 -99.115 ;
        RECT -23.965 -100.805 -23.635 -100.475 ;
        RECT -23.965 -102.165 -23.635 -101.835 ;
        RECT -23.965 -104.885 -23.635 -104.555 ;
        RECT -23.965 -110.325 -23.635 -109.995 ;
        RECT -23.965 -111.685 -23.635 -111.355 ;
        RECT -23.965 -115.765 -23.635 -115.435 ;
        RECT -23.965 -117.125 -23.635 -116.795 ;
        RECT -23.965 -121.205 -23.635 -120.875 ;
        RECT -23.965 -122.565 -23.635 -122.235 ;
        RECT -23.965 -126.645 -23.635 -126.315 ;
        RECT -23.965 -128.005 -23.635 -127.675 ;
        RECT -23.965 -133.445 -23.635 -133.115 ;
        RECT -23.965 -134.805 -23.635 -134.475 ;
        RECT -23.965 -136.165 -23.635 -135.835 ;
        RECT -23.965 -137.525 -23.635 -137.195 ;
        RECT -23.965 -138.885 -23.635 -138.555 ;
        RECT -23.965 -140.245 -23.635 -139.915 ;
        RECT -23.965 -141.605 -23.635 -141.275 ;
        RECT -23.965 -142.965 -23.635 -142.635 ;
        RECT -23.965 -145.685 -23.635 -145.355 ;
        RECT -23.965 -147.045 -23.635 -146.715 ;
        RECT -23.965 -149.765 -23.635 -149.435 ;
        RECT -23.965 -150.825 -23.635 -150.495 ;
        RECT -23.965 -152.485 -23.635 -152.155 ;
        RECT -23.965 -153.845 -23.635 -153.515 ;
        RECT -23.965 -156.09 -23.635 -154.96 ;
        RECT -23.96 -156.205 -23.64 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.605 42.08 -22.275 43.21 ;
        RECT -22.605 40.635 -22.275 40.965 ;
        RECT -22.605 39.275 -22.275 39.605 ;
        RECT -22.605 37.915 -22.275 38.245 ;
        RECT -22.605 36.555 -22.275 36.885 ;
        RECT -22.605 35.195 -22.275 35.525 ;
        RECT -22.605 33.835 -22.275 34.165 ;
        RECT -22.605 32.475 -22.275 32.805 ;
        RECT -22.605 31.115 -22.275 31.445 ;
        RECT -22.605 29.755 -22.275 30.085 ;
        RECT -22.605 28.395 -22.275 28.725 ;
        RECT -22.605 27.035 -22.275 27.365 ;
        RECT -22.605 25.675 -22.275 26.005 ;
        RECT -22.605 24.315 -22.275 24.645 ;
        RECT -22.605 22.955 -22.275 23.285 ;
        RECT -22.605 21.595 -22.275 21.925 ;
        RECT -22.605 20.235 -22.275 20.565 ;
        RECT -22.605 18.875 -22.275 19.205 ;
        RECT -22.605 17.515 -22.275 17.845 ;
        RECT -22.605 16.155 -22.275 16.485 ;
        RECT -22.605 14.795 -22.275 15.125 ;
        RECT -22.605 13.435 -22.275 13.765 ;
        RECT -22.605 12.075 -22.275 12.405 ;
        RECT -22.605 10.715 -22.275 11.045 ;
        RECT -22.605 9.355 -22.275 9.685 ;
        RECT -22.605 7.995 -22.275 8.325 ;
        RECT -22.605 6.635 -22.275 6.965 ;
        RECT -22.605 5.275 -22.275 5.605 ;
        RECT -22.605 3.915 -22.275 4.245 ;
        RECT -22.605 2.555 -22.275 2.885 ;
        RECT -22.605 -1.525 -22.275 -1.195 ;
        RECT -22.605 -2.885 -22.275 -2.555 ;
        RECT -22.605 -4.245 -22.275 -3.915 ;
        RECT -22.605 -5.605 -22.275 -5.275 ;
        RECT -22.605 -6.965 -22.275 -6.635 ;
        RECT -22.605 -8.325 -22.275 -7.995 ;
        RECT -22.605 -9.685 -22.275 -9.355 ;
        RECT -22.605 -11.045 -22.275 -10.715 ;
        RECT -22.605 -12.405 -22.275 -12.075 ;
        RECT -22.605 -13.765 -22.275 -13.435 ;
        RECT -22.605 -15.125 -22.275 -14.795 ;
        RECT -22.605 -16.485 -22.275 -16.155 ;
        RECT -22.605 -17.845 -22.275 -17.515 ;
        RECT -22.605 -19.205 -22.275 -18.875 ;
        RECT -22.605 -24.645 -22.275 -24.315 ;
        RECT -22.605 -26.005 -22.275 -25.675 ;
        RECT -22.605 -27.365 -22.275 -27.035 ;
        RECT -22.605 -28.725 -22.275 -28.395 ;
        RECT -22.605 -30.085 -22.275 -29.755 ;
        RECT -22.605 -31.445 -22.275 -31.115 ;
        RECT -22.605 -32.805 -22.275 -32.475 ;
        RECT -22.605 -34.165 -22.275 -33.835 ;
        RECT -22.605 -35.525 -22.275 -35.195 ;
        RECT -22.605 -36.885 -22.275 -36.555 ;
        RECT -22.605 -38.245 -22.275 -37.915 ;
        RECT -22.605 -39.605 -22.275 -39.275 ;
        RECT -22.605 -40.965 -22.275 -40.635 ;
        RECT -22.605 -45.045 -22.275 -44.715 ;
        RECT -22.605 -46.405 -22.275 -46.075 ;
        RECT -22.605 -47.765 -22.275 -47.435 ;
        RECT -22.605 -49.125 -22.275 -48.795 ;
        RECT -22.605 -50.485 -22.275 -50.155 ;
        RECT -22.605 -51.845 -22.275 -51.515 ;
        RECT -22.605 -53.205 -22.275 -52.875 ;
        RECT -22.605 -54.565 -22.275 -54.235 ;
        RECT -22.605 -55.925 -22.275 -55.595 ;
        RECT -22.605 -57.285 -22.275 -56.955 ;
        RECT -22.605 -58.645 -22.275 -58.315 ;
        RECT -22.605 -60.005 -22.275 -59.675 ;
        RECT -22.605 -61.365 -22.275 -61.035 ;
        RECT -22.605 -62.725 -22.275 -62.395 ;
        RECT -22.605 -64.085 -22.275 -63.755 ;
        RECT -22.605 -65.445 -22.275 -65.115 ;
        RECT -22.605 -66.805 -22.275 -66.475 ;
        RECT -22.605 -68.165 -22.275 -67.835 ;
        RECT -22.605 -69.525 -22.275 -69.195 ;
        RECT -22.605 -70.885 -22.275 -70.555 ;
        RECT -22.605 -72.245 -22.275 -71.915 ;
        RECT -22.605 -73.605 -22.275 -73.275 ;
        RECT -22.605 -74.965 -22.275 -74.635 ;
        RECT -22.605 -76.325 -22.275 -75.995 ;
        RECT -22.605 -77.685 -22.275 -77.355 ;
        RECT -22.605 -79.045 -22.275 -78.715 ;
        RECT -22.605 -80.405 -22.275 -80.075 ;
        RECT -22.605 -81.765 -22.275 -81.435 ;
        RECT -22.605 -83.125 -22.275 -82.795 ;
        RECT -22.605 -84.485 -22.275 -84.155 ;
        RECT -22.605 -85.845 -22.275 -85.515 ;
        RECT -22.605 -87.205 -22.275 -86.875 ;
        RECT -22.605 -88.565 -22.275 -88.235 ;
        RECT -22.605 -89.925 -22.275 -89.595 ;
        RECT -22.605 -91.285 -22.275 -90.955 ;
        RECT -22.605 -92.645 -22.275 -92.315 ;
        RECT -22.605 -98.085 -22.275 -97.755 ;
        RECT -22.605 -99.445 -22.275 -99.115 ;
        RECT -22.605 -100.805 -22.275 -100.475 ;
        RECT -22.605 -102.165 -22.275 -101.835 ;
        RECT -22.605 -104.885 -22.275 -104.555 ;
        RECT -22.605 -110.325 -22.275 -109.995 ;
        RECT -22.605 -111.685 -22.275 -111.355 ;
        RECT -22.605 -115.765 -22.275 -115.435 ;
        RECT -22.605 -117.125 -22.275 -116.795 ;
        RECT -22.605 -118.485 -22.275 -118.155 ;
        RECT -22.605 -121.205 -22.275 -120.875 ;
        RECT -22.605 -122.565 -22.275 -122.235 ;
        RECT -22.605 -126.645 -22.275 -126.315 ;
        RECT -22.605 -128.005 -22.275 -127.675 ;
        RECT -22.605 -133.445 -22.275 -133.115 ;
        RECT -22.605 -134.805 -22.275 -134.475 ;
        RECT -22.605 -136.165 -22.275 -135.835 ;
        RECT -22.605 -137.525 -22.275 -137.195 ;
        RECT -22.605 -138.885 -22.275 -138.555 ;
        RECT -22.605 -140.245 -22.275 -139.915 ;
        RECT -22.605 -141.605 -22.275 -141.275 ;
        RECT -22.605 -142.965 -22.275 -142.635 ;
        RECT -22.605 -145.685 -22.275 -145.355 ;
        RECT -22.605 -149.765 -22.275 -149.435 ;
        RECT -22.605 -152.485 -22.275 -152.155 ;
        RECT -22.605 -153.845 -22.275 -153.515 ;
        RECT -22.605 -156.09 -22.275 -154.96 ;
        RECT -22.6 -156.205 -22.28 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 42.08 -20.915 43.21 ;
        RECT -21.245 40.635 -20.915 40.965 ;
        RECT -21.245 39.275 -20.915 39.605 ;
        RECT -21.245 37.915 -20.915 38.245 ;
        RECT -21.245 36.555 -20.915 36.885 ;
        RECT -21.245 35.195 -20.915 35.525 ;
        RECT -21.245 33.835 -20.915 34.165 ;
        RECT -21.245 32.475 -20.915 32.805 ;
        RECT -21.245 31.115 -20.915 31.445 ;
        RECT -21.245 29.755 -20.915 30.085 ;
        RECT -21.245 28.395 -20.915 28.725 ;
        RECT -21.245 27.035 -20.915 27.365 ;
        RECT -21.245 25.675 -20.915 26.005 ;
        RECT -21.245 24.315 -20.915 24.645 ;
        RECT -21.245 22.955 -20.915 23.285 ;
        RECT -21.245 21.595 -20.915 21.925 ;
        RECT -21.245 20.235 -20.915 20.565 ;
        RECT -21.245 18.875 -20.915 19.205 ;
        RECT -21.245 17.515 -20.915 17.845 ;
        RECT -21.245 16.155 -20.915 16.485 ;
        RECT -21.245 14.795 -20.915 15.125 ;
        RECT -21.245 13.435 -20.915 13.765 ;
        RECT -21.245 12.075 -20.915 12.405 ;
        RECT -21.245 10.715 -20.915 11.045 ;
        RECT -21.245 9.355 -20.915 9.685 ;
        RECT -21.245 7.995 -20.915 8.325 ;
        RECT -21.245 6.635 -20.915 6.965 ;
        RECT -21.245 5.275 -20.915 5.605 ;
        RECT -21.245 3.915 -20.915 4.245 ;
        RECT -21.245 2.555 -20.915 2.885 ;
        RECT -21.245 -1.525 -20.915 -1.195 ;
        RECT -21.245 -2.885 -20.915 -2.555 ;
        RECT -21.245 -4.245 -20.915 -3.915 ;
        RECT -21.245 -6.965 -20.915 -6.635 ;
        RECT -21.245 -8.325 -20.915 -7.995 ;
        RECT -21.245 -12.405 -20.915 -12.075 ;
        RECT -21.245 -13.765 -20.915 -13.435 ;
        RECT -21.245 -16.485 -20.915 -16.155 ;
        RECT -21.245 -24.645 -20.915 -24.315 ;
        RECT -21.245 -26.005 -20.915 -25.675 ;
        RECT -21.245 -28.725 -20.915 -28.395 ;
        RECT -21.245 -30.085 -20.915 -29.755 ;
        RECT -21.245 -32.805 -20.915 -32.475 ;
        RECT -21.245 -35.525 -20.915 -35.195 ;
        RECT -21.245 -38.245 -20.915 -37.915 ;
        RECT -21.245 -45.045 -20.915 -44.715 ;
        RECT -21.245 -46.405 -20.915 -46.075 ;
        RECT -21.245 -49.125 -20.915 -48.795 ;
        RECT -21.245 -50.485 -20.915 -50.155 ;
        RECT -21.245 -53.205 -20.915 -52.875 ;
        RECT -21.245 -54.565 -20.915 -54.235 ;
        RECT -21.245 -57.285 -20.915 -56.955 ;
        RECT -21.245 -58.645 -20.915 -58.315 ;
        RECT -21.245 -61.365 -20.915 -61.035 ;
        RECT -21.24 -62.72 -20.92 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 -99.445 -20.915 -99.115 ;
        RECT -21.245 -100.805 -20.915 -100.475 ;
        RECT -21.245 -102.165 -20.915 -101.835 ;
        RECT -21.245 -104.885 -20.915 -104.555 ;
        RECT -21.245 -110.325 -20.915 -109.995 ;
        RECT -21.245 -115.765 -20.915 -115.435 ;
        RECT -21.245 -118.485 -20.915 -118.155 ;
        RECT -21.245 -121.205 -20.915 -120.875 ;
        RECT -21.245 -122.565 -20.915 -122.235 ;
        RECT -21.245 -126.645 -20.915 -126.315 ;
        RECT -21.245 -128.005 -20.915 -127.675 ;
        RECT -21.245 -133.445 -20.915 -133.115 ;
        RECT -21.245 -134.805 -20.915 -134.475 ;
        RECT -21.245 -136.165 -20.915 -135.835 ;
        RECT -21.245 -137.525 -20.915 -137.195 ;
        RECT -21.245 -138.885 -20.915 -138.555 ;
        RECT -21.245 -140.245 -20.915 -139.915 ;
        RECT -21.245 -141.605 -20.915 -141.275 ;
        RECT -21.245 -142.965 -20.915 -142.635 ;
        RECT -21.245 -145.685 -20.915 -145.355 ;
        RECT -21.245 -149.765 -20.915 -149.435 ;
        RECT -21.245 -150.825 -20.915 -150.495 ;
        RECT -21.245 -152.485 -20.915 -152.155 ;
        RECT -21.245 -153.845 -20.915 -153.515 ;
        RECT -21.245 -156.09 -20.915 -154.96 ;
        RECT -21.24 -156.205 -20.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 6.635 -19.555 6.965 ;
        RECT -19.885 5.275 -19.555 5.605 ;
        RECT -19.885 3.915 -19.555 4.245 ;
        RECT -19.885 2.555 -19.555 2.885 ;
        RECT -19.885 -1.525 -19.555 -1.195 ;
        RECT -19.885 -2.885 -19.555 -2.555 ;
        RECT -19.885 -4.245 -19.555 -3.915 ;
        RECT -19.885 -6.965 -19.555 -6.635 ;
        RECT -19.885 -8.325 -19.555 -7.995 ;
        RECT -19.885 -9.87 -19.555 -9.54 ;
        RECT -19.885 -12.405 -19.555 -12.075 ;
        RECT -19.885 -13.765 -19.555 -13.435 ;
        RECT -19.885 -14.71 -19.555 -14.38 ;
        RECT -19.885 -16.485 -19.555 -16.155 ;
        RECT -19.885 -24.645 -19.555 -24.315 ;
        RECT -19.885 -26.005 -19.555 -25.675 ;
        RECT -19.885 -28.725 -19.555 -28.395 ;
        RECT -19.885 -30.085 -19.555 -29.755 ;
        RECT -19.885 -31.89 -19.555 -31.56 ;
        RECT -19.885 -32.805 -19.555 -32.475 ;
        RECT -19.885 -35.525 -19.555 -35.195 ;
        RECT -19.885 -36.73 -19.555 -36.4 ;
        RECT -19.885 -38.245 -19.555 -37.915 ;
        RECT -19.885 -45.045 -19.555 -44.715 ;
        RECT -19.885 -46.405 -19.555 -46.075 ;
        RECT -19.885 -49.125 -19.555 -48.795 ;
        RECT -19.885 -50.485 -19.555 -50.155 ;
        RECT -19.885 -51.81 -19.555 -51.48 ;
        RECT -19.885 -53.205 -19.555 -52.875 ;
        RECT -19.885 -54.565 -19.555 -54.235 ;
        RECT -19.885 -57.285 -19.555 -56.955 ;
        RECT -19.885 -58.645 -19.555 -58.315 ;
        RECT -19.885 -60.35 -19.555 -60.02 ;
        RECT -19.885 -61.365 -19.555 -61.035 ;
        RECT -19.885 -64.085 -19.555 -63.755 ;
        RECT -19.885 -65.445 -19.555 -65.115 ;
        RECT -19.885 -66.805 -19.555 -66.475 ;
        RECT -19.885 -68.165 -19.555 -67.835 ;
        RECT -19.885 -69.525 -19.555 -69.195 ;
        RECT -19.885 -72.245 -19.555 -71.915 ;
        RECT -19.885 -73.99 -19.555 -73.66 ;
        RECT -19.885 -74.965 -19.555 -74.635 ;
        RECT -19.885 -76.325 -19.555 -75.995 ;
        RECT -19.885 -79.045 -19.555 -78.715 ;
        RECT -19.885 -80.405 -19.555 -80.075 ;
        RECT -19.885 -81.765 -19.555 -81.435 ;
        RECT -19.885 -82.53 -19.555 -82.2 ;
        RECT -19.885 -84.485 -19.555 -84.155 ;
        RECT -19.885 -88.565 -19.555 -88.235 ;
        RECT -19.885 -89.925 -19.555 -89.595 ;
        RECT -19.885 -91.285 -19.555 -90.955 ;
        RECT -19.885 -92.645 -19.555 -92.315 ;
        RECT -19.885 -99.445 -19.555 -99.115 ;
        RECT -19.885 -100.805 -19.555 -100.475 ;
        RECT -19.885 -102.165 -19.555 -101.835 ;
        RECT -19.885 -110.325 -19.555 -109.995 ;
        RECT -19.885 -115.765 -19.555 -115.435 ;
        RECT -19.885 -118.485 -19.555 -118.155 ;
        RECT -19.885 -119.845 -19.555 -119.515 ;
        RECT -19.885 -122.565 -19.555 -122.235 ;
        RECT -19.885 -126.645 -19.555 -126.315 ;
        RECT -19.885 -128.005 -19.555 -127.675 ;
        RECT -19.885 -133.445 -19.555 -133.115 ;
        RECT -19.885 -134.805 -19.555 -134.475 ;
        RECT -19.885 -136.165 -19.555 -135.835 ;
        RECT -19.885 -137.525 -19.555 -137.195 ;
        RECT -19.885 -138.885 -19.555 -138.555 ;
        RECT -19.885 -140.245 -19.555 -139.915 ;
        RECT -19.885 -141.605 -19.555 -141.275 ;
        RECT -19.885 -142.965 -19.555 -142.635 ;
        RECT -19.885 -145.685 -19.555 -145.355 ;
        RECT -19.885 -147.045 -19.555 -146.715 ;
        RECT -19.885 -148.405 -19.555 -148.075 ;
        RECT -19.885 -149.765 -19.555 -149.435 ;
        RECT -19.885 -150.825 -19.555 -150.495 ;
        RECT -19.885 -152.485 -19.555 -152.155 ;
        RECT -19.885 -153.845 -19.555 -153.515 ;
        RECT -19.885 -156.09 -19.555 -154.96 ;
        RECT -19.88 -156.205 -19.56 43.325 ;
        RECT -19.885 42.08 -19.555 43.21 ;
        RECT -19.885 40.635 -19.555 40.965 ;
        RECT -19.885 39.275 -19.555 39.605 ;
        RECT -19.885 37.915 -19.555 38.245 ;
        RECT -19.885 36.555 -19.555 36.885 ;
        RECT -19.885 35.195 -19.555 35.525 ;
        RECT -19.885 33.835 -19.555 34.165 ;
        RECT -19.885 32.475 -19.555 32.805 ;
        RECT -19.885 31.115 -19.555 31.445 ;
        RECT -19.885 29.755 -19.555 30.085 ;
        RECT -19.885 28.395 -19.555 28.725 ;
        RECT -19.885 27.035 -19.555 27.365 ;
        RECT -19.885 25.675 -19.555 26.005 ;
        RECT -19.885 24.315 -19.555 24.645 ;
        RECT -19.885 22.955 -19.555 23.285 ;
        RECT -19.885 21.595 -19.555 21.925 ;
        RECT -19.885 20.235 -19.555 20.565 ;
        RECT -19.885 18.875 -19.555 19.205 ;
        RECT -19.885 17.515 -19.555 17.845 ;
        RECT -19.885 16.155 -19.555 16.485 ;
        RECT -19.885 14.795 -19.555 15.125 ;
        RECT -19.885 13.435 -19.555 13.765 ;
        RECT -19.885 12.075 -19.555 12.405 ;
        RECT -19.885 10.715 -19.555 11.045 ;
        RECT -19.885 9.355 -19.555 9.685 ;
        RECT -19.885 7.995 -19.555 8.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.645 42.08 -41.315 43.21 ;
        RECT -41.645 40.635 -41.315 40.965 ;
        RECT -41.645 39.275 -41.315 39.605 ;
        RECT -41.645 37.915 -41.315 38.245 ;
        RECT -41.645 36.555 -41.315 36.885 ;
        RECT -41.645 35.195 -41.315 35.525 ;
        RECT -41.645 33.835 -41.315 34.165 ;
        RECT -41.645 32.475 -41.315 32.805 ;
        RECT -41.645 31.115 -41.315 31.445 ;
        RECT -41.645 29.755 -41.315 30.085 ;
        RECT -41.645 28.395 -41.315 28.725 ;
        RECT -41.645 27.035 -41.315 27.365 ;
        RECT -41.645 25.675 -41.315 26.005 ;
        RECT -41.645 24.315 -41.315 24.645 ;
        RECT -41.645 23.465 -41.315 23.795 ;
        RECT -41.645 21.415 -41.315 21.745 ;
        RECT -41.645 19.055 -41.315 19.385 ;
        RECT -41.645 17.735 -41.315 18.065 ;
        RECT -41.645 15.545 -41.315 15.875 ;
        RECT -41.645 13.49 -41.315 13.82 ;
        RECT -41.645 12.075 -41.315 12.405 ;
        RECT -41.645 10.715 -41.315 11.045 ;
        RECT -41.645 9.355 -41.315 9.685 ;
        RECT -41.645 7.995 -41.315 8.325 ;
        RECT -41.645 6.635 -41.315 6.965 ;
        RECT -41.645 5.275 -41.315 5.605 ;
        RECT -41.645 3.915 -41.315 4.245 ;
        RECT -41.645 2.555 -41.315 2.885 ;
        RECT -41.645 1.195 -41.315 1.525 ;
        RECT -41.645 -0.165 -41.315 0.165 ;
        RECT -41.645 -1.525 -41.315 -1.195 ;
        RECT -41.645 -2.885 -41.315 -2.555 ;
        RECT -41.645 -4.245 -41.315 -3.915 ;
        RECT -41.645 -5.605 -41.315 -5.275 ;
        RECT -41.645 -6.965 -41.315 -6.635 ;
        RECT -41.645 -8.325 -41.315 -7.995 ;
        RECT -41.645 -9.685 -41.315 -9.355 ;
        RECT -41.645 -11.045 -41.315 -10.715 ;
        RECT -41.645 -12.405 -41.315 -12.075 ;
        RECT -41.645 -13.765 -41.315 -13.435 ;
        RECT -41.645 -15.125 -41.315 -14.795 ;
        RECT -41.645 -16.485 -41.315 -16.155 ;
        RECT -41.645 -17.845 -41.315 -17.515 ;
        RECT -41.645 -19.205 -41.315 -18.875 ;
        RECT -41.645 -21.925 -41.315 -21.595 ;
        RECT -41.645 -23.285 -41.315 -22.955 ;
        RECT -41.645 -24.645 -41.315 -24.315 ;
        RECT -41.645 -26.005 -41.315 -25.675 ;
        RECT -41.645 -27.365 -41.315 -27.035 ;
        RECT -41.645 -28.725 -41.315 -28.395 ;
        RECT -41.645 -30.085 -41.315 -29.755 ;
        RECT -41.645 -31.445 -41.315 -31.115 ;
        RECT -41.645 -32.805 -41.315 -32.475 ;
        RECT -41.645 -34.165 -41.315 -33.835 ;
        RECT -41.645 -35.525 -41.315 -35.195 ;
        RECT -41.645 -36.885 -41.315 -36.555 ;
        RECT -41.645 -38.245 -41.315 -37.915 ;
        RECT -41.645 -39.605 -41.315 -39.275 ;
        RECT -41.645 -40.965 -41.315 -40.635 ;
        RECT -41.645 -42.325 -41.315 -41.995 ;
        RECT -41.645 -43.685 -41.315 -43.355 ;
        RECT -41.645 -45.045 -41.315 -44.715 ;
        RECT -41.645 -46.405 -41.315 -46.075 ;
        RECT -41.645 -47.765 -41.315 -47.435 ;
        RECT -41.645 -49.125 -41.315 -48.795 ;
        RECT -41.645 -50.485 -41.315 -50.155 ;
        RECT -41.645 -51.845 -41.315 -51.515 ;
        RECT -41.645 -53.205 -41.315 -52.875 ;
        RECT -41.645 -54.565 -41.315 -54.235 ;
        RECT -41.645 -55.925 -41.315 -55.595 ;
        RECT -41.645 -57.285 -41.315 -56.955 ;
        RECT -41.645 -58.645 -41.315 -58.315 ;
        RECT -41.645 -60.005 -41.315 -59.675 ;
        RECT -41.645 -61.365 -41.315 -61.035 ;
        RECT -41.645 -62.725 -41.315 -62.395 ;
        RECT -41.645 -64.085 -41.315 -63.755 ;
        RECT -41.645 -66.805 -41.315 -66.475 ;
        RECT -41.645 -68.165 -41.315 -67.835 ;
        RECT -41.645 -69.525 -41.315 -69.195 ;
        RECT -41.645 -70.885 -41.315 -70.555 ;
        RECT -41.645 -72.245 -41.315 -71.915 ;
        RECT -41.645 -73.83 -41.315 -73.5 ;
        RECT -41.645 -74.965 -41.315 -74.635 ;
        RECT -41.645 -77.685 -41.315 -77.355 ;
        RECT -41.645 -79.045 -41.315 -78.715 ;
        RECT -41.645 -80.405 -41.315 -80.075 ;
        RECT -41.645 -81.97 -41.315 -81.64 ;
        RECT -41.645 -83.125 -41.315 -82.795 ;
        RECT -41.645 -84.485 -41.315 -84.155 ;
        RECT -41.645 -85.845 -41.315 -85.515 ;
        RECT -41.645 -89.925 -41.315 -89.595 ;
        RECT -41.645 -91.285 -41.315 -90.955 ;
        RECT -41.645 -92.645 -41.315 -92.315 ;
        RECT -41.645 -98.085 -41.315 -97.755 ;
        RECT -41.645 -99.445 -41.315 -99.115 ;
        RECT -41.645 -100.805 -41.315 -100.475 ;
        RECT -41.645 -102.165 -41.315 -101.835 ;
        RECT -41.645 -103.525 -41.315 -103.195 ;
        RECT -41.645 -104.885 -41.315 -104.555 ;
        RECT -41.645 -106.245 -41.315 -105.915 ;
        RECT -41.645 -107.605 -41.315 -107.275 ;
        RECT -41.645 -108.965 -41.315 -108.635 ;
        RECT -41.645 -110.325 -41.315 -109.995 ;
        RECT -41.645 -111.685 -41.315 -111.355 ;
        RECT -41.645 -113.045 -41.315 -112.715 ;
        RECT -41.645 -114.405 -41.315 -114.075 ;
        RECT -41.645 -115.765 -41.315 -115.435 ;
        RECT -41.645 -117.125 -41.315 -116.795 ;
        RECT -41.645 -118.485 -41.315 -118.155 ;
        RECT -41.645 -119.845 -41.315 -119.515 ;
        RECT -41.645 -121.205 -41.315 -120.875 ;
        RECT -41.645 -122.565 -41.315 -122.235 ;
        RECT -41.645 -123.925 -41.315 -123.595 ;
        RECT -41.645 -125.285 -41.315 -124.955 ;
        RECT -41.645 -126.645 -41.315 -126.315 ;
        RECT -41.645 -128.005 -41.315 -127.675 ;
        RECT -41.645 -129.365 -41.315 -129.035 ;
        RECT -41.645 -130.725 -41.315 -130.395 ;
        RECT -41.645 -132.085 -41.315 -131.755 ;
        RECT -41.645 -133.445 -41.315 -133.115 ;
        RECT -41.645 -134.805 -41.315 -134.475 ;
        RECT -41.645 -136.165 -41.315 -135.835 ;
        RECT -41.645 -137.525 -41.315 -137.195 ;
        RECT -41.645 -138.885 -41.315 -138.555 ;
        RECT -41.645 -140.245 -41.315 -139.915 ;
        RECT -41.645 -141.605 -41.315 -141.275 ;
        RECT -41.645 -142.965 -41.315 -142.635 ;
        RECT -41.645 -145.685 -41.315 -145.355 ;
        RECT -41.645 -149.765 -41.315 -149.435 ;
        RECT -41.645 -152.485 -41.315 -152.155 ;
        RECT -41.645 -153.845 -41.315 -153.515 ;
        RECT -41.645 -156.09 -41.315 -154.96 ;
        RECT -41.64 -156.205 -41.32 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.285 42.08 -39.955 43.21 ;
        RECT -40.285 40.635 -39.955 40.965 ;
        RECT -40.285 39.275 -39.955 39.605 ;
        RECT -40.285 37.915 -39.955 38.245 ;
        RECT -40.285 36.555 -39.955 36.885 ;
        RECT -40.285 35.195 -39.955 35.525 ;
        RECT -40.285 33.835 -39.955 34.165 ;
        RECT -40.285 32.475 -39.955 32.805 ;
        RECT -40.285 31.115 -39.955 31.445 ;
        RECT -40.285 29.755 -39.955 30.085 ;
        RECT -40.285 28.395 -39.955 28.725 ;
        RECT -40.285 27.035 -39.955 27.365 ;
        RECT -40.285 25.675 -39.955 26.005 ;
        RECT -40.285 24.315 -39.955 24.645 ;
        RECT -40.285 12.075 -39.955 12.405 ;
        RECT -40.285 10.715 -39.955 11.045 ;
        RECT -40.285 9.355 -39.955 9.685 ;
        RECT -40.285 7.995 -39.955 8.325 ;
        RECT -40.285 6.635 -39.955 6.965 ;
        RECT -40.285 5.275 -39.955 5.605 ;
        RECT -40.285 3.915 -39.955 4.245 ;
        RECT -40.285 2.555 -39.955 2.885 ;
        RECT -40.285 1.195 -39.955 1.525 ;
        RECT -40.285 -0.165 -39.955 0.165 ;
        RECT -40.285 -1.525 -39.955 -1.195 ;
        RECT -40.285 -2.885 -39.955 -2.555 ;
        RECT -40.285 -4.245 -39.955 -3.915 ;
        RECT -40.285 -5.605 -39.955 -5.275 ;
        RECT -40.285 -6.965 -39.955 -6.635 ;
        RECT -40.285 -8.325 -39.955 -7.995 ;
        RECT -40.285 -9.685 -39.955 -9.355 ;
        RECT -40.285 -11.045 -39.955 -10.715 ;
        RECT -40.285 -12.405 -39.955 -12.075 ;
        RECT -40.285 -13.765 -39.955 -13.435 ;
        RECT -40.285 -15.125 -39.955 -14.795 ;
        RECT -40.285 -16.485 -39.955 -16.155 ;
        RECT -40.285 -17.845 -39.955 -17.515 ;
        RECT -40.285 -19.205 -39.955 -18.875 ;
        RECT -40.285 -21.925 -39.955 -21.595 ;
        RECT -40.285 -24.645 -39.955 -24.315 ;
        RECT -40.285 -26.005 -39.955 -25.675 ;
        RECT -40.285 -27.365 -39.955 -27.035 ;
        RECT -40.285 -28.725 -39.955 -28.395 ;
        RECT -40.285 -30.085 -39.955 -29.755 ;
        RECT -40.285 -31.445 -39.955 -31.115 ;
        RECT -40.285 -32.805 -39.955 -32.475 ;
        RECT -40.285 -34.165 -39.955 -33.835 ;
        RECT -40.285 -35.525 -39.955 -35.195 ;
        RECT -40.285 -36.885 -39.955 -36.555 ;
        RECT -40.285 -38.245 -39.955 -37.915 ;
        RECT -40.285 -39.605 -39.955 -39.275 ;
        RECT -40.285 -40.965 -39.955 -40.635 ;
        RECT -40.285 -42.325 -39.955 -41.995 ;
        RECT -40.285 -43.685 -39.955 -43.355 ;
        RECT -40.285 -45.045 -39.955 -44.715 ;
        RECT -40.285 -46.405 -39.955 -46.075 ;
        RECT -40.285 -47.765 -39.955 -47.435 ;
        RECT -40.285 -49.125 -39.955 -48.795 ;
        RECT -40.285 -50.485 -39.955 -50.155 ;
        RECT -40.285 -51.845 -39.955 -51.515 ;
        RECT -40.285 -53.205 -39.955 -52.875 ;
        RECT -40.285 -54.565 -39.955 -54.235 ;
        RECT -40.285 -55.925 -39.955 -55.595 ;
        RECT -40.285 -57.285 -39.955 -56.955 ;
        RECT -40.285 -58.645 -39.955 -58.315 ;
        RECT -40.285 -60.005 -39.955 -59.675 ;
        RECT -40.285 -61.365 -39.955 -61.035 ;
        RECT -40.285 -62.725 -39.955 -62.395 ;
        RECT -40.285 -64.085 -39.955 -63.755 ;
        RECT -40.285 -66.805 -39.955 -66.475 ;
        RECT -40.285 -68.165 -39.955 -67.835 ;
        RECT -40.285 -69.525 -39.955 -69.195 ;
        RECT -40.285 -70.885 -39.955 -70.555 ;
        RECT -40.285 -72.245 -39.955 -71.915 ;
        RECT -40.285 -73.83 -39.955 -73.5 ;
        RECT -40.285 -74.965 -39.955 -74.635 ;
        RECT -40.285 -77.685 -39.955 -77.355 ;
        RECT -40.285 -79.045 -39.955 -78.715 ;
        RECT -40.285 -80.405 -39.955 -80.075 ;
        RECT -40.285 -81.97 -39.955 -81.64 ;
        RECT -40.285 -83.125 -39.955 -82.795 ;
        RECT -40.285 -84.485 -39.955 -84.155 ;
        RECT -40.285 -85.845 -39.955 -85.515 ;
        RECT -40.28 -87.2 -39.96 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.925 42.08 -38.595 43.21 ;
        RECT -38.925 40.635 -38.595 40.965 ;
        RECT -38.925 39.275 -38.595 39.605 ;
        RECT -38.925 37.915 -38.595 38.245 ;
        RECT -38.925 36.555 -38.595 36.885 ;
        RECT -38.925 35.195 -38.595 35.525 ;
        RECT -38.925 33.835 -38.595 34.165 ;
        RECT -38.925 32.475 -38.595 32.805 ;
        RECT -38.925 31.115 -38.595 31.445 ;
        RECT -38.925 29.755 -38.595 30.085 ;
        RECT -38.925 28.395 -38.595 28.725 ;
        RECT -38.925 27.035 -38.595 27.365 ;
        RECT -38.925 25.675 -38.595 26.005 ;
        RECT -38.925 24.315 -38.595 24.645 ;
        RECT -38.925 22.955 -38.595 23.285 ;
        RECT -38.925 21.595 -38.595 21.925 ;
        RECT -38.925 20.235 -38.595 20.565 ;
        RECT -38.925 18.875 -38.595 19.205 ;
        RECT -38.925 17.515 -38.595 17.845 ;
        RECT -38.925 16.155 -38.595 16.485 ;
        RECT -38.925 14.795 -38.595 15.125 ;
        RECT -38.925 13.435 -38.595 13.765 ;
        RECT -38.925 12.075 -38.595 12.405 ;
        RECT -38.925 10.715 -38.595 11.045 ;
        RECT -38.925 9.355 -38.595 9.685 ;
        RECT -38.925 7.995 -38.595 8.325 ;
        RECT -38.925 6.635 -38.595 6.965 ;
        RECT -38.925 5.275 -38.595 5.605 ;
        RECT -38.925 3.915 -38.595 4.245 ;
        RECT -38.925 2.555 -38.595 2.885 ;
        RECT -38.925 1.195 -38.595 1.525 ;
        RECT -38.925 -1.525 -38.595 -1.195 ;
        RECT -38.925 -2.885 -38.595 -2.555 ;
        RECT -38.925 -4.245 -38.595 -3.915 ;
        RECT -38.925 -5.605 -38.595 -5.275 ;
        RECT -38.925 -6.965 -38.595 -6.635 ;
        RECT -38.925 -8.325 -38.595 -7.995 ;
        RECT -38.925 -9.685 -38.595 -9.355 ;
        RECT -38.925 -11.045 -38.595 -10.715 ;
        RECT -38.925 -12.405 -38.595 -12.075 ;
        RECT -38.925 -13.765 -38.595 -13.435 ;
        RECT -38.925 -15.125 -38.595 -14.795 ;
        RECT -38.925 -16.485 -38.595 -16.155 ;
        RECT -38.925 -17.845 -38.595 -17.515 ;
        RECT -38.925 -19.205 -38.595 -18.875 ;
        RECT -38.925 -24.645 -38.595 -24.315 ;
        RECT -38.925 -26.005 -38.595 -25.675 ;
        RECT -38.925 -27.365 -38.595 -27.035 ;
        RECT -38.925 -28.725 -38.595 -28.395 ;
        RECT -38.925 -30.085 -38.595 -29.755 ;
        RECT -38.925 -31.445 -38.595 -31.115 ;
        RECT -38.925 -32.805 -38.595 -32.475 ;
        RECT -38.925 -34.165 -38.595 -33.835 ;
        RECT -38.925 -35.525 -38.595 -35.195 ;
        RECT -38.925 -36.885 -38.595 -36.555 ;
        RECT -38.925 -38.245 -38.595 -37.915 ;
        RECT -38.925 -39.605 -38.595 -39.275 ;
        RECT -38.925 -40.965 -38.595 -40.635 ;
        RECT -38.925 -42.325 -38.595 -41.995 ;
        RECT -38.925 -43.685 -38.595 -43.355 ;
        RECT -38.925 -45.045 -38.595 -44.715 ;
        RECT -38.925 -46.405 -38.595 -46.075 ;
        RECT -38.925 -47.765 -38.595 -47.435 ;
        RECT -38.925 -49.125 -38.595 -48.795 ;
        RECT -38.925 -50.485 -38.595 -50.155 ;
        RECT -38.925 -51.845 -38.595 -51.515 ;
        RECT -38.925 -53.205 -38.595 -52.875 ;
        RECT -38.925 -54.565 -38.595 -54.235 ;
        RECT -38.925 -55.925 -38.595 -55.595 ;
        RECT -38.925 -57.285 -38.595 -56.955 ;
        RECT -38.925 -58.645 -38.595 -58.315 ;
        RECT -38.925 -60.005 -38.595 -59.675 ;
        RECT -38.925 -61.365 -38.595 -61.035 ;
        RECT -38.925 -62.725 -38.595 -62.395 ;
        RECT -38.925 -64.085 -38.595 -63.755 ;
        RECT -38.925 -66.805 -38.595 -66.475 ;
        RECT -38.925 -68.165 -38.595 -67.835 ;
        RECT -38.925 -69.525 -38.595 -69.195 ;
        RECT -38.925 -70.885 -38.595 -70.555 ;
        RECT -38.925 -72.245 -38.595 -71.915 ;
        RECT -38.925 -73.83 -38.595 -73.5 ;
        RECT -38.925 -74.965 -38.595 -74.635 ;
        RECT -38.925 -77.685 -38.595 -77.355 ;
        RECT -38.925 -79.045 -38.595 -78.715 ;
        RECT -38.925 -80.405 -38.595 -80.075 ;
        RECT -38.925 -81.97 -38.595 -81.64 ;
        RECT -38.925 -83.125 -38.595 -82.795 ;
        RECT -38.925 -84.485 -38.595 -84.155 ;
        RECT -38.925 -85.845 -38.595 -85.515 ;
        RECT -38.925 -89.925 -38.595 -89.595 ;
        RECT -38.925 -91.285 -38.595 -90.955 ;
        RECT -38.925 -92.645 -38.595 -92.315 ;
        RECT -38.925 -98.085 -38.595 -97.755 ;
        RECT -38.925 -99.445 -38.595 -99.115 ;
        RECT -38.925 -100.805 -38.595 -100.475 ;
        RECT -38.925 -102.165 -38.595 -101.835 ;
        RECT -38.925 -103.525 -38.595 -103.195 ;
        RECT -38.925 -104.885 -38.595 -104.555 ;
        RECT -38.925 -107.605 -38.595 -107.275 ;
        RECT -38.925 -108.965 -38.595 -108.635 ;
        RECT -38.925 -110.325 -38.595 -109.995 ;
        RECT -38.925 -111.685 -38.595 -111.355 ;
        RECT -38.925 -113.045 -38.595 -112.715 ;
        RECT -38.925 -114.405 -38.595 -114.075 ;
        RECT -38.925 -115.765 -38.595 -115.435 ;
        RECT -38.925 -117.125 -38.595 -116.795 ;
        RECT -38.925 -118.485 -38.595 -118.155 ;
        RECT -38.925 -119.845 -38.595 -119.515 ;
        RECT -38.925 -121.205 -38.595 -120.875 ;
        RECT -38.925 -122.565 -38.595 -122.235 ;
        RECT -38.925 -125.285 -38.595 -124.955 ;
        RECT -38.925 -126.645 -38.595 -126.315 ;
        RECT -38.925 -128.005 -38.595 -127.675 ;
        RECT -38.925 -130.725 -38.595 -130.395 ;
        RECT -38.925 -132.085 -38.595 -131.755 ;
        RECT -38.925 -133.445 -38.595 -133.115 ;
        RECT -38.925 -134.805 -38.595 -134.475 ;
        RECT -38.925 -136.165 -38.595 -135.835 ;
        RECT -38.925 -137.525 -38.595 -137.195 ;
        RECT -38.925 -138.885 -38.595 -138.555 ;
        RECT -38.925 -140.245 -38.595 -139.915 ;
        RECT -38.925 -141.605 -38.595 -141.275 ;
        RECT -38.92 -141.605 -38.6 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.925 -148.405 -38.595 -148.075 ;
        RECT -38.925 -149.765 -38.595 -149.435 ;
        RECT -38.925 -150.825 -38.595 -150.495 ;
        RECT -38.925 -152.485 -38.595 -152.155 ;
        RECT -38.925 -153.845 -38.595 -153.515 ;
        RECT -38.925 -156.09 -38.595 -154.96 ;
        RECT -38.92 -156.205 -38.6 -147.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.565 42.08 -37.235 43.21 ;
        RECT -37.565 40.635 -37.235 40.965 ;
        RECT -37.565 39.275 -37.235 39.605 ;
        RECT -37.565 37.915 -37.235 38.245 ;
        RECT -37.565 36.555 -37.235 36.885 ;
        RECT -37.565 35.195 -37.235 35.525 ;
        RECT -37.565 33.835 -37.235 34.165 ;
        RECT -37.565 32.475 -37.235 32.805 ;
        RECT -37.565 31.115 -37.235 31.445 ;
        RECT -37.565 29.755 -37.235 30.085 ;
        RECT -37.565 28.395 -37.235 28.725 ;
        RECT -37.565 27.035 -37.235 27.365 ;
        RECT -37.565 25.675 -37.235 26.005 ;
        RECT -37.565 24.315 -37.235 24.645 ;
        RECT -37.565 22.955 -37.235 23.285 ;
        RECT -37.565 21.595 -37.235 21.925 ;
        RECT -37.565 20.235 -37.235 20.565 ;
        RECT -37.565 18.875 -37.235 19.205 ;
        RECT -37.565 17.515 -37.235 17.845 ;
        RECT -37.565 16.155 -37.235 16.485 ;
        RECT -37.565 14.795 -37.235 15.125 ;
        RECT -37.565 13.435 -37.235 13.765 ;
        RECT -37.565 12.075 -37.235 12.405 ;
        RECT -37.565 10.715 -37.235 11.045 ;
        RECT -37.565 9.355 -37.235 9.685 ;
        RECT -37.565 7.995 -37.235 8.325 ;
        RECT -37.565 6.635 -37.235 6.965 ;
        RECT -37.565 5.275 -37.235 5.605 ;
        RECT -37.565 3.915 -37.235 4.245 ;
        RECT -37.565 2.555 -37.235 2.885 ;
        RECT -37.565 -1.525 -37.235 -1.195 ;
        RECT -37.565 -2.885 -37.235 -2.555 ;
        RECT -37.565 -4.245 -37.235 -3.915 ;
        RECT -37.565 -5.605 -37.235 -5.275 ;
        RECT -37.565 -6.965 -37.235 -6.635 ;
        RECT -37.565 -8.325 -37.235 -7.995 ;
        RECT -37.565 -9.685 -37.235 -9.355 ;
        RECT -37.565 -11.045 -37.235 -10.715 ;
        RECT -37.565 -12.405 -37.235 -12.075 ;
        RECT -37.565 -13.765 -37.235 -13.435 ;
        RECT -37.565 -15.125 -37.235 -14.795 ;
        RECT -37.565 -16.485 -37.235 -16.155 ;
        RECT -37.565 -17.845 -37.235 -17.515 ;
        RECT -37.565 -19.205 -37.235 -18.875 ;
        RECT -37.565 -24.645 -37.235 -24.315 ;
        RECT -37.565 -26.005 -37.235 -25.675 ;
        RECT -37.565 -27.365 -37.235 -27.035 ;
        RECT -37.565 -28.725 -37.235 -28.395 ;
        RECT -37.565 -30.085 -37.235 -29.755 ;
        RECT -37.565 -31.445 -37.235 -31.115 ;
        RECT -37.565 -32.805 -37.235 -32.475 ;
        RECT -37.565 -34.165 -37.235 -33.835 ;
        RECT -37.565 -35.525 -37.235 -35.195 ;
        RECT -37.565 -36.885 -37.235 -36.555 ;
        RECT -37.565 -38.245 -37.235 -37.915 ;
        RECT -37.565 -39.605 -37.235 -39.275 ;
        RECT -37.565 -40.965 -37.235 -40.635 ;
        RECT -37.565 -42.325 -37.235 -41.995 ;
        RECT -37.565 -43.685 -37.235 -43.355 ;
        RECT -37.565 -45.045 -37.235 -44.715 ;
        RECT -37.565 -46.405 -37.235 -46.075 ;
        RECT -37.565 -47.765 -37.235 -47.435 ;
        RECT -37.565 -49.125 -37.235 -48.795 ;
        RECT -37.565 -50.485 -37.235 -50.155 ;
        RECT -37.565 -51.845 -37.235 -51.515 ;
        RECT -37.565 -53.205 -37.235 -52.875 ;
        RECT -37.565 -54.565 -37.235 -54.235 ;
        RECT -37.565 -55.925 -37.235 -55.595 ;
        RECT -37.565 -57.285 -37.235 -56.955 ;
        RECT -37.565 -58.645 -37.235 -58.315 ;
        RECT -37.565 -60.005 -37.235 -59.675 ;
        RECT -37.565 -61.365 -37.235 -61.035 ;
        RECT -37.565 -62.725 -37.235 -62.395 ;
        RECT -37.565 -64.085 -37.235 -63.755 ;
        RECT -37.565 -66.805 -37.235 -66.475 ;
        RECT -37.565 -68.165 -37.235 -67.835 ;
        RECT -37.565 -69.525 -37.235 -69.195 ;
        RECT -37.565 -70.885 -37.235 -70.555 ;
        RECT -37.565 -72.245 -37.235 -71.915 ;
        RECT -37.565 -73.83 -37.235 -73.5 ;
        RECT -37.565 -74.965 -37.235 -74.635 ;
        RECT -37.565 -77.685 -37.235 -77.355 ;
        RECT -37.565 -79.045 -37.235 -78.715 ;
        RECT -37.565 -80.405 -37.235 -80.075 ;
        RECT -37.565 -81.97 -37.235 -81.64 ;
        RECT -37.565 -83.125 -37.235 -82.795 ;
        RECT -37.565 -84.485 -37.235 -84.155 ;
        RECT -37.565 -85.845 -37.235 -85.515 ;
        RECT -37.565 -88.565 -37.235 -88.235 ;
        RECT -37.565 -89.925 -37.235 -89.595 ;
        RECT -37.565 -91.285 -37.235 -90.955 ;
        RECT -37.565 -92.645 -37.235 -92.315 ;
        RECT -37.565 -98.085 -37.235 -97.755 ;
        RECT -37.565 -99.445 -37.235 -99.115 ;
        RECT -37.565 -100.805 -37.235 -100.475 ;
        RECT -37.565 -102.165 -37.235 -101.835 ;
        RECT -37.565 -103.525 -37.235 -103.195 ;
        RECT -37.565 -104.885 -37.235 -104.555 ;
        RECT -37.565 -107.605 -37.235 -107.275 ;
        RECT -37.565 -108.965 -37.235 -108.635 ;
        RECT -37.565 -110.325 -37.235 -109.995 ;
        RECT -37.565 -111.685 -37.235 -111.355 ;
        RECT -37.565 -113.045 -37.235 -112.715 ;
        RECT -37.565 -114.405 -37.235 -114.075 ;
        RECT -37.565 -115.765 -37.235 -115.435 ;
        RECT -37.565 -117.125 -37.235 -116.795 ;
        RECT -37.565 -118.485 -37.235 -118.155 ;
        RECT -37.565 -119.845 -37.235 -119.515 ;
        RECT -37.565 -121.205 -37.235 -120.875 ;
        RECT -37.565 -122.565 -37.235 -122.235 ;
        RECT -37.565 -125.285 -37.235 -124.955 ;
        RECT -37.565 -126.645 -37.235 -126.315 ;
        RECT -37.565 -128.005 -37.235 -127.675 ;
        RECT -37.565 -132.085 -37.235 -131.755 ;
        RECT -37.565 -133.445 -37.235 -133.115 ;
        RECT -37.565 -134.805 -37.235 -134.475 ;
        RECT -37.565 -136.165 -37.235 -135.835 ;
        RECT -37.565 -137.525 -37.235 -137.195 ;
        RECT -37.565 -138.885 -37.235 -138.555 ;
        RECT -37.565 -140.245 -37.235 -139.915 ;
        RECT -37.565 -141.605 -37.235 -141.275 ;
        RECT -37.565 -142.965 -37.235 -142.635 ;
        RECT -37.565 -145.685 -37.235 -145.355 ;
        RECT -37.565 -147.045 -37.235 -146.715 ;
        RECT -37.565 -148.405 -37.235 -148.075 ;
        RECT -37.565 -149.765 -37.235 -149.435 ;
        RECT -37.565 -150.825 -37.235 -150.495 ;
        RECT -37.565 -152.485 -37.235 -152.155 ;
        RECT -37.565 -153.845 -37.235 -153.515 ;
        RECT -37.565 -156.09 -37.235 -154.96 ;
        RECT -37.56 -156.205 -37.24 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.205 42.08 -35.875 43.21 ;
        RECT -36.205 40.635 -35.875 40.965 ;
        RECT -36.205 39.275 -35.875 39.605 ;
        RECT -36.205 37.915 -35.875 38.245 ;
        RECT -36.205 36.555 -35.875 36.885 ;
        RECT -36.205 35.195 -35.875 35.525 ;
        RECT -36.205 33.835 -35.875 34.165 ;
        RECT -36.205 32.475 -35.875 32.805 ;
        RECT -36.205 31.115 -35.875 31.445 ;
        RECT -36.205 29.755 -35.875 30.085 ;
        RECT -36.205 28.395 -35.875 28.725 ;
        RECT -36.205 27.035 -35.875 27.365 ;
        RECT -36.205 25.675 -35.875 26.005 ;
        RECT -36.205 24.315 -35.875 24.645 ;
        RECT -36.205 22.955 -35.875 23.285 ;
        RECT -36.205 21.595 -35.875 21.925 ;
        RECT -36.205 20.235 -35.875 20.565 ;
        RECT -36.205 18.875 -35.875 19.205 ;
        RECT -36.205 17.515 -35.875 17.845 ;
        RECT -36.205 16.155 -35.875 16.485 ;
        RECT -36.205 14.795 -35.875 15.125 ;
        RECT -36.205 13.435 -35.875 13.765 ;
        RECT -36.205 12.075 -35.875 12.405 ;
        RECT -36.205 10.715 -35.875 11.045 ;
        RECT -36.205 9.355 -35.875 9.685 ;
        RECT -36.205 7.995 -35.875 8.325 ;
        RECT -36.205 6.635 -35.875 6.965 ;
        RECT -36.205 5.275 -35.875 5.605 ;
        RECT -36.205 3.915 -35.875 4.245 ;
        RECT -36.205 2.555 -35.875 2.885 ;
        RECT -36.205 -1.525 -35.875 -1.195 ;
        RECT -36.205 -2.885 -35.875 -2.555 ;
        RECT -36.205 -4.245 -35.875 -3.915 ;
        RECT -36.205 -5.605 -35.875 -5.275 ;
        RECT -36.205 -6.965 -35.875 -6.635 ;
        RECT -36.205 -8.325 -35.875 -7.995 ;
        RECT -36.205 -9.685 -35.875 -9.355 ;
        RECT -36.205 -11.045 -35.875 -10.715 ;
        RECT -36.205 -12.405 -35.875 -12.075 ;
        RECT -36.205 -13.765 -35.875 -13.435 ;
        RECT -36.205 -15.125 -35.875 -14.795 ;
        RECT -36.205 -16.485 -35.875 -16.155 ;
        RECT -36.205 -17.845 -35.875 -17.515 ;
        RECT -36.205 -19.205 -35.875 -18.875 ;
        RECT -36.205 -24.645 -35.875 -24.315 ;
        RECT -36.205 -26.005 -35.875 -25.675 ;
        RECT -36.205 -27.365 -35.875 -27.035 ;
        RECT -36.205 -28.725 -35.875 -28.395 ;
        RECT -36.205 -30.085 -35.875 -29.755 ;
        RECT -36.205 -31.445 -35.875 -31.115 ;
        RECT -36.205 -32.805 -35.875 -32.475 ;
        RECT -36.205 -34.165 -35.875 -33.835 ;
        RECT -36.205 -35.525 -35.875 -35.195 ;
        RECT -36.205 -36.885 -35.875 -36.555 ;
        RECT -36.205 -38.245 -35.875 -37.915 ;
        RECT -36.205 -39.605 -35.875 -39.275 ;
        RECT -36.205 -40.965 -35.875 -40.635 ;
        RECT -36.205 -42.325 -35.875 -41.995 ;
        RECT -36.205 -43.685 -35.875 -43.355 ;
        RECT -36.205 -45.045 -35.875 -44.715 ;
        RECT -36.205 -46.405 -35.875 -46.075 ;
        RECT -36.205 -47.765 -35.875 -47.435 ;
        RECT -36.205 -49.125 -35.875 -48.795 ;
        RECT -36.205 -50.485 -35.875 -50.155 ;
        RECT -36.205 -51.845 -35.875 -51.515 ;
        RECT -36.205 -53.205 -35.875 -52.875 ;
        RECT -36.205 -54.565 -35.875 -54.235 ;
        RECT -36.205 -55.925 -35.875 -55.595 ;
        RECT -36.205 -57.285 -35.875 -56.955 ;
        RECT -36.205 -58.645 -35.875 -58.315 ;
        RECT -36.205 -60.005 -35.875 -59.675 ;
        RECT -36.205 -61.365 -35.875 -61.035 ;
        RECT -36.205 -62.725 -35.875 -62.395 ;
        RECT -36.205 -64.085 -35.875 -63.755 ;
        RECT -36.205 -66.805 -35.875 -66.475 ;
        RECT -36.205 -68.165 -35.875 -67.835 ;
        RECT -36.205 -69.525 -35.875 -69.195 ;
        RECT -36.205 -70.885 -35.875 -70.555 ;
        RECT -36.205 -72.245 -35.875 -71.915 ;
        RECT -36.205 -73.83 -35.875 -73.5 ;
        RECT -36.205 -74.965 -35.875 -74.635 ;
        RECT -36.205 -77.685 -35.875 -77.355 ;
        RECT -36.205 -79.045 -35.875 -78.715 ;
        RECT -36.205 -80.405 -35.875 -80.075 ;
        RECT -36.205 -81.97 -35.875 -81.64 ;
        RECT -36.205 -83.125 -35.875 -82.795 ;
        RECT -36.205 -84.485 -35.875 -84.155 ;
        RECT -36.205 -85.845 -35.875 -85.515 ;
        RECT -36.2 -87.88 -35.88 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.205 -149.765 -35.875 -149.435 ;
        RECT -36.205 -150.825 -35.875 -150.495 ;
        RECT -36.205 -152.485 -35.875 -152.155 ;
        RECT -36.205 -153.845 -35.875 -153.515 ;
        RECT -36.205 -156.09 -35.875 -154.96 ;
        RECT -36.2 -156.205 -35.88 -149.435 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.845 42.08 -34.515 43.21 ;
        RECT -34.845 40.635 -34.515 40.965 ;
        RECT -34.845 39.275 -34.515 39.605 ;
        RECT -34.845 37.915 -34.515 38.245 ;
        RECT -34.845 36.555 -34.515 36.885 ;
        RECT -34.845 35.195 -34.515 35.525 ;
        RECT -34.845 33.835 -34.515 34.165 ;
        RECT -34.845 32.475 -34.515 32.805 ;
        RECT -34.845 31.115 -34.515 31.445 ;
        RECT -34.845 29.755 -34.515 30.085 ;
        RECT -34.845 28.395 -34.515 28.725 ;
        RECT -34.845 27.035 -34.515 27.365 ;
        RECT -34.845 25.675 -34.515 26.005 ;
        RECT -34.845 24.315 -34.515 24.645 ;
        RECT -34.845 22.955 -34.515 23.285 ;
        RECT -34.845 21.595 -34.515 21.925 ;
        RECT -34.845 20.235 -34.515 20.565 ;
        RECT -34.845 18.875 -34.515 19.205 ;
        RECT -34.845 17.515 -34.515 17.845 ;
        RECT -34.845 16.155 -34.515 16.485 ;
        RECT -34.845 14.795 -34.515 15.125 ;
        RECT -34.845 13.435 -34.515 13.765 ;
        RECT -34.845 12.075 -34.515 12.405 ;
        RECT -34.845 10.715 -34.515 11.045 ;
        RECT -34.845 9.355 -34.515 9.685 ;
        RECT -34.845 7.995 -34.515 8.325 ;
        RECT -34.845 6.635 -34.515 6.965 ;
        RECT -34.845 5.275 -34.515 5.605 ;
        RECT -34.845 3.915 -34.515 4.245 ;
        RECT -34.845 2.555 -34.515 2.885 ;
        RECT -34.845 -1.525 -34.515 -1.195 ;
        RECT -34.845 -2.885 -34.515 -2.555 ;
        RECT -34.845 -4.245 -34.515 -3.915 ;
        RECT -34.845 -5.605 -34.515 -5.275 ;
        RECT -34.845 -6.965 -34.515 -6.635 ;
        RECT -34.845 -8.325 -34.515 -7.995 ;
        RECT -34.845 -9.685 -34.515 -9.355 ;
        RECT -34.845 -11.045 -34.515 -10.715 ;
        RECT -34.845 -12.405 -34.515 -12.075 ;
        RECT -34.845 -13.765 -34.515 -13.435 ;
        RECT -34.845 -15.125 -34.515 -14.795 ;
        RECT -34.845 -16.485 -34.515 -16.155 ;
        RECT -34.845 -17.845 -34.515 -17.515 ;
        RECT -34.845 -19.205 -34.515 -18.875 ;
        RECT -34.845 -24.645 -34.515 -24.315 ;
        RECT -34.845 -26.005 -34.515 -25.675 ;
        RECT -34.845 -27.365 -34.515 -27.035 ;
        RECT -34.845 -28.725 -34.515 -28.395 ;
        RECT -34.845 -30.085 -34.515 -29.755 ;
        RECT -34.845 -31.445 -34.515 -31.115 ;
        RECT -34.845 -32.805 -34.515 -32.475 ;
        RECT -34.845 -34.165 -34.515 -33.835 ;
        RECT -34.845 -35.525 -34.515 -35.195 ;
        RECT -34.845 -36.885 -34.515 -36.555 ;
        RECT -34.845 -38.245 -34.515 -37.915 ;
        RECT -34.845 -39.605 -34.515 -39.275 ;
        RECT -34.845 -40.965 -34.515 -40.635 ;
        RECT -34.845 -42.325 -34.515 -41.995 ;
        RECT -34.845 -43.685 -34.515 -43.355 ;
        RECT -34.845 -45.045 -34.515 -44.715 ;
        RECT -34.845 -46.405 -34.515 -46.075 ;
        RECT -34.845 -47.765 -34.515 -47.435 ;
        RECT -34.845 -49.125 -34.515 -48.795 ;
        RECT -34.845 -50.485 -34.515 -50.155 ;
        RECT -34.845 -51.845 -34.515 -51.515 ;
        RECT -34.845 -53.205 -34.515 -52.875 ;
        RECT -34.845 -54.565 -34.515 -54.235 ;
        RECT -34.845 -55.925 -34.515 -55.595 ;
        RECT -34.845 -57.285 -34.515 -56.955 ;
        RECT -34.845 -58.645 -34.515 -58.315 ;
        RECT -34.845 -60.005 -34.515 -59.675 ;
        RECT -34.845 -61.365 -34.515 -61.035 ;
        RECT -34.845 -62.725 -34.515 -62.395 ;
        RECT -34.845 -64.085 -34.515 -63.755 ;
        RECT -34.845 -66.805 -34.515 -66.475 ;
        RECT -34.845 -68.165 -34.515 -67.835 ;
        RECT -34.845 -69.525 -34.515 -69.195 ;
        RECT -34.845 -70.885 -34.515 -70.555 ;
        RECT -34.845 -72.245 -34.515 -71.915 ;
        RECT -34.845 -73.83 -34.515 -73.5 ;
        RECT -34.845 -74.965 -34.515 -74.635 ;
        RECT -34.845 -77.685 -34.515 -77.355 ;
        RECT -34.845 -79.045 -34.515 -78.715 ;
        RECT -34.845 -80.405 -34.515 -80.075 ;
        RECT -34.845 -81.97 -34.515 -81.64 ;
        RECT -34.845 -83.125 -34.515 -82.795 ;
        RECT -34.845 -84.485 -34.515 -84.155 ;
        RECT -34.845 -85.845 -34.515 -85.515 ;
        RECT -34.84 -87.2 -34.52 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.845 -149.765 -34.515 -149.435 ;
        RECT -34.845 -150.825 -34.515 -150.495 ;
        RECT -34.845 -152.485 -34.515 -152.155 ;
        RECT -34.845 -153.845 -34.515 -153.515 ;
        RECT -34.845 -156.09 -34.515 -154.96 ;
        RECT -34.84 -156.205 -34.52 -147.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.485 42.08 -33.155 43.21 ;
        RECT -33.485 40.635 -33.155 40.965 ;
        RECT -33.485 39.275 -33.155 39.605 ;
        RECT -33.485 37.915 -33.155 38.245 ;
        RECT -33.485 36.555 -33.155 36.885 ;
        RECT -33.485 35.195 -33.155 35.525 ;
        RECT -33.485 33.835 -33.155 34.165 ;
        RECT -33.485 32.475 -33.155 32.805 ;
        RECT -33.485 31.115 -33.155 31.445 ;
        RECT -33.485 29.755 -33.155 30.085 ;
        RECT -33.485 28.395 -33.155 28.725 ;
        RECT -33.485 27.035 -33.155 27.365 ;
        RECT -33.485 25.675 -33.155 26.005 ;
        RECT -33.485 24.315 -33.155 24.645 ;
        RECT -33.485 22.955 -33.155 23.285 ;
        RECT -33.485 21.595 -33.155 21.925 ;
        RECT -33.485 20.235 -33.155 20.565 ;
        RECT -33.485 18.875 -33.155 19.205 ;
        RECT -33.485 17.515 -33.155 17.845 ;
        RECT -33.485 16.155 -33.155 16.485 ;
        RECT -33.485 14.795 -33.155 15.125 ;
        RECT -33.485 13.435 -33.155 13.765 ;
        RECT -33.485 12.075 -33.155 12.405 ;
        RECT -33.485 10.715 -33.155 11.045 ;
        RECT -33.485 9.355 -33.155 9.685 ;
        RECT -33.485 7.995 -33.155 8.325 ;
        RECT -33.485 6.635 -33.155 6.965 ;
        RECT -33.485 5.275 -33.155 5.605 ;
        RECT -33.485 3.915 -33.155 4.245 ;
        RECT -33.485 2.555 -33.155 2.885 ;
        RECT -33.485 -1.525 -33.155 -1.195 ;
        RECT -33.485 -2.885 -33.155 -2.555 ;
        RECT -33.485 -4.245 -33.155 -3.915 ;
        RECT -33.485 -5.605 -33.155 -5.275 ;
        RECT -33.485 -6.965 -33.155 -6.635 ;
        RECT -33.485 -8.325 -33.155 -7.995 ;
        RECT -33.485 -9.685 -33.155 -9.355 ;
        RECT -33.485 -11.045 -33.155 -10.715 ;
        RECT -33.485 -12.405 -33.155 -12.075 ;
        RECT -33.485 -13.765 -33.155 -13.435 ;
        RECT -33.485 -15.125 -33.155 -14.795 ;
        RECT -33.485 -16.485 -33.155 -16.155 ;
        RECT -33.485 -17.845 -33.155 -17.515 ;
        RECT -33.485 -19.205 -33.155 -18.875 ;
        RECT -33.485 -24.645 -33.155 -24.315 ;
        RECT -33.485 -26.005 -33.155 -25.675 ;
        RECT -33.485 -27.365 -33.155 -27.035 ;
        RECT -33.485 -28.725 -33.155 -28.395 ;
        RECT -33.485 -30.085 -33.155 -29.755 ;
        RECT -33.485 -31.445 -33.155 -31.115 ;
        RECT -33.485 -32.805 -33.155 -32.475 ;
        RECT -33.485 -34.165 -33.155 -33.835 ;
        RECT -33.485 -35.525 -33.155 -35.195 ;
        RECT -33.485 -36.885 -33.155 -36.555 ;
        RECT -33.485 -38.245 -33.155 -37.915 ;
        RECT -33.485 -39.605 -33.155 -39.275 ;
        RECT -33.485 -40.965 -33.155 -40.635 ;
        RECT -33.485 -43.685 -33.155 -43.355 ;
        RECT -33.485 -45.045 -33.155 -44.715 ;
        RECT -33.485 -46.405 -33.155 -46.075 ;
        RECT -33.485 -47.765 -33.155 -47.435 ;
        RECT -33.485 -49.125 -33.155 -48.795 ;
        RECT -33.485 -50.485 -33.155 -50.155 ;
        RECT -33.485 -51.845 -33.155 -51.515 ;
        RECT -33.485 -53.205 -33.155 -52.875 ;
        RECT -33.485 -54.565 -33.155 -54.235 ;
        RECT -33.485 -55.925 -33.155 -55.595 ;
        RECT -33.485 -57.285 -33.155 -56.955 ;
        RECT -33.485 -58.645 -33.155 -58.315 ;
        RECT -33.485 -60.005 -33.155 -59.675 ;
        RECT -33.485 -61.365 -33.155 -61.035 ;
        RECT -33.485 -62.725 -33.155 -62.395 ;
        RECT -33.485 -64.085 -33.155 -63.755 ;
        RECT -33.485 -66.805 -33.155 -66.475 ;
        RECT -33.485 -68.165 -33.155 -67.835 ;
        RECT -33.485 -69.525 -33.155 -69.195 ;
        RECT -33.485 -70.885 -33.155 -70.555 ;
        RECT -33.485 -72.245 -33.155 -71.915 ;
        RECT -33.485 -73.83 -33.155 -73.5 ;
        RECT -33.485 -74.965 -33.155 -74.635 ;
        RECT -33.485 -77.685 -33.155 -77.355 ;
        RECT -33.485 -79.045 -33.155 -78.715 ;
        RECT -33.485 -80.405 -33.155 -80.075 ;
        RECT -33.485 -81.97 -33.155 -81.64 ;
        RECT -33.485 -83.125 -33.155 -82.795 ;
        RECT -33.485 -84.485 -33.155 -84.155 ;
        RECT -33.485 -85.845 -33.155 -85.515 ;
        RECT -33.485 -88.565 -33.155 -88.235 ;
        RECT -33.485 -89.925 -33.155 -89.595 ;
        RECT -33.485 -91.285 -33.155 -90.955 ;
        RECT -33.485 -92.645 -33.155 -92.315 ;
        RECT -33.485 -98.085 -33.155 -97.755 ;
        RECT -33.485 -100.805 -33.155 -100.475 ;
        RECT -33.485 -102.165 -33.155 -101.835 ;
        RECT -33.485 -103.525 -33.155 -103.195 ;
        RECT -33.485 -104.885 -33.155 -104.555 ;
        RECT -33.485 -107.605 -33.155 -107.275 ;
        RECT -33.485 -108.965 -33.155 -108.635 ;
        RECT -33.485 -110.325 -33.155 -109.995 ;
        RECT -33.485 -111.685 -33.155 -111.355 ;
        RECT -33.485 -113.045 -33.155 -112.715 ;
        RECT -33.485 -115.765 -33.155 -115.435 ;
        RECT -33.485 -117.125 -33.155 -116.795 ;
        RECT -33.485 -118.485 -33.155 -118.155 ;
        RECT -33.485 -119.845 -33.155 -119.515 ;
        RECT -33.485 -121.205 -33.155 -120.875 ;
        RECT -33.485 -122.565 -33.155 -122.235 ;
        RECT -33.485 -125.285 -33.155 -124.955 ;
        RECT -33.485 -126.645 -33.155 -126.315 ;
        RECT -33.485 -128.005 -33.155 -127.675 ;
        RECT -33.485 -132.085 -33.155 -131.755 ;
        RECT -33.485 -133.445 -33.155 -133.115 ;
        RECT -33.485 -134.805 -33.155 -134.475 ;
        RECT -33.485 -136.165 -33.155 -135.835 ;
        RECT -33.485 -137.525 -33.155 -137.195 ;
        RECT -33.485 -138.885 -33.155 -138.555 ;
        RECT -33.485 -140.245 -33.155 -139.915 ;
        RECT -33.485 -141.605 -33.155 -141.275 ;
        RECT -33.485 -142.965 -33.155 -142.635 ;
        RECT -33.485 -145.685 -33.155 -145.355 ;
        RECT -33.485 -149.765 -33.155 -149.435 ;
        RECT -33.485 -150.825 -33.155 -150.495 ;
        RECT -33.485 -152.485 -33.155 -152.155 ;
        RECT -33.485 -153.845 -33.155 -153.515 ;
        RECT -33.485 -156.09 -33.155 -154.96 ;
        RECT -33.48 -156.205 -33.16 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.125 24.315 -31.795 24.645 ;
        RECT -32.125 22.955 -31.795 23.285 ;
        RECT -32.125 21.595 -31.795 21.925 ;
        RECT -32.125 20.235 -31.795 20.565 ;
        RECT -32.125 18.875 -31.795 19.205 ;
        RECT -32.125 17.515 -31.795 17.845 ;
        RECT -32.125 16.155 -31.795 16.485 ;
        RECT -32.125 14.795 -31.795 15.125 ;
        RECT -32.125 13.435 -31.795 13.765 ;
        RECT -32.125 12.075 -31.795 12.405 ;
        RECT -32.125 10.715 -31.795 11.045 ;
        RECT -32.125 9.355 -31.795 9.685 ;
        RECT -32.125 7.995 -31.795 8.325 ;
        RECT -32.125 6.635 -31.795 6.965 ;
        RECT -32.125 5.275 -31.795 5.605 ;
        RECT -32.125 3.915 -31.795 4.245 ;
        RECT -32.125 2.555 -31.795 2.885 ;
        RECT -32.125 -1.525 -31.795 -1.195 ;
        RECT -32.125 -2.885 -31.795 -2.555 ;
        RECT -32.125 -4.245 -31.795 -3.915 ;
        RECT -32.125 -5.605 -31.795 -5.275 ;
        RECT -32.125 -6.965 -31.795 -6.635 ;
        RECT -32.125 -8.325 -31.795 -7.995 ;
        RECT -32.125 -9.685 -31.795 -9.355 ;
        RECT -32.125 -11.045 -31.795 -10.715 ;
        RECT -32.125 -12.405 -31.795 -12.075 ;
        RECT -32.125 -13.765 -31.795 -13.435 ;
        RECT -32.125 -15.125 -31.795 -14.795 ;
        RECT -32.125 -16.485 -31.795 -16.155 ;
        RECT -32.125 -17.845 -31.795 -17.515 ;
        RECT -32.125 -19.205 -31.795 -18.875 ;
        RECT -32.125 -24.645 -31.795 -24.315 ;
        RECT -32.125 -26.005 -31.795 -25.675 ;
        RECT -32.125 -27.365 -31.795 -27.035 ;
        RECT -32.125 -28.725 -31.795 -28.395 ;
        RECT -32.125 -30.085 -31.795 -29.755 ;
        RECT -32.125 -31.445 -31.795 -31.115 ;
        RECT -32.125 -32.805 -31.795 -32.475 ;
        RECT -32.125 -34.165 -31.795 -33.835 ;
        RECT -32.125 -35.525 -31.795 -35.195 ;
        RECT -32.125 -36.885 -31.795 -36.555 ;
        RECT -32.125 -38.245 -31.795 -37.915 ;
        RECT -32.125 -39.605 -31.795 -39.275 ;
        RECT -32.125 -40.965 -31.795 -40.635 ;
        RECT -32.125 -43.685 -31.795 -43.355 ;
        RECT -32.125 -45.045 -31.795 -44.715 ;
        RECT -32.125 -46.405 -31.795 -46.075 ;
        RECT -32.125 -47.765 -31.795 -47.435 ;
        RECT -32.125 -49.125 -31.795 -48.795 ;
        RECT -32.125 -50.485 -31.795 -50.155 ;
        RECT -32.125 -51.845 -31.795 -51.515 ;
        RECT -32.125 -53.205 -31.795 -52.875 ;
        RECT -32.125 -54.565 -31.795 -54.235 ;
        RECT -32.125 -55.925 -31.795 -55.595 ;
        RECT -32.125 -57.285 -31.795 -56.955 ;
        RECT -32.125 -58.645 -31.795 -58.315 ;
        RECT -32.125 -60.005 -31.795 -59.675 ;
        RECT -32.125 -61.365 -31.795 -61.035 ;
        RECT -32.125 -62.725 -31.795 -62.395 ;
        RECT -32.125 -64.085 -31.795 -63.755 ;
        RECT -32.125 -66.805 -31.795 -66.475 ;
        RECT -32.125 -68.165 -31.795 -67.835 ;
        RECT -32.125 -69.525 -31.795 -69.195 ;
        RECT -32.125 -70.885 -31.795 -70.555 ;
        RECT -32.125 -72.245 -31.795 -71.915 ;
        RECT -32.125 -73.83 -31.795 -73.5 ;
        RECT -32.125 -74.965 -31.795 -74.635 ;
        RECT -32.125 -77.685 -31.795 -77.355 ;
        RECT -32.125 -79.045 -31.795 -78.715 ;
        RECT -32.125 -80.405 -31.795 -80.075 ;
        RECT -32.125 -81.97 -31.795 -81.64 ;
        RECT -32.125 -83.125 -31.795 -82.795 ;
        RECT -32.125 -84.485 -31.795 -84.155 ;
        RECT -32.125 -85.845 -31.795 -85.515 ;
        RECT -32.125 -88.565 -31.795 -88.235 ;
        RECT -32.125 -89.925 -31.795 -89.595 ;
        RECT -32.125 -91.285 -31.795 -90.955 ;
        RECT -32.125 -92.645 -31.795 -92.315 ;
        RECT -32.125 -98.085 -31.795 -97.755 ;
        RECT -32.125 -100.805 -31.795 -100.475 ;
        RECT -32.125 -102.165 -31.795 -101.835 ;
        RECT -32.125 -103.525 -31.795 -103.195 ;
        RECT -32.125 -104.885 -31.795 -104.555 ;
        RECT -32.125 -107.605 -31.795 -107.275 ;
        RECT -32.125 -108.965 -31.795 -108.635 ;
        RECT -32.125 -110.325 -31.795 -109.995 ;
        RECT -32.125 -111.685 -31.795 -111.355 ;
        RECT -32.125 -115.765 -31.795 -115.435 ;
        RECT -32.125 -117.125 -31.795 -116.795 ;
        RECT -32.125 -118.485 -31.795 -118.155 ;
        RECT -32.125 -119.845 -31.795 -119.515 ;
        RECT -32.125 -121.205 -31.795 -120.875 ;
        RECT -32.125 -122.565 -31.795 -122.235 ;
        RECT -32.125 -125.285 -31.795 -124.955 ;
        RECT -32.125 -126.645 -31.795 -126.315 ;
        RECT -32.125 -128.005 -31.795 -127.675 ;
        RECT -32.125 -132.085 -31.795 -131.755 ;
        RECT -32.125 -133.445 -31.795 -133.115 ;
        RECT -32.125 -134.805 -31.795 -134.475 ;
        RECT -32.125 -136.165 -31.795 -135.835 ;
        RECT -32.125 -137.525 -31.795 -137.195 ;
        RECT -32.125 -138.885 -31.795 -138.555 ;
        RECT -32.125 -140.245 -31.795 -139.915 ;
        RECT -32.125 -141.605 -31.795 -141.275 ;
        RECT -32.125 -142.965 -31.795 -142.635 ;
        RECT -32.125 -145.685 -31.795 -145.355 ;
        RECT -32.125 -147.045 -31.795 -146.715 ;
        RECT -32.125 -148.405 -31.795 -148.075 ;
        RECT -32.125 -149.765 -31.795 -149.435 ;
        RECT -32.125 -150.825 -31.795 -150.495 ;
        RECT -32.125 -152.485 -31.795 -152.155 ;
        RECT -32.125 -153.845 -31.795 -153.515 ;
        RECT -32.125 -156.09 -31.795 -154.96 ;
        RECT -32.12 -156.205 -31.8 43.325 ;
        RECT -32.125 42.08 -31.795 43.21 ;
        RECT -32.125 40.635 -31.795 40.965 ;
        RECT -32.125 39.275 -31.795 39.605 ;
        RECT -32.125 37.915 -31.795 38.245 ;
        RECT -32.125 36.555 -31.795 36.885 ;
        RECT -32.125 35.195 -31.795 35.525 ;
        RECT -32.125 33.835 -31.795 34.165 ;
        RECT -32.125 32.475 -31.795 32.805 ;
        RECT -32.125 31.115 -31.795 31.445 ;
        RECT -32.125 29.755 -31.795 30.085 ;
        RECT -32.125 28.395 -31.795 28.725 ;
        RECT -32.125 27.035 -31.795 27.365 ;
        RECT -32.125 25.675 -31.795 26.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.525 42.08 -52.195 43.21 ;
        RECT -52.525 40.635 -52.195 40.965 ;
        RECT -52.525 39.275 -52.195 39.605 ;
        RECT -52.525 37.915 -52.195 38.245 ;
        RECT -52.525 36.555 -52.195 36.885 ;
        RECT -52.525 35.195 -52.195 35.525 ;
        RECT -52.525 33.835 -52.195 34.165 ;
        RECT -52.525 32.475 -52.195 32.805 ;
        RECT -52.525 31.115 -52.195 31.445 ;
        RECT -52.525 29.755 -52.195 30.085 ;
        RECT -52.525 28.395 -52.195 28.725 ;
        RECT -52.525 27.035 -52.195 27.365 ;
        RECT -52.525 25.675 -52.195 26.005 ;
        RECT -52.525 24.315 -52.195 24.645 ;
        RECT -52.525 23.465 -52.195 23.795 ;
        RECT -52.525 21.415 -52.195 21.745 ;
        RECT -52.525 19.055 -52.195 19.385 ;
        RECT -52.525 17.735 -52.195 18.065 ;
        RECT -52.525 15.545 -52.195 15.875 ;
        RECT -52.525 13.49 -52.195 13.82 ;
        RECT -52.525 12.075 -52.195 12.405 ;
        RECT -52.525 10.715 -52.195 11.045 ;
        RECT -52.525 9.355 -52.195 9.685 ;
        RECT -52.525 7.995 -52.195 8.325 ;
        RECT -52.525 6.635 -52.195 6.965 ;
        RECT -52.525 5.275 -52.195 5.605 ;
        RECT -52.525 3.915 -52.195 4.245 ;
        RECT -52.525 2.555 -52.195 2.885 ;
        RECT -52.525 -0.165 -52.195 0.165 ;
        RECT -52.525 -1.525 -52.195 -1.195 ;
        RECT -52.525 -2.885 -52.195 -2.555 ;
        RECT -52.525 -4.245 -52.195 -3.915 ;
        RECT -52.525 -5.605 -52.195 -5.275 ;
        RECT -52.525 -6.965 -52.195 -6.635 ;
        RECT -52.525 -8.325 -52.195 -7.995 ;
        RECT -52.525 -9.685 -52.195 -9.355 ;
        RECT -52.525 -11.045 -52.195 -10.715 ;
        RECT -52.525 -12.405 -52.195 -12.075 ;
        RECT -52.525 -13.765 -52.195 -13.435 ;
        RECT -52.525 -15.125 -52.195 -14.795 ;
        RECT -52.525 -16.485 -52.195 -16.155 ;
        RECT -52.525 -17.845 -52.195 -17.515 ;
        RECT -52.525 -19.205 -52.195 -18.875 ;
        RECT -52.525 -20.565 -52.195 -20.235 ;
        RECT -52.525 -21.925 -52.195 -21.595 ;
        RECT -52.525 -23.285 -52.195 -22.955 ;
        RECT -52.525 -24.645 -52.195 -24.315 ;
        RECT -52.525 -26.005 -52.195 -25.675 ;
        RECT -52.525 -27.365 -52.195 -27.035 ;
        RECT -52.525 -28.725 -52.195 -28.395 ;
        RECT -52.525 -30.085 -52.195 -29.755 ;
        RECT -52.525 -31.445 -52.195 -31.115 ;
        RECT -52.525 -32.805 -52.195 -32.475 ;
        RECT -52.525 -34.165 -52.195 -33.835 ;
        RECT -52.525 -35.525 -52.195 -35.195 ;
        RECT -52.525 -36.885 -52.195 -36.555 ;
        RECT -52.525 -38.245 -52.195 -37.915 ;
        RECT -52.525 -39.605 -52.195 -39.275 ;
        RECT -52.525 -40.965 -52.195 -40.635 ;
        RECT -52.525 -42.325 -52.195 -41.995 ;
        RECT -52.525 -43.685 -52.195 -43.355 ;
        RECT -52.525 -45.045 -52.195 -44.715 ;
        RECT -52.525 -46.405 -52.195 -46.075 ;
        RECT -52.525 -47.765 -52.195 -47.435 ;
        RECT -52.525 -49.125 -52.195 -48.795 ;
        RECT -52.525 -50.485 -52.195 -50.155 ;
        RECT -52.525 -51.845 -52.195 -51.515 ;
        RECT -52.525 -53.205 -52.195 -52.875 ;
        RECT -52.525 -54.565 -52.195 -54.235 ;
        RECT -52.525 -55.925 -52.195 -55.595 ;
        RECT -52.525 -57.285 -52.195 -56.955 ;
        RECT -52.525 -58.645 -52.195 -58.315 ;
        RECT -52.525 -60.005 -52.195 -59.675 ;
        RECT -52.525 -61.365 -52.195 -61.035 ;
        RECT -52.525 -62.725 -52.195 -62.395 ;
        RECT -52.525 -64.085 -52.195 -63.755 ;
        RECT -52.525 -65.445 -52.195 -65.115 ;
        RECT -52.525 -66.805 -52.195 -66.475 ;
        RECT -52.525 -68.165 -52.195 -67.835 ;
        RECT -52.525 -69.525 -52.195 -69.195 ;
        RECT -52.525 -70.885 -52.195 -70.555 ;
        RECT -52.525 -72.245 -52.195 -71.915 ;
        RECT -52.525 -73.605 -52.195 -73.275 ;
        RECT -52.525 -74.965 -52.195 -74.635 ;
        RECT -52.525 -76.325 -52.195 -75.995 ;
        RECT -52.525 -77.685 -52.195 -77.355 ;
        RECT -52.525 -79.045 -52.195 -78.715 ;
        RECT -52.525 -80.405 -52.195 -80.075 ;
        RECT -52.525 -81.765 -52.195 -81.435 ;
        RECT -52.525 -83.125 -52.195 -82.795 ;
        RECT -52.525 -84.485 -52.195 -84.155 ;
        RECT -52.525 -85.845 -52.195 -85.515 ;
        RECT -52.525 -87.205 -52.195 -86.875 ;
        RECT -52.525 -88.565 -52.195 -88.235 ;
        RECT -52.525 -89.925 -52.195 -89.595 ;
        RECT -52.525 -91.285 -52.195 -90.955 ;
        RECT -52.525 -92.645 -52.195 -92.315 ;
        RECT -52.525 -94.005 -52.195 -93.675 ;
        RECT -52.525 -95.365 -52.195 -95.035 ;
        RECT -52.525 -96.725 -52.195 -96.395 ;
        RECT -52.525 -98.085 -52.195 -97.755 ;
        RECT -52.525 -99.445 -52.195 -99.115 ;
        RECT -52.525 -100.805 -52.195 -100.475 ;
        RECT -52.525 -102.165 -52.195 -101.835 ;
        RECT -52.525 -103.525 -52.195 -103.195 ;
        RECT -52.525 -104.885 -52.195 -104.555 ;
        RECT -52.525 -106.245 -52.195 -105.915 ;
        RECT -52.525 -107.605 -52.195 -107.275 ;
        RECT -52.525 -108.965 -52.195 -108.635 ;
        RECT -52.525 -110.325 -52.195 -109.995 ;
        RECT -52.525 -111.685 -52.195 -111.355 ;
        RECT -52.525 -113.045 -52.195 -112.715 ;
        RECT -52.525 -114.405 -52.195 -114.075 ;
        RECT -52.525 -115.765 -52.195 -115.435 ;
        RECT -52.525 -117.125 -52.195 -116.795 ;
        RECT -52.525 -118.485 -52.195 -118.155 ;
        RECT -52.525 -119.845 -52.195 -119.515 ;
        RECT -52.525 -121.205 -52.195 -120.875 ;
        RECT -52.525 -122.565 -52.195 -122.235 ;
        RECT -52.525 -123.925 -52.195 -123.595 ;
        RECT -52.525 -125.285 -52.195 -124.955 ;
        RECT -52.525 -126.645 -52.195 -126.315 ;
        RECT -52.525 -128.005 -52.195 -127.675 ;
        RECT -52.525 -129.365 -52.195 -129.035 ;
        RECT -52.525 -130.725 -52.195 -130.395 ;
        RECT -52.525 -132.085 -52.195 -131.755 ;
        RECT -52.525 -133.445 -52.195 -133.115 ;
        RECT -52.525 -134.805 -52.195 -134.475 ;
        RECT -52.525 -136.165 -52.195 -135.835 ;
        RECT -52.525 -137.525 -52.195 -137.195 ;
        RECT -52.525 -138.885 -52.195 -138.555 ;
        RECT -52.525 -140.245 -52.195 -139.915 ;
        RECT -52.525 -141.605 -52.195 -141.275 ;
        RECT -52.525 -142.965 -52.195 -142.635 ;
        RECT -52.525 -145.685 -52.195 -145.355 ;
        RECT -52.525 -147.045 -52.195 -146.715 ;
        RECT -52.52 -147.045 -52.2 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.165 42.08 -50.835 43.21 ;
        RECT -51.165 40.635 -50.835 40.965 ;
        RECT -51.165 39.275 -50.835 39.605 ;
        RECT -51.165 37.915 -50.835 38.245 ;
        RECT -51.165 36.555 -50.835 36.885 ;
        RECT -51.165 35.195 -50.835 35.525 ;
        RECT -51.165 33.835 -50.835 34.165 ;
        RECT -51.165 32.475 -50.835 32.805 ;
        RECT -51.165 31.115 -50.835 31.445 ;
        RECT -51.165 29.755 -50.835 30.085 ;
        RECT -51.165 28.395 -50.835 28.725 ;
        RECT -51.165 27.035 -50.835 27.365 ;
        RECT -51.165 25.675 -50.835 26.005 ;
        RECT -51.165 24.315 -50.835 24.645 ;
        RECT -51.16 24.315 -50.84 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.165 12.075 -50.835 12.405 ;
        RECT -51.165 10.715 -50.835 11.045 ;
        RECT -51.165 9.355 -50.835 9.685 ;
        RECT -51.165 7.995 -50.835 8.325 ;
        RECT -51.165 3.915 -50.835 4.245 ;
        RECT -51.165 2.555 -50.835 2.885 ;
        RECT -51.165 -0.165 -50.835 0.165 ;
        RECT -51.165 -1.525 -50.835 -1.195 ;
        RECT -51.165 -2.885 -50.835 -2.555 ;
        RECT -51.165 -4.245 -50.835 -3.915 ;
        RECT -51.165 -5.605 -50.835 -5.275 ;
        RECT -51.165 -6.965 -50.835 -6.635 ;
        RECT -51.165 -8.325 -50.835 -7.995 ;
        RECT -51.165 -9.685 -50.835 -9.355 ;
        RECT -51.165 -11.045 -50.835 -10.715 ;
        RECT -51.165 -12.405 -50.835 -12.075 ;
        RECT -51.165 -13.765 -50.835 -13.435 ;
        RECT -51.165 -15.125 -50.835 -14.795 ;
        RECT -51.165 -16.485 -50.835 -16.155 ;
        RECT -51.165 -17.845 -50.835 -17.515 ;
        RECT -51.165 -19.205 -50.835 -18.875 ;
        RECT -51.165 -20.565 -50.835 -20.235 ;
        RECT -51.165 -21.925 -50.835 -21.595 ;
        RECT -51.165 -23.285 -50.835 -22.955 ;
        RECT -51.165 -24.645 -50.835 -24.315 ;
        RECT -51.165 -26.005 -50.835 -25.675 ;
        RECT -51.165 -27.365 -50.835 -27.035 ;
        RECT -51.165 -28.725 -50.835 -28.395 ;
        RECT -51.165 -30.085 -50.835 -29.755 ;
        RECT -51.165 -31.445 -50.835 -31.115 ;
        RECT -51.165 -32.805 -50.835 -32.475 ;
        RECT -51.165 -34.165 -50.835 -33.835 ;
        RECT -51.165 -35.525 -50.835 -35.195 ;
        RECT -51.165 -36.885 -50.835 -36.555 ;
        RECT -51.165 -38.245 -50.835 -37.915 ;
        RECT -51.165 -39.605 -50.835 -39.275 ;
        RECT -51.165 -40.965 -50.835 -40.635 ;
        RECT -51.165 -42.325 -50.835 -41.995 ;
        RECT -51.165 -43.685 -50.835 -43.355 ;
        RECT -51.165 -45.045 -50.835 -44.715 ;
        RECT -51.165 -46.405 -50.835 -46.075 ;
        RECT -51.165 -47.765 -50.835 -47.435 ;
        RECT -51.165 -49.125 -50.835 -48.795 ;
        RECT -51.165 -50.485 -50.835 -50.155 ;
        RECT -51.165 -51.845 -50.835 -51.515 ;
        RECT -51.165 -53.205 -50.835 -52.875 ;
        RECT -51.165 -54.565 -50.835 -54.235 ;
        RECT -51.165 -55.925 -50.835 -55.595 ;
        RECT -51.165 -57.285 -50.835 -56.955 ;
        RECT -51.165 -58.645 -50.835 -58.315 ;
        RECT -51.165 -60.005 -50.835 -59.675 ;
        RECT -51.165 -61.365 -50.835 -61.035 ;
        RECT -51.165 -62.725 -50.835 -62.395 ;
        RECT -51.165 -64.085 -50.835 -63.755 ;
        RECT -51.165 -65.445 -50.835 -65.115 ;
        RECT -51.165 -66.805 -50.835 -66.475 ;
        RECT -51.165 -68.165 -50.835 -67.835 ;
        RECT -51.165 -69.525 -50.835 -69.195 ;
        RECT -51.165 -70.885 -50.835 -70.555 ;
        RECT -51.165 -72.245 -50.835 -71.915 ;
        RECT -51.165 -73.605 -50.835 -73.275 ;
        RECT -51.165 -74.965 -50.835 -74.635 ;
        RECT -51.165 -76.325 -50.835 -75.995 ;
        RECT -51.165 -77.685 -50.835 -77.355 ;
        RECT -51.165 -79.045 -50.835 -78.715 ;
        RECT -51.165 -80.405 -50.835 -80.075 ;
        RECT -51.165 -81.765 -50.835 -81.435 ;
        RECT -51.165 -83.125 -50.835 -82.795 ;
        RECT -51.165 -84.485 -50.835 -84.155 ;
        RECT -51.165 -85.845 -50.835 -85.515 ;
        RECT -51.165 -87.205 -50.835 -86.875 ;
        RECT -51.165 -88.565 -50.835 -88.235 ;
        RECT -51.165 -89.925 -50.835 -89.595 ;
        RECT -51.165 -91.285 -50.835 -90.955 ;
        RECT -51.165 -92.645 -50.835 -92.315 ;
        RECT -51.165 -94.005 -50.835 -93.675 ;
        RECT -51.165 -95.365 -50.835 -95.035 ;
        RECT -51.165 -98.085 -50.835 -97.755 ;
        RECT -51.165 -99.445 -50.835 -99.115 ;
        RECT -51.165 -100.805 -50.835 -100.475 ;
        RECT -51.165 -102.165 -50.835 -101.835 ;
        RECT -51.165 -103.525 -50.835 -103.195 ;
        RECT -51.165 -104.885 -50.835 -104.555 ;
        RECT -51.165 -106.245 -50.835 -105.915 ;
        RECT -51.165 -107.605 -50.835 -107.275 ;
        RECT -51.165 -108.965 -50.835 -108.635 ;
        RECT -51.165 -110.325 -50.835 -109.995 ;
        RECT -51.165 -111.685 -50.835 -111.355 ;
        RECT -51.165 -113.045 -50.835 -112.715 ;
        RECT -51.165 -114.405 -50.835 -114.075 ;
        RECT -51.165 -115.765 -50.835 -115.435 ;
        RECT -51.165 -117.125 -50.835 -116.795 ;
        RECT -51.165 -118.485 -50.835 -118.155 ;
        RECT -51.165 -119.845 -50.835 -119.515 ;
        RECT -51.165 -121.205 -50.835 -120.875 ;
        RECT -51.165 -122.565 -50.835 -122.235 ;
        RECT -51.165 -123.925 -50.835 -123.595 ;
        RECT -51.165 -125.285 -50.835 -124.955 ;
        RECT -51.165 -126.645 -50.835 -126.315 ;
        RECT -51.165 -128.005 -50.835 -127.675 ;
        RECT -51.165 -129.365 -50.835 -129.035 ;
        RECT -51.165 -130.725 -50.835 -130.395 ;
        RECT -51.165 -132.085 -50.835 -131.755 ;
        RECT -51.165 -133.445 -50.835 -133.115 ;
        RECT -51.165 -134.805 -50.835 -134.475 ;
        RECT -51.165 -136.165 -50.835 -135.835 ;
        RECT -51.165 -137.525 -50.835 -137.195 ;
        RECT -51.165 -138.885 -50.835 -138.555 ;
        RECT -51.165 -140.245 -50.835 -139.915 ;
        RECT -51.165 -141.605 -50.835 -141.275 ;
        RECT -51.165 -142.965 -50.835 -142.635 ;
        RECT -51.165 -145.685 -50.835 -145.355 ;
        RECT -51.165 -148.405 -50.835 -148.075 ;
        RECT -51.165 -149.765 -50.835 -149.435 ;
        RECT -51.165 -150.825 -50.835 -150.495 ;
        RECT -51.165 -152.485 -50.835 -152.155 ;
        RECT -51.165 -153.845 -50.835 -153.515 ;
        RECT -51.165 -156.09 -50.835 -154.96 ;
        RECT -51.16 -156.205 -50.84 12.405 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.805 42.08 -49.475 43.21 ;
        RECT -49.805 40.635 -49.475 40.965 ;
        RECT -49.805 39.275 -49.475 39.605 ;
        RECT -49.805 37.915 -49.475 38.245 ;
        RECT -49.805 36.555 -49.475 36.885 ;
        RECT -49.805 35.195 -49.475 35.525 ;
        RECT -49.805 33.835 -49.475 34.165 ;
        RECT -49.805 32.475 -49.475 32.805 ;
        RECT -49.805 31.115 -49.475 31.445 ;
        RECT -49.805 29.755 -49.475 30.085 ;
        RECT -49.805 28.395 -49.475 28.725 ;
        RECT -49.805 27.035 -49.475 27.365 ;
        RECT -49.805 25.675 -49.475 26.005 ;
        RECT -49.805 24.315 -49.475 24.645 ;
        RECT -49.8 24.315 -49.48 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.805 12.075 -49.475 12.405 ;
        RECT -49.805 10.715 -49.475 11.045 ;
        RECT -49.805 9.355 -49.475 9.685 ;
        RECT -49.805 7.995 -49.475 8.325 ;
        RECT -49.805 3.915 -49.475 4.245 ;
        RECT -49.805 2.555 -49.475 2.885 ;
        RECT -49.805 -0.165 -49.475 0.165 ;
        RECT -49.805 -1.525 -49.475 -1.195 ;
        RECT -49.805 -2.885 -49.475 -2.555 ;
        RECT -49.805 -4.245 -49.475 -3.915 ;
        RECT -49.805 -5.605 -49.475 -5.275 ;
        RECT -49.805 -6.965 -49.475 -6.635 ;
        RECT -49.805 -8.325 -49.475 -7.995 ;
        RECT -49.805 -9.685 -49.475 -9.355 ;
        RECT -49.805 -11.045 -49.475 -10.715 ;
        RECT -49.805 -12.405 -49.475 -12.075 ;
        RECT -49.805 -13.765 -49.475 -13.435 ;
        RECT -49.805 -15.125 -49.475 -14.795 ;
        RECT -49.805 -16.485 -49.475 -16.155 ;
        RECT -49.805 -17.845 -49.475 -17.515 ;
        RECT -49.805 -19.205 -49.475 -18.875 ;
        RECT -49.805 -20.565 -49.475 -20.235 ;
        RECT -49.805 -21.925 -49.475 -21.595 ;
        RECT -49.805 -23.285 -49.475 -22.955 ;
        RECT -49.805 -24.645 -49.475 -24.315 ;
        RECT -49.805 -26.005 -49.475 -25.675 ;
        RECT -49.805 -27.365 -49.475 -27.035 ;
        RECT -49.805 -28.725 -49.475 -28.395 ;
        RECT -49.805 -30.085 -49.475 -29.755 ;
        RECT -49.805 -31.445 -49.475 -31.115 ;
        RECT -49.805 -32.805 -49.475 -32.475 ;
        RECT -49.805 -34.165 -49.475 -33.835 ;
        RECT -49.805 -35.525 -49.475 -35.195 ;
        RECT -49.805 -36.885 -49.475 -36.555 ;
        RECT -49.805 -38.245 -49.475 -37.915 ;
        RECT -49.805 -39.605 -49.475 -39.275 ;
        RECT -49.805 -40.965 -49.475 -40.635 ;
        RECT -49.805 -42.325 -49.475 -41.995 ;
        RECT -49.805 -43.685 -49.475 -43.355 ;
        RECT -49.805 -45.045 -49.475 -44.715 ;
        RECT -49.805 -46.405 -49.475 -46.075 ;
        RECT -49.805 -47.765 -49.475 -47.435 ;
        RECT -49.805 -49.125 -49.475 -48.795 ;
        RECT -49.805 -50.485 -49.475 -50.155 ;
        RECT -49.805 -51.845 -49.475 -51.515 ;
        RECT -49.805 -53.205 -49.475 -52.875 ;
        RECT -49.805 -54.565 -49.475 -54.235 ;
        RECT -49.805 -55.925 -49.475 -55.595 ;
        RECT -49.805 -57.285 -49.475 -56.955 ;
        RECT -49.805 -58.645 -49.475 -58.315 ;
        RECT -49.805 -60.005 -49.475 -59.675 ;
        RECT -49.805 -61.365 -49.475 -61.035 ;
        RECT -49.805 -62.725 -49.475 -62.395 ;
        RECT -49.805 -64.085 -49.475 -63.755 ;
        RECT -49.805 -65.445 -49.475 -65.115 ;
        RECT -49.805 -66.805 -49.475 -66.475 ;
        RECT -49.805 -68.165 -49.475 -67.835 ;
        RECT -49.805 -69.525 -49.475 -69.195 ;
        RECT -49.805 -70.885 -49.475 -70.555 ;
        RECT -49.805 -72.245 -49.475 -71.915 ;
        RECT -49.805 -73.605 -49.475 -73.275 ;
        RECT -49.805 -74.965 -49.475 -74.635 ;
        RECT -49.805 -76.325 -49.475 -75.995 ;
        RECT -49.805 -77.685 -49.475 -77.355 ;
        RECT -49.805 -79.045 -49.475 -78.715 ;
        RECT -49.805 -80.405 -49.475 -80.075 ;
        RECT -49.805 -81.765 -49.475 -81.435 ;
        RECT -49.805 -83.125 -49.475 -82.795 ;
        RECT -49.805 -84.485 -49.475 -84.155 ;
        RECT -49.805 -85.845 -49.475 -85.515 ;
        RECT -49.805 -87.205 -49.475 -86.875 ;
        RECT -49.805 -88.565 -49.475 -88.235 ;
        RECT -49.805 -89.925 -49.475 -89.595 ;
        RECT -49.805 -91.285 -49.475 -90.955 ;
        RECT -49.805 -92.645 -49.475 -92.315 ;
        RECT -49.805 -94.005 -49.475 -93.675 ;
        RECT -49.805 -95.365 -49.475 -95.035 ;
        RECT -49.805 -98.085 -49.475 -97.755 ;
        RECT -49.805 -99.445 -49.475 -99.115 ;
        RECT -49.805 -100.805 -49.475 -100.475 ;
        RECT -49.805 -102.165 -49.475 -101.835 ;
        RECT -49.805 -103.525 -49.475 -103.195 ;
        RECT -49.805 -104.885 -49.475 -104.555 ;
        RECT -49.805 -106.245 -49.475 -105.915 ;
        RECT -49.805 -107.605 -49.475 -107.275 ;
        RECT -49.805 -108.965 -49.475 -108.635 ;
        RECT -49.805 -110.325 -49.475 -109.995 ;
        RECT -49.805 -111.685 -49.475 -111.355 ;
        RECT -49.805 -113.045 -49.475 -112.715 ;
        RECT -49.805 -114.405 -49.475 -114.075 ;
        RECT -49.805 -115.765 -49.475 -115.435 ;
        RECT -49.805 -117.125 -49.475 -116.795 ;
        RECT -49.805 -118.485 -49.475 -118.155 ;
        RECT -49.805 -119.845 -49.475 -119.515 ;
        RECT -49.805 -121.205 -49.475 -120.875 ;
        RECT -49.805 -122.565 -49.475 -122.235 ;
        RECT -49.805 -123.925 -49.475 -123.595 ;
        RECT -49.805 -125.285 -49.475 -124.955 ;
        RECT -49.805 -126.645 -49.475 -126.315 ;
        RECT -49.805 -128.005 -49.475 -127.675 ;
        RECT -49.805 -129.365 -49.475 -129.035 ;
        RECT -49.805 -130.725 -49.475 -130.395 ;
        RECT -49.805 -132.085 -49.475 -131.755 ;
        RECT -49.805 -133.445 -49.475 -133.115 ;
        RECT -49.805 -134.805 -49.475 -134.475 ;
        RECT -49.805 -136.165 -49.475 -135.835 ;
        RECT -49.805 -137.525 -49.475 -137.195 ;
        RECT -49.805 -138.885 -49.475 -138.555 ;
        RECT -49.805 -140.245 -49.475 -139.915 ;
        RECT -49.805 -141.605 -49.475 -141.275 ;
        RECT -49.805 -142.965 -49.475 -142.635 ;
        RECT -49.805 -145.685 -49.475 -145.355 ;
        RECT -49.805 -148.405 -49.475 -148.075 ;
        RECT -49.805 -149.765 -49.475 -149.435 ;
        RECT -49.805 -150.825 -49.475 -150.495 ;
        RECT -49.805 -152.485 -49.475 -152.155 ;
        RECT -49.805 -153.845 -49.475 -153.515 ;
        RECT -49.805 -156.09 -49.475 -154.96 ;
        RECT -49.8 -156.205 -49.48 12.405 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 42.08 -48.115 43.21 ;
        RECT -48.445 40.635 -48.115 40.965 ;
        RECT -48.445 39.275 -48.115 39.605 ;
        RECT -48.445 37.915 -48.115 38.245 ;
        RECT -48.445 36.555 -48.115 36.885 ;
        RECT -48.445 35.195 -48.115 35.525 ;
        RECT -48.445 33.835 -48.115 34.165 ;
        RECT -48.445 32.475 -48.115 32.805 ;
        RECT -48.445 31.115 -48.115 31.445 ;
        RECT -48.445 29.755 -48.115 30.085 ;
        RECT -48.445 28.395 -48.115 28.725 ;
        RECT -48.445 27.035 -48.115 27.365 ;
        RECT -48.445 25.675 -48.115 26.005 ;
        RECT -48.445 24.315 -48.115 24.645 ;
        RECT -48.44 24.315 -48.12 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 12.075 -48.115 12.405 ;
        RECT -48.445 10.715 -48.115 11.045 ;
        RECT -48.445 9.355 -48.115 9.685 ;
        RECT -48.445 7.995 -48.115 8.325 ;
        RECT -48.445 3.915 -48.115 4.245 ;
        RECT -48.445 2.555 -48.115 2.885 ;
        RECT -48.445 -0.165 -48.115 0.165 ;
        RECT -48.445 -1.525 -48.115 -1.195 ;
        RECT -48.445 -2.885 -48.115 -2.555 ;
        RECT -48.445 -4.245 -48.115 -3.915 ;
        RECT -48.445 -5.605 -48.115 -5.275 ;
        RECT -48.445 -6.965 -48.115 -6.635 ;
        RECT -48.445 -8.325 -48.115 -7.995 ;
        RECT -48.445 -9.685 -48.115 -9.355 ;
        RECT -48.445 -11.045 -48.115 -10.715 ;
        RECT -48.445 -12.405 -48.115 -12.075 ;
        RECT -48.445 -13.765 -48.115 -13.435 ;
        RECT -48.445 -15.125 -48.115 -14.795 ;
        RECT -48.445 -16.485 -48.115 -16.155 ;
        RECT -48.445 -17.845 -48.115 -17.515 ;
        RECT -48.445 -19.205 -48.115 -18.875 ;
        RECT -48.445 -20.565 -48.115 -20.235 ;
        RECT -48.445 -21.925 -48.115 -21.595 ;
        RECT -48.445 -23.285 -48.115 -22.955 ;
        RECT -48.445 -24.645 -48.115 -24.315 ;
        RECT -48.445 -26.005 -48.115 -25.675 ;
        RECT -48.445 -27.365 -48.115 -27.035 ;
        RECT -48.445 -28.725 -48.115 -28.395 ;
        RECT -48.445 -30.085 -48.115 -29.755 ;
        RECT -48.445 -31.445 -48.115 -31.115 ;
        RECT -48.445 -32.805 -48.115 -32.475 ;
        RECT -48.445 -34.165 -48.115 -33.835 ;
        RECT -48.445 -35.525 -48.115 -35.195 ;
        RECT -48.445 -36.885 -48.115 -36.555 ;
        RECT -48.445 -38.245 -48.115 -37.915 ;
        RECT -48.445 -39.605 -48.115 -39.275 ;
        RECT -48.445 -40.965 -48.115 -40.635 ;
        RECT -48.445 -42.325 -48.115 -41.995 ;
        RECT -48.445 -43.685 -48.115 -43.355 ;
        RECT -48.445 -45.045 -48.115 -44.715 ;
        RECT -48.445 -46.405 -48.115 -46.075 ;
        RECT -48.445 -47.765 -48.115 -47.435 ;
        RECT -48.445 -49.125 -48.115 -48.795 ;
        RECT -48.445 -50.485 -48.115 -50.155 ;
        RECT -48.445 -51.845 -48.115 -51.515 ;
        RECT -48.445 -53.205 -48.115 -52.875 ;
        RECT -48.445 -54.565 -48.115 -54.235 ;
        RECT -48.445 -55.925 -48.115 -55.595 ;
        RECT -48.445 -57.285 -48.115 -56.955 ;
        RECT -48.445 -58.645 -48.115 -58.315 ;
        RECT -48.445 -60.005 -48.115 -59.675 ;
        RECT -48.445 -61.365 -48.115 -61.035 ;
        RECT -48.445 -62.725 -48.115 -62.395 ;
        RECT -48.445 -64.085 -48.115 -63.755 ;
        RECT -48.445 -65.445 -48.115 -65.115 ;
        RECT -48.445 -66.805 -48.115 -66.475 ;
        RECT -48.445 -68.165 -48.115 -67.835 ;
        RECT -48.445 -69.525 -48.115 -69.195 ;
        RECT -48.445 -70.885 -48.115 -70.555 ;
        RECT -48.445 -72.245 -48.115 -71.915 ;
        RECT -48.445 -73.605 -48.115 -73.275 ;
        RECT -48.445 -74.965 -48.115 -74.635 ;
        RECT -48.445 -76.325 -48.115 -75.995 ;
        RECT -48.445 -77.685 -48.115 -77.355 ;
        RECT -48.445 -79.045 -48.115 -78.715 ;
        RECT -48.445 -80.405 -48.115 -80.075 ;
        RECT -48.445 -81.765 -48.115 -81.435 ;
        RECT -48.445 -83.125 -48.115 -82.795 ;
        RECT -48.445 -84.485 -48.115 -84.155 ;
        RECT -48.445 -85.845 -48.115 -85.515 ;
        RECT -48.445 -87.205 -48.115 -86.875 ;
        RECT -48.44 -87.88 -48.12 12.405 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 -149.765 -48.115 -149.435 ;
        RECT -48.445 -150.825 -48.115 -150.495 ;
        RECT -48.445 -152.485 -48.115 -152.155 ;
        RECT -48.445 -153.845 -48.115 -153.515 ;
        RECT -48.445 -156.09 -48.115 -154.96 ;
        RECT -48.44 -156.205 -48.12 -149.435 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.085 42.08 -46.755 43.21 ;
        RECT -47.085 40.635 -46.755 40.965 ;
        RECT -47.085 39.275 -46.755 39.605 ;
        RECT -47.085 37.915 -46.755 38.245 ;
        RECT -47.085 36.555 -46.755 36.885 ;
        RECT -47.085 35.195 -46.755 35.525 ;
        RECT -47.085 33.835 -46.755 34.165 ;
        RECT -47.085 32.475 -46.755 32.805 ;
        RECT -47.085 31.115 -46.755 31.445 ;
        RECT -47.085 29.755 -46.755 30.085 ;
        RECT -47.085 28.395 -46.755 28.725 ;
        RECT -47.085 27.035 -46.755 27.365 ;
        RECT -47.085 25.675 -46.755 26.005 ;
        RECT -47.085 24.315 -46.755 24.645 ;
        RECT -47.08 24.315 -46.76 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.085 12.075 -46.755 12.405 ;
        RECT -47.085 10.715 -46.755 11.045 ;
        RECT -47.085 9.355 -46.755 9.685 ;
        RECT -47.085 7.995 -46.755 8.325 ;
        RECT -47.085 3.915 -46.755 4.245 ;
        RECT -47.085 2.555 -46.755 2.885 ;
        RECT -47.085 -0.165 -46.755 0.165 ;
        RECT -47.085 -1.525 -46.755 -1.195 ;
        RECT -47.085 -2.885 -46.755 -2.555 ;
        RECT -47.085 -4.245 -46.755 -3.915 ;
        RECT -47.085 -5.605 -46.755 -5.275 ;
        RECT -47.085 -6.965 -46.755 -6.635 ;
        RECT -47.085 -8.325 -46.755 -7.995 ;
        RECT -47.085 -9.685 -46.755 -9.355 ;
        RECT -47.085 -11.045 -46.755 -10.715 ;
        RECT -47.085 -12.405 -46.755 -12.075 ;
        RECT -47.085 -13.765 -46.755 -13.435 ;
        RECT -47.085 -15.125 -46.755 -14.795 ;
        RECT -47.085 -16.485 -46.755 -16.155 ;
        RECT -47.085 -17.845 -46.755 -17.515 ;
        RECT -47.085 -19.205 -46.755 -18.875 ;
        RECT -47.085 -20.565 -46.755 -20.235 ;
        RECT -47.085 -21.925 -46.755 -21.595 ;
        RECT -47.085 -23.285 -46.755 -22.955 ;
        RECT -47.085 -24.645 -46.755 -24.315 ;
        RECT -47.085 -26.005 -46.755 -25.675 ;
        RECT -47.085 -27.365 -46.755 -27.035 ;
        RECT -47.085 -28.725 -46.755 -28.395 ;
        RECT -47.085 -30.085 -46.755 -29.755 ;
        RECT -47.085 -31.445 -46.755 -31.115 ;
        RECT -47.085 -32.805 -46.755 -32.475 ;
        RECT -47.085 -34.165 -46.755 -33.835 ;
        RECT -47.085 -35.525 -46.755 -35.195 ;
        RECT -47.085 -36.885 -46.755 -36.555 ;
        RECT -47.085 -38.245 -46.755 -37.915 ;
        RECT -47.085 -39.605 -46.755 -39.275 ;
        RECT -47.085 -40.965 -46.755 -40.635 ;
        RECT -47.085 -42.325 -46.755 -41.995 ;
        RECT -47.085 -43.685 -46.755 -43.355 ;
        RECT -47.085 -45.045 -46.755 -44.715 ;
        RECT -47.085 -46.405 -46.755 -46.075 ;
        RECT -47.085 -47.765 -46.755 -47.435 ;
        RECT -47.085 -49.125 -46.755 -48.795 ;
        RECT -47.085 -50.485 -46.755 -50.155 ;
        RECT -47.085 -51.845 -46.755 -51.515 ;
        RECT -47.085 -53.205 -46.755 -52.875 ;
        RECT -47.085 -54.565 -46.755 -54.235 ;
        RECT -47.085 -55.925 -46.755 -55.595 ;
        RECT -47.085 -57.285 -46.755 -56.955 ;
        RECT -47.085 -58.645 -46.755 -58.315 ;
        RECT -47.085 -60.005 -46.755 -59.675 ;
        RECT -47.085 -61.365 -46.755 -61.035 ;
        RECT -47.085 -62.725 -46.755 -62.395 ;
        RECT -47.085 -64.085 -46.755 -63.755 ;
        RECT -47.085 -66.805 -46.755 -66.475 ;
        RECT -47.085 -68.165 -46.755 -67.835 ;
        RECT -47.085 -69.525 -46.755 -69.195 ;
        RECT -47.085 -70.885 -46.755 -70.555 ;
        RECT -47.085 -72.245 -46.755 -71.915 ;
        RECT -47.085 -74.965 -46.755 -74.635 ;
        RECT -47.085 -77.685 -46.755 -77.355 ;
        RECT -47.085 -79.045 -46.755 -78.715 ;
        RECT -47.085 -80.405 -46.755 -80.075 ;
        RECT -47.085 -83.125 -46.755 -82.795 ;
        RECT -47.085 -84.485 -46.755 -84.155 ;
        RECT -47.085 -85.845 -46.755 -85.515 ;
        RECT -47.085 -89.925 -46.755 -89.595 ;
        RECT -47.085 -91.285 -46.755 -90.955 ;
        RECT -47.085 -92.645 -46.755 -92.315 ;
        RECT -47.085 -94.005 -46.755 -93.675 ;
        RECT -47.085 -98.085 -46.755 -97.755 ;
        RECT -47.085 -99.445 -46.755 -99.115 ;
        RECT -47.085 -100.805 -46.755 -100.475 ;
        RECT -47.085 -102.165 -46.755 -101.835 ;
        RECT -47.085 -103.525 -46.755 -103.195 ;
        RECT -47.085 -104.885 -46.755 -104.555 ;
        RECT -47.085 -106.245 -46.755 -105.915 ;
        RECT -47.085 -107.605 -46.755 -107.275 ;
        RECT -47.085 -108.965 -46.755 -108.635 ;
        RECT -47.085 -110.325 -46.755 -109.995 ;
        RECT -47.085 -111.685 -46.755 -111.355 ;
        RECT -47.085 -113.045 -46.755 -112.715 ;
        RECT -47.085 -114.405 -46.755 -114.075 ;
        RECT -47.085 -115.765 -46.755 -115.435 ;
        RECT -47.085 -117.125 -46.755 -116.795 ;
        RECT -47.085 -118.485 -46.755 -118.155 ;
        RECT -47.085 -119.845 -46.755 -119.515 ;
        RECT -47.085 -121.205 -46.755 -120.875 ;
        RECT -47.085 -122.565 -46.755 -122.235 ;
        RECT -47.085 -123.925 -46.755 -123.595 ;
        RECT -47.085 -125.285 -46.755 -124.955 ;
        RECT -47.085 -126.645 -46.755 -126.315 ;
        RECT -47.085 -128.005 -46.755 -127.675 ;
        RECT -47.085 -129.365 -46.755 -129.035 ;
        RECT -47.085 -130.725 -46.755 -130.395 ;
        RECT -47.085 -132.085 -46.755 -131.755 ;
        RECT -47.085 -133.445 -46.755 -133.115 ;
        RECT -47.085 -134.805 -46.755 -134.475 ;
        RECT -47.085 -136.165 -46.755 -135.835 ;
        RECT -47.085 -137.525 -46.755 -137.195 ;
        RECT -47.085 -138.885 -46.755 -138.555 ;
        RECT -47.085 -140.245 -46.755 -139.915 ;
        RECT -47.085 -141.605 -46.755 -141.275 ;
        RECT -47.085 -142.965 -46.755 -142.635 ;
        RECT -47.085 -145.685 -46.755 -145.355 ;
        RECT -47.085 -149.765 -46.755 -149.435 ;
        RECT -47.085 -150.825 -46.755 -150.495 ;
        RECT -47.085 -152.485 -46.755 -152.155 ;
        RECT -47.085 -153.845 -46.755 -153.515 ;
        RECT -47.085 -156.09 -46.755 -154.96 ;
        RECT -47.08 -156.205 -46.76 12.405 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.725 42.08 -45.395 43.21 ;
        RECT -45.725 40.635 -45.395 40.965 ;
        RECT -45.725 39.275 -45.395 39.605 ;
        RECT -45.725 37.915 -45.395 38.245 ;
        RECT -45.725 36.555 -45.395 36.885 ;
        RECT -45.725 35.195 -45.395 35.525 ;
        RECT -45.725 33.835 -45.395 34.165 ;
        RECT -45.725 32.475 -45.395 32.805 ;
        RECT -45.725 31.115 -45.395 31.445 ;
        RECT -45.725 29.755 -45.395 30.085 ;
        RECT -45.725 28.395 -45.395 28.725 ;
        RECT -45.725 27.035 -45.395 27.365 ;
        RECT -45.725 25.675 -45.395 26.005 ;
        RECT -45.725 24.315 -45.395 24.645 ;
        RECT -45.72 24.315 -45.4 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.725 12.075 -45.395 12.405 ;
        RECT -45.725 10.715 -45.395 11.045 ;
        RECT -45.725 9.355 -45.395 9.685 ;
        RECT -45.725 7.995 -45.395 8.325 ;
        RECT -45.725 3.915 -45.395 4.245 ;
        RECT -45.725 2.555 -45.395 2.885 ;
        RECT -45.725 -0.165 -45.395 0.165 ;
        RECT -45.725 -1.525 -45.395 -1.195 ;
        RECT -45.725 -2.885 -45.395 -2.555 ;
        RECT -45.725 -4.245 -45.395 -3.915 ;
        RECT -45.725 -5.605 -45.395 -5.275 ;
        RECT -45.725 -6.965 -45.395 -6.635 ;
        RECT -45.725 -8.325 -45.395 -7.995 ;
        RECT -45.725 -9.685 -45.395 -9.355 ;
        RECT -45.725 -11.045 -45.395 -10.715 ;
        RECT -45.725 -12.405 -45.395 -12.075 ;
        RECT -45.725 -13.765 -45.395 -13.435 ;
        RECT -45.725 -15.125 -45.395 -14.795 ;
        RECT -45.725 -16.485 -45.395 -16.155 ;
        RECT -45.725 -17.845 -45.395 -17.515 ;
        RECT -45.725 -19.205 -45.395 -18.875 ;
        RECT -45.725 -20.565 -45.395 -20.235 ;
        RECT -45.725 -21.925 -45.395 -21.595 ;
        RECT -45.725 -23.285 -45.395 -22.955 ;
        RECT -45.725 -24.645 -45.395 -24.315 ;
        RECT -45.725 -26.005 -45.395 -25.675 ;
        RECT -45.725 -27.365 -45.395 -27.035 ;
        RECT -45.725 -28.725 -45.395 -28.395 ;
        RECT -45.725 -30.085 -45.395 -29.755 ;
        RECT -45.725 -31.445 -45.395 -31.115 ;
        RECT -45.725 -32.805 -45.395 -32.475 ;
        RECT -45.725 -34.165 -45.395 -33.835 ;
        RECT -45.725 -35.525 -45.395 -35.195 ;
        RECT -45.725 -36.885 -45.395 -36.555 ;
        RECT -45.725 -38.245 -45.395 -37.915 ;
        RECT -45.725 -39.605 -45.395 -39.275 ;
        RECT -45.725 -40.965 -45.395 -40.635 ;
        RECT -45.725 -42.325 -45.395 -41.995 ;
        RECT -45.725 -43.685 -45.395 -43.355 ;
        RECT -45.725 -45.045 -45.395 -44.715 ;
        RECT -45.725 -46.405 -45.395 -46.075 ;
        RECT -45.725 -47.765 -45.395 -47.435 ;
        RECT -45.725 -49.125 -45.395 -48.795 ;
        RECT -45.725 -50.485 -45.395 -50.155 ;
        RECT -45.725 -51.845 -45.395 -51.515 ;
        RECT -45.725 -53.205 -45.395 -52.875 ;
        RECT -45.725 -54.565 -45.395 -54.235 ;
        RECT -45.725 -55.925 -45.395 -55.595 ;
        RECT -45.725 -57.285 -45.395 -56.955 ;
        RECT -45.725 -58.645 -45.395 -58.315 ;
        RECT -45.725 -60.005 -45.395 -59.675 ;
        RECT -45.725 -61.365 -45.395 -61.035 ;
        RECT -45.725 -62.725 -45.395 -62.395 ;
        RECT -45.725 -64.085 -45.395 -63.755 ;
        RECT -45.725 -66.805 -45.395 -66.475 ;
        RECT -45.725 -68.165 -45.395 -67.835 ;
        RECT -45.725 -69.525 -45.395 -69.195 ;
        RECT -45.725 -70.885 -45.395 -70.555 ;
        RECT -45.725 -72.245 -45.395 -71.915 ;
        RECT -45.725 -73.83 -45.395 -73.5 ;
        RECT -45.725 -74.965 -45.395 -74.635 ;
        RECT -45.725 -77.685 -45.395 -77.355 ;
        RECT -45.725 -79.045 -45.395 -78.715 ;
        RECT -45.725 -80.405 -45.395 -80.075 ;
        RECT -45.725 -81.97 -45.395 -81.64 ;
        RECT -45.725 -83.125 -45.395 -82.795 ;
        RECT -45.725 -84.485 -45.395 -84.155 ;
        RECT -45.725 -85.845 -45.395 -85.515 ;
        RECT -45.725 -89.925 -45.395 -89.595 ;
        RECT -45.725 -91.285 -45.395 -90.955 ;
        RECT -45.725 -92.645 -45.395 -92.315 ;
        RECT -45.725 -94.005 -45.395 -93.675 ;
        RECT -45.725 -98.085 -45.395 -97.755 ;
        RECT -45.725 -99.445 -45.395 -99.115 ;
        RECT -45.725 -100.805 -45.395 -100.475 ;
        RECT -45.725 -102.165 -45.395 -101.835 ;
        RECT -45.725 -103.525 -45.395 -103.195 ;
        RECT -45.725 -104.885 -45.395 -104.555 ;
        RECT -45.725 -106.245 -45.395 -105.915 ;
        RECT -45.725 -107.605 -45.395 -107.275 ;
        RECT -45.725 -108.965 -45.395 -108.635 ;
        RECT -45.725 -110.325 -45.395 -109.995 ;
        RECT -45.725 -111.685 -45.395 -111.355 ;
        RECT -45.725 -113.045 -45.395 -112.715 ;
        RECT -45.725 -114.405 -45.395 -114.075 ;
        RECT -45.725 -115.765 -45.395 -115.435 ;
        RECT -45.725 -117.125 -45.395 -116.795 ;
        RECT -45.725 -118.485 -45.395 -118.155 ;
        RECT -45.725 -119.845 -45.395 -119.515 ;
        RECT -45.725 -121.205 -45.395 -120.875 ;
        RECT -45.725 -122.565 -45.395 -122.235 ;
        RECT -45.725 -123.925 -45.395 -123.595 ;
        RECT -45.725 -125.285 -45.395 -124.955 ;
        RECT -45.725 -126.645 -45.395 -126.315 ;
        RECT -45.725 -128.005 -45.395 -127.675 ;
        RECT -45.725 -129.365 -45.395 -129.035 ;
        RECT -45.725 -130.725 -45.395 -130.395 ;
        RECT -45.725 -132.085 -45.395 -131.755 ;
        RECT -45.725 -133.445 -45.395 -133.115 ;
        RECT -45.725 -134.805 -45.395 -134.475 ;
        RECT -45.725 -136.165 -45.395 -135.835 ;
        RECT -45.725 -137.525 -45.395 -137.195 ;
        RECT -45.725 -138.885 -45.395 -138.555 ;
        RECT -45.725 -140.245 -45.395 -139.915 ;
        RECT -45.725 -141.605 -45.395 -141.275 ;
        RECT -45.72 -141.605 -45.4 12.405 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.725 -148.405 -45.395 -148.075 ;
        RECT -45.725 -149.765 -45.395 -149.435 ;
        RECT -45.725 -150.825 -45.395 -150.495 ;
        RECT -45.725 -152.485 -45.395 -152.155 ;
        RECT -45.725 -153.845 -45.395 -153.515 ;
        RECT -45.725 -156.09 -45.395 -154.96 ;
        RECT -45.72 -156.205 -45.4 -147.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.365 42.08 -44.035 43.21 ;
        RECT -44.365 40.635 -44.035 40.965 ;
        RECT -44.365 39.275 -44.035 39.605 ;
        RECT -44.365 37.915 -44.035 38.245 ;
        RECT -44.365 36.555 -44.035 36.885 ;
        RECT -44.365 35.195 -44.035 35.525 ;
        RECT -44.365 33.835 -44.035 34.165 ;
        RECT -44.365 32.475 -44.035 32.805 ;
        RECT -44.365 31.115 -44.035 31.445 ;
        RECT -44.365 29.755 -44.035 30.085 ;
        RECT -44.365 28.395 -44.035 28.725 ;
        RECT -44.365 27.035 -44.035 27.365 ;
        RECT -44.365 25.675 -44.035 26.005 ;
        RECT -44.365 24.315 -44.035 24.645 ;
        RECT -44.365 23.465 -44.035 23.795 ;
        RECT -44.365 21.415 -44.035 21.745 ;
        RECT -44.365 19.055 -44.035 19.385 ;
        RECT -44.365 17.735 -44.035 18.065 ;
        RECT -44.365 15.545 -44.035 15.875 ;
        RECT -44.365 13.49 -44.035 13.82 ;
        RECT -44.365 12.075 -44.035 12.405 ;
        RECT -44.365 10.715 -44.035 11.045 ;
        RECT -44.365 9.355 -44.035 9.685 ;
        RECT -44.365 7.995 -44.035 8.325 ;
        RECT -44.365 6.635 -44.035 6.965 ;
        RECT -44.365 5.275 -44.035 5.605 ;
        RECT -44.365 3.915 -44.035 4.245 ;
        RECT -44.365 2.555 -44.035 2.885 ;
        RECT -44.365 1.195 -44.035 1.525 ;
        RECT -44.365 -0.165 -44.035 0.165 ;
        RECT -44.365 -1.525 -44.035 -1.195 ;
        RECT -44.365 -2.885 -44.035 -2.555 ;
        RECT -44.365 -4.245 -44.035 -3.915 ;
        RECT -44.365 -5.605 -44.035 -5.275 ;
        RECT -44.365 -6.965 -44.035 -6.635 ;
        RECT -44.365 -8.325 -44.035 -7.995 ;
        RECT -44.365 -9.685 -44.035 -9.355 ;
        RECT -44.365 -11.045 -44.035 -10.715 ;
        RECT -44.365 -12.405 -44.035 -12.075 ;
        RECT -44.365 -13.765 -44.035 -13.435 ;
        RECT -44.365 -15.125 -44.035 -14.795 ;
        RECT -44.365 -16.485 -44.035 -16.155 ;
        RECT -44.365 -17.845 -44.035 -17.515 ;
        RECT -44.365 -19.205 -44.035 -18.875 ;
        RECT -44.365 -20.565 -44.035 -20.235 ;
        RECT -44.365 -21.925 -44.035 -21.595 ;
        RECT -44.365 -23.285 -44.035 -22.955 ;
        RECT -44.365 -24.645 -44.035 -24.315 ;
        RECT -44.365 -26.005 -44.035 -25.675 ;
        RECT -44.365 -27.365 -44.035 -27.035 ;
        RECT -44.365 -28.725 -44.035 -28.395 ;
        RECT -44.365 -30.085 -44.035 -29.755 ;
        RECT -44.365 -31.445 -44.035 -31.115 ;
        RECT -44.365 -32.805 -44.035 -32.475 ;
        RECT -44.365 -34.165 -44.035 -33.835 ;
        RECT -44.365 -35.525 -44.035 -35.195 ;
        RECT -44.365 -36.885 -44.035 -36.555 ;
        RECT -44.365 -38.245 -44.035 -37.915 ;
        RECT -44.365 -39.605 -44.035 -39.275 ;
        RECT -44.365 -40.965 -44.035 -40.635 ;
        RECT -44.365 -42.325 -44.035 -41.995 ;
        RECT -44.365 -43.685 -44.035 -43.355 ;
        RECT -44.365 -45.045 -44.035 -44.715 ;
        RECT -44.365 -46.405 -44.035 -46.075 ;
        RECT -44.365 -47.765 -44.035 -47.435 ;
        RECT -44.365 -49.125 -44.035 -48.795 ;
        RECT -44.365 -50.485 -44.035 -50.155 ;
        RECT -44.365 -51.845 -44.035 -51.515 ;
        RECT -44.365 -53.205 -44.035 -52.875 ;
        RECT -44.365 -54.565 -44.035 -54.235 ;
        RECT -44.365 -55.925 -44.035 -55.595 ;
        RECT -44.365 -57.285 -44.035 -56.955 ;
        RECT -44.365 -58.645 -44.035 -58.315 ;
        RECT -44.365 -60.005 -44.035 -59.675 ;
        RECT -44.365 -61.365 -44.035 -61.035 ;
        RECT -44.365 -62.725 -44.035 -62.395 ;
        RECT -44.365 -64.085 -44.035 -63.755 ;
        RECT -44.365 -66.805 -44.035 -66.475 ;
        RECT -44.365 -68.165 -44.035 -67.835 ;
        RECT -44.365 -69.525 -44.035 -69.195 ;
        RECT -44.365 -70.885 -44.035 -70.555 ;
        RECT -44.365 -72.245 -44.035 -71.915 ;
        RECT -44.365 -73.83 -44.035 -73.5 ;
        RECT -44.365 -74.965 -44.035 -74.635 ;
        RECT -44.365 -77.685 -44.035 -77.355 ;
        RECT -44.365 -79.045 -44.035 -78.715 ;
        RECT -44.365 -80.405 -44.035 -80.075 ;
        RECT -44.365 -81.97 -44.035 -81.64 ;
        RECT -44.365 -83.125 -44.035 -82.795 ;
        RECT -44.365 -84.485 -44.035 -84.155 ;
        RECT -44.365 -85.845 -44.035 -85.515 ;
        RECT -44.365 -89.925 -44.035 -89.595 ;
        RECT -44.365 -91.285 -44.035 -90.955 ;
        RECT -44.365 -92.645 -44.035 -92.315 ;
        RECT -44.365 -98.085 -44.035 -97.755 ;
        RECT -44.365 -99.445 -44.035 -99.115 ;
        RECT -44.365 -100.805 -44.035 -100.475 ;
        RECT -44.365 -102.165 -44.035 -101.835 ;
        RECT -44.365 -103.525 -44.035 -103.195 ;
        RECT -44.365 -104.885 -44.035 -104.555 ;
        RECT -44.365 -106.245 -44.035 -105.915 ;
        RECT -44.365 -107.605 -44.035 -107.275 ;
        RECT -44.365 -108.965 -44.035 -108.635 ;
        RECT -44.365 -110.325 -44.035 -109.995 ;
        RECT -44.365 -111.685 -44.035 -111.355 ;
        RECT -44.365 -113.045 -44.035 -112.715 ;
        RECT -44.365 -114.405 -44.035 -114.075 ;
        RECT -44.365 -115.765 -44.035 -115.435 ;
        RECT -44.365 -117.125 -44.035 -116.795 ;
        RECT -44.365 -118.485 -44.035 -118.155 ;
        RECT -44.365 -119.845 -44.035 -119.515 ;
        RECT -44.365 -121.205 -44.035 -120.875 ;
        RECT -44.365 -122.565 -44.035 -122.235 ;
        RECT -44.365 -123.925 -44.035 -123.595 ;
        RECT -44.365 -125.285 -44.035 -124.955 ;
        RECT -44.365 -126.645 -44.035 -126.315 ;
        RECT -44.365 -128.005 -44.035 -127.675 ;
        RECT -44.365 -129.365 -44.035 -129.035 ;
        RECT -44.365 -130.725 -44.035 -130.395 ;
        RECT -44.365 -132.085 -44.035 -131.755 ;
        RECT -44.365 -133.445 -44.035 -133.115 ;
        RECT -44.365 -134.805 -44.035 -134.475 ;
        RECT -44.365 -136.165 -44.035 -135.835 ;
        RECT -44.365 -137.525 -44.035 -137.195 ;
        RECT -44.365 -138.885 -44.035 -138.555 ;
        RECT -44.365 -140.245 -44.035 -139.915 ;
        RECT -44.365 -141.605 -44.035 -141.275 ;
        RECT -44.365 -142.965 -44.035 -142.635 ;
        RECT -44.365 -145.685 -44.035 -145.355 ;
        RECT -44.365 -147.045 -44.035 -146.715 ;
        RECT -44.365 -148.405 -44.035 -148.075 ;
        RECT -44.365 -149.765 -44.035 -149.435 ;
        RECT -44.365 -150.825 -44.035 -150.495 ;
        RECT -44.365 -152.485 -44.035 -152.155 ;
        RECT -44.365 -153.845 -44.035 -153.515 ;
        RECT -44.365 -156.09 -44.035 -154.96 ;
        RECT -44.36 -156.205 -44.04 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.005 -92.645 -42.675 -92.315 ;
        RECT -43.005 -98.085 -42.675 -97.755 ;
        RECT -43.005 -99.445 -42.675 -99.115 ;
        RECT -43.005 -100.805 -42.675 -100.475 ;
        RECT -43.005 -102.165 -42.675 -101.835 ;
        RECT -43.005 -103.525 -42.675 -103.195 ;
        RECT -43.005 -104.885 -42.675 -104.555 ;
        RECT -43.005 -106.245 -42.675 -105.915 ;
        RECT -43.005 -107.605 -42.675 -107.275 ;
        RECT -43.005 -108.965 -42.675 -108.635 ;
        RECT -43.005 -110.325 -42.675 -109.995 ;
        RECT -43.005 -111.685 -42.675 -111.355 ;
        RECT -43.005 -113.045 -42.675 -112.715 ;
        RECT -43.005 -114.405 -42.675 -114.075 ;
        RECT -43.005 -115.765 -42.675 -115.435 ;
        RECT -43.005 -117.125 -42.675 -116.795 ;
        RECT -43.005 -118.485 -42.675 -118.155 ;
        RECT -43.005 -119.845 -42.675 -119.515 ;
        RECT -43.005 -121.205 -42.675 -120.875 ;
        RECT -43.005 -122.565 -42.675 -122.235 ;
        RECT -43.005 -123.925 -42.675 -123.595 ;
        RECT -43.005 -125.285 -42.675 -124.955 ;
        RECT -43.005 -126.645 -42.675 -126.315 ;
        RECT -43.005 -128.005 -42.675 -127.675 ;
        RECT -43.005 -129.365 -42.675 -129.035 ;
        RECT -43.005 -130.725 -42.675 -130.395 ;
        RECT -43.005 -132.085 -42.675 -131.755 ;
        RECT -43.005 -133.445 -42.675 -133.115 ;
        RECT -43.005 -134.805 -42.675 -134.475 ;
        RECT -43.005 -136.165 -42.675 -135.835 ;
        RECT -43.005 -137.525 -42.675 -137.195 ;
        RECT -43.005 -138.885 -42.675 -138.555 ;
        RECT -43.005 -140.245 -42.675 -139.915 ;
        RECT -43.005 -141.605 -42.675 -141.275 ;
        RECT -43.005 -142.965 -42.675 -142.635 ;
        RECT -43.005 -145.685 -42.675 -145.355 ;
        RECT -43.005 -147.045 -42.675 -146.715 ;
        RECT -43.005 -148.405 -42.675 -148.075 ;
        RECT -43.005 -149.765 -42.675 -149.435 ;
        RECT -43.005 -150.825 -42.675 -150.495 ;
        RECT -43.005 -152.485 -42.675 -152.155 ;
        RECT -43.005 -153.845 -42.675 -153.515 ;
        RECT -43.005 -156.09 -42.675 -154.96 ;
        RECT -43 -156.205 -42.68 43.325 ;
        RECT -43.005 42.08 -42.675 43.21 ;
        RECT -43.005 40.635 -42.675 40.965 ;
        RECT -43.005 39.275 -42.675 39.605 ;
        RECT -43.005 37.915 -42.675 38.245 ;
        RECT -43.005 36.555 -42.675 36.885 ;
        RECT -43.005 35.195 -42.675 35.525 ;
        RECT -43.005 33.835 -42.675 34.165 ;
        RECT -43.005 32.475 -42.675 32.805 ;
        RECT -43.005 31.115 -42.675 31.445 ;
        RECT -43.005 29.755 -42.675 30.085 ;
        RECT -43.005 28.395 -42.675 28.725 ;
        RECT -43.005 27.035 -42.675 27.365 ;
        RECT -43.005 25.675 -42.675 26.005 ;
        RECT -43.005 24.315 -42.675 24.645 ;
        RECT -43.005 23.465 -42.675 23.795 ;
        RECT -43.005 21.415 -42.675 21.745 ;
        RECT -43.005 19.055 -42.675 19.385 ;
        RECT -43.005 17.735 -42.675 18.065 ;
        RECT -43.005 15.545 -42.675 15.875 ;
        RECT -43.005 13.49 -42.675 13.82 ;
        RECT -43.005 12.075 -42.675 12.405 ;
        RECT -43.005 10.715 -42.675 11.045 ;
        RECT -43.005 9.355 -42.675 9.685 ;
        RECT -43.005 7.995 -42.675 8.325 ;
        RECT -43.005 6.635 -42.675 6.965 ;
        RECT -43.005 5.275 -42.675 5.605 ;
        RECT -43.005 3.915 -42.675 4.245 ;
        RECT -43.005 2.555 -42.675 2.885 ;
        RECT -43.005 1.195 -42.675 1.525 ;
        RECT -43.005 -0.165 -42.675 0.165 ;
        RECT -43.005 -1.525 -42.675 -1.195 ;
        RECT -43.005 -2.885 -42.675 -2.555 ;
        RECT -43.005 -4.245 -42.675 -3.915 ;
        RECT -43.005 -5.605 -42.675 -5.275 ;
        RECT -43.005 -6.965 -42.675 -6.635 ;
        RECT -43.005 -8.325 -42.675 -7.995 ;
        RECT -43.005 -9.685 -42.675 -9.355 ;
        RECT -43.005 -11.045 -42.675 -10.715 ;
        RECT -43.005 -12.405 -42.675 -12.075 ;
        RECT -43.005 -13.765 -42.675 -13.435 ;
        RECT -43.005 -15.125 -42.675 -14.795 ;
        RECT -43.005 -16.485 -42.675 -16.155 ;
        RECT -43.005 -17.845 -42.675 -17.515 ;
        RECT -43.005 -19.205 -42.675 -18.875 ;
        RECT -43.005 -21.925 -42.675 -21.595 ;
        RECT -43.005 -23.285 -42.675 -22.955 ;
        RECT -43.005 -24.645 -42.675 -24.315 ;
        RECT -43.005 -26.005 -42.675 -25.675 ;
        RECT -43.005 -27.365 -42.675 -27.035 ;
        RECT -43.005 -28.725 -42.675 -28.395 ;
        RECT -43.005 -30.085 -42.675 -29.755 ;
        RECT -43.005 -31.445 -42.675 -31.115 ;
        RECT -43.005 -32.805 -42.675 -32.475 ;
        RECT -43.005 -34.165 -42.675 -33.835 ;
        RECT -43.005 -35.525 -42.675 -35.195 ;
        RECT -43.005 -36.885 -42.675 -36.555 ;
        RECT -43.005 -38.245 -42.675 -37.915 ;
        RECT -43.005 -39.605 -42.675 -39.275 ;
        RECT -43.005 -40.965 -42.675 -40.635 ;
        RECT -43.005 -42.325 -42.675 -41.995 ;
        RECT -43.005 -43.685 -42.675 -43.355 ;
        RECT -43.005 -45.045 -42.675 -44.715 ;
        RECT -43.005 -46.405 -42.675 -46.075 ;
        RECT -43.005 -47.765 -42.675 -47.435 ;
        RECT -43.005 -49.125 -42.675 -48.795 ;
        RECT -43.005 -50.485 -42.675 -50.155 ;
        RECT -43.005 -51.845 -42.675 -51.515 ;
        RECT -43.005 -53.205 -42.675 -52.875 ;
        RECT -43.005 -54.565 -42.675 -54.235 ;
        RECT -43.005 -55.925 -42.675 -55.595 ;
        RECT -43.005 -57.285 -42.675 -56.955 ;
        RECT -43.005 -58.645 -42.675 -58.315 ;
        RECT -43.005 -60.005 -42.675 -59.675 ;
        RECT -43.005 -61.365 -42.675 -61.035 ;
        RECT -43.005 -62.725 -42.675 -62.395 ;
        RECT -43.005 -64.085 -42.675 -63.755 ;
        RECT -43.005 -66.805 -42.675 -66.475 ;
        RECT -43.005 -68.165 -42.675 -67.835 ;
        RECT -43.005 -69.525 -42.675 -69.195 ;
        RECT -43.005 -70.885 -42.675 -70.555 ;
        RECT -43.005 -72.245 -42.675 -71.915 ;
        RECT -43.005 -73.83 -42.675 -73.5 ;
        RECT -43.005 -74.965 -42.675 -74.635 ;
        RECT -43.005 -77.685 -42.675 -77.355 ;
        RECT -43.005 -79.045 -42.675 -78.715 ;
        RECT -43.005 -80.405 -42.675 -80.075 ;
        RECT -43.005 -81.97 -42.675 -81.64 ;
        RECT -43.005 -83.125 -42.675 -82.795 ;
        RECT -43.005 -84.485 -42.675 -84.155 ;
        RECT -43.005 -85.845 -42.675 -85.515 ;
        RECT -43.005 -89.925 -42.675 -89.595 ;
        RECT -43.005 -91.285 -42.675 -90.955 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.605 42.08 -56.275 43.21 ;
        RECT -56.605 40.635 -56.275 40.965 ;
        RECT -56.605 39.275 -56.275 39.605 ;
        RECT -56.605 37.915 -56.275 38.245 ;
        RECT -56.605 36.555 -56.275 36.885 ;
        RECT -56.605 35.195 -56.275 35.525 ;
        RECT -56.605 33.835 -56.275 34.165 ;
        RECT -56.605 32.475 -56.275 32.805 ;
        RECT -56.605 31.115 -56.275 31.445 ;
        RECT -56.605 29.755 -56.275 30.085 ;
        RECT -56.605 28.395 -56.275 28.725 ;
        RECT -56.605 27.035 -56.275 27.365 ;
        RECT -56.605 25.675 -56.275 26.005 ;
        RECT -56.605 24.315 -56.275 24.645 ;
        RECT -56.605 23.465 -56.275 23.795 ;
        RECT -56.605 21.415 -56.275 21.745 ;
        RECT -56.605 19.055 -56.275 19.385 ;
        RECT -56.605 17.735 -56.275 18.065 ;
        RECT -56.605 15.545 -56.275 15.875 ;
        RECT -56.605 13.49 -56.275 13.82 ;
        RECT -56.605 12.075 -56.275 12.405 ;
        RECT -56.605 10.715 -56.275 11.045 ;
        RECT -56.605 9.355 -56.275 9.685 ;
        RECT -56.605 7.995 -56.275 8.325 ;
        RECT -56.605 6.635 -56.275 6.965 ;
        RECT -56.605 5.275 -56.275 5.605 ;
        RECT -56.605 3.915 -56.275 4.245 ;
        RECT -56.605 2.555 -56.275 2.885 ;
        RECT -56.605 1.195 -56.275 1.525 ;
        RECT -56.605 -0.165 -56.275 0.165 ;
        RECT -56.605 -1.525 -56.275 -1.195 ;
        RECT -56.605 -2.885 -56.275 -2.555 ;
        RECT -56.605 -4.245 -56.275 -3.915 ;
        RECT -56.605 -5.605 -56.275 -5.275 ;
        RECT -56.605 -6.965 -56.275 -6.635 ;
        RECT -56.605 -8.325 -56.275 -7.995 ;
        RECT -56.605 -9.685 -56.275 -9.355 ;
        RECT -56.605 -11.045 -56.275 -10.715 ;
        RECT -56.605 -12.405 -56.275 -12.075 ;
        RECT -56.605 -13.765 -56.275 -13.435 ;
        RECT -56.605 -15.125 -56.275 -14.795 ;
        RECT -56.605 -16.485 -56.275 -16.155 ;
        RECT -56.605 -17.845 -56.275 -17.515 ;
        RECT -56.605 -19.205 -56.275 -18.875 ;
        RECT -56.605 -20.565 -56.275 -20.235 ;
        RECT -56.605 -21.925 -56.275 -21.595 ;
        RECT -56.605 -23.285 -56.275 -22.955 ;
        RECT -56.605 -24.645 -56.275 -24.315 ;
        RECT -56.605 -26.005 -56.275 -25.675 ;
        RECT -56.605 -27.365 -56.275 -27.035 ;
        RECT -56.605 -28.725 -56.275 -28.395 ;
        RECT -56.605 -30.085 -56.275 -29.755 ;
        RECT -56.605 -31.445 -56.275 -31.115 ;
        RECT -56.605 -32.805 -56.275 -32.475 ;
        RECT -56.605 -34.165 -56.275 -33.835 ;
        RECT -56.605 -35.525 -56.275 -35.195 ;
        RECT -56.605 -36.885 -56.275 -36.555 ;
        RECT -56.605 -38.245 -56.275 -37.915 ;
        RECT -56.605 -39.605 -56.275 -39.275 ;
        RECT -56.605 -40.965 -56.275 -40.635 ;
        RECT -56.605 -42.325 -56.275 -41.995 ;
        RECT -56.605 -43.685 -56.275 -43.355 ;
        RECT -56.605 -45.045 -56.275 -44.715 ;
        RECT -56.605 -46.405 -56.275 -46.075 ;
        RECT -56.605 -47.765 -56.275 -47.435 ;
        RECT -56.605 -49.125 -56.275 -48.795 ;
        RECT -56.605 -50.485 -56.275 -50.155 ;
        RECT -56.605 -51.845 -56.275 -51.515 ;
        RECT -56.605 -53.205 -56.275 -52.875 ;
        RECT -56.605 -54.565 -56.275 -54.235 ;
        RECT -56.605 -55.925 -56.275 -55.595 ;
        RECT -56.605 -57.285 -56.275 -56.955 ;
        RECT -56.605 -58.645 -56.275 -58.315 ;
        RECT -56.605 -60.005 -56.275 -59.675 ;
        RECT -56.605 -61.365 -56.275 -61.035 ;
        RECT -56.605 -62.725 -56.275 -62.395 ;
        RECT -56.605 -64.085 -56.275 -63.755 ;
        RECT -56.605 -65.445 -56.275 -65.115 ;
        RECT -56.605 -66.805 -56.275 -66.475 ;
        RECT -56.605 -68.165 -56.275 -67.835 ;
        RECT -56.605 -69.525 -56.275 -69.195 ;
        RECT -56.605 -70.885 -56.275 -70.555 ;
        RECT -56.605 -72.245 -56.275 -71.915 ;
        RECT -56.605 -73.605 -56.275 -73.275 ;
        RECT -56.605 -74.965 -56.275 -74.635 ;
        RECT -56.605 -76.325 -56.275 -75.995 ;
        RECT -56.605 -77.685 -56.275 -77.355 ;
        RECT -56.605 -79.045 -56.275 -78.715 ;
        RECT -56.605 -80.405 -56.275 -80.075 ;
        RECT -56.605 -81.765 -56.275 -81.435 ;
        RECT -56.605 -83.125 -56.275 -82.795 ;
        RECT -56.605 -84.485 -56.275 -84.155 ;
        RECT -56.605 -85.845 -56.275 -85.515 ;
        RECT -56.605 -87.205 -56.275 -86.875 ;
        RECT -56.605 -88.565 -56.275 -88.235 ;
        RECT -56.605 -89.925 -56.275 -89.595 ;
        RECT -56.605 -91.285 -56.275 -90.955 ;
        RECT -56.605 -92.645 -56.275 -92.315 ;
        RECT -56.605 -94.005 -56.275 -93.675 ;
        RECT -56.605 -95.365 -56.275 -95.035 ;
        RECT -56.605 -96.725 -56.275 -96.395 ;
        RECT -56.605 -98.085 -56.275 -97.755 ;
        RECT -56.605 -99.445 -56.275 -99.115 ;
        RECT -56.605 -100.805 -56.275 -100.475 ;
        RECT -56.605 -102.165 -56.275 -101.835 ;
        RECT -56.605 -103.525 -56.275 -103.195 ;
        RECT -56.605 -104.885 -56.275 -104.555 ;
        RECT -56.605 -106.245 -56.275 -105.915 ;
        RECT -56.605 -107.605 -56.275 -107.275 ;
        RECT -56.605 -108.965 -56.275 -108.635 ;
        RECT -56.605 -110.325 -56.275 -109.995 ;
        RECT -56.605 -111.685 -56.275 -111.355 ;
        RECT -56.605 -113.045 -56.275 -112.715 ;
        RECT -56.605 -114.405 -56.275 -114.075 ;
        RECT -56.605 -115.765 -56.275 -115.435 ;
        RECT -56.605 -117.125 -56.275 -116.795 ;
        RECT -56.605 -118.485 -56.275 -118.155 ;
        RECT -56.605 -119.845 -56.275 -119.515 ;
        RECT -56.605 -121.205 -56.275 -120.875 ;
        RECT -56.605 -122.565 -56.275 -122.235 ;
        RECT -56.605 -123.925 -56.275 -123.595 ;
        RECT -56.605 -125.285 -56.275 -124.955 ;
        RECT -56.605 -126.645 -56.275 -126.315 ;
        RECT -56.605 -128.005 -56.275 -127.675 ;
        RECT -56.605 -129.365 -56.275 -129.035 ;
        RECT -56.605 -130.725 -56.275 -130.395 ;
        RECT -56.605 -132.085 -56.275 -131.755 ;
        RECT -56.605 -133.445 -56.275 -133.115 ;
        RECT -56.605 -134.805 -56.275 -134.475 ;
        RECT -56.605 -136.165 -56.275 -135.835 ;
        RECT -56.605 -137.525 -56.275 -137.195 ;
        RECT -56.605 -138.885 -56.275 -138.555 ;
        RECT -56.605 -140.245 -56.275 -139.915 ;
        RECT -56.605 -141.605 -56.275 -141.275 ;
        RECT -56.605 -142.965 -56.275 -142.635 ;
        RECT -56.605 -144.325 -56.275 -143.995 ;
        RECT -56.605 -145.685 -56.275 -145.355 ;
        RECT -56.605 -147.045 -56.275 -146.715 ;
        RECT -56.605 -148.405 -56.275 -148.075 ;
        RECT -56.605 -149.765 -56.275 -149.435 ;
        RECT -56.605 -151.125 -56.275 -150.795 ;
        RECT -56.605 -152.485 -56.275 -152.155 ;
        RECT -56.605 -153.845 -56.275 -153.515 ;
        RECT -56.605 -156.09 -56.275 -154.96 ;
        RECT -56.6 -156.205 -56.28 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.245 42.08 -54.915 43.21 ;
        RECT -55.245 40.635 -54.915 40.965 ;
        RECT -55.245 39.275 -54.915 39.605 ;
        RECT -55.245 37.915 -54.915 38.245 ;
        RECT -55.245 36.555 -54.915 36.885 ;
        RECT -55.245 35.195 -54.915 35.525 ;
        RECT -55.245 33.835 -54.915 34.165 ;
        RECT -55.245 32.475 -54.915 32.805 ;
        RECT -55.245 31.115 -54.915 31.445 ;
        RECT -55.245 29.755 -54.915 30.085 ;
        RECT -55.245 28.395 -54.915 28.725 ;
        RECT -55.245 27.035 -54.915 27.365 ;
        RECT -55.245 25.675 -54.915 26.005 ;
        RECT -55.245 24.315 -54.915 24.645 ;
        RECT -55.245 23.465 -54.915 23.795 ;
        RECT -55.245 21.415 -54.915 21.745 ;
        RECT -55.245 19.055 -54.915 19.385 ;
        RECT -55.245 17.735 -54.915 18.065 ;
        RECT -55.245 15.545 -54.915 15.875 ;
        RECT -55.245 13.49 -54.915 13.82 ;
        RECT -55.245 12.075 -54.915 12.405 ;
        RECT -55.245 10.715 -54.915 11.045 ;
        RECT -55.245 9.355 -54.915 9.685 ;
        RECT -55.245 7.995 -54.915 8.325 ;
        RECT -55.245 6.635 -54.915 6.965 ;
        RECT -55.245 5.275 -54.915 5.605 ;
        RECT -55.245 3.915 -54.915 4.245 ;
        RECT -55.245 2.555 -54.915 2.885 ;
        RECT -55.245 1.195 -54.915 1.525 ;
        RECT -55.245 -0.165 -54.915 0.165 ;
        RECT -55.245 -1.525 -54.915 -1.195 ;
        RECT -55.245 -2.885 -54.915 -2.555 ;
        RECT -55.245 -4.245 -54.915 -3.915 ;
        RECT -55.245 -5.605 -54.915 -5.275 ;
        RECT -55.245 -6.965 -54.915 -6.635 ;
        RECT -55.245 -8.325 -54.915 -7.995 ;
        RECT -55.245 -9.685 -54.915 -9.355 ;
        RECT -55.245 -11.045 -54.915 -10.715 ;
        RECT -55.245 -12.405 -54.915 -12.075 ;
        RECT -55.245 -13.765 -54.915 -13.435 ;
        RECT -55.245 -15.125 -54.915 -14.795 ;
        RECT -55.245 -16.485 -54.915 -16.155 ;
        RECT -55.245 -17.845 -54.915 -17.515 ;
        RECT -55.245 -19.205 -54.915 -18.875 ;
        RECT -55.245 -20.565 -54.915 -20.235 ;
        RECT -55.245 -21.925 -54.915 -21.595 ;
        RECT -55.245 -23.285 -54.915 -22.955 ;
        RECT -55.245 -24.645 -54.915 -24.315 ;
        RECT -55.245 -26.005 -54.915 -25.675 ;
        RECT -55.245 -27.365 -54.915 -27.035 ;
        RECT -55.245 -28.725 -54.915 -28.395 ;
        RECT -55.245 -30.085 -54.915 -29.755 ;
        RECT -55.245 -31.445 -54.915 -31.115 ;
        RECT -55.245 -32.805 -54.915 -32.475 ;
        RECT -55.245 -34.165 -54.915 -33.835 ;
        RECT -55.245 -35.525 -54.915 -35.195 ;
        RECT -55.245 -36.885 -54.915 -36.555 ;
        RECT -55.245 -38.245 -54.915 -37.915 ;
        RECT -55.245 -39.605 -54.915 -39.275 ;
        RECT -55.245 -40.965 -54.915 -40.635 ;
        RECT -55.245 -42.325 -54.915 -41.995 ;
        RECT -55.245 -43.685 -54.915 -43.355 ;
        RECT -55.245 -45.045 -54.915 -44.715 ;
        RECT -55.245 -46.405 -54.915 -46.075 ;
        RECT -55.245 -47.765 -54.915 -47.435 ;
        RECT -55.245 -49.125 -54.915 -48.795 ;
        RECT -55.245 -50.485 -54.915 -50.155 ;
        RECT -55.245 -51.845 -54.915 -51.515 ;
        RECT -55.245 -53.205 -54.915 -52.875 ;
        RECT -55.245 -54.565 -54.915 -54.235 ;
        RECT -55.245 -55.925 -54.915 -55.595 ;
        RECT -55.245 -57.285 -54.915 -56.955 ;
        RECT -55.245 -58.645 -54.915 -58.315 ;
        RECT -55.245 -60.005 -54.915 -59.675 ;
        RECT -55.245 -61.365 -54.915 -61.035 ;
        RECT -55.245 -62.725 -54.915 -62.395 ;
        RECT -55.245 -64.085 -54.915 -63.755 ;
        RECT -55.245 -65.445 -54.915 -65.115 ;
        RECT -55.245 -66.805 -54.915 -66.475 ;
        RECT -55.245 -68.165 -54.915 -67.835 ;
        RECT -55.245 -69.525 -54.915 -69.195 ;
        RECT -55.245 -70.885 -54.915 -70.555 ;
        RECT -55.245 -72.245 -54.915 -71.915 ;
        RECT -55.245 -73.605 -54.915 -73.275 ;
        RECT -55.245 -74.965 -54.915 -74.635 ;
        RECT -55.245 -76.325 -54.915 -75.995 ;
        RECT -55.245 -77.685 -54.915 -77.355 ;
        RECT -55.245 -79.045 -54.915 -78.715 ;
        RECT -55.245 -80.405 -54.915 -80.075 ;
        RECT -55.245 -81.765 -54.915 -81.435 ;
        RECT -55.245 -83.125 -54.915 -82.795 ;
        RECT -55.245 -84.485 -54.915 -84.155 ;
        RECT -55.245 -85.845 -54.915 -85.515 ;
        RECT -55.245 -87.205 -54.915 -86.875 ;
        RECT -55.245 -88.565 -54.915 -88.235 ;
        RECT -55.245 -89.925 -54.915 -89.595 ;
        RECT -55.245 -91.285 -54.915 -90.955 ;
        RECT -55.245 -92.645 -54.915 -92.315 ;
        RECT -55.245 -94.005 -54.915 -93.675 ;
        RECT -55.245 -95.365 -54.915 -95.035 ;
        RECT -55.245 -96.725 -54.915 -96.395 ;
        RECT -55.245 -98.085 -54.915 -97.755 ;
        RECT -55.245 -99.445 -54.915 -99.115 ;
        RECT -55.245 -100.805 -54.915 -100.475 ;
        RECT -55.245 -102.165 -54.915 -101.835 ;
        RECT -55.245 -103.525 -54.915 -103.195 ;
        RECT -55.245 -104.885 -54.915 -104.555 ;
        RECT -55.245 -106.245 -54.915 -105.915 ;
        RECT -55.245 -107.605 -54.915 -107.275 ;
        RECT -55.245 -108.965 -54.915 -108.635 ;
        RECT -55.245 -110.325 -54.915 -109.995 ;
        RECT -55.245 -111.685 -54.915 -111.355 ;
        RECT -55.245 -113.045 -54.915 -112.715 ;
        RECT -55.245 -114.405 -54.915 -114.075 ;
        RECT -55.245 -115.765 -54.915 -115.435 ;
        RECT -55.245 -117.125 -54.915 -116.795 ;
        RECT -55.245 -118.485 -54.915 -118.155 ;
        RECT -55.245 -119.845 -54.915 -119.515 ;
        RECT -55.245 -121.205 -54.915 -120.875 ;
        RECT -55.245 -122.565 -54.915 -122.235 ;
        RECT -55.245 -123.925 -54.915 -123.595 ;
        RECT -55.245 -125.285 -54.915 -124.955 ;
        RECT -55.245 -126.645 -54.915 -126.315 ;
        RECT -55.245 -128.005 -54.915 -127.675 ;
        RECT -55.245 -129.365 -54.915 -129.035 ;
        RECT -55.245 -130.725 -54.915 -130.395 ;
        RECT -55.245 -132.085 -54.915 -131.755 ;
        RECT -55.245 -133.445 -54.915 -133.115 ;
        RECT -55.245 -134.805 -54.915 -134.475 ;
        RECT -55.245 -136.165 -54.915 -135.835 ;
        RECT -55.245 -137.525 -54.915 -137.195 ;
        RECT -55.245 -138.885 -54.915 -138.555 ;
        RECT -55.245 -140.245 -54.915 -139.915 ;
        RECT -55.245 -141.605 -54.915 -141.275 ;
        RECT -55.245 -142.965 -54.915 -142.635 ;
        RECT -55.245 -144.325 -54.915 -143.995 ;
        RECT -55.245 -145.685 -54.915 -145.355 ;
        RECT -55.245 -147.045 -54.915 -146.715 ;
        RECT -55.245 -148.405 -54.915 -148.075 ;
        RECT -55.245 -149.765 -54.915 -149.435 ;
        RECT -55.245 -151.125 -54.915 -150.795 ;
        RECT -55.245 -152.485 -54.915 -152.155 ;
        RECT -55.245 -153.845 -54.915 -153.515 ;
        RECT -55.245 -156.09 -54.915 -154.96 ;
        RECT -55.24 -156.205 -54.92 43.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.885 -51.845 -53.555 -51.515 ;
        RECT -53.885 -53.205 -53.555 -52.875 ;
        RECT -53.885 -54.565 -53.555 -54.235 ;
        RECT -53.885 -55.925 -53.555 -55.595 ;
        RECT -53.885 -57.285 -53.555 -56.955 ;
        RECT -53.885 -58.645 -53.555 -58.315 ;
        RECT -53.885 -60.005 -53.555 -59.675 ;
        RECT -53.885 -61.365 -53.555 -61.035 ;
        RECT -53.885 -62.725 -53.555 -62.395 ;
        RECT -53.885 -64.085 -53.555 -63.755 ;
        RECT -53.885 -65.445 -53.555 -65.115 ;
        RECT -53.885 -66.805 -53.555 -66.475 ;
        RECT -53.885 -68.165 -53.555 -67.835 ;
        RECT -53.885 -69.525 -53.555 -69.195 ;
        RECT -53.885 -70.885 -53.555 -70.555 ;
        RECT -53.885 -72.245 -53.555 -71.915 ;
        RECT -53.885 -73.605 -53.555 -73.275 ;
        RECT -53.885 -74.965 -53.555 -74.635 ;
        RECT -53.885 -76.325 -53.555 -75.995 ;
        RECT -53.885 -77.685 -53.555 -77.355 ;
        RECT -53.885 -79.045 -53.555 -78.715 ;
        RECT -53.885 -80.405 -53.555 -80.075 ;
        RECT -53.885 -81.765 -53.555 -81.435 ;
        RECT -53.885 -83.125 -53.555 -82.795 ;
        RECT -53.885 -84.485 -53.555 -84.155 ;
        RECT -53.885 -85.845 -53.555 -85.515 ;
        RECT -53.885 -87.205 -53.555 -86.875 ;
        RECT -53.885 -88.565 -53.555 -88.235 ;
        RECT -53.885 -89.925 -53.555 -89.595 ;
        RECT -53.885 -91.285 -53.555 -90.955 ;
        RECT -53.885 -92.645 -53.555 -92.315 ;
        RECT -53.885 -94.005 -53.555 -93.675 ;
        RECT -53.885 -95.365 -53.555 -95.035 ;
        RECT -53.885 -96.725 -53.555 -96.395 ;
        RECT -53.885 -98.085 -53.555 -97.755 ;
        RECT -53.885 -99.445 -53.555 -99.115 ;
        RECT -53.885 -100.805 -53.555 -100.475 ;
        RECT -53.885 -102.165 -53.555 -101.835 ;
        RECT -53.885 -103.525 -53.555 -103.195 ;
        RECT -53.885 -104.885 -53.555 -104.555 ;
        RECT -53.885 -106.245 -53.555 -105.915 ;
        RECT -53.885 -107.605 -53.555 -107.275 ;
        RECT -53.885 -108.965 -53.555 -108.635 ;
        RECT -53.885 -110.325 -53.555 -109.995 ;
        RECT -53.885 -111.685 -53.555 -111.355 ;
        RECT -53.885 -113.045 -53.555 -112.715 ;
        RECT -53.885 -114.405 -53.555 -114.075 ;
        RECT -53.885 -115.765 -53.555 -115.435 ;
        RECT -53.885 -117.125 -53.555 -116.795 ;
        RECT -53.885 -118.485 -53.555 -118.155 ;
        RECT -53.885 -119.845 -53.555 -119.515 ;
        RECT -53.885 -121.205 -53.555 -120.875 ;
        RECT -53.885 -122.565 -53.555 -122.235 ;
        RECT -53.885 -123.925 -53.555 -123.595 ;
        RECT -53.885 -125.285 -53.555 -124.955 ;
        RECT -53.885 -126.645 -53.555 -126.315 ;
        RECT -53.885 -128.005 -53.555 -127.675 ;
        RECT -53.885 -129.365 -53.555 -129.035 ;
        RECT -53.885 -130.725 -53.555 -130.395 ;
        RECT -53.885 -132.085 -53.555 -131.755 ;
        RECT -53.885 -133.445 -53.555 -133.115 ;
        RECT -53.885 -134.805 -53.555 -134.475 ;
        RECT -53.885 -136.165 -53.555 -135.835 ;
        RECT -53.885 -137.525 -53.555 -137.195 ;
        RECT -53.885 -138.885 -53.555 -138.555 ;
        RECT -53.885 -140.245 -53.555 -139.915 ;
        RECT -53.885 -141.605 -53.555 -141.275 ;
        RECT -53.885 -142.965 -53.555 -142.635 ;
        RECT -53.885 -145.685 -53.555 -145.355 ;
        RECT -53.885 -147.045 -53.555 -146.715 ;
        RECT -53.885 -148.405 -53.555 -148.075 ;
        RECT -53.885 -149.765 -53.555 -149.435 ;
        RECT -53.885 -152.485 -53.555 -152.155 ;
        RECT -53.885 -153.845 -53.555 -153.515 ;
        RECT -53.885 -156.09 -53.555 -154.96 ;
        RECT -53.88 -156.205 -53.56 43.325 ;
        RECT -53.885 42.08 -53.555 43.21 ;
        RECT -53.885 40.635 -53.555 40.965 ;
        RECT -53.885 39.275 -53.555 39.605 ;
        RECT -53.885 37.915 -53.555 38.245 ;
        RECT -53.885 36.555 -53.555 36.885 ;
        RECT -53.885 35.195 -53.555 35.525 ;
        RECT -53.885 33.835 -53.555 34.165 ;
        RECT -53.885 32.475 -53.555 32.805 ;
        RECT -53.885 31.115 -53.555 31.445 ;
        RECT -53.885 29.755 -53.555 30.085 ;
        RECT -53.885 28.395 -53.555 28.725 ;
        RECT -53.885 27.035 -53.555 27.365 ;
        RECT -53.885 25.675 -53.555 26.005 ;
        RECT -53.885 24.315 -53.555 24.645 ;
        RECT -53.885 23.465 -53.555 23.795 ;
        RECT -53.885 21.415 -53.555 21.745 ;
        RECT -53.885 19.055 -53.555 19.385 ;
        RECT -53.885 17.735 -53.555 18.065 ;
        RECT -53.885 15.545 -53.555 15.875 ;
        RECT -53.885 13.49 -53.555 13.82 ;
        RECT -53.885 12.075 -53.555 12.405 ;
        RECT -53.885 10.715 -53.555 11.045 ;
        RECT -53.885 9.355 -53.555 9.685 ;
        RECT -53.885 7.995 -53.555 8.325 ;
        RECT -53.885 6.635 -53.555 6.965 ;
        RECT -53.885 5.275 -53.555 5.605 ;
        RECT -53.885 3.915 -53.555 4.245 ;
        RECT -53.885 2.555 -53.555 2.885 ;
        RECT -53.885 1.195 -53.555 1.525 ;
        RECT -53.885 -0.165 -53.555 0.165 ;
        RECT -53.885 -1.525 -53.555 -1.195 ;
        RECT -53.885 -2.885 -53.555 -2.555 ;
        RECT -53.885 -4.245 -53.555 -3.915 ;
        RECT -53.885 -5.605 -53.555 -5.275 ;
        RECT -53.885 -6.965 -53.555 -6.635 ;
        RECT -53.885 -8.325 -53.555 -7.995 ;
        RECT -53.885 -9.685 -53.555 -9.355 ;
        RECT -53.885 -11.045 -53.555 -10.715 ;
        RECT -53.885 -12.405 -53.555 -12.075 ;
        RECT -53.885 -13.765 -53.555 -13.435 ;
        RECT -53.885 -15.125 -53.555 -14.795 ;
        RECT -53.885 -16.485 -53.555 -16.155 ;
        RECT -53.885 -17.845 -53.555 -17.515 ;
        RECT -53.885 -19.205 -53.555 -18.875 ;
        RECT -53.885 -20.565 -53.555 -20.235 ;
        RECT -53.885 -21.925 -53.555 -21.595 ;
        RECT -53.885 -23.285 -53.555 -22.955 ;
        RECT -53.885 -24.645 -53.555 -24.315 ;
        RECT -53.885 -26.005 -53.555 -25.675 ;
        RECT -53.885 -27.365 -53.555 -27.035 ;
        RECT -53.885 -28.725 -53.555 -28.395 ;
        RECT -53.885 -30.085 -53.555 -29.755 ;
        RECT -53.885 -31.445 -53.555 -31.115 ;
        RECT -53.885 -32.805 -53.555 -32.475 ;
        RECT -53.885 -34.165 -53.555 -33.835 ;
        RECT -53.885 -35.525 -53.555 -35.195 ;
        RECT -53.885 -36.885 -53.555 -36.555 ;
        RECT -53.885 -38.245 -53.555 -37.915 ;
        RECT -53.885 -39.605 -53.555 -39.275 ;
        RECT -53.885 -40.965 -53.555 -40.635 ;
        RECT -53.885 -42.325 -53.555 -41.995 ;
        RECT -53.885 -43.685 -53.555 -43.355 ;
        RECT -53.885 -45.045 -53.555 -44.715 ;
        RECT -53.885 -46.405 -53.555 -46.075 ;
        RECT -53.885 -47.765 -53.555 -47.435 ;
        RECT -53.885 -49.125 -53.555 -48.795 ;
        RECT -53.885 -50.485 -53.555 -50.155 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -21.92 -159.085 -21.6 -158.765 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -28.04 -159.085 -27.72 -158.765 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -34.16 -159.085 -33.84 -158.765 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -40.28 -159.085 -39.96 -158.765 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -46.4 -159.085 -46.08 -158.765 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -52.52 -159.085 -52.2 -158.765 ;
    END
  END addr[5]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -9.68 -159.085 -9.36 -158.765 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.6 -159.085 6 -158.685 ;
    END
  END din[0]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 11.7 -159.085 12.1 -158.685 ;
    END
  END din[1]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 17.8 -159.085 18.2 -158.685 ;
    END
  END din[2]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 23.9 -159.085 24.3 -158.685 ;
    END
  END din[3]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4 -159.085 4.4 -158.685 ;
    END
  END dout[0]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 10.1 -159.085 10.5 -158.685 ;
    END
  END dout[1]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 16.2 -159.085 16.6 -158.685 ;
    END
  END dout[2]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 22.3 -159.085 22.7 -158.685 ;
    END
  END dout[3]
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -15.8 -159.085 -15.48 -158.765 ;
    END
  END we
  PIN wmask[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 6.4 -159.085 6.8 -158.685 ;
    END
  END wmask[0]
  PIN wmask[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 18.6 -159.085 19 -158.685 ;
    END
  END wmask[1]
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -61.96 -159.085 42.145 46.205 ;
    LAYER met2 SPACING 0.14 ;
      RECT -61.96 -159.085 42.145 46.205 ;
    LAYER met3 SPACING 0.3 ;
      RECT 0.515 -35.525 0.845 -35.195 ;
      RECT 0.52 -44.365 0.84 -35.195 ;
      RECT 0.515 -44.365 0.845 -44.035 ;
      RECT -0.165 -34.165 0.165 -33.835 ;
      RECT -0.16 -41.645 0.16 -33.835 ;
      RECT -0.165 -41.645 0.165 -41.315 ;
      RECT -9.005 -9.005 -8.675 -8.675 ;
      RECT -9 -96.725 -8.68 -8.675 ;
      RECT -9.005 -11.045 -8.675 -10.715 ;
      RECT -9.005 -96.725 -8.675 -96.395 ;
      RECT -9.685 -142.285 -9.355 -141.955 ;
      RECT -9.68 -158.275 -9.36 -141.955 ;
      RECT -9.685 -86.525 -9.355 -86.195 ;
      RECT -9.68 -133.445 -9.36 -86.195 ;
      RECT -9.685 -133.445 -9.355 -133.115 ;
      RECT -9.685 -19.205 -9.355 -18.875 ;
      RECT -9.68 -76.325 -9.36 -18.875 ;
      RECT -9.685 -76.325 -9.355 -75.995 ;
      RECT -11.045 -142.965 -10.715 -142.635 ;
      RECT -11.04 -147.725 -10.72 -142.635 ;
      RECT -11.045 -147.725 -10.715 -147.395 ;
      RECT -13.085 -19.885 -12.755 -19.555 ;
      RECT -13.08 -83.805 -12.76 -19.555 ;
      RECT -13.085 -83.805 -12.755 -83.475 ;
      RECT -13.765 -20.565 -13.435 -20.235 ;
      RECT -13.76 -76.325 -13.44 -20.235 ;
      RECT -13.765 -76.325 -13.435 -75.995 ;
      RECT -14.445 -142.285 -14.115 -141.955 ;
      RECT -14.44 -147.045 -14.12 -141.955 ;
      RECT -14.445 -147.045 -14.115 -146.715 ;
      RECT -14.445 -85.23 -14.115 -84.9 ;
      RECT -14.44 -87.885 -14.12 -84.9 ;
      RECT -14.445 -87.885 -14.115 -87.555 ;
      RECT -14.445 -39.43 -14.115 -39.1 ;
      RECT -14.44 -41.645 -14.12 -39.1 ;
      RECT -14.445 -41.645 -14.115 -41.315 ;
      RECT -14.445 -17.41 -14.115 -17.08 ;
      RECT -14.44 -19.885 -14.12 -17.08 ;
      RECT -14.445 -19.885 -14.115 -19.555 ;
      RECT -15.125 -85.71 -14.795 -85.38 ;
      RECT -15.12 -88.565 -14.8 -85.38 ;
      RECT -15.125 -88.565 -14.795 -88.235 ;
      RECT -15.125 -39.91 -14.795 -39.58 ;
      RECT -15.12 -42.325 -14.8 -39.58 ;
      RECT -15.125 -42.325 -14.795 -41.995 ;
      RECT -15.125 -17.89 -14.795 -17.56 ;
      RECT -15.12 -20.565 -14.8 -17.56 ;
      RECT -15.125 -20.565 -14.795 -20.235 ;
      RECT -15.8 -158.275 -15.48 -147.4 ;
      RECT -15.805 -147.85 -15.475 -147.52 ;
      RECT -15.805 -86.19 -15.475 -85.86 ;
      RECT -15.8 -89.245 -15.48 -85.86 ;
      RECT -15.805 -89.245 -15.475 -88.915 ;
      RECT -15.805 -40.39 -15.475 -40.06 ;
      RECT -15.8 -43.005 -15.48 -40.06 ;
      RECT -15.805 -43.005 -15.475 -42.675 ;
      RECT -15.805 -18.37 -15.475 -18.04 ;
      RECT -15.8 -21.245 -15.48 -18.04 ;
      RECT -15.805 -21.245 -15.475 -20.915 ;
      RECT -16.485 -86.67 -16.155 -86.34 ;
      RECT -16.48 -149.085 -16.16 -86.34 ;
      RECT -16.485 -149.085 -16.155 -148.755 ;
      RECT -16.485 -40.87 -16.155 -40.54 ;
      RECT -16.48 -43.685 -16.16 -40.54 ;
      RECT -16.485 -43.685 -16.155 -43.355 ;
      RECT -16.485 -18.85 -16.155 -18.52 ;
      RECT -16.48 -21.925 -16.16 -18.52 ;
      RECT -16.485 -21.925 -16.155 -21.595 ;
      RECT -17.165 -89.245 -16.835 -88.915 ;
      RECT -17.16 -147.045 -16.84 -88.915 ;
      RECT -17.165 -147.045 -16.835 -146.715 ;
      RECT -18.525 -88.565 -18.195 -88.235 ;
      RECT -18.52 -149.085 -18.2 -88.235 ;
      RECT -18.525 -149.085 -18.195 -148.755 ;
      RECT -19.205 -32.805 -18.875 -32.475 ;
      RECT -19.2 -96.045 -18.88 -32.475 ;
      RECT -19.205 -96.045 -18.875 -95.715 ;
      RECT -20.565 -142.285 -20.235 -141.955 ;
      RECT -20.56 -147.045 -20.24 -141.955 ;
      RECT -20.565 -147.045 -20.235 -146.715 ;
      RECT -21.245 -63.405 -20.915 -63.075 ;
      RECT -21.24 -94.685 -20.92 -63.075 ;
      RECT -21.245 -94.685 -20.915 -94.355 ;
      RECT -21.92 -158.275 -21.6 -147.4 ;
      RECT -21.925 -147.85 -21.595 -147.52 ;
      RECT -23.285 -87.885 -22.955 -87.555 ;
      RECT -23.28 -147.045 -22.96 -87.555 ;
      RECT -23.285 -147.045 -22.955 -146.715 ;
      RECT -26.685 -142.285 -26.355 -141.955 ;
      RECT -26.68 -147.045 -26.36 -141.955 ;
      RECT -26.685 -147.045 -26.355 -146.715 ;
      RECT -28.04 -158.275 -27.72 -147.4 ;
      RECT -28.045 -147.85 -27.715 -147.52 ;
      RECT -29.405 -87.885 -29.075 -87.555 ;
      RECT -29.4 -147.045 -29.08 -87.555 ;
      RECT -29.405 -147.045 -29.075 -146.715 ;
      RECT -30.085 -88.565 -29.755 -88.235 ;
      RECT -30.08 -149.085 -29.76 -88.235 ;
      RECT -30.085 -149.085 -29.755 -148.755 ;
      RECT -32.805 -142.285 -32.475 -141.955 ;
      RECT -32.8 -147.045 -32.48 -141.955 ;
      RECT -32.805 -147.045 -32.475 -146.715 ;
      RECT -34.16 -158.275 -33.84 -147.4 ;
      RECT -34.165 -147.85 -33.835 -147.52 ;
      RECT -34.845 -87.885 -34.515 -87.555 ;
      RECT -34.84 -147.045 -34.52 -87.555 ;
      RECT -34.845 -147.045 -34.515 -146.715 ;
      RECT -36.205 -88.565 -35.875 -88.235 ;
      RECT -36.2 -149.085 -35.88 -88.235 ;
      RECT -36.205 -149.085 -35.875 -148.755 ;
      RECT -38.925 -142.285 -38.595 -141.955 ;
      RECT -38.92 -147.045 -38.6 -141.955 ;
      RECT -38.925 -147.045 -38.595 -146.715 ;
      RECT -40.28 -158.275 -39.96 -147.4 ;
      RECT -40.285 -147.85 -39.955 -147.52 ;
      RECT -40.285 -87.885 -39.955 -87.555 ;
      RECT -40.28 -147.045 -39.96 -87.555 ;
      RECT -40.285 -147.045 -39.955 -146.715 ;
      RECT -42.325 -88.565 -41.995 -88.235 ;
      RECT -42.32 -149.085 -42 -88.235 ;
      RECT -42.325 -149.085 -41.995 -148.755 ;
      RECT -46 18.18 -44.72 18.77 ;
      RECT -45.04 -94.005 -44.72 18.77 ;
      RECT -45.045 -94.005 -44.715 -93.675 ;
      RECT -45.725 -142.285 -45.395 -141.955 ;
      RECT -45.72 -147.045 -45.4 -141.955 ;
      RECT -45.725 -147.045 -45.395 -146.715 ;
      RECT -46.4 -158.275 -46.08 -147.4 ;
      RECT -46.405 -147.85 -46.075 -147.52 ;
      RECT -46.405 -87.885 -46.075 -87.555 ;
      RECT -46.4 -147.045 -46.08 -87.555 ;
      RECT -46.405 -147.045 -46.075 -146.715 ;
      RECT -47.765 -87.205 -47.435 -86.875 ;
      RECT -47.76 -95.365 -47.44 -86.875 ;
      RECT -47.765 -95.365 -47.435 -95.035 ;
      RECT -48.445 -88.565 -48.115 -88.235 ;
      RECT -48.44 -149.085 -48.12 -88.235 ;
      RECT -48.445 -149.085 -48.115 -148.755 ;
      RECT -49.125 -142.285 -48.795 -141.955 ;
      RECT -49.12 -147.045 -48.8 -141.955 ;
      RECT -49.125 -147.045 -48.795 -146.715 ;
      RECT -51.845 1.875 -51.515 2.205 ;
      RECT -51.84 -9.005 -51.52 2.205 ;
      RECT -51.845 -9.005 -51.515 -8.675 ;
      RECT -52.52 -158.275 -52.2 -147.4 ;
      RECT -52.525 -147.85 -52.195 -147.52 ;
      RECT 25.5 -80.215 25.9 -20.12 ;
      RECT 24.7 -79.355 25.1 -20.12 ;
      RECT 23.9 -158.195 24.3 -79.445 ;
      RECT 23.1 -63.5 23.5 -48.905 ;
      RECT 23.1 -45.08 23.5 -15.74 ;
      RECT 22.3 -158.195 22.7 -73.605 ;
      RECT 22.3 -64 22.7 -49.36 ;
      RECT 22.3 -45.51 22.7 -12.47 ;
      RECT 20.2 -87.06 20.6 -20.12 ;
      RECT 19.4 -80.215 19.8 -20.12 ;
      RECT 18.6 -158.195 19 -87.15 ;
      RECT 18.6 -79.355 19 -20.12 ;
      RECT 17.8 -158.195 18.2 -79.445 ;
      RECT 17 -63.5 17.4 -48.905 ;
      RECT 17 -45.08 17.4 -15.74 ;
      RECT 16.2 -158.195 16.6 -73.605 ;
      RECT 16.2 -64 16.6 -49.36 ;
      RECT 16.2 -45.51 16.6 -12.47 ;
      RECT 13.3 -80.215 13.7 -20.12 ;
      RECT 12.5 -79.355 12.9 -20.12 ;
      RECT 11.7 -158.195 12.1 -79.445 ;
      RECT 10.9 -63.5 11.3 -48.905 ;
      RECT 10.9 -45.08 11.3 -15.74 ;
      RECT 10.1 -158.195 10.5 -73.605 ;
      RECT 10.1 -64 10.5 -49.36 ;
      RECT 10.1 -45.51 10.5 -12.47 ;
      RECT 8 -87.06 8.4 -20.12 ;
      RECT 7.2 -80.215 7.6 -20.12 ;
      RECT 6.4 -158.195 6.8 -87.15 ;
      RECT 6.4 -79.355 6.8 -20.12 ;
      RECT 5.6 -158.195 6 -79.445 ;
      RECT 4.8 -63.5 5.2 -48.905 ;
      RECT 4.8 -45.08 5.2 -15.74 ;
      RECT 4 -158.195 4.4 -73.605 ;
      RECT 4 -64 4.4 -49.36 ;
      RECT 4 -45.51 4.4 -12.47 ;
  END
END sram22_64x4m4w2

END LIBRARY
