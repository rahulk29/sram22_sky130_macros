VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 
MACRO sram22_64x24m4w8
    CLASS BLOCK  ;
    FOREIGN sram22_64x24m4w8   ;
    SIZE 298.440 BY 191.000 ;
    SYMMETRY X Y R90 ;
    PIN dout[0] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 138.470 0.000 138.610 0.140 ; 
        END 
    END dout[0] 
    PIN dout[1] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 144.570 0.000 144.710 0.140 ; 
        END 
    END dout[1] 
    PIN dout[2] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 150.670 0.000 150.810 0.140 ; 
        END 
    END dout[2] 
    PIN dout[3] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 156.770 0.000 156.910 0.140 ; 
        END 
    END dout[3] 
    PIN dout[4] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 162.870 0.000 163.010 0.140 ; 
        END 
    END dout[4] 
    PIN dout[5] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 168.970 0.000 169.110 0.140 ; 
        END 
    END dout[5] 
    PIN dout[6] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 175.070 0.000 175.210 0.140 ; 
        END 
    END dout[6] 
    PIN dout[7] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 181.170 0.000 181.310 0.140 ; 
        END 
    END dout[7] 
    PIN dout[8] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 187.270 0.000 187.410 0.140 ; 
        END 
    END dout[8] 
    PIN dout[9] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 193.370 0.000 193.510 0.140 ; 
        END 
    END dout[9] 
    PIN dout[10] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 199.470 0.000 199.610 0.140 ; 
        END 
    END dout[10] 
    PIN dout[11] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 205.570 0.000 205.710 0.140 ; 
        END 
    END dout[11] 
    PIN dout[12] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 211.670 0.000 211.810 0.140 ; 
        END 
    END dout[12] 
    PIN dout[13] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 217.770 0.000 217.910 0.140 ; 
        END 
    END dout[13] 
    PIN dout[14] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 223.870 0.000 224.010 0.140 ; 
        END 
    END dout[14] 
    PIN dout[15] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 229.970 0.000 230.110 0.140 ; 
        END 
    END dout[15] 
    PIN dout[16] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 236.070 0.000 236.210 0.140 ; 
        END 
    END dout[16] 
    PIN dout[17] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 242.170 0.000 242.310 0.140 ; 
        END 
    END dout[17] 
    PIN dout[18] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 248.270 0.000 248.410 0.140 ; 
        END 
    END dout[18] 
    PIN dout[19] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 254.370 0.000 254.510 0.140 ; 
        END 
    END dout[19] 
    PIN dout[20] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 260.470 0.000 260.610 0.140 ; 
        END 
    END dout[20] 
    PIN dout[21] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 266.570 0.000 266.710 0.140 ; 
        END 
    END dout[21] 
    PIN dout[22] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 272.670 0.000 272.810 0.140 ; 
        END 
    END dout[22] 
    PIN dout[23] 
        DIRECTION OUTPUT ; 
        ANTENNADIFFAREA 0.448000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 0.950300 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 7.107200 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 278.770 0.000 278.910 0.140 ; 
        END 
    END dout[23] 
    PIN din[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 138.050 0.000 138.190 0.140 ; 
        END 
    END din[0] 
    PIN din[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 144.150 0.000 144.290 0.140 ; 
        END 
    END din[1] 
    PIN din[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 150.250 0.000 150.390 0.140 ; 
        END 
    END din[2] 
    PIN din[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 156.350 0.000 156.490 0.140 ; 
        END 
    END din[3] 
    PIN din[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 162.450 0.000 162.590 0.140 ; 
        END 
    END din[4] 
    PIN din[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 168.550 0.000 168.690 0.140 ; 
        END 
    END din[5] 
    PIN din[6] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 174.650 0.000 174.790 0.140 ; 
        END 
    END din[6] 
    PIN din[7] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 180.750 0.000 180.890 0.140 ; 
        END 
    END din[7] 
    PIN din[8] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 186.850 0.000 186.990 0.140 ; 
        END 
    END din[8] 
    PIN din[9] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 192.950 0.000 193.090 0.140 ; 
        END 
    END din[9] 
    PIN din[10] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 199.050 0.000 199.190 0.140 ; 
        END 
    END din[10] 
    PIN din[11] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 205.150 0.000 205.290 0.140 ; 
        END 
    END din[11] 
    PIN din[12] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 211.250 0.000 211.390 0.140 ; 
        END 
    END din[12] 
    PIN din[13] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 217.350 0.000 217.490 0.140 ; 
        END 
    END din[13] 
    PIN din[14] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 223.450 0.000 223.590 0.140 ; 
        END 
    END din[14] 
    PIN din[15] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 229.550 0.000 229.690 0.140 ; 
        END 
    END din[15] 
    PIN din[16] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 235.650 0.000 235.790 0.140 ; 
        END 
    END din[16] 
    PIN din[17] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 241.750 0.000 241.890 0.140 ; 
        END 
    END din[17] 
    PIN din[18] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 247.850 0.000 247.990 0.140 ; 
        END 
    END din[18] 
    PIN din[19] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 253.950 0.000 254.090 0.140 ; 
        END 
    END din[19] 
    PIN din[20] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 260.050 0.000 260.190 0.140 ; 
        END 
    END din[20] 
    PIN din[21] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 266.150 0.000 266.290 0.140 ; 
        END 
    END din[21] 
    PIN din[22] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 272.250 0.000 272.390 0.140 ; 
        END 
    END din[22] 
    PIN din[23] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 5.238500 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 6.828800 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 278.350 0.000 278.490 0.140 ; 
        END 
    END din[23] 
    PIN wmask[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.048900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 137.700 0.000 137.840 0.140 ; 
        END 
    END wmask[0] 
    PIN wmask[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.048900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 186.500 0.000 186.640 0.140 ; 
        END 
    END wmask[1] 
    PIN wmask[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met2 ;
        ANTENNAPARTIALMETALAREA 3.048900 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 0.278400 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 235.300 0.000 235.440 0.140 ; 
        END 
    END wmask[2] 
    PIN addr[0] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 96.360 0.000 96.680 0.320 ; 
        END 
    END addr[0] 
    PIN addr[1] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 90.240 0.000 90.560 0.320 ; 
        END 
    END addr[1] 
    PIN addr[2] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 84.120 0.000 84.440 0.320 ; 
        END 
    END addr[2] 
    PIN addr[3] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 78.000 0.000 78.320 0.320 ; 
        END 
    END addr[3] 
    PIN addr[4] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 71.880 0.000 72.200 0.320 ; 
        END 
    END addr[4] 
    PIN addr[5] 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 65.760 0.000 66.080 0.320 ; 
        END 
    END addr[5] 
    PIN we 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 108.600 0.000 108.920 0.320 ; 
        END 
    END we 
    PIN ce 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 0.126000 LAYER met1 ;
        ANTENNAPARTIALMETALAREA 3.880700 LAYER met1 ;
        PORT 
            LAYER met1 ;
                RECT 102.480 0.000 102.800 0.320 ; 
        END 
    END ce 
    PIN clk 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 17.019000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 111.320 0.000 111.640 0.320 ; 
        END 
    END clk 
    PIN rstb 
        DIRECTION INPUT ; 
        ANTENNAGATEAREA 20.925000 LAYER met2 ;
        PORT 
            LAYER met1 ;
                RECT 112.000 0.000 112.320 0.320 ; 
        END 
    END rstb 
    PIN vdd 
        DIRECTION INOUT ; 
        USE POWER ; 
        PORT 
            LAYER met2 ;
                RECT 0.160 5.920 137.480 6.240 ; 
                RECT 139.200 5.920 143.600 6.240 ; 
                RECT 145.320 5.920 149.720 6.240 ; 
                RECT 151.440 5.920 155.840 6.240 ; 
                RECT 157.560 5.920 161.960 6.240 ; 
                RECT 163.680 5.920 168.080 6.240 ; 
                RECT 169.800 5.920 174.200 6.240 ; 
                RECT 175.920 5.920 180.320 6.240 ; 
                RECT 182.040 5.920 186.440 6.240 ; 
                RECT 188.160 5.920 192.560 6.240 ; 
                RECT 194.280 5.920 198.680 6.240 ; 
                RECT 200.400 5.920 204.800 6.240 ; 
                RECT 206.520 5.920 210.920 6.240 ; 
                RECT 212.640 5.920 217.040 6.240 ; 
                RECT 218.760 5.920 223.160 6.240 ; 
                RECT 224.880 5.920 229.280 6.240 ; 
                RECT 231.000 5.920 235.400 6.240 ; 
                RECT 237.120 5.920 241.520 6.240 ; 
                RECT 243.240 5.920 247.640 6.240 ; 
                RECT 249.360 5.920 253.760 6.240 ; 
                RECT 255.480 5.920 259.880 6.240 ; 
                RECT 261.600 5.920 266.000 6.240 ; 
                RECT 267.720 5.920 272.120 6.240 ; 
                RECT 273.840 5.920 278.240 6.240 ; 
                RECT 279.280 5.920 298.280 6.240 ; 
                RECT 0.160 7.280 298.280 7.600 ; 
                RECT 0.160 8.640 298.280 8.960 ; 
                RECT 0.160 10.000 110.960 10.320 ; 
                RECT 133.760 10.000 298.280 10.320 ; 
                RECT 0.160 11.360 298.280 11.680 ; 
                RECT 0.160 12.720 298.280 13.040 ; 
                RECT 0.160 14.080 62.000 14.400 ; 
                RECT 112.680 14.080 298.280 14.400 ; 
                RECT 0.160 15.440 298.280 15.760 ; 
                RECT 0.160 16.800 298.280 17.120 ; 
                RECT 0.160 18.160 62.000 18.480 ; 
                RECT 112.000 18.160 298.280 18.480 ; 
                RECT 0.160 19.520 298.280 19.840 ; 
                RECT 0.160 20.880 127.280 21.200 ; 
                RECT 288.120 20.880 298.280 21.200 ; 
                RECT 0.160 22.240 127.280 22.560 ; 
                RECT 288.120 22.240 298.280 22.560 ; 
                RECT 0.160 23.600 127.280 23.920 ; 
                RECT 288.120 23.600 298.280 23.920 ; 
                RECT 0.160 24.960 127.280 25.280 ; 
                RECT 288.120 24.960 298.280 25.280 ; 
                RECT 0.160 26.320 127.280 26.640 ; 
                RECT 288.120 26.320 298.280 26.640 ; 
                RECT 0.160 27.680 127.280 28.000 ; 
                RECT 288.120 27.680 298.280 28.000 ; 
                RECT 0.160 29.040 127.280 29.360 ; 
                RECT 288.120 29.040 298.280 29.360 ; 
                RECT 0.160 30.400 127.280 30.720 ; 
                RECT 288.120 30.400 298.280 30.720 ; 
                RECT 0.160 31.760 79.000 32.080 ; 
                RECT 89.560 31.760 127.280 32.080 ; 
                RECT 288.120 31.760 298.280 32.080 ; 
                RECT 0.160 33.120 77.640 33.440 ; 
                RECT 95.680 33.120 127.280 33.440 ; 
                RECT 288.120 33.120 298.280 33.440 ; 
                RECT 0.160 34.480 57.920 34.800 ; 
                RECT 112.680 34.480 127.280 34.800 ; 
                RECT 288.120 34.480 298.280 34.800 ; 
                RECT 0.160 35.840 57.240 36.160 ; 
                RECT 108.600 35.840 127.280 36.160 ; 
                RECT 288.120 35.840 298.280 36.160 ; 
                RECT 0.160 37.200 127.280 37.520 ; 
                RECT 288.120 37.200 298.280 37.520 ; 
                RECT 0.160 38.560 126.600 38.880 ; 
                RECT 288.120 38.560 298.280 38.880 ; 
                RECT 0.160 39.920 127.280 40.240 ; 
                RECT 288.120 39.920 298.280 40.240 ; 
                RECT 0.160 41.280 127.280 41.600 ; 
                RECT 288.120 41.280 298.280 41.600 ; 
                RECT 0.160 42.640 53.840 42.960 ; 
                RECT 64.400 42.640 127.280 42.960 ; 
                RECT 288.120 42.640 298.280 42.960 ; 
                RECT 0.160 44.000 55.200 44.320 ; 
                RECT 61.000 44.000 68.120 44.320 ; 
                RECT 71.200 44.000 127.280 44.320 ; 
                RECT 288.120 44.000 298.280 44.320 ; 
                RECT 0.160 45.360 56.560 45.680 ; 
                RECT 59.640 45.360 127.280 45.680 ; 
                RECT 288.120 45.360 298.280 45.680 ; 
                RECT 0.160 46.720 127.280 47.040 ; 
                RECT 288.120 46.720 298.280 47.040 ; 
                RECT 0.160 48.080 62.680 48.400 ; 
                RECT 71.200 48.080 104.160 48.400 ; 
                RECT 110.640 48.080 127.280 48.400 ; 
                RECT 288.120 48.080 298.280 48.400 ; 
                RECT 0.160 49.440 55.200 49.760 ; 
                RECT 64.400 49.440 104.160 49.760 ; 
                RECT 110.640 49.440 127.280 49.760 ; 
                RECT 288.120 49.440 298.280 49.760 ; 
                RECT 0.160 50.800 59.280 51.120 ; 
                RECT 63.720 50.800 104.160 51.120 ; 
                RECT 288.120 50.800 298.280 51.120 ; 
                RECT 0.160 52.160 104.160 52.480 ; 
                RECT 110.640 52.160 127.280 52.480 ; 
                RECT 288.120 52.160 298.280 52.480 ; 
                RECT 0.160 53.520 55.200 53.840 ; 
                RECT 64.400 53.520 127.280 53.840 ; 
                RECT 288.120 53.520 298.280 53.840 ; 
                RECT 0.160 54.880 62.000 55.200 ; 
                RECT 70.520 54.880 127.280 55.200 ; 
                RECT 288.120 54.880 298.280 55.200 ; 
                RECT 0.160 56.240 127.280 56.560 ; 
                RECT 288.120 56.240 298.280 56.560 ; 
                RECT 0.160 57.600 62.680 57.920 ; 
                RECT 68.480 57.600 89.200 57.920 ; 
                RECT 109.960 57.600 127.280 57.920 ; 
                RECT 288.120 57.600 298.280 57.920 ; 
                RECT 0.160 58.960 65.400 59.280 ; 
                RECT 71.200 58.960 78.320 59.280 ; 
                RECT 83.440 58.960 89.200 59.280 ; 
                RECT 109.960 58.960 127.280 59.280 ; 
                RECT 288.120 58.960 298.280 59.280 ; 
                RECT 0.160 60.320 59.280 60.640 ; 
                RECT 64.400 60.320 79.680 60.640 ; 
                RECT 82.080 60.320 89.200 60.640 ; 
                RECT 119.480 60.320 127.280 60.640 ; 
                RECT 288.120 60.320 298.280 60.640 ; 
                RECT 0.160 61.680 89.200 62.000 ; 
                RECT 119.480 61.680 127.280 62.000 ; 
                RECT 288.120 61.680 298.280 62.000 ; 
                RECT 0.160 63.040 53.160 63.360 ; 
                RECT 75.960 63.040 89.200 63.360 ; 
                RECT 118.120 63.040 127.280 63.360 ; 
                RECT 288.120 63.040 298.280 63.360 ; 
                RECT 0.160 64.400 62.680 64.720 ; 
                RECT 71.200 64.400 89.200 64.720 ; 
                RECT 119.480 64.400 127.280 64.720 ; 
                RECT 288.120 64.400 298.280 64.720 ; 
                RECT 0.160 65.760 62.000 66.080 ; 
                RECT 64.400 65.760 71.520 66.080 ; 
                RECT 78.000 65.760 89.200 66.080 ; 
                RECT 119.480 65.760 127.280 66.080 ; 
                RECT 288.120 65.760 298.280 66.080 ; 
                RECT 0.160 67.120 53.840 67.440 ; 
                RECT 67.120 67.120 89.200 67.440 ; 
                RECT 109.960 67.120 127.280 67.440 ; 
                RECT 288.120 67.120 298.280 67.440 ; 
                RECT 0.160 68.480 62.000 68.800 ; 
                RECT 71.200 68.480 89.200 68.800 ; 
                RECT 122.200 68.480 127.280 68.800 ; 
                RECT 288.120 68.480 298.280 68.800 ; 
                RECT 0.160 69.840 59.960 70.160 ; 
                RECT 63.720 69.840 89.200 70.160 ; 
                RECT 120.840 69.840 127.280 70.160 ; 
                RECT 288.120 69.840 298.280 70.160 ; 
                RECT 0.160 71.200 55.200 71.520 ; 
                RECT 59.640 71.200 62.680 71.520 ; 
                RECT 71.200 71.200 89.200 71.520 ; 
                RECT 122.200 71.200 127.280 71.520 ; 
                RECT 288.120 71.200 298.280 71.520 ; 
                RECT 0.160 72.560 57.920 72.880 ; 
                RECT 61.680 72.560 89.200 72.880 ; 
                RECT 122.200 72.560 127.280 72.880 ; 
                RECT 288.120 72.560 298.280 72.880 ; 
                RECT 0.160 73.920 55.200 74.240 ; 
                RECT 58.280 73.920 89.200 74.240 ; 
                RECT 122.200 73.920 127.280 74.240 ; 
                RECT 288.120 73.920 298.280 74.240 ; 
                RECT 0.160 75.280 59.280 75.600 ; 
                RECT 64.400 75.280 89.200 75.600 ; 
                RECT 120.840 75.280 127.280 75.600 ; 
                RECT 288.120 75.280 298.280 75.600 ; 
                RECT 0.160 76.640 55.200 76.960 ; 
                RECT 71.200 76.640 89.200 76.960 ; 
                RECT 109.960 76.640 127.280 76.960 ; 
                RECT 288.120 76.640 298.280 76.960 ; 
                RECT 0.160 78.000 63.360 78.320 ; 
                RECT 67.120 78.000 89.200 78.320 ; 
                RECT 123.560 78.000 127.280 78.320 ; 
                RECT 288.120 78.000 298.280 78.320 ; 
                RECT 0.160 79.360 62.000 79.680 ; 
                RECT 65.080 79.360 89.200 79.680 ; 
                RECT 124.920 79.360 127.280 79.680 ; 
                RECT 288.120 79.360 298.280 79.680 ; 
                RECT 0.160 80.720 62.680 81.040 ; 
                RECT 67.120 80.720 89.200 81.040 ; 
                RECT 124.920 80.720 127.280 81.040 ; 
                RECT 288.120 80.720 298.280 81.040 ; 
                RECT 0.160 82.080 53.840 82.400 ; 
                RECT 61.000 82.080 89.200 82.400 ; 
                RECT 123.560 82.080 127.280 82.400 ; 
                RECT 288.120 82.080 298.280 82.400 ; 
                RECT 0.160 83.440 53.840 83.760 ; 
                RECT 64.400 83.440 89.200 83.760 ; 
                RECT 124.920 83.440 127.280 83.760 ; 
                RECT 288.120 83.440 298.280 83.760 ; 
                RECT 0.160 84.800 56.560 85.120 ; 
                RECT 63.720 84.800 89.200 85.120 ; 
                RECT 109.960 84.800 127.280 85.120 ; 
                RECT 288.120 84.800 298.280 85.120 ; 
                RECT 0.160 86.160 62.000 86.480 ; 
                RECT 65.080 86.160 89.200 86.480 ; 
                RECT 288.120 86.160 298.280 86.480 ; 
                RECT 0.160 87.520 58.600 87.840 ; 
                RECT 71.200 87.520 89.200 87.840 ; 
                RECT 288.120 87.520 298.280 87.840 ; 
                RECT 0.160 88.880 89.200 89.200 ; 
                RECT 288.120 88.880 298.280 89.200 ; 
                RECT 0.160 90.240 49.760 90.560 ; 
                RECT 67.120 90.240 89.200 90.560 ; 
                RECT 288.120 90.240 298.280 90.560 ; 
                RECT 0.160 91.600 89.200 91.920 ; 
                RECT 288.120 91.600 298.280 91.920 ; 
                RECT 0.160 92.960 89.200 93.280 ; 
                RECT 109.960 92.960 127.280 93.280 ; 
                RECT 288.120 92.960 298.280 93.280 ; 
                RECT 0.160 94.320 127.280 94.640 ; 
                RECT 288.120 94.320 298.280 94.640 ; 
                RECT 0.160 95.680 65.400 96.000 ; 
                RECT 73.240 95.680 127.280 96.000 ; 
                RECT 288.120 95.680 298.280 96.000 ; 
                RECT 0.160 97.040 68.800 97.360 ; 
                RECT 71.200 97.040 127.280 97.360 ; 
                RECT 288.120 97.040 298.280 97.360 ; 
                RECT 0.160 98.400 127.280 98.720 ; 
                RECT 288.120 98.400 298.280 98.720 ; 
                RECT 0.160 99.760 53.160 100.080 ; 
                RECT 58.280 99.760 76.960 100.080 ; 
                RECT 86.840 99.760 89.200 100.080 ; 
                RECT 110.640 99.760 127.280 100.080 ; 
                RECT 288.120 99.760 298.280 100.080 ; 
                RECT 0.160 101.120 89.200 101.440 ; 
                RECT 110.640 101.120 127.280 101.440 ; 
                RECT 288.120 101.120 298.280 101.440 ; 
                RECT 0.160 102.480 89.200 102.800 ; 
                RECT 110.640 102.480 127.280 102.800 ; 
                RECT 288.120 102.480 298.280 102.800 ; 
                RECT 0.160 103.840 89.200 104.160 ; 
                RECT 110.640 103.840 127.280 104.160 ; 
                RECT 288.120 103.840 298.280 104.160 ; 
                RECT 0.160 105.200 62.000 105.520 ; 
                RECT 70.520 105.200 89.200 105.520 ; 
                RECT 110.640 105.200 127.280 105.520 ; 
                RECT 288.120 105.200 298.280 105.520 ; 
                RECT 0.160 106.560 89.200 106.880 ; 
                RECT 110.640 106.560 127.280 106.880 ; 
                RECT 288.120 106.560 298.280 106.880 ; 
                RECT 0.160 107.920 89.200 108.240 ; 
                RECT 110.640 107.920 127.280 108.240 ; 
                RECT 288.120 107.920 298.280 108.240 ; 
                RECT 0.160 109.280 55.200 109.600 ; 
                RECT 60.320 109.280 89.200 109.600 ; 
                RECT 288.120 109.280 298.280 109.600 ; 
                RECT 0.160 110.640 89.200 110.960 ; 
                RECT 110.640 110.640 124.560 110.960 ; 
                RECT 288.120 110.640 298.280 110.960 ; 
                RECT 0.160 112.000 89.200 112.320 ; 
                RECT 110.640 112.000 121.840 112.320 ; 
                RECT 288.120 112.000 298.280 112.320 ; 
                RECT 0.160 113.360 89.200 113.680 ; 
                RECT 110.640 113.360 119.120 113.680 ; 
                RECT 288.120 113.360 298.280 113.680 ; 
                RECT 0.160 114.720 32.080 115.040 ; 
                RECT 50.120 114.720 57.920 115.040 ; 
                RECT 61.000 114.720 89.200 115.040 ; 
                RECT 110.640 114.720 116.400 115.040 ; 
                RECT 288.120 114.720 298.280 115.040 ; 
                RECT 0.160 116.080 32.080 116.400 ; 
                RECT 50.120 116.080 55.200 116.400 ; 
                RECT 58.280 116.080 89.200 116.400 ; 
                RECT 110.640 116.080 127.280 116.400 ; 
                RECT 288.120 116.080 298.280 116.400 ; 
                RECT 0.160 117.440 32.080 117.760 ; 
                RECT 50.120 117.440 89.200 117.760 ; 
                RECT 110.640 117.440 127.280 117.760 ; 
                RECT 288.120 117.440 298.280 117.760 ; 
                RECT 0.160 118.800 32.080 119.120 ; 
                RECT 50.120 118.800 127.280 119.120 ; 
                RECT 288.120 118.800 298.280 119.120 ; 
                RECT 0.160 120.160 32.080 120.480 ; 
                RECT 50.800 120.160 127.280 120.480 ; 
                RECT 288.120 120.160 298.280 120.480 ; 
                RECT 0.160 121.520 32.080 121.840 ; 
                RECT 50.120 121.520 127.280 121.840 ; 
                RECT 288.120 121.520 298.280 121.840 ; 
                RECT 0.160 122.880 32.080 123.200 ; 
                RECT 50.120 122.880 127.280 123.200 ; 
                RECT 288.120 122.880 298.280 123.200 ; 
                RECT 0.160 124.240 32.080 124.560 ; 
                RECT 50.120 124.240 89.200 124.560 ; 
                RECT 109.960 124.240 117.760 124.560 ; 
                RECT 288.120 124.240 298.280 124.560 ; 
                RECT 0.160 125.600 32.080 125.920 ; 
                RECT 50.120 125.600 56.560 125.920 ; 
                RECT 61.000 125.600 89.200 125.920 ; 
                RECT 109.960 125.600 120.480 125.920 ; 
                RECT 288.120 125.600 298.280 125.920 ; 
                RECT 0.160 126.960 89.200 127.280 ; 
                RECT 109.960 126.960 123.200 127.280 ; 
                RECT 288.120 126.960 298.280 127.280 ; 
                RECT 0.160 128.320 89.200 128.640 ; 
                RECT 109.960 128.320 125.920 128.640 ; 
                RECT 288.120 128.320 298.280 128.640 ; 
                RECT 0.160 129.680 59.280 130.000 ; 
                RECT 65.080 129.680 89.200 130.000 ; 
                RECT 288.120 129.680 298.280 130.000 ; 
                RECT 0.160 131.040 15.760 131.360 ; 
                RECT 31.760 131.040 38.200 131.360 ; 
                RECT 45.360 131.040 89.200 131.360 ; 
                RECT 109.960 131.040 127.280 131.360 ; 
                RECT 288.120 131.040 298.280 131.360 ; 
                RECT 0.160 132.400 15.760 132.720 ; 
                RECT 50.120 132.400 89.200 132.720 ; 
                RECT 109.960 132.400 127.280 132.720 ; 
                RECT 288.120 132.400 298.280 132.720 ; 
                RECT 0.160 133.760 15.760 134.080 ; 
                RECT 50.120 133.760 89.200 134.080 ; 
                RECT 288.120 133.760 298.280 134.080 ; 
                RECT 0.160 135.120 15.760 135.440 ; 
                RECT 31.760 135.120 38.200 135.440 ; 
                RECT 45.360 135.120 53.840 135.440 ; 
                RECT 63.720 135.120 89.200 135.440 ; 
                RECT 109.960 135.120 113.680 135.440 ; 
                RECT 288.120 135.120 298.280 135.440 ; 
                RECT 0.160 136.480 16.440 136.800 ; 
                RECT 44.680 136.480 89.200 136.800 ; 
                RECT 109.960 136.480 298.280 136.800 ; 
                RECT 0.160 137.840 44.320 138.160 ; 
                RECT 86.160 137.840 298.280 138.160 ; 
                RECT 0.160 139.200 124.560 139.520 ; 
                RECT 290.840 139.200 298.280 139.520 ; 
                RECT 0.160 140.560 124.560 140.880 ; 
                RECT 290.840 140.560 298.280 140.880 ; 
                RECT 0.160 141.920 124.560 142.240 ; 
                RECT 290.840 141.920 298.280 142.240 ; 
                RECT 0.160 143.280 23.240 143.600 ; 
                RECT 30.400 143.280 32.080 143.600 ; 
                RECT 40.600 143.280 70.160 143.600 ; 
                RECT 290.840 143.280 298.280 143.600 ; 
                RECT 0.160 144.640 21.200 144.960 ; 
                RECT 31.760 144.640 33.440 144.960 ; 
                RECT 39.920 144.640 51.120 144.960 ; 
                RECT 52.160 144.640 70.160 144.960 ; 
                RECT 290.840 144.640 298.280 144.960 ; 
                RECT 0.160 146.000 21.200 146.320 ; 
                RECT 31.760 146.000 51.120 146.320 ; 
                RECT 54.880 146.000 70.160 146.320 ; 
                RECT 290.840 146.000 298.280 146.320 ; 
                RECT 0.160 147.360 21.200 147.680 ; 
                RECT 31.760 147.360 51.120 147.680 ; 
                RECT 55.560 147.360 70.160 147.680 ; 
                RECT 290.840 147.360 298.280 147.680 ; 
                RECT 0.160 148.720 51.120 149.040 ; 
                RECT 56.240 148.720 70.160 149.040 ; 
                RECT 290.840 148.720 298.280 149.040 ; 
                RECT 0.160 150.080 21.200 150.400 ; 
                RECT 31.760 150.080 51.120 150.400 ; 
                RECT 52.160 150.080 70.160 150.400 ; 
                RECT 290.840 150.080 298.280 150.400 ; 
                RECT 0.160 151.440 21.200 151.760 ; 
                RECT 31.760 151.440 70.160 151.760 ; 
                RECT 290.840 151.440 298.280 151.760 ; 
                RECT 0.160 152.800 70.160 153.120 ; 
                RECT 290.840 152.800 298.280 153.120 ; 
                RECT 0.160 154.160 70.160 154.480 ; 
                RECT 290.840 154.160 298.280 154.480 ; 
                RECT 0.160 155.520 14.400 155.840 ; 
                RECT 17.480 155.520 70.160 155.840 ; 
                RECT 290.840 155.520 298.280 155.840 ; 
                RECT 0.160 156.880 70.160 157.200 ; 
                RECT 290.840 156.880 298.280 157.200 ; 
                RECT 0.160 158.240 13.720 158.560 ; 
                RECT 17.480 158.240 30.720 158.560 ; 
                RECT 33.800 158.240 70.160 158.560 ; 
                RECT 290.840 158.240 298.280 158.560 ; 
                RECT 0.160 159.600 13.040 159.920 ; 
                RECT 17.480 159.600 30.720 159.920 ; 
                RECT 40.600 159.600 70.160 159.920 ; 
                RECT 290.840 159.600 298.280 159.920 ; 
                RECT 0.160 160.960 12.360 161.280 ; 
                RECT 17.480 160.960 30.720 161.280 ; 
                RECT 39.240 160.960 51.120 161.280 ; 
                RECT 52.160 160.960 70.160 161.280 ; 
                RECT 290.840 160.960 298.280 161.280 ; 
                RECT 0.160 162.320 51.120 162.640 ; 
                RECT 52.840 162.320 70.160 162.640 ; 
                RECT 290.840 162.320 298.280 162.640 ; 
                RECT 0.160 163.680 11.680 164.000 ; 
                RECT 17.480 163.680 30.720 164.000 ; 
                RECT 35.840 163.680 51.120 164.000 ; 
                RECT 53.520 163.680 70.160 164.000 ; 
                RECT 290.840 163.680 298.280 164.000 ; 
                RECT 0.160 165.040 11.000 165.360 ; 
                RECT 17.480 165.040 51.120 165.360 ; 
                RECT 54.200 165.040 70.160 165.360 ; 
                RECT 290.840 165.040 298.280 165.360 ; 
                RECT 0.160 166.400 10.320 166.720 ; 
                RECT 17.480 166.400 51.120 166.720 ; 
                RECT 54.200 166.400 70.160 166.720 ; 
                RECT 290.840 166.400 298.280 166.720 ; 
                RECT 0.160 167.760 9.640 168.080 ; 
                RECT 17.480 167.760 70.160 168.080 ; 
                RECT 290.840 167.760 298.280 168.080 ; 
                RECT 0.160 169.120 70.160 169.440 ; 
                RECT 290.840 169.120 298.280 169.440 ; 
                RECT 0.160 170.480 70.160 170.800 ; 
                RECT 290.840 170.480 298.280 170.800 ; 
                RECT 0.160 171.840 70.160 172.160 ; 
                RECT 290.840 171.840 298.280 172.160 ; 
                RECT 0.160 173.200 70.160 173.520 ; 
                RECT 290.840 173.200 298.280 173.520 ; 
                RECT 0.160 174.560 70.160 174.880 ; 
                RECT 290.840 174.560 298.280 174.880 ; 
                RECT 0.160 175.920 70.160 176.240 ; 
                RECT 290.840 175.920 298.280 176.240 ; 
                RECT 0.160 177.280 124.560 177.600 ; 
                RECT 290.840 177.280 298.280 177.600 ; 
                RECT 0.160 178.640 124.560 178.960 ; 
                RECT 290.840 178.640 298.280 178.960 ; 
                RECT 0.160 180.000 124.560 180.320 ; 
                RECT 290.840 180.000 298.280 180.320 ; 
                RECT 0.160 181.360 298.280 181.680 ; 
                RECT 0.160 182.720 298.280 183.040 ; 
                RECT 0.160 184.080 298.280 184.400 ; 
                RECT 0.160 185.440 298.280 185.760 ; 
                RECT 0.160 0.160 298.280 1.520 ; 
                RECT 0.160 189.480 298.280 190.840 ; 
                RECT 128.700 42.275 134.500 43.645 ; 
                RECT 280.600 42.275 286.400 43.645 ; 
                RECT 128.700 47.315 134.500 48.685 ; 
                RECT 280.600 47.315 286.400 48.685 ; 
                RECT 128.700 52.415 134.500 53.835 ; 
                RECT 280.600 52.415 286.400 53.835 ; 
                RECT 128.700 57.585 134.500 59.005 ; 
                RECT 280.600 57.585 286.400 59.005 ; 
                RECT 128.700 95.445 286.400 95.735 ; 
                RECT 128.700 117.700 286.400 118.570 ; 
                RECT 128.700 65.770 286.400 67.570 ; 
                RECT 128.700 77.240 286.400 78.040 ; 
                RECT 128.700 85.140 286.400 85.940 ; 
                RECT 128.700 132.025 286.400 132.825 ; 
                RECT 128.700 91.365 286.400 92.165 ; 
                RECT 128.700 80.250 286.400 81.050 ; 
                RECT 128.700 26.520 286.400 28.320 ; 
                RECT 77.290 142.995 79.210 176.175 ; 
                RECT 81.130 142.995 83.050 176.175 ; 
                RECT 100.235 142.995 102.155 176.175 ; 
                RECT 104.075 142.995 105.995 176.175 ; 
                RECT 107.915 142.995 109.835 176.175 ; 
                RECT 111.755 142.995 113.675 176.175 ; 
                RECT 115.595 142.995 117.515 176.175 ; 
                RECT 119.435 142.995 121.355 176.175 ; 
                RECT 92.345 58.260 94.265 93.660 ; 
                RECT 98.975 58.260 100.725 93.660 ; 
                RECT 107.155 58.260 109.075 93.660 ; 
                RECT 92.970 123.880 94.890 136.360 ; 
                RECT 99.945 123.880 101.865 136.360 ; 
                RECT 107.565 123.880 109.485 136.360 ; 
                RECT 93.615 99.660 95.535 117.880 ; 
                RECT 100.675 99.660 102.425 117.880 ; 
                RECT 107.780 99.660 109.700 117.880 ; 
                RECT 107.800 48.680 109.720 52.260 ; 
                RECT 22.230 145.265 31.390 146.015 ; 
                RECT 22.230 149.890 31.390 151.640 ; 
                RECT 33.090 133.050 49.130 133.850 ; 
                RECT 16.290 133.760 31.130 135.450 ; 
        END 
    END vdd 
    PIN vss 
        DIRECTION INOUT ; 
        USE GROUND ; 
        PORT 
            LAYER met2 ;
                RECT 2.880 5.240 137.480 5.560 ; 
                RECT 139.200 5.240 143.600 5.560 ; 
                RECT 145.320 5.240 149.720 5.560 ; 
                RECT 151.440 5.240 155.840 5.560 ; 
                RECT 157.560 5.240 161.960 5.560 ; 
                RECT 163.680 5.240 168.080 5.560 ; 
                RECT 169.800 5.240 174.200 5.560 ; 
                RECT 175.920 5.240 180.320 5.560 ; 
                RECT 182.040 5.240 186.440 5.560 ; 
                RECT 188.160 5.240 192.560 5.560 ; 
                RECT 194.280 5.240 198.680 5.560 ; 
                RECT 200.400 5.240 204.800 5.560 ; 
                RECT 206.520 5.240 210.920 5.560 ; 
                RECT 212.640 5.240 217.040 5.560 ; 
                RECT 218.760 5.240 223.160 5.560 ; 
                RECT 224.880 5.240 229.280 5.560 ; 
                RECT 231.000 5.240 235.400 5.560 ; 
                RECT 237.120 5.240 241.520 5.560 ; 
                RECT 243.240 5.240 247.640 5.560 ; 
                RECT 249.360 5.240 253.760 5.560 ; 
                RECT 255.480 5.240 259.880 5.560 ; 
                RECT 261.600 5.240 266.000 5.560 ; 
                RECT 267.720 5.240 272.120 5.560 ; 
                RECT 273.840 5.240 278.240 5.560 ; 
                RECT 279.280 5.240 295.560 5.560 ; 
                RECT 2.880 6.600 295.560 6.920 ; 
                RECT 2.880 7.960 295.560 8.280 ; 
                RECT 2.880 9.320 111.640 9.640 ; 
                RECT 133.080 9.320 295.560 9.640 ; 
                RECT 2.880 10.680 295.560 11.000 ; 
                RECT 2.880 12.040 295.560 12.360 ; 
                RECT 2.880 13.400 62.000 13.720 ; 
                RECT 112.680 13.400 295.560 13.720 ; 
                RECT 2.880 14.760 295.560 15.080 ; 
                RECT 2.880 16.120 295.560 16.440 ; 
                RECT 2.880 17.480 62.000 17.800 ; 
                RECT 112.000 17.480 295.560 17.800 ; 
                RECT 2.880 18.840 295.560 19.160 ; 
                RECT 2.880 20.200 127.280 20.520 ; 
                RECT 288.120 20.200 295.560 20.520 ; 
                RECT 2.880 21.560 127.280 21.880 ; 
                RECT 288.120 21.560 295.560 21.880 ; 
                RECT 2.880 22.920 127.280 23.240 ; 
                RECT 288.120 22.920 295.560 23.240 ; 
                RECT 2.880 24.280 127.280 24.600 ; 
                RECT 288.120 24.280 295.560 24.600 ; 
                RECT 2.880 25.640 127.280 25.960 ; 
                RECT 288.120 25.640 295.560 25.960 ; 
                RECT 2.880 27.000 127.280 27.320 ; 
                RECT 288.120 27.000 295.560 27.320 ; 
                RECT 2.880 28.360 127.280 28.680 ; 
                RECT 288.120 28.360 295.560 28.680 ; 
                RECT 2.880 29.720 127.280 30.040 ; 
                RECT 288.120 29.720 295.560 30.040 ; 
                RECT 2.880 31.080 79.680 31.400 ; 
                RECT 90.920 31.080 127.280 31.400 ; 
                RECT 288.120 31.080 295.560 31.400 ; 
                RECT 2.880 32.440 78.320 32.760 ; 
                RECT 97.040 32.440 127.280 32.760 ; 
                RECT 288.120 32.440 295.560 32.760 ; 
                RECT 2.880 33.800 55.200 34.120 ; 
                RECT 112.000 33.800 127.280 34.120 ; 
                RECT 288.120 33.800 295.560 34.120 ; 
                RECT 2.880 35.160 56.560 35.480 ; 
                RECT 102.480 35.160 127.280 35.480 ; 
                RECT 288.120 35.160 295.560 35.480 ; 
                RECT 2.880 36.520 127.280 36.840 ; 
                RECT 288.120 36.520 295.560 36.840 ; 
                RECT 2.880 37.880 126.600 38.200 ; 
                RECT 288.120 37.880 295.560 38.200 ; 
                RECT 2.880 39.240 127.280 39.560 ; 
                RECT 288.120 39.240 295.560 39.560 ; 
                RECT 2.880 40.600 127.280 40.920 ; 
                RECT 288.120 40.600 295.560 40.920 ; 
                RECT 2.880 41.960 53.840 42.280 ; 
                RECT 64.400 41.960 127.280 42.280 ; 
                RECT 288.120 41.960 295.560 42.280 ; 
                RECT 2.880 43.320 55.200 43.640 ; 
                RECT 56.920 43.320 127.280 43.640 ; 
                RECT 288.120 43.320 295.560 43.640 ; 
                RECT 2.880 44.680 56.560 45.000 ; 
                RECT 61.000 44.680 68.120 45.000 ; 
                RECT 71.200 44.680 127.280 45.000 ; 
                RECT 288.120 44.680 295.560 45.000 ; 
                RECT 2.880 46.040 56.560 46.360 ; 
                RECT 59.640 46.040 127.280 46.360 ; 
                RECT 288.120 46.040 295.560 46.360 ; 
                RECT 2.880 47.400 62.680 47.720 ; 
                RECT 71.200 47.400 127.280 47.720 ; 
                RECT 288.120 47.400 295.560 47.720 ; 
                RECT 2.880 48.760 57.920 49.080 ; 
                RECT 64.400 48.760 104.160 49.080 ; 
                RECT 110.640 48.760 127.280 49.080 ; 
                RECT 288.120 48.760 295.560 49.080 ; 
                RECT 2.880 50.120 55.200 50.440 ; 
                RECT 64.400 50.120 104.160 50.440 ; 
                RECT 288.120 50.120 295.560 50.440 ; 
                RECT 2.880 51.480 76.280 51.800 ; 
                RECT 101.120 51.480 104.160 51.800 ; 
                RECT 110.640 51.480 127.280 51.800 ; 
                RECT 288.120 51.480 295.560 51.800 ; 
                RECT 2.880 52.840 55.200 53.160 ; 
                RECT 64.400 52.840 127.280 53.160 ; 
                RECT 288.120 52.840 295.560 53.160 ; 
                RECT 2.880 54.200 62.680 54.520 ; 
                RECT 70.520 54.200 127.280 54.520 ; 
                RECT 288.120 54.200 295.560 54.520 ; 
                RECT 2.880 55.560 62.000 55.880 ; 
                RECT 64.400 55.560 127.280 55.880 ; 
                RECT 288.120 55.560 295.560 55.880 ; 
                RECT 2.880 56.920 127.280 57.240 ; 
                RECT 288.120 56.920 295.560 57.240 ; 
                RECT 2.880 58.280 62.680 58.600 ; 
                RECT 71.200 58.280 77.640 58.600 ; 
                RECT 83.440 58.280 89.200 58.600 ; 
                RECT 109.960 58.280 127.280 58.600 ; 
                RECT 288.120 58.280 295.560 58.600 ; 
                RECT 2.880 59.640 59.280 59.960 ; 
                RECT 64.400 59.640 79.000 59.960 ; 
                RECT 82.760 59.640 89.200 59.960 ; 
                RECT 119.480 59.640 127.280 59.960 ; 
                RECT 288.120 59.640 295.560 59.960 ; 
                RECT 2.880 61.000 62.000 61.320 ; 
                RECT 64.400 61.000 89.200 61.320 ; 
                RECT 118.120 61.000 127.280 61.320 ; 
                RECT 288.120 61.000 295.560 61.320 ; 
                RECT 2.880 62.360 89.200 62.680 ; 
                RECT 119.480 62.360 127.280 62.680 ; 
                RECT 288.120 62.360 295.560 62.680 ; 
                RECT 2.880 63.720 53.160 64.040 ; 
                RECT 75.960 63.720 89.200 64.040 ; 
                RECT 119.480 63.720 127.280 64.040 ; 
                RECT 288.120 63.720 295.560 64.040 ; 
                RECT 2.880 65.080 71.520 65.400 ; 
                RECT 77.320 65.080 89.200 65.400 ; 
                RECT 109.960 65.080 127.280 65.400 ; 
                RECT 288.120 65.080 295.560 65.400 ; 
                RECT 2.880 66.440 62.000 66.760 ; 
                RECT 64.400 66.440 74.240 66.760 ; 
                RECT 78.000 66.440 89.200 66.760 ; 
                RECT 118.120 66.440 127.280 66.760 ; 
                RECT 288.120 66.440 295.560 66.760 ; 
                RECT 2.880 67.800 53.840 68.120 ; 
                RECT 67.120 67.800 89.200 68.120 ; 
                RECT 109.960 67.800 127.280 68.120 ; 
                RECT 288.120 67.800 295.560 68.120 ; 
                RECT 2.880 69.160 62.000 69.480 ; 
                RECT 71.200 69.160 89.200 69.480 ; 
                RECT 122.200 69.160 127.280 69.480 ; 
                RECT 288.120 69.160 295.560 69.480 ; 
                RECT 2.880 70.520 59.960 70.840 ; 
                RECT 71.200 70.520 89.200 70.840 ; 
                RECT 122.200 70.520 127.280 70.840 ; 
                RECT 288.120 70.520 295.560 70.840 ; 
                RECT 2.880 71.880 55.200 72.200 ; 
                RECT 61.680 71.880 89.200 72.200 ; 
                RECT 122.200 71.880 127.280 72.200 ; 
                RECT 288.120 71.880 295.560 72.200 ; 
                RECT 2.880 73.240 89.200 73.560 ; 
                RECT 120.840 73.240 127.280 73.560 ; 
                RECT 288.120 73.240 295.560 73.560 ; 
                RECT 2.880 74.600 55.200 74.920 ; 
                RECT 58.280 74.600 89.200 74.920 ; 
                RECT 122.200 74.600 127.280 74.920 ; 
                RECT 288.120 74.600 295.560 74.920 ; 
                RECT 2.880 75.960 55.200 76.280 ; 
                RECT 64.400 75.960 89.200 76.280 ; 
                RECT 109.960 75.960 127.280 76.280 ; 
                RECT 288.120 75.960 295.560 76.280 ; 
                RECT 2.880 77.320 59.280 77.640 ; 
                RECT 71.200 77.320 89.200 77.640 ; 
                RECT 124.920 77.320 127.280 77.640 ; 
                RECT 288.120 77.320 295.560 77.640 ; 
                RECT 2.880 78.680 62.000 79.000 ; 
                RECT 67.120 78.680 89.200 79.000 ; 
                RECT 124.920 78.680 127.280 79.000 ; 
                RECT 288.120 78.680 295.560 79.000 ; 
                RECT 2.880 80.040 62.680 80.360 ; 
                RECT 67.120 80.040 89.200 80.360 ; 
                RECT 123.560 80.040 127.280 80.360 ; 
                RECT 288.120 80.040 295.560 80.360 ; 
                RECT 2.880 81.400 89.200 81.720 ; 
                RECT 124.920 81.400 127.280 81.720 ; 
                RECT 288.120 81.400 295.560 81.720 ; 
                RECT 2.880 82.760 53.840 83.080 ; 
                RECT 61.000 82.760 89.200 83.080 ; 
                RECT 124.920 82.760 127.280 83.080 ; 
                RECT 288.120 82.760 295.560 83.080 ; 
                RECT 2.880 84.120 53.840 84.440 ; 
                RECT 64.400 84.120 89.200 84.440 ; 
                RECT 123.560 84.120 127.280 84.440 ; 
                RECT 288.120 84.120 295.560 84.440 ; 
                RECT 2.880 85.480 62.000 85.800 ; 
                RECT 65.080 85.480 89.200 85.800 ; 
                RECT 288.120 85.480 295.560 85.800 ; 
                RECT 2.880 86.840 89.200 87.160 ; 
                RECT 288.120 86.840 295.560 87.160 ; 
                RECT 2.880 88.200 58.600 88.520 ; 
                RECT 71.200 88.200 89.200 88.520 ; 
                RECT 288.120 88.200 295.560 88.520 ; 
                RECT 2.880 89.560 49.760 89.880 ; 
                RECT 63.720 89.560 89.200 89.880 ; 
                RECT 288.120 89.560 295.560 89.880 ; 
                RECT 2.880 90.920 59.960 91.240 ; 
                RECT 67.120 90.920 89.200 91.240 ; 
                RECT 109.960 90.920 127.280 91.240 ; 
                RECT 288.120 90.920 295.560 91.240 ; 
                RECT 2.880 92.280 89.200 92.600 ; 
                RECT 288.120 92.280 295.560 92.600 ; 
                RECT 2.880 93.640 89.200 93.960 ; 
                RECT 109.960 93.640 127.280 93.960 ; 
                RECT 288.120 93.640 295.560 93.960 ; 
                RECT 2.880 95.000 65.400 95.320 ; 
                RECT 73.240 95.000 127.280 95.320 ; 
                RECT 288.120 95.000 295.560 95.320 ; 
                RECT 2.880 96.360 127.280 96.680 ; 
                RECT 288.120 96.360 295.560 96.680 ; 
                RECT 2.880 97.720 68.800 98.040 ; 
                RECT 71.200 97.720 127.280 98.040 ; 
                RECT 288.120 97.720 295.560 98.040 ; 
                RECT 2.880 99.080 55.200 99.400 ; 
                RECT 58.280 99.080 89.200 99.400 ; 
                RECT 110.640 99.080 127.280 99.400 ; 
                RECT 288.120 99.080 295.560 99.400 ; 
                RECT 2.880 100.440 53.160 100.760 ; 
                RECT 56.920 100.440 89.200 100.760 ; 
                RECT 110.640 100.440 127.280 100.760 ; 
                RECT 288.120 100.440 295.560 100.760 ; 
                RECT 2.880 101.800 89.200 102.120 ; 
                RECT 110.640 101.800 127.280 102.120 ; 
                RECT 288.120 101.800 295.560 102.120 ; 
                RECT 2.880 103.160 89.200 103.480 ; 
                RECT 110.640 103.160 127.280 103.480 ; 
                RECT 288.120 103.160 295.560 103.480 ; 
                RECT 2.880 104.520 89.200 104.840 ; 
                RECT 110.640 104.520 127.280 104.840 ; 
                RECT 288.120 104.520 295.560 104.840 ; 
                RECT 2.880 105.880 62.000 106.200 ; 
                RECT 70.520 105.880 89.200 106.200 ; 
                RECT 110.640 105.880 127.280 106.200 ; 
                RECT 288.120 105.880 295.560 106.200 ; 
                RECT 2.880 107.240 89.200 107.560 ; 
                RECT 110.640 107.240 127.280 107.560 ; 
                RECT 288.120 107.240 295.560 107.560 ; 
                RECT 2.880 108.600 55.200 108.920 ; 
                RECT 60.320 108.600 89.200 108.920 ; 
                RECT 110.640 108.600 127.280 108.920 ; 
                RECT 288.120 108.600 295.560 108.920 ; 
                RECT 2.880 109.960 89.200 110.280 ; 
                RECT 288.120 109.960 295.560 110.280 ; 
                RECT 2.880 111.320 89.200 111.640 ; 
                RECT 110.640 111.320 124.560 111.640 ; 
                RECT 288.120 111.320 295.560 111.640 ; 
                RECT 2.880 112.680 89.200 113.000 ; 
                RECT 110.640 112.680 121.840 113.000 ; 
                RECT 288.120 112.680 295.560 113.000 ; 
                RECT 2.880 114.040 57.920 114.360 ; 
                RECT 61.000 114.040 89.200 114.360 ; 
                RECT 110.640 114.040 116.400 114.360 ; 
                RECT 288.120 114.040 295.560 114.360 ; 
                RECT 2.880 115.400 32.080 115.720 ; 
                RECT 50.120 115.400 55.200 115.720 ; 
                RECT 58.280 115.400 89.200 115.720 ; 
                RECT 110.640 115.400 116.400 115.720 ; 
                RECT 288.120 115.400 295.560 115.720 ; 
                RECT 2.880 116.760 32.080 117.080 ; 
                RECT 50.120 116.760 89.200 117.080 ; 
                RECT 110.640 116.760 127.280 117.080 ; 
                RECT 288.120 116.760 295.560 117.080 ; 
                RECT 2.880 118.120 32.080 118.440 ; 
                RECT 50.120 118.120 89.200 118.440 ; 
                RECT 110.640 118.120 127.280 118.440 ; 
                RECT 288.120 118.120 295.560 118.440 ; 
                RECT 2.880 119.480 32.080 119.800 ; 
                RECT 50.800 119.480 127.280 119.800 ; 
                RECT 288.120 119.480 295.560 119.800 ; 
                RECT 2.880 120.840 32.080 121.160 ; 
                RECT 50.120 120.840 127.280 121.160 ; 
                RECT 288.120 120.840 295.560 121.160 ; 
                RECT 2.880 122.200 32.080 122.520 ; 
                RECT 50.120 122.200 127.280 122.520 ; 
                RECT 288.120 122.200 295.560 122.520 ; 
                RECT 2.880 123.560 32.080 123.880 ; 
                RECT 50.120 123.560 89.200 123.880 ; 
                RECT 109.960 123.560 117.760 123.880 ; 
                RECT 288.120 123.560 295.560 123.880 ; 
                RECT 2.880 124.920 32.080 125.240 ; 
                RECT 50.120 124.920 56.560 125.240 ; 
                RECT 61.000 124.920 89.200 125.240 ; 
                RECT 109.960 124.920 117.760 125.240 ; 
                RECT 288.120 124.920 295.560 125.240 ; 
                RECT 2.880 126.280 32.080 126.600 ; 
                RECT 50.120 126.280 89.200 126.600 ; 
                RECT 109.960 126.280 120.480 126.600 ; 
                RECT 288.120 126.280 295.560 126.600 ; 
                RECT 2.880 127.640 89.200 127.960 ; 
                RECT 109.960 127.640 123.200 127.960 ; 
                RECT 288.120 127.640 295.560 127.960 ; 
                RECT 2.880 129.000 89.200 129.320 ; 
                RECT 288.120 129.000 295.560 129.320 ; 
                RECT 2.880 130.360 15.760 130.680 ; 
                RECT 31.760 130.360 59.280 130.680 ; 
                RECT 65.080 130.360 89.200 130.680 ; 
                RECT 288.120 130.360 295.560 130.680 ; 
                RECT 2.880 131.720 15.760 132.040 ; 
                RECT 31.760 131.720 38.200 132.040 ; 
                RECT 45.360 131.720 89.200 132.040 ; 
                RECT 109.960 131.720 127.280 132.040 ; 
                RECT 288.120 131.720 295.560 132.040 ; 
                RECT 2.880 133.080 15.760 133.400 ; 
                RECT 50.120 133.080 89.200 133.400 ; 
                RECT 109.960 133.080 127.280 133.400 ; 
                RECT 288.120 133.080 295.560 133.400 ; 
                RECT 2.880 134.440 15.760 134.760 ; 
                RECT 31.760 134.440 89.200 134.760 ; 
                RECT 288.120 134.440 295.560 134.760 ; 
                RECT 2.880 135.800 15.760 136.120 ; 
                RECT 45.360 135.800 53.840 136.120 ; 
                RECT 63.720 135.800 89.200 136.120 ; 
                RECT 109.960 135.800 127.280 136.120 ; 
                RECT 288.120 135.800 295.560 136.120 ; 
                RECT 2.880 137.160 38.200 137.480 ; 
                RECT 58.280 137.160 295.560 137.480 ; 
                RECT 2.880 138.520 28.680 138.840 ; 
                RECT 56.920 138.520 295.560 138.840 ; 
                RECT 2.880 139.880 124.560 140.200 ; 
                RECT 290.840 139.880 295.560 140.200 ; 
                RECT 2.880 141.240 124.560 141.560 ; 
                RECT 290.840 141.240 295.560 141.560 ; 
                RECT 2.880 142.600 23.240 142.920 ; 
                RECT 30.400 142.600 70.160 142.920 ; 
                RECT 290.840 142.600 295.560 142.920 ; 
                RECT 2.880 143.960 21.200 144.280 ; 
                RECT 40.600 143.960 70.160 144.280 ; 
                RECT 290.840 143.960 295.560 144.280 ; 
                RECT 2.880 145.320 21.200 145.640 ; 
                RECT 39.240 145.320 51.120 145.640 ; 
                RECT 52.160 145.320 70.160 145.640 ; 
                RECT 290.840 145.320 295.560 145.640 ; 
                RECT 2.880 146.680 51.120 147.000 ; 
                RECT 52.160 146.680 70.160 147.000 ; 
                RECT 290.840 146.680 295.560 147.000 ; 
                RECT 2.880 148.040 21.200 148.360 ; 
                RECT 31.760 148.040 51.120 148.360 ; 
                RECT 55.560 148.040 70.160 148.360 ; 
                RECT 290.840 148.040 295.560 148.360 ; 
                RECT 2.880 149.400 21.200 149.720 ; 
                RECT 31.760 149.400 51.120 149.720 ; 
                RECT 56.240 149.400 70.160 149.720 ; 
                RECT 290.840 149.400 295.560 149.720 ; 
                RECT 2.880 150.760 21.200 151.080 ; 
                RECT 31.760 150.760 51.120 151.080 ; 
                RECT 56.240 150.760 70.160 151.080 ; 
                RECT 290.840 150.760 295.560 151.080 ; 
                RECT 2.880 152.120 70.160 152.440 ; 
                RECT 290.840 152.120 295.560 152.440 ; 
                RECT 2.880 153.480 70.160 153.800 ; 
                RECT 290.840 153.480 295.560 153.800 ; 
                RECT 2.880 154.840 70.160 155.160 ; 
                RECT 290.840 154.840 295.560 155.160 ; 
                RECT 2.880 156.200 14.400 156.520 ; 
                RECT 17.480 156.200 30.720 156.520 ; 
                RECT 33.120 156.200 70.160 156.520 ; 
                RECT 290.840 156.200 295.560 156.520 ; 
                RECT 2.880 157.560 13.720 157.880 ; 
                RECT 17.480 157.560 70.160 157.880 ; 
                RECT 290.840 157.560 295.560 157.880 ; 
                RECT 2.880 158.920 13.040 159.240 ; 
                RECT 17.480 158.920 34.800 159.240 ; 
                RECT 40.600 158.920 70.160 159.240 ; 
                RECT 290.840 158.920 295.560 159.240 ; 
                RECT 2.880 160.280 12.360 160.600 ; 
                RECT 17.480 160.280 36.160 160.600 ; 
                RECT 39.920 160.280 70.160 160.600 ; 
                RECT 290.840 160.280 295.560 160.600 ; 
                RECT 2.880 161.640 51.120 161.960 ; 
                RECT 52.840 161.640 70.160 161.960 ; 
                RECT 290.840 161.640 295.560 161.960 ; 
                RECT 2.880 163.000 11.680 163.320 ; 
                RECT 17.480 163.000 51.120 163.320 ; 
                RECT 53.520 163.000 70.160 163.320 ; 
                RECT 290.840 163.000 295.560 163.320 ; 
                RECT 2.880 164.360 51.120 164.680 ; 
                RECT 54.200 164.360 70.160 164.680 ; 
                RECT 290.840 164.360 295.560 164.680 ; 
                RECT 2.880 165.720 11.000 166.040 ; 
                RECT 17.480 165.720 30.720 166.040 ; 
                RECT 36.520 165.720 51.120 166.040 ; 
                RECT 52.160 165.720 70.160 166.040 ; 
                RECT 290.840 165.720 295.560 166.040 ; 
                RECT 2.880 167.080 10.320 167.400 ; 
                RECT 17.480 167.080 30.720 167.400 ; 
                RECT 37.200 167.080 51.120 167.400 ; 
                RECT 54.200 167.080 70.160 167.400 ; 
                RECT 290.840 167.080 295.560 167.400 ; 
                RECT 2.880 168.440 9.640 168.760 ; 
                RECT 17.480 168.440 30.720 168.760 ; 
                RECT 37.880 168.440 70.160 168.760 ; 
                RECT 290.840 168.440 295.560 168.760 ; 
                RECT 2.880 169.800 70.160 170.120 ; 
                RECT 290.840 169.800 295.560 170.120 ; 
                RECT 2.880 171.160 70.160 171.480 ; 
                RECT 290.840 171.160 295.560 171.480 ; 
                RECT 2.880 172.520 70.160 172.840 ; 
                RECT 290.840 172.520 295.560 172.840 ; 
                RECT 2.880 173.880 70.160 174.200 ; 
                RECT 290.840 173.880 295.560 174.200 ; 
                RECT 2.880 175.240 70.160 175.560 ; 
                RECT 290.840 175.240 295.560 175.560 ; 
                RECT 2.880 176.600 124.560 176.920 ; 
                RECT 290.840 176.600 295.560 176.920 ; 
                RECT 2.880 177.960 124.560 178.280 ; 
                RECT 290.840 177.960 295.560 178.280 ; 
                RECT 2.880 179.320 124.560 179.640 ; 
                RECT 290.840 179.320 295.560 179.640 ; 
                RECT 2.880 180.680 295.560 181.000 ; 
                RECT 2.880 182.040 295.560 182.360 ; 
                RECT 2.880 183.400 295.560 183.720 ; 
                RECT 2.880 184.760 295.560 185.080 ; 
                RECT 2.880 2.880 295.560 4.240 ; 
                RECT 2.880 186.760 295.560 188.120 ; 
                RECT 128.700 39.630 134.500 40.750 ; 
                RECT 280.600 39.630 286.400 40.750 ; 
                RECT 128.700 45.420 134.500 46.040 ; 
                RECT 280.600 45.420 286.400 46.040 ; 
                RECT 128.700 50.470 134.500 51.110 ; 
                RECT 280.600 50.470 286.400 51.110 ; 
                RECT 128.700 55.640 134.500 56.280 ; 
                RECT 280.600 55.640 286.400 56.280 ; 
                RECT 128.700 83.250 286.400 84.050 ; 
                RECT 128.700 121.980 286.400 122.225 ; 
                RECT 128.700 86.460 286.400 87.260 ; 
                RECT 128.700 108.005 286.400 108.295 ; 
                RECT 128.700 81.570 286.400 82.370 ; 
                RECT 128.700 69.510 286.400 71.310 ; 
                RECT 128.700 78.560 286.400 79.360 ; 
                RECT 128.700 89.645 286.400 90.445 ; 
                RECT 128.700 30.260 286.400 32.060 ; 
                RECT 70.910 142.995 72.830 176.175 ; 
                RECT 89.080 142.995 91.000 176.175 ; 
                RECT 92.920 142.995 94.840 176.175 ; 
                RECT 89.720 58.260 90.610 93.660 ; 
                RECT 96.480 58.260 97.370 93.660 ; 
                RECT 103.025 58.260 104.345 93.660 ; 
                RECT 89.805 123.880 90.915 136.360 ; 
                RECT 97.320 123.880 98.210 136.360 ; 
                RECT 104.185 123.880 105.295 136.360 ; 
                RECT 90.235 99.660 91.345 117.880 ; 
                RECT 98.180 99.660 99.070 117.880 ; 
                RECT 104.615 99.660 105.725 117.880 ; 
                RECT 104.635 48.680 105.745 52.260 ; 
                RECT 22.230 144.060 31.390 144.430 ; 
                RECT 22.230 147.395 31.390 148.285 ; 
                RECT 16.290 130.420 31.130 131.090 ; 
                RECT 16.290 131.720 31.130 132.730 ; 
        END 
    END vss 
    OBS 
        LAYER met1 ;
            RECT 0.000 0.000 298.440 191.000 ; 
        LAYER met2 ;
            RECT 0.000 0.000 298.440 191.000 ; 
    END 
END sram22_64x24m4w8 
END LIBRARY 

