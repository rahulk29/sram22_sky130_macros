VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram22_1024x32m8w32
  CLASS BLOCK ;
  ORIGIN 86.345 184.925 ;
  FOREIGN sram22_1024x32m8w32 -86.345 -184.925 ;
  SIZE 452.85 BY 430.37 ;
  SYMMETRY X Y R90 ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met3 ;
        RECT 357.515 244.04 357.845 245.17 ;
        RECT 357.515 239.875 357.845 240.205 ;
        RECT 357.515 238.515 357.845 238.845 ;
        RECT 357.515 237.155 357.845 237.485 ;
        RECT 357.515 235.17 357.845 235.5 ;
        RECT 357.515 232.995 357.845 233.325 ;
        RECT 357.515 231.415 357.845 231.745 ;
        RECT 357.515 230.565 357.845 230.895 ;
        RECT 357.515 228.255 357.845 228.585 ;
        RECT 357.515 227.405 357.845 227.735 ;
        RECT 357.515 225.095 357.845 225.425 ;
        RECT 357.515 224.245 357.845 224.575 ;
        RECT 357.515 221.935 357.845 222.265 ;
        RECT 357.515 221.085 357.845 221.415 ;
        RECT 357.515 218.775 357.845 219.105 ;
        RECT 357.515 217.195 357.845 217.525 ;
        RECT 357.515 216.345 357.845 216.675 ;
        RECT 357.515 214.035 357.845 214.365 ;
        RECT 357.515 213.185 357.845 213.515 ;
        RECT 357.515 210.875 357.845 211.205 ;
        RECT 357.515 210.025 357.845 210.355 ;
        RECT 357.515 207.715 357.845 208.045 ;
        RECT 357.515 206.865 357.845 207.195 ;
        RECT 357.515 204.555 357.845 204.885 ;
        RECT 357.515 202.975 357.845 203.305 ;
        RECT 357.515 202.125 357.845 202.455 ;
        RECT 357.515 199.815 357.845 200.145 ;
        RECT 357.515 198.965 357.845 199.295 ;
        RECT 357.515 196.655 357.845 196.985 ;
        RECT 357.515 195.805 357.845 196.135 ;
        RECT 357.515 193.495 357.845 193.825 ;
        RECT 357.515 192.645 357.845 192.975 ;
        RECT 357.515 190.335 357.845 190.665 ;
        RECT 357.515 188.755 357.845 189.085 ;
        RECT 357.515 187.905 357.845 188.235 ;
        RECT 357.515 185.595 357.845 185.925 ;
        RECT 357.515 184.745 357.845 185.075 ;
        RECT 357.515 182.435 357.845 182.765 ;
        RECT 357.515 181.585 357.845 181.915 ;
        RECT 357.515 179.275 357.845 179.605 ;
        RECT 357.515 178.425 357.845 178.755 ;
        RECT 357.515 176.115 357.845 176.445 ;
        RECT 357.515 174.535 357.845 174.865 ;
        RECT 357.515 173.685 357.845 174.015 ;
        RECT 357.515 171.375 357.845 171.705 ;
        RECT 357.515 170.525 357.845 170.855 ;
        RECT 357.515 168.215 357.845 168.545 ;
        RECT 357.515 167.365 357.845 167.695 ;
        RECT 357.515 165.055 357.845 165.385 ;
        RECT 357.515 164.205 357.845 164.535 ;
        RECT 357.515 161.895 357.845 162.225 ;
        RECT 357.515 160.315 357.845 160.645 ;
        RECT 357.515 159.465 357.845 159.795 ;
        RECT 357.515 157.155 357.845 157.485 ;
        RECT 357.515 156.305 357.845 156.635 ;
        RECT 357.515 153.995 357.845 154.325 ;
        RECT 357.515 153.145 357.845 153.475 ;
        RECT 357.515 150.835 357.845 151.165 ;
        RECT 357.515 149.985 357.845 150.315 ;
        RECT 357.515 147.675 357.845 148.005 ;
        RECT 357.515 146.095 357.845 146.425 ;
        RECT 357.515 145.245 357.845 145.575 ;
        RECT 357.515 142.935 357.845 143.265 ;
        RECT 357.515 142.085 357.845 142.415 ;
        RECT 357.515 139.775 357.845 140.105 ;
        RECT 357.515 138.925 357.845 139.255 ;
        RECT 357.515 136.615 357.845 136.945 ;
        RECT 357.515 135.765 357.845 136.095 ;
        RECT 357.515 133.455 357.845 133.785 ;
        RECT 357.515 131.875 357.845 132.205 ;
        RECT 357.515 131.025 357.845 131.355 ;
        RECT 357.515 128.715 357.845 129.045 ;
        RECT 357.515 127.865 357.845 128.195 ;
        RECT 357.515 125.555 357.845 125.885 ;
        RECT 357.515 124.705 357.845 125.035 ;
        RECT 357.515 122.395 357.845 122.725 ;
        RECT 357.515 121.545 357.845 121.875 ;
        RECT 357.515 119.235 357.845 119.565 ;
        RECT 357.515 117.655 357.845 117.985 ;
        RECT 357.515 116.805 357.845 117.135 ;
        RECT 357.515 114.495 357.845 114.825 ;
        RECT 357.515 113.645 357.845 113.975 ;
        RECT 357.515 111.335 357.845 111.665 ;
        RECT 357.515 110.485 357.845 110.815 ;
        RECT 357.515 108.175 357.845 108.505 ;
        RECT 357.515 107.325 357.845 107.655 ;
        RECT 357.515 105.015 357.845 105.345 ;
        RECT 357.515 103.435 357.845 103.765 ;
        RECT 357.515 102.585 357.845 102.915 ;
        RECT 357.515 100.275 357.845 100.605 ;
        RECT 357.515 99.425 357.845 99.755 ;
        RECT 357.515 97.115 357.845 97.445 ;
        RECT 357.515 96.265 357.845 96.595 ;
        RECT 357.515 93.955 357.845 94.285 ;
        RECT 357.515 93.105 357.845 93.435 ;
        RECT 357.515 90.795 357.845 91.125 ;
        RECT 357.515 89.215 357.845 89.545 ;
        RECT 357.515 88.365 357.845 88.695 ;
        RECT 357.515 86.055 357.845 86.385 ;
        RECT 357.515 85.205 357.845 85.535 ;
        RECT 357.515 82.895 357.845 83.225 ;
        RECT 357.515 82.045 357.845 82.375 ;
        RECT 357.515 79.735 357.845 80.065 ;
        RECT 357.515 78.885 357.845 79.215 ;
        RECT 357.515 76.575 357.845 76.905 ;
        RECT 357.515 74.995 357.845 75.325 ;
        RECT 357.515 74.145 357.845 74.475 ;
        RECT 357.515 71.835 357.845 72.165 ;
        RECT 357.515 70.985 357.845 71.315 ;
        RECT 357.515 68.675 357.845 69.005 ;
        RECT 357.515 67.825 357.845 68.155 ;
        RECT 357.515 65.515 357.845 65.845 ;
        RECT 357.515 64.665 357.845 64.995 ;
        RECT 357.515 62.355 357.845 62.685 ;
        RECT 357.515 60.775 357.845 61.105 ;
        RECT 357.515 59.925 357.845 60.255 ;
        RECT 357.515 57.615 357.845 57.945 ;
        RECT 357.515 56.765 357.845 57.095 ;
        RECT 357.515 54.455 357.845 54.785 ;
        RECT 357.515 53.605 357.845 53.935 ;
        RECT 357.515 51.295 357.845 51.625 ;
        RECT 357.515 50.445 357.845 50.775 ;
        RECT 357.515 48.135 357.845 48.465 ;
        RECT 357.515 46.555 357.845 46.885 ;
        RECT 357.515 45.705 357.845 46.035 ;
        RECT 357.515 43.395 357.845 43.725 ;
        RECT 357.515 42.545 357.845 42.875 ;
        RECT 357.515 40.235 357.845 40.565 ;
        RECT 357.515 39.385 357.845 39.715 ;
        RECT 357.515 37.075 357.845 37.405 ;
        RECT 357.515 36.225 357.845 36.555 ;
        RECT 357.515 33.915 357.845 34.245 ;
        RECT 357.515 32.335 357.845 32.665 ;
        RECT 357.515 31.485 357.845 31.815 ;
        RECT 357.515 29.175 357.845 29.505 ;
        RECT 357.515 28.325 357.845 28.655 ;
        RECT 357.515 26.015 357.845 26.345 ;
        RECT 357.515 25.165 357.845 25.495 ;
        RECT 357.515 22.855 357.845 23.185 ;
        RECT 357.515 22.005 357.845 22.335 ;
        RECT 357.515 19.695 357.845 20.025 ;
        RECT 357.515 18.115 357.845 18.445 ;
        RECT 357.515 17.265 357.845 17.595 ;
        RECT 357.515 14.955 357.845 15.285 ;
        RECT 357.515 14.105 357.845 14.435 ;
        RECT 357.515 11.795 357.845 12.125 ;
        RECT 357.515 10.945 357.845 11.275 ;
        RECT 357.515 8.635 357.845 8.965 ;
        RECT 357.515 7.785 357.845 8.115 ;
        RECT 357.515 5.475 357.845 5.805 ;
        RECT 357.515 3.895 357.845 4.225 ;
        RECT 357.515 3.045 357.845 3.375 ;
        RECT 357.515 0.87 357.845 1.2 ;
        RECT 357.515 -0.845 357.845 -0.515 ;
        RECT 357.515 -2.205 357.845 -1.875 ;
        RECT 357.515 -3.565 357.845 -3.235 ;
        RECT 357.515 -4.925 357.845 -4.595 ;
        RECT 357.515 -6.285 357.845 -5.955 ;
        RECT 357.515 -7.645 357.845 -7.315 ;
        RECT 357.515 -9.005 357.845 -8.675 ;
        RECT 357.515 -10.365 357.845 -10.035 ;
        RECT 357.515 -11.725 357.845 -11.395 ;
        RECT 357.515 -13.085 357.845 -12.755 ;
        RECT 357.515 -14.445 357.845 -14.115 ;
        RECT 357.515 -15.805 357.845 -15.475 ;
        RECT 357.515 -17.165 357.845 -16.835 ;
        RECT 357.515 -18.525 357.845 -18.195 ;
        RECT 357.515 -19.885 357.845 -19.555 ;
        RECT 357.515 -21.245 357.845 -20.915 ;
        RECT 357.515 -22.605 357.845 -22.275 ;
        RECT 357.515 -23.965 357.845 -23.635 ;
        RECT 357.515 -25.325 357.845 -24.995 ;
        RECT 357.515 -26.685 357.845 -26.355 ;
        RECT 357.515 -28.045 357.845 -27.715 ;
        RECT 357.515 -29.405 357.845 -29.075 ;
        RECT 357.515 -30.765 357.845 -30.435 ;
        RECT 357.515 -32.125 357.845 -31.795 ;
        RECT 357.515 -33.485 357.845 -33.155 ;
        RECT 357.515 -34.845 357.845 -34.515 ;
        RECT 357.515 -36.205 357.845 -35.875 ;
        RECT 357.515 -37.565 357.845 -37.235 ;
        RECT 357.515 -38.925 357.845 -38.595 ;
        RECT 357.515 -40.285 357.845 -39.955 ;
        RECT 357.515 -41.645 357.845 -41.315 ;
        RECT 357.515 -43.005 357.845 -42.675 ;
        RECT 357.515 -44.365 357.845 -44.035 ;
        RECT 357.515 -45.725 357.845 -45.395 ;
        RECT 357.515 -47.085 357.845 -46.755 ;
        RECT 357.515 -48.445 357.845 -48.115 ;
        RECT 357.515 -49.805 357.845 -49.475 ;
        RECT 357.515 -51.165 357.845 -50.835 ;
        RECT 357.515 -52.525 357.845 -52.195 ;
        RECT 357.515 -53.885 357.845 -53.555 ;
        RECT 357.515 -55.245 357.845 -54.915 ;
        RECT 357.515 -56.605 357.845 -56.275 ;
        RECT 357.515 -57.965 357.845 -57.635 ;
        RECT 357.515 -59.325 357.845 -58.995 ;
        RECT 357.515 -60.685 357.845 -60.355 ;
        RECT 357.515 -62.045 357.845 -61.715 ;
        RECT 357.515 -63.405 357.845 -63.075 ;
        RECT 357.515 -64.765 357.845 -64.435 ;
        RECT 357.515 -66.125 357.845 -65.795 ;
        RECT 357.515 -67.485 357.845 -67.155 ;
        RECT 357.515 -68.845 357.845 -68.515 ;
        RECT 357.515 -70.205 357.845 -69.875 ;
        RECT 357.515 -71.565 357.845 -71.235 ;
        RECT 357.515 -72.925 357.845 -72.595 ;
        RECT 357.515 -74.285 357.845 -73.955 ;
        RECT 357.515 -75.645 357.845 -75.315 ;
        RECT 357.515 -77.005 357.845 -76.675 ;
        RECT 357.515 -78.365 357.845 -78.035 ;
        RECT 357.515 -79.725 357.845 -79.395 ;
        RECT 357.515 -81.085 357.845 -80.755 ;
        RECT 357.515 -82.445 357.845 -82.115 ;
        RECT 357.515 -83.805 357.845 -83.475 ;
        RECT 357.515 -85.165 357.845 -84.835 ;
        RECT 357.515 -86.525 357.845 -86.195 ;
        RECT 357.515 -87.885 357.845 -87.555 ;
        RECT 357.515 -89.245 357.845 -88.915 ;
        RECT 357.515 -90.605 357.845 -90.275 ;
        RECT 357.515 -91.965 357.845 -91.635 ;
        RECT 357.515 -93.325 357.845 -92.995 ;
        RECT 357.515 -94.685 357.845 -94.355 ;
        RECT 357.515 -96.045 357.845 -95.715 ;
        RECT 357.515 -97.405 357.845 -97.075 ;
        RECT 357.515 -98.765 357.845 -98.435 ;
        RECT 357.515 -100.125 357.845 -99.795 ;
        RECT 357.515 -101.485 357.845 -101.155 ;
        RECT 357.515 -102.845 357.845 -102.515 ;
        RECT 357.515 -104.205 357.845 -103.875 ;
        RECT 357.515 -105.565 357.845 -105.235 ;
        RECT 357.515 -106.925 357.845 -106.595 ;
        RECT 357.515 -108.285 357.845 -107.955 ;
        RECT 357.515 -109.645 357.845 -109.315 ;
        RECT 357.515 -111.005 357.845 -110.675 ;
        RECT 357.515 -112.365 357.845 -112.035 ;
        RECT 357.515 -113.725 357.845 -113.395 ;
        RECT 357.515 -115.085 357.845 -114.755 ;
        RECT 357.515 -116.445 357.845 -116.115 ;
        RECT 357.515 -117.805 357.845 -117.475 ;
        RECT 357.515 -119.165 357.845 -118.835 ;
        RECT 357.515 -120.525 357.845 -120.195 ;
        RECT 357.515 -121.885 357.845 -121.555 ;
        RECT 357.515 -123.245 357.845 -122.915 ;
        RECT 357.515 -124.605 357.845 -124.275 ;
        RECT 357.515 -125.965 357.845 -125.635 ;
        RECT 357.515 -127.325 357.845 -126.995 ;
        RECT 357.515 -128.685 357.845 -128.355 ;
        RECT 357.515 -130.045 357.845 -129.715 ;
        RECT 357.515 -131.405 357.845 -131.075 ;
        RECT 357.515 -132.765 357.845 -132.435 ;
        RECT 357.515 -134.125 357.845 -133.795 ;
        RECT 357.515 -135.485 357.845 -135.155 ;
        RECT 357.515 -136.845 357.845 -136.515 ;
        RECT 357.515 -138.205 357.845 -137.875 ;
        RECT 357.515 -139.565 357.845 -139.235 ;
        RECT 357.515 -140.925 357.845 -140.595 ;
        RECT 357.515 -142.285 357.845 -141.955 ;
        RECT 357.515 -143.645 357.845 -143.315 ;
        RECT 357.515 -145.005 357.845 -144.675 ;
        RECT 357.515 -146.365 357.845 -146.035 ;
        RECT 357.515 -147.725 357.845 -147.395 ;
        RECT 357.515 -149.085 357.845 -148.755 ;
        RECT 357.515 -150.445 357.845 -150.115 ;
        RECT 357.515 -151.805 357.845 -151.475 ;
        RECT 357.515 -153.165 357.845 -152.835 ;
        RECT 357.515 -154.525 357.845 -154.195 ;
        RECT 357.515 -155.885 357.845 -155.555 ;
        RECT 357.515 -157.245 357.845 -156.915 ;
        RECT 357.515 -158.605 357.845 -158.275 ;
        RECT 357.515 -159.965 357.845 -159.635 ;
        RECT 357.515 -161.325 357.845 -160.995 ;
        RECT 357.515 -162.685 357.845 -162.355 ;
        RECT 357.515 -164.045 357.845 -163.715 ;
        RECT 357.515 -165.405 357.845 -165.075 ;
        RECT 357.515 -166.765 357.845 -166.435 ;
        RECT 357.515 -168.125 357.845 -167.795 ;
        RECT 357.515 -169.485 357.845 -169.155 ;
        RECT 357.515 -170.845 357.845 -170.515 ;
        RECT 357.515 -172.205 357.845 -171.875 ;
        RECT 357.515 -173.565 357.845 -173.235 ;
        RECT 357.515 -174.925 357.845 -174.595 ;
        RECT 357.515 -176.285 357.845 -175.955 ;
        RECT 357.515 -177.645 357.845 -177.315 ;
        RECT 357.515 -179.005 357.845 -178.675 ;
        RECT 357.515 -184.65 357.845 -183.52 ;
        RECT 357.52 -184.765 357.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.875 244.04 359.205 245.17 ;
        RECT 358.875 239.875 359.205 240.205 ;
        RECT 358.875 238.515 359.205 238.845 ;
        RECT 358.875 237.155 359.205 237.485 ;
        RECT 358.875 235.17 359.205 235.5 ;
        RECT 358.875 232.995 359.205 233.325 ;
        RECT 358.875 231.415 359.205 231.745 ;
        RECT 358.875 230.565 359.205 230.895 ;
        RECT 358.875 228.255 359.205 228.585 ;
        RECT 358.875 227.405 359.205 227.735 ;
        RECT 358.875 225.095 359.205 225.425 ;
        RECT 358.875 224.245 359.205 224.575 ;
        RECT 358.875 221.935 359.205 222.265 ;
        RECT 358.875 221.085 359.205 221.415 ;
        RECT 358.875 218.775 359.205 219.105 ;
        RECT 358.875 217.195 359.205 217.525 ;
        RECT 358.875 216.345 359.205 216.675 ;
        RECT 358.875 214.035 359.205 214.365 ;
        RECT 358.875 213.185 359.205 213.515 ;
        RECT 358.875 210.875 359.205 211.205 ;
        RECT 358.875 210.025 359.205 210.355 ;
        RECT 358.875 207.715 359.205 208.045 ;
        RECT 358.875 206.865 359.205 207.195 ;
        RECT 358.875 204.555 359.205 204.885 ;
        RECT 358.875 202.975 359.205 203.305 ;
        RECT 358.875 202.125 359.205 202.455 ;
        RECT 358.875 199.815 359.205 200.145 ;
        RECT 358.875 198.965 359.205 199.295 ;
        RECT 358.875 196.655 359.205 196.985 ;
        RECT 358.875 195.805 359.205 196.135 ;
        RECT 358.875 193.495 359.205 193.825 ;
        RECT 358.875 192.645 359.205 192.975 ;
        RECT 358.875 190.335 359.205 190.665 ;
        RECT 358.875 188.755 359.205 189.085 ;
        RECT 358.875 187.905 359.205 188.235 ;
        RECT 358.875 185.595 359.205 185.925 ;
        RECT 358.875 184.745 359.205 185.075 ;
        RECT 358.875 182.435 359.205 182.765 ;
        RECT 358.875 181.585 359.205 181.915 ;
        RECT 358.875 179.275 359.205 179.605 ;
        RECT 358.875 178.425 359.205 178.755 ;
        RECT 358.875 176.115 359.205 176.445 ;
        RECT 358.875 174.535 359.205 174.865 ;
        RECT 358.875 173.685 359.205 174.015 ;
        RECT 358.875 171.375 359.205 171.705 ;
        RECT 358.875 170.525 359.205 170.855 ;
        RECT 358.875 168.215 359.205 168.545 ;
        RECT 358.875 167.365 359.205 167.695 ;
        RECT 358.875 165.055 359.205 165.385 ;
        RECT 358.875 164.205 359.205 164.535 ;
        RECT 358.875 161.895 359.205 162.225 ;
        RECT 358.875 160.315 359.205 160.645 ;
        RECT 358.875 159.465 359.205 159.795 ;
        RECT 358.875 157.155 359.205 157.485 ;
        RECT 358.875 156.305 359.205 156.635 ;
        RECT 358.875 153.995 359.205 154.325 ;
        RECT 358.875 153.145 359.205 153.475 ;
        RECT 358.875 150.835 359.205 151.165 ;
        RECT 358.875 149.985 359.205 150.315 ;
        RECT 358.875 147.675 359.205 148.005 ;
        RECT 358.875 146.095 359.205 146.425 ;
        RECT 358.875 145.245 359.205 145.575 ;
        RECT 358.875 142.935 359.205 143.265 ;
        RECT 358.875 142.085 359.205 142.415 ;
        RECT 358.875 139.775 359.205 140.105 ;
        RECT 358.875 138.925 359.205 139.255 ;
        RECT 358.875 136.615 359.205 136.945 ;
        RECT 358.875 135.765 359.205 136.095 ;
        RECT 358.875 133.455 359.205 133.785 ;
        RECT 358.875 131.875 359.205 132.205 ;
        RECT 358.875 131.025 359.205 131.355 ;
        RECT 358.875 128.715 359.205 129.045 ;
        RECT 358.875 127.865 359.205 128.195 ;
        RECT 358.875 125.555 359.205 125.885 ;
        RECT 358.875 124.705 359.205 125.035 ;
        RECT 358.875 122.395 359.205 122.725 ;
        RECT 358.875 121.545 359.205 121.875 ;
        RECT 358.875 119.235 359.205 119.565 ;
        RECT 358.875 117.655 359.205 117.985 ;
        RECT 358.875 116.805 359.205 117.135 ;
        RECT 358.875 114.495 359.205 114.825 ;
        RECT 358.875 113.645 359.205 113.975 ;
        RECT 358.875 111.335 359.205 111.665 ;
        RECT 358.875 110.485 359.205 110.815 ;
        RECT 358.875 108.175 359.205 108.505 ;
        RECT 358.875 107.325 359.205 107.655 ;
        RECT 358.875 105.015 359.205 105.345 ;
        RECT 358.875 103.435 359.205 103.765 ;
        RECT 358.875 102.585 359.205 102.915 ;
        RECT 358.875 100.275 359.205 100.605 ;
        RECT 358.875 99.425 359.205 99.755 ;
        RECT 358.875 97.115 359.205 97.445 ;
        RECT 358.875 96.265 359.205 96.595 ;
        RECT 358.875 93.955 359.205 94.285 ;
        RECT 358.875 93.105 359.205 93.435 ;
        RECT 358.875 90.795 359.205 91.125 ;
        RECT 358.875 89.215 359.205 89.545 ;
        RECT 358.875 88.365 359.205 88.695 ;
        RECT 358.875 86.055 359.205 86.385 ;
        RECT 358.875 85.205 359.205 85.535 ;
        RECT 358.875 82.895 359.205 83.225 ;
        RECT 358.875 82.045 359.205 82.375 ;
        RECT 358.875 79.735 359.205 80.065 ;
        RECT 358.875 78.885 359.205 79.215 ;
        RECT 358.875 76.575 359.205 76.905 ;
        RECT 358.875 74.995 359.205 75.325 ;
        RECT 358.875 74.145 359.205 74.475 ;
        RECT 358.875 71.835 359.205 72.165 ;
        RECT 358.875 70.985 359.205 71.315 ;
        RECT 358.875 68.675 359.205 69.005 ;
        RECT 358.875 67.825 359.205 68.155 ;
        RECT 358.875 65.515 359.205 65.845 ;
        RECT 358.875 64.665 359.205 64.995 ;
        RECT 358.875 62.355 359.205 62.685 ;
        RECT 358.875 60.775 359.205 61.105 ;
        RECT 358.875 59.925 359.205 60.255 ;
        RECT 358.875 57.615 359.205 57.945 ;
        RECT 358.875 56.765 359.205 57.095 ;
        RECT 358.875 54.455 359.205 54.785 ;
        RECT 358.875 53.605 359.205 53.935 ;
        RECT 358.875 51.295 359.205 51.625 ;
        RECT 358.875 50.445 359.205 50.775 ;
        RECT 358.875 48.135 359.205 48.465 ;
        RECT 358.875 46.555 359.205 46.885 ;
        RECT 358.875 45.705 359.205 46.035 ;
        RECT 358.875 43.395 359.205 43.725 ;
        RECT 358.875 42.545 359.205 42.875 ;
        RECT 358.875 40.235 359.205 40.565 ;
        RECT 358.875 39.385 359.205 39.715 ;
        RECT 358.875 37.075 359.205 37.405 ;
        RECT 358.875 36.225 359.205 36.555 ;
        RECT 358.875 33.915 359.205 34.245 ;
        RECT 358.875 32.335 359.205 32.665 ;
        RECT 358.875 31.485 359.205 31.815 ;
        RECT 358.875 29.175 359.205 29.505 ;
        RECT 358.875 28.325 359.205 28.655 ;
        RECT 358.875 26.015 359.205 26.345 ;
        RECT 358.875 25.165 359.205 25.495 ;
        RECT 358.875 22.855 359.205 23.185 ;
        RECT 358.875 22.005 359.205 22.335 ;
        RECT 358.875 19.695 359.205 20.025 ;
        RECT 358.875 18.115 359.205 18.445 ;
        RECT 358.875 17.265 359.205 17.595 ;
        RECT 358.875 14.955 359.205 15.285 ;
        RECT 358.875 14.105 359.205 14.435 ;
        RECT 358.875 11.795 359.205 12.125 ;
        RECT 358.875 10.945 359.205 11.275 ;
        RECT 358.875 8.635 359.205 8.965 ;
        RECT 358.875 7.785 359.205 8.115 ;
        RECT 358.875 5.475 359.205 5.805 ;
        RECT 358.875 3.895 359.205 4.225 ;
        RECT 358.875 3.045 359.205 3.375 ;
        RECT 358.875 0.87 359.205 1.2 ;
        RECT 358.875 -0.845 359.205 -0.515 ;
        RECT 358.875 -2.205 359.205 -1.875 ;
        RECT 358.875 -3.565 359.205 -3.235 ;
        RECT 358.875 -4.925 359.205 -4.595 ;
        RECT 358.875 -6.285 359.205 -5.955 ;
        RECT 358.875 -7.645 359.205 -7.315 ;
        RECT 358.875 -9.005 359.205 -8.675 ;
        RECT 358.875 -10.365 359.205 -10.035 ;
        RECT 358.875 -11.725 359.205 -11.395 ;
        RECT 358.875 -13.085 359.205 -12.755 ;
        RECT 358.875 -14.445 359.205 -14.115 ;
        RECT 358.875 -15.805 359.205 -15.475 ;
        RECT 358.875 -17.165 359.205 -16.835 ;
        RECT 358.875 -18.525 359.205 -18.195 ;
        RECT 358.875 -19.885 359.205 -19.555 ;
        RECT 358.875 -21.245 359.205 -20.915 ;
        RECT 358.875 -22.605 359.205 -22.275 ;
        RECT 358.875 -23.965 359.205 -23.635 ;
        RECT 358.875 -25.325 359.205 -24.995 ;
        RECT 358.875 -26.685 359.205 -26.355 ;
        RECT 358.875 -28.045 359.205 -27.715 ;
        RECT 358.875 -29.405 359.205 -29.075 ;
        RECT 358.875 -30.765 359.205 -30.435 ;
        RECT 358.875 -32.125 359.205 -31.795 ;
        RECT 358.875 -33.485 359.205 -33.155 ;
        RECT 358.875 -34.845 359.205 -34.515 ;
        RECT 358.875 -36.205 359.205 -35.875 ;
        RECT 358.875 -37.565 359.205 -37.235 ;
        RECT 358.875 -38.925 359.205 -38.595 ;
        RECT 358.875 -40.285 359.205 -39.955 ;
        RECT 358.875 -41.645 359.205 -41.315 ;
        RECT 358.875 -43.005 359.205 -42.675 ;
        RECT 358.875 -44.365 359.205 -44.035 ;
        RECT 358.875 -45.725 359.205 -45.395 ;
        RECT 358.875 -47.085 359.205 -46.755 ;
        RECT 358.875 -48.445 359.205 -48.115 ;
        RECT 358.875 -49.805 359.205 -49.475 ;
        RECT 358.875 -51.165 359.205 -50.835 ;
        RECT 358.875 -52.525 359.205 -52.195 ;
        RECT 358.875 -53.885 359.205 -53.555 ;
        RECT 358.875 -55.245 359.205 -54.915 ;
        RECT 358.875 -56.605 359.205 -56.275 ;
        RECT 358.875 -57.965 359.205 -57.635 ;
        RECT 358.875 -59.325 359.205 -58.995 ;
        RECT 358.875 -60.685 359.205 -60.355 ;
        RECT 358.875 -62.045 359.205 -61.715 ;
        RECT 358.875 -63.405 359.205 -63.075 ;
        RECT 358.875 -64.765 359.205 -64.435 ;
        RECT 358.875 -66.125 359.205 -65.795 ;
        RECT 358.875 -67.485 359.205 -67.155 ;
        RECT 358.875 -68.845 359.205 -68.515 ;
        RECT 358.875 -70.205 359.205 -69.875 ;
        RECT 358.875 -71.565 359.205 -71.235 ;
        RECT 358.875 -72.925 359.205 -72.595 ;
        RECT 358.875 -74.285 359.205 -73.955 ;
        RECT 358.875 -75.645 359.205 -75.315 ;
        RECT 358.875 -77.005 359.205 -76.675 ;
        RECT 358.875 -78.365 359.205 -78.035 ;
        RECT 358.875 -79.725 359.205 -79.395 ;
        RECT 358.875 -81.085 359.205 -80.755 ;
        RECT 358.875 -82.445 359.205 -82.115 ;
        RECT 358.875 -83.805 359.205 -83.475 ;
        RECT 358.875 -85.165 359.205 -84.835 ;
        RECT 358.875 -86.525 359.205 -86.195 ;
        RECT 358.875 -87.885 359.205 -87.555 ;
        RECT 358.875 -89.245 359.205 -88.915 ;
        RECT 358.875 -90.605 359.205 -90.275 ;
        RECT 358.875 -91.965 359.205 -91.635 ;
        RECT 358.875 -93.325 359.205 -92.995 ;
        RECT 358.875 -94.685 359.205 -94.355 ;
        RECT 358.875 -96.045 359.205 -95.715 ;
        RECT 358.875 -97.405 359.205 -97.075 ;
        RECT 358.875 -98.765 359.205 -98.435 ;
        RECT 358.875 -100.125 359.205 -99.795 ;
        RECT 358.875 -101.485 359.205 -101.155 ;
        RECT 358.875 -102.845 359.205 -102.515 ;
        RECT 358.875 -104.205 359.205 -103.875 ;
        RECT 358.875 -105.565 359.205 -105.235 ;
        RECT 358.875 -106.925 359.205 -106.595 ;
        RECT 358.875 -108.285 359.205 -107.955 ;
        RECT 358.875 -109.645 359.205 -109.315 ;
        RECT 358.875 -111.005 359.205 -110.675 ;
        RECT 358.875 -112.365 359.205 -112.035 ;
        RECT 358.875 -113.725 359.205 -113.395 ;
        RECT 358.875 -115.085 359.205 -114.755 ;
        RECT 358.875 -116.445 359.205 -116.115 ;
        RECT 358.875 -117.805 359.205 -117.475 ;
        RECT 358.875 -119.165 359.205 -118.835 ;
        RECT 358.875 -120.525 359.205 -120.195 ;
        RECT 358.875 -121.885 359.205 -121.555 ;
        RECT 358.875 -123.245 359.205 -122.915 ;
        RECT 358.875 -124.605 359.205 -124.275 ;
        RECT 358.875 -125.965 359.205 -125.635 ;
        RECT 358.875 -127.325 359.205 -126.995 ;
        RECT 358.875 -128.685 359.205 -128.355 ;
        RECT 358.875 -130.045 359.205 -129.715 ;
        RECT 358.875 -131.405 359.205 -131.075 ;
        RECT 358.875 -132.765 359.205 -132.435 ;
        RECT 358.875 -134.125 359.205 -133.795 ;
        RECT 358.875 -135.485 359.205 -135.155 ;
        RECT 358.875 -136.845 359.205 -136.515 ;
        RECT 358.875 -138.205 359.205 -137.875 ;
        RECT 358.875 -139.565 359.205 -139.235 ;
        RECT 358.875 -140.925 359.205 -140.595 ;
        RECT 358.875 -142.285 359.205 -141.955 ;
        RECT 358.875 -143.645 359.205 -143.315 ;
        RECT 358.875 -145.005 359.205 -144.675 ;
        RECT 358.875 -146.365 359.205 -146.035 ;
        RECT 358.875 -147.725 359.205 -147.395 ;
        RECT 358.875 -149.085 359.205 -148.755 ;
        RECT 358.875 -150.445 359.205 -150.115 ;
        RECT 358.875 -151.805 359.205 -151.475 ;
        RECT 358.875 -153.165 359.205 -152.835 ;
        RECT 358.875 -154.525 359.205 -154.195 ;
        RECT 358.875 -155.885 359.205 -155.555 ;
        RECT 358.875 -157.245 359.205 -156.915 ;
        RECT 358.875 -158.605 359.205 -158.275 ;
        RECT 358.875 -159.965 359.205 -159.635 ;
        RECT 358.875 -161.325 359.205 -160.995 ;
        RECT 358.875 -162.685 359.205 -162.355 ;
        RECT 358.875 -164.045 359.205 -163.715 ;
        RECT 358.875 -165.405 359.205 -165.075 ;
        RECT 358.875 -166.765 359.205 -166.435 ;
        RECT 358.875 -168.125 359.205 -167.795 ;
        RECT 358.875 -169.485 359.205 -169.155 ;
        RECT 358.875 -170.845 359.205 -170.515 ;
        RECT 358.875 -172.205 359.205 -171.875 ;
        RECT 358.875 -173.565 359.205 -173.235 ;
        RECT 358.875 -174.925 359.205 -174.595 ;
        RECT 358.875 -176.285 359.205 -175.955 ;
        RECT 358.875 -177.645 359.205 -177.315 ;
        RECT 358.875 -179.005 359.205 -178.675 ;
        RECT 358.875 -184.65 359.205 -183.52 ;
        RECT 358.88 -184.765 359.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.235 244.04 360.565 245.17 ;
        RECT 360.235 239.875 360.565 240.205 ;
        RECT 360.235 238.515 360.565 238.845 ;
        RECT 360.235 237.155 360.565 237.485 ;
        RECT 360.235 235.17 360.565 235.5 ;
        RECT 360.235 232.995 360.565 233.325 ;
        RECT 360.235 231.415 360.565 231.745 ;
        RECT 360.235 230.565 360.565 230.895 ;
        RECT 360.235 228.255 360.565 228.585 ;
        RECT 360.235 227.405 360.565 227.735 ;
        RECT 360.235 225.095 360.565 225.425 ;
        RECT 360.235 224.245 360.565 224.575 ;
        RECT 360.235 221.935 360.565 222.265 ;
        RECT 360.235 221.085 360.565 221.415 ;
        RECT 360.235 218.775 360.565 219.105 ;
        RECT 360.235 217.195 360.565 217.525 ;
        RECT 360.235 216.345 360.565 216.675 ;
        RECT 360.235 214.035 360.565 214.365 ;
        RECT 360.235 213.185 360.565 213.515 ;
        RECT 360.235 210.875 360.565 211.205 ;
        RECT 360.235 210.025 360.565 210.355 ;
        RECT 360.235 207.715 360.565 208.045 ;
        RECT 360.235 206.865 360.565 207.195 ;
        RECT 360.235 204.555 360.565 204.885 ;
        RECT 360.235 202.975 360.565 203.305 ;
        RECT 360.235 202.125 360.565 202.455 ;
        RECT 360.235 199.815 360.565 200.145 ;
        RECT 360.235 198.965 360.565 199.295 ;
        RECT 360.235 196.655 360.565 196.985 ;
        RECT 360.235 195.805 360.565 196.135 ;
        RECT 360.235 193.495 360.565 193.825 ;
        RECT 360.235 192.645 360.565 192.975 ;
        RECT 360.235 190.335 360.565 190.665 ;
        RECT 360.235 188.755 360.565 189.085 ;
        RECT 360.235 187.905 360.565 188.235 ;
        RECT 360.235 185.595 360.565 185.925 ;
        RECT 360.235 184.745 360.565 185.075 ;
        RECT 360.235 182.435 360.565 182.765 ;
        RECT 360.235 181.585 360.565 181.915 ;
        RECT 360.235 179.275 360.565 179.605 ;
        RECT 360.235 178.425 360.565 178.755 ;
        RECT 360.235 176.115 360.565 176.445 ;
        RECT 360.235 174.535 360.565 174.865 ;
        RECT 360.235 173.685 360.565 174.015 ;
        RECT 360.235 171.375 360.565 171.705 ;
        RECT 360.235 170.525 360.565 170.855 ;
        RECT 360.235 168.215 360.565 168.545 ;
        RECT 360.235 167.365 360.565 167.695 ;
        RECT 360.235 165.055 360.565 165.385 ;
        RECT 360.235 164.205 360.565 164.535 ;
        RECT 360.235 161.895 360.565 162.225 ;
        RECT 360.235 160.315 360.565 160.645 ;
        RECT 360.235 159.465 360.565 159.795 ;
        RECT 360.235 157.155 360.565 157.485 ;
        RECT 360.235 156.305 360.565 156.635 ;
        RECT 360.235 153.995 360.565 154.325 ;
        RECT 360.235 153.145 360.565 153.475 ;
        RECT 360.235 150.835 360.565 151.165 ;
        RECT 360.235 149.985 360.565 150.315 ;
        RECT 360.235 147.675 360.565 148.005 ;
        RECT 360.235 146.095 360.565 146.425 ;
        RECT 360.235 145.245 360.565 145.575 ;
        RECT 360.235 142.935 360.565 143.265 ;
        RECT 360.235 142.085 360.565 142.415 ;
        RECT 360.235 139.775 360.565 140.105 ;
        RECT 360.235 138.925 360.565 139.255 ;
        RECT 360.235 136.615 360.565 136.945 ;
        RECT 360.235 135.765 360.565 136.095 ;
        RECT 360.235 133.455 360.565 133.785 ;
        RECT 360.235 131.875 360.565 132.205 ;
        RECT 360.235 131.025 360.565 131.355 ;
        RECT 360.235 128.715 360.565 129.045 ;
        RECT 360.235 127.865 360.565 128.195 ;
        RECT 360.235 125.555 360.565 125.885 ;
        RECT 360.235 124.705 360.565 125.035 ;
        RECT 360.235 122.395 360.565 122.725 ;
        RECT 360.235 121.545 360.565 121.875 ;
        RECT 360.235 119.235 360.565 119.565 ;
        RECT 360.235 117.655 360.565 117.985 ;
        RECT 360.235 116.805 360.565 117.135 ;
        RECT 360.235 114.495 360.565 114.825 ;
        RECT 360.235 113.645 360.565 113.975 ;
        RECT 360.235 111.335 360.565 111.665 ;
        RECT 360.235 110.485 360.565 110.815 ;
        RECT 360.235 108.175 360.565 108.505 ;
        RECT 360.235 107.325 360.565 107.655 ;
        RECT 360.235 105.015 360.565 105.345 ;
        RECT 360.235 103.435 360.565 103.765 ;
        RECT 360.235 102.585 360.565 102.915 ;
        RECT 360.235 100.275 360.565 100.605 ;
        RECT 360.235 99.425 360.565 99.755 ;
        RECT 360.235 97.115 360.565 97.445 ;
        RECT 360.235 96.265 360.565 96.595 ;
        RECT 360.235 93.955 360.565 94.285 ;
        RECT 360.235 93.105 360.565 93.435 ;
        RECT 360.235 90.795 360.565 91.125 ;
        RECT 360.235 89.215 360.565 89.545 ;
        RECT 360.235 88.365 360.565 88.695 ;
        RECT 360.235 86.055 360.565 86.385 ;
        RECT 360.235 85.205 360.565 85.535 ;
        RECT 360.235 82.895 360.565 83.225 ;
        RECT 360.235 82.045 360.565 82.375 ;
        RECT 360.235 79.735 360.565 80.065 ;
        RECT 360.235 78.885 360.565 79.215 ;
        RECT 360.235 76.575 360.565 76.905 ;
        RECT 360.235 74.995 360.565 75.325 ;
        RECT 360.235 74.145 360.565 74.475 ;
        RECT 360.235 71.835 360.565 72.165 ;
        RECT 360.235 70.985 360.565 71.315 ;
        RECT 360.235 68.675 360.565 69.005 ;
        RECT 360.235 67.825 360.565 68.155 ;
        RECT 360.235 65.515 360.565 65.845 ;
        RECT 360.235 64.665 360.565 64.995 ;
        RECT 360.235 62.355 360.565 62.685 ;
        RECT 360.235 60.775 360.565 61.105 ;
        RECT 360.235 59.925 360.565 60.255 ;
        RECT 360.235 57.615 360.565 57.945 ;
        RECT 360.235 56.765 360.565 57.095 ;
        RECT 360.235 54.455 360.565 54.785 ;
        RECT 360.235 53.605 360.565 53.935 ;
        RECT 360.235 51.295 360.565 51.625 ;
        RECT 360.235 50.445 360.565 50.775 ;
        RECT 360.235 48.135 360.565 48.465 ;
        RECT 360.235 46.555 360.565 46.885 ;
        RECT 360.235 45.705 360.565 46.035 ;
        RECT 360.235 43.395 360.565 43.725 ;
        RECT 360.235 42.545 360.565 42.875 ;
        RECT 360.235 40.235 360.565 40.565 ;
        RECT 360.235 39.385 360.565 39.715 ;
        RECT 360.235 37.075 360.565 37.405 ;
        RECT 360.235 36.225 360.565 36.555 ;
        RECT 360.235 33.915 360.565 34.245 ;
        RECT 360.235 32.335 360.565 32.665 ;
        RECT 360.235 31.485 360.565 31.815 ;
        RECT 360.235 29.175 360.565 29.505 ;
        RECT 360.235 28.325 360.565 28.655 ;
        RECT 360.235 26.015 360.565 26.345 ;
        RECT 360.235 25.165 360.565 25.495 ;
        RECT 360.235 22.855 360.565 23.185 ;
        RECT 360.235 22.005 360.565 22.335 ;
        RECT 360.235 19.695 360.565 20.025 ;
        RECT 360.235 18.115 360.565 18.445 ;
        RECT 360.235 17.265 360.565 17.595 ;
        RECT 360.235 14.955 360.565 15.285 ;
        RECT 360.235 14.105 360.565 14.435 ;
        RECT 360.235 11.795 360.565 12.125 ;
        RECT 360.235 10.945 360.565 11.275 ;
        RECT 360.235 8.635 360.565 8.965 ;
        RECT 360.235 7.785 360.565 8.115 ;
        RECT 360.235 5.475 360.565 5.805 ;
        RECT 360.235 3.895 360.565 4.225 ;
        RECT 360.235 3.045 360.565 3.375 ;
        RECT 360.235 0.87 360.565 1.2 ;
        RECT 360.235 -0.845 360.565 -0.515 ;
        RECT 360.235 -2.205 360.565 -1.875 ;
        RECT 360.235 -3.565 360.565 -3.235 ;
        RECT 360.235 -4.925 360.565 -4.595 ;
        RECT 360.235 -6.285 360.565 -5.955 ;
        RECT 360.235 -7.645 360.565 -7.315 ;
        RECT 360.235 -9.005 360.565 -8.675 ;
        RECT 360.235 -10.365 360.565 -10.035 ;
        RECT 360.235 -11.725 360.565 -11.395 ;
        RECT 360.235 -13.085 360.565 -12.755 ;
        RECT 360.235 -14.445 360.565 -14.115 ;
        RECT 360.235 -15.805 360.565 -15.475 ;
        RECT 360.235 -17.165 360.565 -16.835 ;
        RECT 360.235 -18.525 360.565 -18.195 ;
        RECT 360.235 -19.885 360.565 -19.555 ;
        RECT 360.235 -21.245 360.565 -20.915 ;
        RECT 360.235 -22.605 360.565 -22.275 ;
        RECT 360.235 -23.965 360.565 -23.635 ;
        RECT 360.235 -25.325 360.565 -24.995 ;
        RECT 360.235 -26.685 360.565 -26.355 ;
        RECT 360.235 -28.045 360.565 -27.715 ;
        RECT 360.235 -29.405 360.565 -29.075 ;
        RECT 360.235 -30.765 360.565 -30.435 ;
        RECT 360.235 -32.125 360.565 -31.795 ;
        RECT 360.235 -33.485 360.565 -33.155 ;
        RECT 360.235 -34.845 360.565 -34.515 ;
        RECT 360.235 -36.205 360.565 -35.875 ;
        RECT 360.235 -37.565 360.565 -37.235 ;
        RECT 360.235 -38.925 360.565 -38.595 ;
        RECT 360.235 -40.285 360.565 -39.955 ;
        RECT 360.235 -41.645 360.565 -41.315 ;
        RECT 360.235 -43.005 360.565 -42.675 ;
        RECT 360.235 -44.365 360.565 -44.035 ;
        RECT 360.235 -45.725 360.565 -45.395 ;
        RECT 360.235 -47.085 360.565 -46.755 ;
        RECT 360.235 -48.445 360.565 -48.115 ;
        RECT 360.235 -49.805 360.565 -49.475 ;
        RECT 360.235 -51.165 360.565 -50.835 ;
        RECT 360.235 -52.525 360.565 -52.195 ;
        RECT 360.235 -53.885 360.565 -53.555 ;
        RECT 360.235 -55.245 360.565 -54.915 ;
        RECT 360.235 -56.605 360.565 -56.275 ;
        RECT 360.235 -57.965 360.565 -57.635 ;
        RECT 360.235 -59.325 360.565 -58.995 ;
        RECT 360.235 -60.685 360.565 -60.355 ;
        RECT 360.235 -62.045 360.565 -61.715 ;
        RECT 360.235 -63.405 360.565 -63.075 ;
        RECT 360.235 -64.765 360.565 -64.435 ;
        RECT 360.235 -66.125 360.565 -65.795 ;
        RECT 360.235 -67.485 360.565 -67.155 ;
        RECT 360.235 -68.845 360.565 -68.515 ;
        RECT 360.235 -70.205 360.565 -69.875 ;
        RECT 360.235 -71.565 360.565 -71.235 ;
        RECT 360.235 -72.925 360.565 -72.595 ;
        RECT 360.235 -74.285 360.565 -73.955 ;
        RECT 360.235 -75.645 360.565 -75.315 ;
        RECT 360.235 -77.005 360.565 -76.675 ;
        RECT 360.235 -78.365 360.565 -78.035 ;
        RECT 360.235 -79.725 360.565 -79.395 ;
        RECT 360.235 -81.085 360.565 -80.755 ;
        RECT 360.235 -82.445 360.565 -82.115 ;
        RECT 360.235 -83.805 360.565 -83.475 ;
        RECT 360.235 -85.165 360.565 -84.835 ;
        RECT 360.235 -86.525 360.565 -86.195 ;
        RECT 360.235 -87.885 360.565 -87.555 ;
        RECT 360.235 -89.245 360.565 -88.915 ;
        RECT 360.235 -90.605 360.565 -90.275 ;
        RECT 360.235 -91.965 360.565 -91.635 ;
        RECT 360.235 -93.325 360.565 -92.995 ;
        RECT 360.235 -94.685 360.565 -94.355 ;
        RECT 360.235 -96.045 360.565 -95.715 ;
        RECT 360.235 -97.405 360.565 -97.075 ;
        RECT 360.235 -98.765 360.565 -98.435 ;
        RECT 360.235 -100.125 360.565 -99.795 ;
        RECT 360.235 -101.485 360.565 -101.155 ;
        RECT 360.235 -102.845 360.565 -102.515 ;
        RECT 360.235 -104.205 360.565 -103.875 ;
        RECT 360.235 -105.565 360.565 -105.235 ;
        RECT 360.235 -106.925 360.565 -106.595 ;
        RECT 360.235 -108.285 360.565 -107.955 ;
        RECT 360.235 -109.645 360.565 -109.315 ;
        RECT 360.235 -111.005 360.565 -110.675 ;
        RECT 360.235 -112.365 360.565 -112.035 ;
        RECT 360.235 -113.725 360.565 -113.395 ;
        RECT 360.235 -115.085 360.565 -114.755 ;
        RECT 360.235 -116.445 360.565 -116.115 ;
        RECT 360.235 -117.805 360.565 -117.475 ;
        RECT 360.235 -119.165 360.565 -118.835 ;
        RECT 360.235 -120.525 360.565 -120.195 ;
        RECT 360.235 -121.885 360.565 -121.555 ;
        RECT 360.235 -123.245 360.565 -122.915 ;
        RECT 360.235 -124.605 360.565 -124.275 ;
        RECT 360.235 -125.965 360.565 -125.635 ;
        RECT 360.235 -127.325 360.565 -126.995 ;
        RECT 360.235 -128.685 360.565 -128.355 ;
        RECT 360.235 -130.045 360.565 -129.715 ;
        RECT 360.235 -131.405 360.565 -131.075 ;
        RECT 360.235 -132.765 360.565 -132.435 ;
        RECT 360.235 -134.125 360.565 -133.795 ;
        RECT 360.235 -135.485 360.565 -135.155 ;
        RECT 360.235 -136.845 360.565 -136.515 ;
        RECT 360.235 -138.205 360.565 -137.875 ;
        RECT 360.235 -139.565 360.565 -139.235 ;
        RECT 360.235 -140.925 360.565 -140.595 ;
        RECT 360.235 -142.285 360.565 -141.955 ;
        RECT 360.235 -143.645 360.565 -143.315 ;
        RECT 360.235 -145.005 360.565 -144.675 ;
        RECT 360.235 -146.365 360.565 -146.035 ;
        RECT 360.235 -147.725 360.565 -147.395 ;
        RECT 360.235 -149.085 360.565 -148.755 ;
        RECT 360.235 -150.445 360.565 -150.115 ;
        RECT 360.235 -151.805 360.565 -151.475 ;
        RECT 360.235 -153.165 360.565 -152.835 ;
        RECT 360.235 -154.525 360.565 -154.195 ;
        RECT 360.235 -155.885 360.565 -155.555 ;
        RECT 360.235 -157.245 360.565 -156.915 ;
        RECT 360.235 -158.605 360.565 -158.275 ;
        RECT 360.235 -159.965 360.565 -159.635 ;
        RECT 360.235 -161.325 360.565 -160.995 ;
        RECT 360.235 -162.685 360.565 -162.355 ;
        RECT 360.235 -164.045 360.565 -163.715 ;
        RECT 360.235 -165.405 360.565 -165.075 ;
        RECT 360.235 -166.765 360.565 -166.435 ;
        RECT 360.235 -168.125 360.565 -167.795 ;
        RECT 360.235 -169.485 360.565 -169.155 ;
        RECT 360.235 -170.845 360.565 -170.515 ;
        RECT 360.235 -172.205 360.565 -171.875 ;
        RECT 360.235 -173.565 360.565 -173.235 ;
        RECT 360.235 -174.925 360.565 -174.595 ;
        RECT 360.235 -176.285 360.565 -175.955 ;
        RECT 360.235 -177.645 360.565 -177.315 ;
        RECT 360.235 -179.005 360.565 -178.675 ;
        RECT 360.235 -184.65 360.565 -183.52 ;
        RECT 360.24 -184.765 360.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.475 244.04 338.805 245.17 ;
        RECT 338.475 239.875 338.805 240.205 ;
        RECT 338.475 238.515 338.805 238.845 ;
        RECT 338.475 237.155 338.805 237.485 ;
        RECT 338.48 237.155 338.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.475 -0.845 338.805 -0.515 ;
        RECT 338.475 -2.205 338.805 -1.875 ;
        RECT 338.475 -3.565 338.805 -3.235 ;
        RECT 338.48 -3.565 338.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 338.475 -96.045 338.805 -95.715 ;
        RECT 338.475 -97.405 338.805 -97.075 ;
        RECT 338.475 -98.765 338.805 -98.435 ;
        RECT 338.475 -100.125 338.805 -99.795 ;
        RECT 338.475 -101.485 338.805 -101.155 ;
        RECT 338.475 -102.845 338.805 -102.515 ;
        RECT 338.475 -104.205 338.805 -103.875 ;
        RECT 338.475 -105.565 338.805 -105.235 ;
        RECT 338.475 -106.925 338.805 -106.595 ;
        RECT 338.475 -108.285 338.805 -107.955 ;
        RECT 338.475 -109.645 338.805 -109.315 ;
        RECT 338.475 -111.005 338.805 -110.675 ;
        RECT 338.475 -112.365 338.805 -112.035 ;
        RECT 338.475 -113.725 338.805 -113.395 ;
        RECT 338.475 -115.085 338.805 -114.755 ;
        RECT 338.475 -116.445 338.805 -116.115 ;
        RECT 338.475 -117.805 338.805 -117.475 ;
        RECT 338.475 -119.165 338.805 -118.835 ;
        RECT 338.475 -120.525 338.805 -120.195 ;
        RECT 338.475 -121.885 338.805 -121.555 ;
        RECT 338.475 -123.245 338.805 -122.915 ;
        RECT 338.475 -124.605 338.805 -124.275 ;
        RECT 338.475 -125.965 338.805 -125.635 ;
        RECT 338.475 -127.325 338.805 -126.995 ;
        RECT 338.475 -128.685 338.805 -128.355 ;
        RECT 338.475 -130.045 338.805 -129.715 ;
        RECT 338.475 -131.405 338.805 -131.075 ;
        RECT 338.475 -132.765 338.805 -132.435 ;
        RECT 338.475 -134.125 338.805 -133.795 ;
        RECT 338.475 -135.485 338.805 -135.155 ;
        RECT 338.475 -136.845 338.805 -136.515 ;
        RECT 338.475 -138.205 338.805 -137.875 ;
        RECT 338.475 -139.565 338.805 -139.235 ;
        RECT 338.475 -140.925 338.805 -140.595 ;
        RECT 338.475 -142.285 338.805 -141.955 ;
        RECT 338.475 -143.645 338.805 -143.315 ;
        RECT 338.475 -145.005 338.805 -144.675 ;
        RECT 338.475 -146.365 338.805 -146.035 ;
        RECT 338.475 -147.725 338.805 -147.395 ;
        RECT 338.475 -149.085 338.805 -148.755 ;
        RECT 338.475 -150.445 338.805 -150.115 ;
        RECT 338.475 -151.805 338.805 -151.475 ;
        RECT 338.475 -153.165 338.805 -152.835 ;
        RECT 338.475 -154.525 338.805 -154.195 ;
        RECT 338.475 -155.885 338.805 -155.555 ;
        RECT 338.475 -157.245 338.805 -156.915 ;
        RECT 338.475 -158.605 338.805 -158.275 ;
        RECT 338.475 -159.965 338.805 -159.635 ;
        RECT 338.475 -161.325 338.805 -160.995 ;
        RECT 338.475 -162.685 338.805 -162.355 ;
        RECT 338.475 -164.045 338.805 -163.715 ;
        RECT 338.475 -165.405 338.805 -165.075 ;
        RECT 338.475 -166.765 338.805 -166.435 ;
        RECT 338.475 -168.125 338.805 -167.795 ;
        RECT 338.475 -169.485 338.805 -169.155 ;
        RECT 338.475 -170.845 338.805 -170.515 ;
        RECT 338.475 -172.205 338.805 -171.875 ;
        RECT 338.475 -173.565 338.805 -173.235 ;
        RECT 338.475 -174.925 338.805 -174.595 ;
        RECT 338.475 -176.285 338.805 -175.955 ;
        RECT 338.475 -177.645 338.805 -177.315 ;
        RECT 338.475 -179.005 338.805 -178.675 ;
        RECT 338.475 -184.65 338.805 -183.52 ;
        RECT 338.48 -184.765 338.8 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.835 244.04 340.165 245.17 ;
        RECT 339.835 239.875 340.165 240.205 ;
        RECT 339.835 238.515 340.165 238.845 ;
        RECT 339.835 237.155 340.165 237.485 ;
        RECT 339.84 237.155 340.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.835 -0.845 340.165 -0.515 ;
        RECT 339.835 -2.205 340.165 -1.875 ;
        RECT 339.835 -3.565 340.165 -3.235 ;
        RECT 339.84 -3.565 340.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.835 -96.045 340.165 -95.715 ;
        RECT 339.835 -97.405 340.165 -97.075 ;
        RECT 339.835 -98.765 340.165 -98.435 ;
        RECT 339.835 -100.125 340.165 -99.795 ;
        RECT 339.835 -101.485 340.165 -101.155 ;
        RECT 339.835 -102.845 340.165 -102.515 ;
        RECT 339.835 -104.205 340.165 -103.875 ;
        RECT 339.835 -105.565 340.165 -105.235 ;
        RECT 339.835 -106.925 340.165 -106.595 ;
        RECT 339.835 -108.285 340.165 -107.955 ;
        RECT 339.835 -109.645 340.165 -109.315 ;
        RECT 339.835 -111.005 340.165 -110.675 ;
        RECT 339.835 -112.365 340.165 -112.035 ;
        RECT 339.835 -113.725 340.165 -113.395 ;
        RECT 339.835 -115.085 340.165 -114.755 ;
        RECT 339.835 -116.445 340.165 -116.115 ;
        RECT 339.835 -117.805 340.165 -117.475 ;
        RECT 339.835 -119.165 340.165 -118.835 ;
        RECT 339.835 -120.525 340.165 -120.195 ;
        RECT 339.835 -121.885 340.165 -121.555 ;
        RECT 339.835 -123.245 340.165 -122.915 ;
        RECT 339.835 -124.605 340.165 -124.275 ;
        RECT 339.835 -125.965 340.165 -125.635 ;
        RECT 339.835 -127.325 340.165 -126.995 ;
        RECT 339.835 -128.685 340.165 -128.355 ;
        RECT 339.835 -130.045 340.165 -129.715 ;
        RECT 339.835 -131.405 340.165 -131.075 ;
        RECT 339.835 -132.765 340.165 -132.435 ;
        RECT 339.835 -134.125 340.165 -133.795 ;
        RECT 339.835 -135.485 340.165 -135.155 ;
        RECT 339.835 -136.845 340.165 -136.515 ;
        RECT 339.835 -138.205 340.165 -137.875 ;
        RECT 339.835 -139.565 340.165 -139.235 ;
        RECT 339.835 -140.925 340.165 -140.595 ;
        RECT 339.835 -142.285 340.165 -141.955 ;
        RECT 339.835 -143.645 340.165 -143.315 ;
        RECT 339.835 -145.005 340.165 -144.675 ;
        RECT 339.835 -146.365 340.165 -146.035 ;
        RECT 339.835 -147.725 340.165 -147.395 ;
        RECT 339.835 -149.085 340.165 -148.755 ;
        RECT 339.835 -150.445 340.165 -150.115 ;
        RECT 339.835 -151.805 340.165 -151.475 ;
        RECT 339.835 -153.165 340.165 -152.835 ;
        RECT 339.835 -154.525 340.165 -154.195 ;
        RECT 339.835 -155.885 340.165 -155.555 ;
        RECT 339.835 -157.245 340.165 -156.915 ;
        RECT 339.835 -158.605 340.165 -158.275 ;
        RECT 339.835 -159.965 340.165 -159.635 ;
        RECT 339.835 -161.325 340.165 -160.995 ;
        RECT 339.835 -162.685 340.165 -162.355 ;
        RECT 339.835 -164.045 340.165 -163.715 ;
        RECT 339.835 -165.405 340.165 -165.075 ;
        RECT 339.835 -166.765 340.165 -166.435 ;
        RECT 339.835 -168.125 340.165 -167.795 ;
        RECT 339.835 -169.485 340.165 -169.155 ;
        RECT 339.835 -170.845 340.165 -170.515 ;
        RECT 339.835 -172.205 340.165 -171.875 ;
        RECT 339.835 -173.565 340.165 -173.235 ;
        RECT 339.835 -174.925 340.165 -174.595 ;
        RECT 339.835 -176.285 340.165 -175.955 ;
        RECT 339.835 -177.645 340.165 -177.315 ;
        RECT 339.835 -179.005 340.165 -178.675 ;
        RECT 339.835 -184.65 340.165 -183.52 ;
        RECT 339.84 -184.765 340.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.56 -98.075 340.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.195 244.04 341.525 245.17 ;
        RECT 341.195 239.875 341.525 240.205 ;
        RECT 341.195 238.515 341.525 238.845 ;
        RECT 341.195 237.155 341.525 237.485 ;
        RECT 341.2 237.155 341.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.195 -98.765 341.525 -98.435 ;
        RECT 341.195 -100.125 341.525 -99.795 ;
        RECT 341.195 -101.485 341.525 -101.155 ;
        RECT 341.195 -102.845 341.525 -102.515 ;
        RECT 341.195 -104.205 341.525 -103.875 ;
        RECT 341.195 -105.565 341.525 -105.235 ;
        RECT 341.195 -106.925 341.525 -106.595 ;
        RECT 341.195 -108.285 341.525 -107.955 ;
        RECT 341.195 -109.645 341.525 -109.315 ;
        RECT 341.195 -111.005 341.525 -110.675 ;
        RECT 341.195 -112.365 341.525 -112.035 ;
        RECT 341.195 -113.725 341.525 -113.395 ;
        RECT 341.195 -115.085 341.525 -114.755 ;
        RECT 341.195 -116.445 341.525 -116.115 ;
        RECT 341.195 -117.805 341.525 -117.475 ;
        RECT 341.195 -119.165 341.525 -118.835 ;
        RECT 341.195 -120.525 341.525 -120.195 ;
        RECT 341.195 -121.885 341.525 -121.555 ;
        RECT 341.195 -123.245 341.525 -122.915 ;
        RECT 341.195 -124.605 341.525 -124.275 ;
        RECT 341.195 -125.965 341.525 -125.635 ;
        RECT 341.195 -127.325 341.525 -126.995 ;
        RECT 341.195 -128.685 341.525 -128.355 ;
        RECT 341.195 -130.045 341.525 -129.715 ;
        RECT 341.195 -131.405 341.525 -131.075 ;
        RECT 341.195 -132.765 341.525 -132.435 ;
        RECT 341.195 -134.125 341.525 -133.795 ;
        RECT 341.195 -135.485 341.525 -135.155 ;
        RECT 341.195 -136.845 341.525 -136.515 ;
        RECT 341.195 -138.205 341.525 -137.875 ;
        RECT 341.195 -139.565 341.525 -139.235 ;
        RECT 341.195 -140.925 341.525 -140.595 ;
        RECT 341.195 -142.285 341.525 -141.955 ;
        RECT 341.195 -143.645 341.525 -143.315 ;
        RECT 341.195 -145.005 341.525 -144.675 ;
        RECT 341.195 -146.365 341.525 -146.035 ;
        RECT 341.195 -147.725 341.525 -147.395 ;
        RECT 341.195 -149.085 341.525 -148.755 ;
        RECT 341.195 -150.445 341.525 -150.115 ;
        RECT 341.195 -151.805 341.525 -151.475 ;
        RECT 341.195 -153.165 341.525 -152.835 ;
        RECT 341.195 -154.525 341.525 -154.195 ;
        RECT 341.195 -155.885 341.525 -155.555 ;
        RECT 341.195 -157.245 341.525 -156.915 ;
        RECT 341.195 -158.605 341.525 -158.275 ;
        RECT 341.195 -159.965 341.525 -159.635 ;
        RECT 341.195 -161.325 341.525 -160.995 ;
        RECT 341.195 -162.685 341.525 -162.355 ;
        RECT 341.195 -164.045 341.525 -163.715 ;
        RECT 341.195 -165.405 341.525 -165.075 ;
        RECT 341.195 -166.765 341.525 -166.435 ;
        RECT 341.195 -168.125 341.525 -167.795 ;
        RECT 341.195 -169.485 341.525 -169.155 ;
        RECT 341.195 -170.845 341.525 -170.515 ;
        RECT 341.195 -172.205 341.525 -171.875 ;
        RECT 341.195 -173.565 341.525 -173.235 ;
        RECT 341.195 -174.925 341.525 -174.595 ;
        RECT 341.195 -176.285 341.525 -175.955 ;
        RECT 341.195 -177.645 341.525 -177.315 ;
        RECT 341.195 -179.005 341.525 -178.675 ;
        RECT 341.195 -184.65 341.525 -183.52 ;
        RECT 341.2 -184.765 341.52 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.555 244.04 342.885 245.17 ;
        RECT 342.555 239.875 342.885 240.205 ;
        RECT 342.555 238.515 342.885 238.845 ;
        RECT 342.555 237.155 342.885 237.485 ;
        RECT 342.56 237.155 342.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 342.555 -0.845 342.885 -0.515 ;
        RECT 342.555 -2.205 342.885 -1.875 ;
        RECT 342.555 -3.565 342.885 -3.235 ;
        RECT 342.56 -3.565 342.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.915 244.04 344.245 245.17 ;
        RECT 343.915 239.875 344.245 240.205 ;
        RECT 343.915 238.515 344.245 238.845 ;
        RECT 343.915 237.155 344.245 237.485 ;
        RECT 343.92 237.155 344.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.915 -0.845 344.245 -0.515 ;
        RECT 343.915 -2.205 344.245 -1.875 ;
        RECT 343.915 -3.565 344.245 -3.235 ;
        RECT 343.92 -3.565 344.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.275 244.04 345.605 245.17 ;
        RECT 345.275 239.875 345.605 240.205 ;
        RECT 345.275 238.515 345.605 238.845 ;
        RECT 345.275 237.155 345.605 237.485 ;
        RECT 345.28 237.155 345.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.275 -0.845 345.605 -0.515 ;
        RECT 345.275 -2.205 345.605 -1.875 ;
        RECT 345.275 -3.565 345.605 -3.235 ;
        RECT 345.28 -3.565 345.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.275 -96.045 345.605 -95.715 ;
        RECT 345.275 -97.405 345.605 -97.075 ;
        RECT 345.275 -98.765 345.605 -98.435 ;
        RECT 345.275 -100.125 345.605 -99.795 ;
        RECT 345.275 -101.485 345.605 -101.155 ;
        RECT 345.275 -102.845 345.605 -102.515 ;
        RECT 345.275 -104.205 345.605 -103.875 ;
        RECT 345.275 -105.565 345.605 -105.235 ;
        RECT 345.275 -106.925 345.605 -106.595 ;
        RECT 345.275 -108.285 345.605 -107.955 ;
        RECT 345.275 -109.645 345.605 -109.315 ;
        RECT 345.275 -111.005 345.605 -110.675 ;
        RECT 345.275 -112.365 345.605 -112.035 ;
        RECT 345.275 -113.725 345.605 -113.395 ;
        RECT 345.275 -115.085 345.605 -114.755 ;
        RECT 345.275 -116.445 345.605 -116.115 ;
        RECT 345.275 -117.805 345.605 -117.475 ;
        RECT 345.275 -119.165 345.605 -118.835 ;
        RECT 345.275 -120.525 345.605 -120.195 ;
        RECT 345.275 -121.885 345.605 -121.555 ;
        RECT 345.275 -123.245 345.605 -122.915 ;
        RECT 345.275 -124.605 345.605 -124.275 ;
        RECT 345.275 -125.965 345.605 -125.635 ;
        RECT 345.275 -127.325 345.605 -126.995 ;
        RECT 345.275 -128.685 345.605 -128.355 ;
        RECT 345.275 -130.045 345.605 -129.715 ;
        RECT 345.275 -131.405 345.605 -131.075 ;
        RECT 345.275 -132.765 345.605 -132.435 ;
        RECT 345.275 -134.125 345.605 -133.795 ;
        RECT 345.275 -135.485 345.605 -135.155 ;
        RECT 345.275 -136.845 345.605 -136.515 ;
        RECT 345.275 -138.205 345.605 -137.875 ;
        RECT 345.275 -139.565 345.605 -139.235 ;
        RECT 345.275 -140.925 345.605 -140.595 ;
        RECT 345.275 -142.285 345.605 -141.955 ;
        RECT 345.275 -143.645 345.605 -143.315 ;
        RECT 345.275 -145.005 345.605 -144.675 ;
        RECT 345.275 -146.365 345.605 -146.035 ;
        RECT 345.275 -147.725 345.605 -147.395 ;
        RECT 345.275 -149.085 345.605 -148.755 ;
        RECT 345.275 -150.445 345.605 -150.115 ;
        RECT 345.275 -151.805 345.605 -151.475 ;
        RECT 345.275 -153.165 345.605 -152.835 ;
        RECT 345.275 -154.525 345.605 -154.195 ;
        RECT 345.275 -155.885 345.605 -155.555 ;
        RECT 345.275 -157.245 345.605 -156.915 ;
        RECT 345.275 -158.605 345.605 -158.275 ;
        RECT 345.275 -159.965 345.605 -159.635 ;
        RECT 345.275 -161.325 345.605 -160.995 ;
        RECT 345.275 -162.685 345.605 -162.355 ;
        RECT 345.275 -164.045 345.605 -163.715 ;
        RECT 345.275 -165.405 345.605 -165.075 ;
        RECT 345.275 -166.765 345.605 -166.435 ;
        RECT 345.275 -168.125 345.605 -167.795 ;
        RECT 345.275 -169.485 345.605 -169.155 ;
        RECT 345.275 -170.845 345.605 -170.515 ;
        RECT 345.275 -172.205 345.605 -171.875 ;
        RECT 345.275 -173.565 345.605 -173.235 ;
        RECT 345.275 -174.925 345.605 -174.595 ;
        RECT 345.275 -176.285 345.605 -175.955 ;
        RECT 345.275 -177.645 345.605 -177.315 ;
        RECT 345.275 -179.005 345.605 -178.675 ;
        RECT 345.275 -184.65 345.605 -183.52 ;
        RECT 345.28 -184.765 345.6 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.635 244.04 346.965 245.17 ;
        RECT 346.635 239.875 346.965 240.205 ;
        RECT 346.635 238.515 346.965 238.845 ;
        RECT 346.635 237.155 346.965 237.485 ;
        RECT 346.64 237.155 346.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.635 -0.845 346.965 -0.515 ;
        RECT 346.635 -2.205 346.965 -1.875 ;
        RECT 346.635 -3.565 346.965 -3.235 ;
        RECT 346.64 -3.565 346.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 346.635 -96.045 346.965 -95.715 ;
        RECT 346.635 -97.405 346.965 -97.075 ;
        RECT 346.635 -98.765 346.965 -98.435 ;
        RECT 346.635 -100.125 346.965 -99.795 ;
        RECT 346.635 -101.485 346.965 -101.155 ;
        RECT 346.635 -102.845 346.965 -102.515 ;
        RECT 346.635 -104.205 346.965 -103.875 ;
        RECT 346.635 -105.565 346.965 -105.235 ;
        RECT 346.635 -106.925 346.965 -106.595 ;
        RECT 346.635 -108.285 346.965 -107.955 ;
        RECT 346.635 -109.645 346.965 -109.315 ;
        RECT 346.635 -111.005 346.965 -110.675 ;
        RECT 346.635 -112.365 346.965 -112.035 ;
        RECT 346.635 -113.725 346.965 -113.395 ;
        RECT 346.635 -115.085 346.965 -114.755 ;
        RECT 346.635 -116.445 346.965 -116.115 ;
        RECT 346.635 -117.805 346.965 -117.475 ;
        RECT 346.635 -119.165 346.965 -118.835 ;
        RECT 346.635 -120.525 346.965 -120.195 ;
        RECT 346.635 -121.885 346.965 -121.555 ;
        RECT 346.635 -123.245 346.965 -122.915 ;
        RECT 346.635 -124.605 346.965 -124.275 ;
        RECT 346.635 -125.965 346.965 -125.635 ;
        RECT 346.635 -127.325 346.965 -126.995 ;
        RECT 346.635 -128.685 346.965 -128.355 ;
        RECT 346.635 -130.045 346.965 -129.715 ;
        RECT 346.635 -131.405 346.965 -131.075 ;
        RECT 346.635 -132.765 346.965 -132.435 ;
        RECT 346.635 -134.125 346.965 -133.795 ;
        RECT 346.635 -135.485 346.965 -135.155 ;
        RECT 346.635 -136.845 346.965 -136.515 ;
        RECT 346.635 -138.205 346.965 -137.875 ;
        RECT 346.635 -139.565 346.965 -139.235 ;
        RECT 346.635 -140.925 346.965 -140.595 ;
        RECT 346.635 -142.285 346.965 -141.955 ;
        RECT 346.635 -143.645 346.965 -143.315 ;
        RECT 346.635 -145.005 346.965 -144.675 ;
        RECT 346.635 -146.365 346.965 -146.035 ;
        RECT 346.635 -147.725 346.965 -147.395 ;
        RECT 346.635 -149.085 346.965 -148.755 ;
        RECT 346.635 -150.445 346.965 -150.115 ;
        RECT 346.635 -151.805 346.965 -151.475 ;
        RECT 346.635 -153.165 346.965 -152.835 ;
        RECT 346.635 -154.525 346.965 -154.195 ;
        RECT 346.635 -155.885 346.965 -155.555 ;
        RECT 346.635 -157.245 346.965 -156.915 ;
        RECT 346.635 -158.605 346.965 -158.275 ;
        RECT 346.635 -159.965 346.965 -159.635 ;
        RECT 346.635 -161.325 346.965 -160.995 ;
        RECT 346.635 -162.685 346.965 -162.355 ;
        RECT 346.635 -164.045 346.965 -163.715 ;
        RECT 346.635 -165.405 346.965 -165.075 ;
        RECT 346.635 -166.765 346.965 -166.435 ;
        RECT 346.635 -168.125 346.965 -167.795 ;
        RECT 346.635 -169.485 346.965 -169.155 ;
        RECT 346.635 -170.845 346.965 -170.515 ;
        RECT 346.635 -172.205 346.965 -171.875 ;
        RECT 346.635 -173.565 346.965 -173.235 ;
        RECT 346.635 -174.925 346.965 -174.595 ;
        RECT 346.635 -176.285 346.965 -175.955 ;
        RECT 346.635 -177.645 346.965 -177.315 ;
        RECT 346.635 -179.005 346.965 -178.675 ;
        RECT 346.635 -184.65 346.965 -183.52 ;
        RECT 346.64 -184.765 346.96 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.995 244.04 348.325 245.17 ;
        RECT 347.995 239.875 348.325 240.205 ;
        RECT 347.995 238.515 348.325 238.845 ;
        RECT 347.995 237.155 348.325 237.485 ;
        RECT 348 237.155 348.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.995 -0.845 348.325 -0.515 ;
        RECT 347.995 -2.205 348.325 -1.875 ;
        RECT 347.995 -3.565 348.325 -3.235 ;
        RECT 348 -3.565 348.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.995 -96.045 348.325 -95.715 ;
        RECT 347.995 -97.405 348.325 -97.075 ;
        RECT 347.995 -98.765 348.325 -98.435 ;
        RECT 347.995 -100.125 348.325 -99.795 ;
        RECT 347.995 -101.485 348.325 -101.155 ;
        RECT 347.995 -102.845 348.325 -102.515 ;
        RECT 347.995 -104.205 348.325 -103.875 ;
        RECT 347.995 -105.565 348.325 -105.235 ;
        RECT 347.995 -106.925 348.325 -106.595 ;
        RECT 347.995 -108.285 348.325 -107.955 ;
        RECT 347.995 -109.645 348.325 -109.315 ;
        RECT 347.995 -111.005 348.325 -110.675 ;
        RECT 347.995 -112.365 348.325 -112.035 ;
        RECT 347.995 -113.725 348.325 -113.395 ;
        RECT 347.995 -115.085 348.325 -114.755 ;
        RECT 347.995 -116.445 348.325 -116.115 ;
        RECT 347.995 -117.805 348.325 -117.475 ;
        RECT 347.995 -119.165 348.325 -118.835 ;
        RECT 347.995 -120.525 348.325 -120.195 ;
        RECT 347.995 -121.885 348.325 -121.555 ;
        RECT 347.995 -123.245 348.325 -122.915 ;
        RECT 347.995 -124.605 348.325 -124.275 ;
        RECT 347.995 -125.965 348.325 -125.635 ;
        RECT 347.995 -127.325 348.325 -126.995 ;
        RECT 347.995 -128.685 348.325 -128.355 ;
        RECT 347.995 -130.045 348.325 -129.715 ;
        RECT 347.995 -131.405 348.325 -131.075 ;
        RECT 347.995 -132.765 348.325 -132.435 ;
        RECT 347.995 -134.125 348.325 -133.795 ;
        RECT 347.995 -135.485 348.325 -135.155 ;
        RECT 347.995 -136.845 348.325 -136.515 ;
        RECT 347.995 -138.205 348.325 -137.875 ;
        RECT 347.995 -139.565 348.325 -139.235 ;
        RECT 347.995 -140.925 348.325 -140.595 ;
        RECT 347.995 -142.285 348.325 -141.955 ;
        RECT 347.995 -143.645 348.325 -143.315 ;
        RECT 347.995 -145.005 348.325 -144.675 ;
        RECT 347.995 -146.365 348.325 -146.035 ;
        RECT 347.995 -147.725 348.325 -147.395 ;
        RECT 347.995 -149.085 348.325 -148.755 ;
        RECT 347.995 -150.445 348.325 -150.115 ;
        RECT 347.995 -151.805 348.325 -151.475 ;
        RECT 347.995 -153.165 348.325 -152.835 ;
        RECT 347.995 -154.525 348.325 -154.195 ;
        RECT 347.995 -155.885 348.325 -155.555 ;
        RECT 347.995 -157.245 348.325 -156.915 ;
        RECT 347.995 -158.605 348.325 -158.275 ;
        RECT 347.995 -159.965 348.325 -159.635 ;
        RECT 347.995 -161.325 348.325 -160.995 ;
        RECT 347.995 -162.685 348.325 -162.355 ;
        RECT 347.995 -164.045 348.325 -163.715 ;
        RECT 347.995 -165.405 348.325 -165.075 ;
        RECT 347.995 -166.765 348.325 -166.435 ;
        RECT 347.995 -168.125 348.325 -167.795 ;
        RECT 347.995 -169.485 348.325 -169.155 ;
        RECT 347.995 -170.845 348.325 -170.515 ;
        RECT 347.995 -172.205 348.325 -171.875 ;
        RECT 347.995 -173.565 348.325 -173.235 ;
        RECT 347.995 -174.925 348.325 -174.595 ;
        RECT 347.995 -176.285 348.325 -175.955 ;
        RECT 347.995 -177.645 348.325 -177.315 ;
        RECT 347.995 -179.005 348.325 -178.675 ;
        RECT 347.995 -184.65 348.325 -183.52 ;
        RECT 348 -184.765 348.32 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.355 244.04 349.685 245.17 ;
        RECT 349.355 239.875 349.685 240.205 ;
        RECT 349.355 238.515 349.685 238.845 ;
        RECT 349.355 237.155 349.685 237.485 ;
        RECT 349.36 237.155 349.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.355 -0.845 349.685 -0.515 ;
        RECT 349.355 -2.205 349.685 -1.875 ;
        RECT 349.355 -3.565 349.685 -3.235 ;
        RECT 349.36 -3.565 349.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 349.355 -96.045 349.685 -95.715 ;
        RECT 349.355 -97.405 349.685 -97.075 ;
        RECT 349.355 -98.765 349.685 -98.435 ;
        RECT 349.355 -100.125 349.685 -99.795 ;
        RECT 349.355 -101.485 349.685 -101.155 ;
        RECT 349.355 -102.845 349.685 -102.515 ;
        RECT 349.355 -104.205 349.685 -103.875 ;
        RECT 349.355 -105.565 349.685 -105.235 ;
        RECT 349.355 -106.925 349.685 -106.595 ;
        RECT 349.355 -108.285 349.685 -107.955 ;
        RECT 349.355 -109.645 349.685 -109.315 ;
        RECT 349.355 -111.005 349.685 -110.675 ;
        RECT 349.355 -112.365 349.685 -112.035 ;
        RECT 349.355 -113.725 349.685 -113.395 ;
        RECT 349.355 -115.085 349.685 -114.755 ;
        RECT 349.355 -116.445 349.685 -116.115 ;
        RECT 349.355 -117.805 349.685 -117.475 ;
        RECT 349.355 -119.165 349.685 -118.835 ;
        RECT 349.355 -120.525 349.685 -120.195 ;
        RECT 349.355 -121.885 349.685 -121.555 ;
        RECT 349.355 -123.245 349.685 -122.915 ;
        RECT 349.355 -124.605 349.685 -124.275 ;
        RECT 349.355 -125.965 349.685 -125.635 ;
        RECT 349.355 -127.325 349.685 -126.995 ;
        RECT 349.355 -128.685 349.685 -128.355 ;
        RECT 349.355 -130.045 349.685 -129.715 ;
        RECT 349.355 -131.405 349.685 -131.075 ;
        RECT 349.355 -132.765 349.685 -132.435 ;
        RECT 349.355 -134.125 349.685 -133.795 ;
        RECT 349.355 -135.485 349.685 -135.155 ;
        RECT 349.355 -136.845 349.685 -136.515 ;
        RECT 349.355 -138.205 349.685 -137.875 ;
        RECT 349.355 -139.565 349.685 -139.235 ;
        RECT 349.355 -140.925 349.685 -140.595 ;
        RECT 349.355 -142.285 349.685 -141.955 ;
        RECT 349.355 -143.645 349.685 -143.315 ;
        RECT 349.355 -145.005 349.685 -144.675 ;
        RECT 349.355 -146.365 349.685 -146.035 ;
        RECT 349.355 -147.725 349.685 -147.395 ;
        RECT 349.355 -149.085 349.685 -148.755 ;
        RECT 349.355 -150.445 349.685 -150.115 ;
        RECT 349.355 -151.805 349.685 -151.475 ;
        RECT 349.355 -153.165 349.685 -152.835 ;
        RECT 349.355 -154.525 349.685 -154.195 ;
        RECT 349.355 -155.885 349.685 -155.555 ;
        RECT 349.355 -157.245 349.685 -156.915 ;
        RECT 349.355 -158.605 349.685 -158.275 ;
        RECT 349.355 -159.965 349.685 -159.635 ;
        RECT 349.355 -161.325 349.685 -160.995 ;
        RECT 349.355 -162.685 349.685 -162.355 ;
        RECT 349.355 -164.045 349.685 -163.715 ;
        RECT 349.355 -165.405 349.685 -165.075 ;
        RECT 349.355 -166.765 349.685 -166.435 ;
        RECT 349.355 -168.125 349.685 -167.795 ;
        RECT 349.355 -169.485 349.685 -169.155 ;
        RECT 349.355 -170.845 349.685 -170.515 ;
        RECT 349.355 -172.205 349.685 -171.875 ;
        RECT 349.355 -173.565 349.685 -173.235 ;
        RECT 349.355 -174.925 349.685 -174.595 ;
        RECT 349.355 -176.285 349.685 -175.955 ;
        RECT 349.355 -177.645 349.685 -177.315 ;
        RECT 349.355 -179.005 349.685 -178.675 ;
        RECT 349.355 -184.65 349.685 -183.52 ;
        RECT 349.36 -184.765 349.68 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.715 244.04 351.045 245.17 ;
        RECT 350.715 239.875 351.045 240.205 ;
        RECT 350.715 238.515 351.045 238.845 ;
        RECT 350.715 237.155 351.045 237.485 ;
        RECT 350.72 237.155 351.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.715 -0.845 351.045 -0.515 ;
        RECT 350.715 -2.205 351.045 -1.875 ;
        RECT 350.715 -3.565 351.045 -3.235 ;
        RECT 350.72 -3.565 351.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.715 -96.045 351.045 -95.715 ;
        RECT 350.715 -97.405 351.045 -97.075 ;
        RECT 350.715 -98.765 351.045 -98.435 ;
        RECT 350.715 -100.125 351.045 -99.795 ;
        RECT 350.715 -101.485 351.045 -101.155 ;
        RECT 350.715 -102.845 351.045 -102.515 ;
        RECT 350.715 -104.205 351.045 -103.875 ;
        RECT 350.715 -105.565 351.045 -105.235 ;
        RECT 350.715 -106.925 351.045 -106.595 ;
        RECT 350.715 -108.285 351.045 -107.955 ;
        RECT 350.715 -109.645 351.045 -109.315 ;
        RECT 350.715 -111.005 351.045 -110.675 ;
        RECT 350.715 -112.365 351.045 -112.035 ;
        RECT 350.715 -113.725 351.045 -113.395 ;
        RECT 350.715 -115.085 351.045 -114.755 ;
        RECT 350.715 -116.445 351.045 -116.115 ;
        RECT 350.715 -117.805 351.045 -117.475 ;
        RECT 350.715 -119.165 351.045 -118.835 ;
        RECT 350.715 -120.525 351.045 -120.195 ;
        RECT 350.715 -121.885 351.045 -121.555 ;
        RECT 350.715 -123.245 351.045 -122.915 ;
        RECT 350.715 -124.605 351.045 -124.275 ;
        RECT 350.715 -125.965 351.045 -125.635 ;
        RECT 350.715 -127.325 351.045 -126.995 ;
        RECT 350.715 -128.685 351.045 -128.355 ;
        RECT 350.715 -130.045 351.045 -129.715 ;
        RECT 350.715 -131.405 351.045 -131.075 ;
        RECT 350.715 -132.765 351.045 -132.435 ;
        RECT 350.715 -134.125 351.045 -133.795 ;
        RECT 350.715 -135.485 351.045 -135.155 ;
        RECT 350.715 -136.845 351.045 -136.515 ;
        RECT 350.715 -138.205 351.045 -137.875 ;
        RECT 350.715 -139.565 351.045 -139.235 ;
        RECT 350.715 -140.925 351.045 -140.595 ;
        RECT 350.715 -142.285 351.045 -141.955 ;
        RECT 350.715 -143.645 351.045 -143.315 ;
        RECT 350.715 -145.005 351.045 -144.675 ;
        RECT 350.715 -146.365 351.045 -146.035 ;
        RECT 350.715 -147.725 351.045 -147.395 ;
        RECT 350.715 -149.085 351.045 -148.755 ;
        RECT 350.715 -150.445 351.045 -150.115 ;
        RECT 350.715 -151.805 351.045 -151.475 ;
        RECT 350.715 -153.165 351.045 -152.835 ;
        RECT 350.715 -154.525 351.045 -154.195 ;
        RECT 350.715 -155.885 351.045 -155.555 ;
        RECT 350.715 -157.245 351.045 -156.915 ;
        RECT 350.715 -158.605 351.045 -158.275 ;
        RECT 350.715 -159.965 351.045 -159.635 ;
        RECT 350.715 -161.325 351.045 -160.995 ;
        RECT 350.715 -162.685 351.045 -162.355 ;
        RECT 350.715 -164.045 351.045 -163.715 ;
        RECT 350.715 -165.405 351.045 -165.075 ;
        RECT 350.715 -166.765 351.045 -166.435 ;
        RECT 350.715 -168.125 351.045 -167.795 ;
        RECT 350.715 -169.485 351.045 -169.155 ;
        RECT 350.715 -170.845 351.045 -170.515 ;
        RECT 350.715 -172.205 351.045 -171.875 ;
        RECT 350.715 -173.565 351.045 -173.235 ;
        RECT 350.715 -174.925 351.045 -174.595 ;
        RECT 350.715 -176.285 351.045 -175.955 ;
        RECT 350.715 -177.645 351.045 -177.315 ;
        RECT 350.715 -179.005 351.045 -178.675 ;
        RECT 350.715 -184.65 351.045 -183.52 ;
        RECT 350.72 -184.765 351.04 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.075 244.04 352.405 245.17 ;
        RECT 352.075 239.875 352.405 240.205 ;
        RECT 352.075 238.515 352.405 238.845 ;
        RECT 352.075 237.155 352.405 237.485 ;
        RECT 352.08 237.155 352.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.075 -98.765 352.405 -98.435 ;
        RECT 352.075 -100.125 352.405 -99.795 ;
        RECT 352.075 -101.485 352.405 -101.155 ;
        RECT 352.075 -102.845 352.405 -102.515 ;
        RECT 352.075 -104.205 352.405 -103.875 ;
        RECT 352.075 -105.565 352.405 -105.235 ;
        RECT 352.075 -106.925 352.405 -106.595 ;
        RECT 352.075 -108.285 352.405 -107.955 ;
        RECT 352.075 -109.645 352.405 -109.315 ;
        RECT 352.075 -111.005 352.405 -110.675 ;
        RECT 352.075 -112.365 352.405 -112.035 ;
        RECT 352.075 -113.725 352.405 -113.395 ;
        RECT 352.075 -115.085 352.405 -114.755 ;
        RECT 352.075 -116.445 352.405 -116.115 ;
        RECT 352.075 -117.805 352.405 -117.475 ;
        RECT 352.075 -119.165 352.405 -118.835 ;
        RECT 352.075 -120.525 352.405 -120.195 ;
        RECT 352.075 -121.885 352.405 -121.555 ;
        RECT 352.075 -123.245 352.405 -122.915 ;
        RECT 352.075 -124.605 352.405 -124.275 ;
        RECT 352.075 -125.965 352.405 -125.635 ;
        RECT 352.075 -127.325 352.405 -126.995 ;
        RECT 352.075 -128.685 352.405 -128.355 ;
        RECT 352.075 -130.045 352.405 -129.715 ;
        RECT 352.075 -131.405 352.405 -131.075 ;
        RECT 352.075 -132.765 352.405 -132.435 ;
        RECT 352.075 -134.125 352.405 -133.795 ;
        RECT 352.075 -135.485 352.405 -135.155 ;
        RECT 352.075 -136.845 352.405 -136.515 ;
        RECT 352.075 -138.205 352.405 -137.875 ;
        RECT 352.075 -139.565 352.405 -139.235 ;
        RECT 352.075 -140.925 352.405 -140.595 ;
        RECT 352.075 -142.285 352.405 -141.955 ;
        RECT 352.075 -143.645 352.405 -143.315 ;
        RECT 352.075 -145.005 352.405 -144.675 ;
        RECT 352.075 -146.365 352.405 -146.035 ;
        RECT 352.075 -147.725 352.405 -147.395 ;
        RECT 352.075 -149.085 352.405 -148.755 ;
        RECT 352.075 -150.445 352.405 -150.115 ;
        RECT 352.075 -151.805 352.405 -151.475 ;
        RECT 352.075 -153.165 352.405 -152.835 ;
        RECT 352.075 -154.525 352.405 -154.195 ;
        RECT 352.075 -155.885 352.405 -155.555 ;
        RECT 352.075 -157.245 352.405 -156.915 ;
        RECT 352.075 -158.605 352.405 -158.275 ;
        RECT 352.075 -159.965 352.405 -159.635 ;
        RECT 352.075 -161.325 352.405 -160.995 ;
        RECT 352.075 -162.685 352.405 -162.355 ;
        RECT 352.075 -164.045 352.405 -163.715 ;
        RECT 352.075 -165.405 352.405 -165.075 ;
        RECT 352.075 -166.765 352.405 -166.435 ;
        RECT 352.075 -168.125 352.405 -167.795 ;
        RECT 352.075 -169.485 352.405 -169.155 ;
        RECT 352.075 -170.845 352.405 -170.515 ;
        RECT 352.075 -172.205 352.405 -171.875 ;
        RECT 352.075 -173.565 352.405 -173.235 ;
        RECT 352.075 -174.925 352.405 -174.595 ;
        RECT 352.075 -176.285 352.405 -175.955 ;
        RECT 352.075 -177.645 352.405 -177.315 ;
        RECT 352.075 -179.005 352.405 -178.675 ;
        RECT 352.075 -184.65 352.405 -183.52 ;
        RECT 352.08 -184.765 352.4 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.11 -98.075 352.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.435 244.04 353.765 245.17 ;
        RECT 353.435 239.875 353.765 240.205 ;
        RECT 353.435 238.515 353.765 238.845 ;
        RECT 353.435 237.155 353.765 237.485 ;
        RECT 353.44 237.155 353.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.435 -0.845 353.765 -0.515 ;
        RECT 353.435 -2.205 353.765 -1.875 ;
        RECT 353.435 -3.565 353.765 -3.235 ;
        RECT 353.44 -3.565 353.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 353.435 -96.045 353.765 -95.715 ;
        RECT 353.435 -97.405 353.765 -97.075 ;
        RECT 353.435 -98.765 353.765 -98.435 ;
        RECT 353.435 -100.125 353.765 -99.795 ;
        RECT 353.435 -101.485 353.765 -101.155 ;
        RECT 353.435 -102.845 353.765 -102.515 ;
        RECT 353.435 -104.205 353.765 -103.875 ;
        RECT 353.435 -105.565 353.765 -105.235 ;
        RECT 353.435 -106.925 353.765 -106.595 ;
        RECT 353.435 -108.285 353.765 -107.955 ;
        RECT 353.435 -109.645 353.765 -109.315 ;
        RECT 353.435 -111.005 353.765 -110.675 ;
        RECT 353.435 -112.365 353.765 -112.035 ;
        RECT 353.435 -113.725 353.765 -113.395 ;
        RECT 353.435 -115.085 353.765 -114.755 ;
        RECT 353.435 -116.445 353.765 -116.115 ;
        RECT 353.435 -117.805 353.765 -117.475 ;
        RECT 353.435 -119.165 353.765 -118.835 ;
        RECT 353.435 -120.525 353.765 -120.195 ;
        RECT 353.435 -121.885 353.765 -121.555 ;
        RECT 353.435 -123.245 353.765 -122.915 ;
        RECT 353.435 -124.605 353.765 -124.275 ;
        RECT 353.435 -125.965 353.765 -125.635 ;
        RECT 353.435 -127.325 353.765 -126.995 ;
        RECT 353.435 -128.685 353.765 -128.355 ;
        RECT 353.435 -130.045 353.765 -129.715 ;
        RECT 353.435 -131.405 353.765 -131.075 ;
        RECT 353.435 -132.765 353.765 -132.435 ;
        RECT 353.435 -134.125 353.765 -133.795 ;
        RECT 353.435 -135.485 353.765 -135.155 ;
        RECT 353.435 -136.845 353.765 -136.515 ;
        RECT 353.435 -138.205 353.765 -137.875 ;
        RECT 353.435 -139.565 353.765 -139.235 ;
        RECT 353.435 -140.925 353.765 -140.595 ;
        RECT 353.435 -142.285 353.765 -141.955 ;
        RECT 353.435 -143.645 353.765 -143.315 ;
        RECT 353.435 -145.005 353.765 -144.675 ;
        RECT 353.435 -146.365 353.765 -146.035 ;
        RECT 353.435 -147.725 353.765 -147.395 ;
        RECT 353.435 -149.085 353.765 -148.755 ;
        RECT 353.435 -150.445 353.765 -150.115 ;
        RECT 353.435 -151.805 353.765 -151.475 ;
        RECT 353.435 -153.165 353.765 -152.835 ;
        RECT 353.435 -154.525 353.765 -154.195 ;
        RECT 353.435 -155.885 353.765 -155.555 ;
        RECT 353.435 -157.245 353.765 -156.915 ;
        RECT 353.435 -158.605 353.765 -158.275 ;
        RECT 353.435 -159.965 353.765 -159.635 ;
        RECT 353.435 -161.325 353.765 -160.995 ;
        RECT 353.435 -162.685 353.765 -162.355 ;
        RECT 353.435 -164.045 353.765 -163.715 ;
        RECT 353.435 -165.405 353.765 -165.075 ;
        RECT 353.435 -166.765 353.765 -166.435 ;
        RECT 353.435 -168.125 353.765 -167.795 ;
        RECT 353.435 -169.485 353.765 -169.155 ;
        RECT 353.435 -170.845 353.765 -170.515 ;
        RECT 353.435 -172.205 353.765 -171.875 ;
        RECT 353.435 -173.565 353.765 -173.235 ;
        RECT 353.435 -174.925 353.765 -174.595 ;
        RECT 353.435 -176.285 353.765 -175.955 ;
        RECT 353.435 -177.645 353.765 -177.315 ;
        RECT 353.435 -179.005 353.765 -178.675 ;
        RECT 353.435 -184.65 353.765 -183.52 ;
        RECT 353.44 -184.765 353.76 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.795 244.04 355.125 245.17 ;
        RECT 354.795 239.875 355.125 240.205 ;
        RECT 354.795 238.515 355.125 238.845 ;
        RECT 354.795 237.155 355.125 237.485 ;
        RECT 354.8 237.155 355.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.795 -0.845 355.125 -0.515 ;
        RECT 354.795 -2.205 355.125 -1.875 ;
        RECT 354.795 -3.565 355.125 -3.235 ;
        RECT 354.8 -3.565 355.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.795 -96.045 355.125 -95.715 ;
        RECT 354.795 -97.405 355.125 -97.075 ;
        RECT 354.795 -98.765 355.125 -98.435 ;
        RECT 354.795 -100.125 355.125 -99.795 ;
        RECT 354.795 -101.485 355.125 -101.155 ;
        RECT 354.795 -102.845 355.125 -102.515 ;
        RECT 354.795 -104.205 355.125 -103.875 ;
        RECT 354.795 -105.565 355.125 -105.235 ;
        RECT 354.795 -106.925 355.125 -106.595 ;
        RECT 354.795 -108.285 355.125 -107.955 ;
        RECT 354.795 -109.645 355.125 -109.315 ;
        RECT 354.795 -111.005 355.125 -110.675 ;
        RECT 354.795 -112.365 355.125 -112.035 ;
        RECT 354.795 -113.725 355.125 -113.395 ;
        RECT 354.795 -115.085 355.125 -114.755 ;
        RECT 354.795 -116.445 355.125 -116.115 ;
        RECT 354.795 -117.805 355.125 -117.475 ;
        RECT 354.795 -119.165 355.125 -118.835 ;
        RECT 354.795 -120.525 355.125 -120.195 ;
        RECT 354.795 -121.885 355.125 -121.555 ;
        RECT 354.795 -123.245 355.125 -122.915 ;
        RECT 354.795 -124.605 355.125 -124.275 ;
        RECT 354.795 -125.965 355.125 -125.635 ;
        RECT 354.795 -127.325 355.125 -126.995 ;
        RECT 354.795 -128.685 355.125 -128.355 ;
        RECT 354.795 -130.045 355.125 -129.715 ;
        RECT 354.795 -131.405 355.125 -131.075 ;
        RECT 354.795 -132.765 355.125 -132.435 ;
        RECT 354.795 -134.125 355.125 -133.795 ;
        RECT 354.795 -135.485 355.125 -135.155 ;
        RECT 354.795 -136.845 355.125 -136.515 ;
        RECT 354.795 -138.205 355.125 -137.875 ;
        RECT 354.795 -139.565 355.125 -139.235 ;
        RECT 354.795 -140.925 355.125 -140.595 ;
        RECT 354.795 -142.285 355.125 -141.955 ;
        RECT 354.795 -143.645 355.125 -143.315 ;
        RECT 354.795 -145.005 355.125 -144.675 ;
        RECT 354.795 -146.365 355.125 -146.035 ;
        RECT 354.795 -147.725 355.125 -147.395 ;
        RECT 354.795 -149.085 355.125 -148.755 ;
        RECT 354.795 -150.445 355.125 -150.115 ;
        RECT 354.795 -151.805 355.125 -151.475 ;
        RECT 354.795 -153.165 355.125 -152.835 ;
        RECT 354.795 -154.525 355.125 -154.195 ;
        RECT 354.795 -155.885 355.125 -155.555 ;
        RECT 354.795 -157.245 355.125 -156.915 ;
        RECT 354.795 -158.605 355.125 -158.275 ;
        RECT 354.795 -159.965 355.125 -159.635 ;
        RECT 354.795 -161.325 355.125 -160.995 ;
        RECT 354.795 -162.685 355.125 -162.355 ;
        RECT 354.795 -164.045 355.125 -163.715 ;
        RECT 354.795 -165.405 355.125 -165.075 ;
        RECT 354.795 -166.765 355.125 -166.435 ;
        RECT 354.795 -168.125 355.125 -167.795 ;
        RECT 354.795 -169.485 355.125 -169.155 ;
        RECT 354.795 -170.845 355.125 -170.515 ;
        RECT 354.795 -172.205 355.125 -171.875 ;
        RECT 354.795 -173.565 355.125 -173.235 ;
        RECT 354.795 -174.925 355.125 -174.595 ;
        RECT 354.795 -176.285 355.125 -175.955 ;
        RECT 354.795 -177.645 355.125 -177.315 ;
        RECT 354.795 -179.005 355.125 -178.675 ;
        RECT 354.795 -184.65 355.125 -183.52 ;
        RECT 354.8 -184.765 355.12 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 356.155 22.005 356.485 22.335 ;
        RECT 356.155 19.695 356.485 20.025 ;
        RECT 356.155 18.115 356.485 18.445 ;
        RECT 356.155 17.265 356.485 17.595 ;
        RECT 356.155 14.955 356.485 15.285 ;
        RECT 356.155 14.105 356.485 14.435 ;
        RECT 356.155 11.795 356.485 12.125 ;
        RECT 356.155 10.945 356.485 11.275 ;
        RECT 356.155 8.635 356.485 8.965 ;
        RECT 356.155 7.785 356.485 8.115 ;
        RECT 356.155 5.475 356.485 5.805 ;
        RECT 356.155 3.895 356.485 4.225 ;
        RECT 356.155 3.045 356.485 3.375 ;
        RECT 356.155 0.87 356.485 1.2 ;
        RECT 356.155 -0.845 356.485 -0.515 ;
        RECT 356.155 -2.205 356.485 -1.875 ;
        RECT 356.155 -3.565 356.485 -3.235 ;
        RECT 356.155 -4.925 356.485 -4.595 ;
        RECT 356.155 -6.285 356.485 -5.955 ;
        RECT 356.155 -7.645 356.485 -7.315 ;
        RECT 356.155 -9.005 356.485 -8.675 ;
        RECT 356.155 -10.365 356.485 -10.035 ;
        RECT 356.155 -11.725 356.485 -11.395 ;
        RECT 356.155 -13.085 356.485 -12.755 ;
        RECT 356.155 -14.445 356.485 -14.115 ;
        RECT 356.155 -15.805 356.485 -15.475 ;
        RECT 356.155 -17.165 356.485 -16.835 ;
        RECT 356.155 -18.525 356.485 -18.195 ;
        RECT 356.155 -19.885 356.485 -19.555 ;
        RECT 356.155 -21.245 356.485 -20.915 ;
        RECT 356.155 -22.605 356.485 -22.275 ;
        RECT 356.155 -23.965 356.485 -23.635 ;
        RECT 356.155 -25.325 356.485 -24.995 ;
        RECT 356.155 -26.685 356.485 -26.355 ;
        RECT 356.155 -28.045 356.485 -27.715 ;
        RECT 356.155 -29.405 356.485 -29.075 ;
        RECT 356.155 -30.765 356.485 -30.435 ;
        RECT 356.155 -32.125 356.485 -31.795 ;
        RECT 356.155 -33.485 356.485 -33.155 ;
        RECT 356.155 -34.845 356.485 -34.515 ;
        RECT 356.155 -36.205 356.485 -35.875 ;
        RECT 356.155 -37.565 356.485 -37.235 ;
        RECT 356.155 -38.925 356.485 -38.595 ;
        RECT 356.155 -40.285 356.485 -39.955 ;
        RECT 356.155 -41.645 356.485 -41.315 ;
        RECT 356.155 -43.005 356.485 -42.675 ;
        RECT 356.155 -44.365 356.485 -44.035 ;
        RECT 356.155 -45.725 356.485 -45.395 ;
        RECT 356.155 -47.085 356.485 -46.755 ;
        RECT 356.155 -48.445 356.485 -48.115 ;
        RECT 356.155 -49.805 356.485 -49.475 ;
        RECT 356.155 -51.165 356.485 -50.835 ;
        RECT 356.155 -52.525 356.485 -52.195 ;
        RECT 356.155 -53.885 356.485 -53.555 ;
        RECT 356.155 -55.245 356.485 -54.915 ;
        RECT 356.155 -56.605 356.485 -56.275 ;
        RECT 356.155 -57.965 356.485 -57.635 ;
        RECT 356.155 -59.325 356.485 -58.995 ;
        RECT 356.155 -60.685 356.485 -60.355 ;
        RECT 356.155 -62.045 356.485 -61.715 ;
        RECT 356.155 -63.405 356.485 -63.075 ;
        RECT 356.155 -64.765 356.485 -64.435 ;
        RECT 356.155 -66.125 356.485 -65.795 ;
        RECT 356.155 -67.485 356.485 -67.155 ;
        RECT 356.155 -68.845 356.485 -68.515 ;
        RECT 356.155 -70.205 356.485 -69.875 ;
        RECT 356.155 -71.565 356.485 -71.235 ;
        RECT 356.155 -72.925 356.485 -72.595 ;
        RECT 356.155 -74.285 356.485 -73.955 ;
        RECT 356.155 -75.645 356.485 -75.315 ;
        RECT 356.155 -77.005 356.485 -76.675 ;
        RECT 356.155 -78.365 356.485 -78.035 ;
        RECT 356.155 -79.725 356.485 -79.395 ;
        RECT 356.155 -81.085 356.485 -80.755 ;
        RECT 356.155 -82.445 356.485 -82.115 ;
        RECT 356.155 -83.805 356.485 -83.475 ;
        RECT 356.155 -85.165 356.485 -84.835 ;
        RECT 356.155 -86.525 356.485 -86.195 ;
        RECT 356.155 -87.885 356.485 -87.555 ;
        RECT 356.155 -89.245 356.485 -88.915 ;
        RECT 356.155 -90.605 356.485 -90.275 ;
        RECT 356.155 -91.965 356.485 -91.635 ;
        RECT 356.155 -93.325 356.485 -92.995 ;
        RECT 356.155 -94.685 356.485 -94.355 ;
        RECT 356.155 -96.045 356.485 -95.715 ;
        RECT 356.155 -97.405 356.485 -97.075 ;
        RECT 356.155 -98.765 356.485 -98.435 ;
        RECT 356.155 -100.125 356.485 -99.795 ;
        RECT 356.155 -101.485 356.485 -101.155 ;
        RECT 356.155 -102.845 356.485 -102.515 ;
        RECT 356.155 -104.205 356.485 -103.875 ;
        RECT 356.155 -105.565 356.485 -105.235 ;
        RECT 356.155 -106.925 356.485 -106.595 ;
        RECT 356.155 -108.285 356.485 -107.955 ;
        RECT 356.155 -109.645 356.485 -109.315 ;
        RECT 356.155 -111.005 356.485 -110.675 ;
        RECT 356.155 -112.365 356.485 -112.035 ;
        RECT 356.155 -113.725 356.485 -113.395 ;
        RECT 356.155 -115.085 356.485 -114.755 ;
        RECT 356.155 -116.445 356.485 -116.115 ;
        RECT 356.155 -117.805 356.485 -117.475 ;
        RECT 356.155 -119.165 356.485 -118.835 ;
        RECT 356.155 -120.525 356.485 -120.195 ;
        RECT 356.155 -121.885 356.485 -121.555 ;
        RECT 356.155 -123.245 356.485 -122.915 ;
        RECT 356.155 -124.605 356.485 -124.275 ;
        RECT 356.155 -125.965 356.485 -125.635 ;
        RECT 356.155 -127.325 356.485 -126.995 ;
        RECT 356.155 -128.685 356.485 -128.355 ;
        RECT 356.155 -130.045 356.485 -129.715 ;
        RECT 356.155 -131.405 356.485 -131.075 ;
        RECT 356.155 -132.765 356.485 -132.435 ;
        RECT 356.155 -134.125 356.485 -133.795 ;
        RECT 356.155 -135.485 356.485 -135.155 ;
        RECT 356.155 -136.845 356.485 -136.515 ;
        RECT 356.155 -138.205 356.485 -137.875 ;
        RECT 356.155 -139.565 356.485 -139.235 ;
        RECT 356.155 -140.925 356.485 -140.595 ;
        RECT 356.155 -142.285 356.485 -141.955 ;
        RECT 356.155 -143.645 356.485 -143.315 ;
        RECT 356.155 -145.005 356.485 -144.675 ;
        RECT 356.155 -146.365 356.485 -146.035 ;
        RECT 356.155 -147.725 356.485 -147.395 ;
        RECT 356.155 -149.085 356.485 -148.755 ;
        RECT 356.155 -150.445 356.485 -150.115 ;
        RECT 356.155 -151.805 356.485 -151.475 ;
        RECT 356.155 -153.165 356.485 -152.835 ;
        RECT 356.155 -154.525 356.485 -154.195 ;
        RECT 356.155 -155.885 356.485 -155.555 ;
        RECT 356.155 -157.245 356.485 -156.915 ;
        RECT 356.155 -158.605 356.485 -158.275 ;
        RECT 356.155 -159.965 356.485 -159.635 ;
        RECT 356.155 -161.325 356.485 -160.995 ;
        RECT 356.155 -162.685 356.485 -162.355 ;
        RECT 356.155 -164.045 356.485 -163.715 ;
        RECT 356.155 -165.405 356.485 -165.075 ;
        RECT 356.155 -166.765 356.485 -166.435 ;
        RECT 356.155 -168.125 356.485 -167.795 ;
        RECT 356.155 -169.485 356.485 -169.155 ;
        RECT 356.155 -170.845 356.485 -170.515 ;
        RECT 356.155 -172.205 356.485 -171.875 ;
        RECT 356.155 -173.565 356.485 -173.235 ;
        RECT 356.155 -174.925 356.485 -174.595 ;
        RECT 356.155 -176.285 356.485 -175.955 ;
        RECT 356.155 -177.645 356.485 -177.315 ;
        RECT 356.155 -179.005 356.485 -178.675 ;
        RECT 356.155 -184.65 356.485 -183.52 ;
        RECT 356.16 -184.765 356.48 245.285 ;
        RECT 356.155 244.04 356.485 245.17 ;
        RECT 356.155 239.875 356.485 240.205 ;
        RECT 356.155 238.515 356.485 238.845 ;
        RECT 356.155 237.155 356.485 237.485 ;
        RECT 356.155 235.17 356.485 235.5 ;
        RECT 356.155 232.995 356.485 233.325 ;
        RECT 356.155 231.415 356.485 231.745 ;
        RECT 356.155 230.565 356.485 230.895 ;
        RECT 356.155 228.255 356.485 228.585 ;
        RECT 356.155 227.405 356.485 227.735 ;
        RECT 356.155 225.095 356.485 225.425 ;
        RECT 356.155 224.245 356.485 224.575 ;
        RECT 356.155 221.935 356.485 222.265 ;
        RECT 356.155 221.085 356.485 221.415 ;
        RECT 356.155 218.775 356.485 219.105 ;
        RECT 356.155 217.195 356.485 217.525 ;
        RECT 356.155 216.345 356.485 216.675 ;
        RECT 356.155 214.035 356.485 214.365 ;
        RECT 356.155 213.185 356.485 213.515 ;
        RECT 356.155 210.875 356.485 211.205 ;
        RECT 356.155 210.025 356.485 210.355 ;
        RECT 356.155 207.715 356.485 208.045 ;
        RECT 356.155 206.865 356.485 207.195 ;
        RECT 356.155 204.555 356.485 204.885 ;
        RECT 356.155 202.975 356.485 203.305 ;
        RECT 356.155 202.125 356.485 202.455 ;
        RECT 356.155 199.815 356.485 200.145 ;
        RECT 356.155 198.965 356.485 199.295 ;
        RECT 356.155 196.655 356.485 196.985 ;
        RECT 356.155 195.805 356.485 196.135 ;
        RECT 356.155 193.495 356.485 193.825 ;
        RECT 356.155 192.645 356.485 192.975 ;
        RECT 356.155 190.335 356.485 190.665 ;
        RECT 356.155 188.755 356.485 189.085 ;
        RECT 356.155 187.905 356.485 188.235 ;
        RECT 356.155 185.595 356.485 185.925 ;
        RECT 356.155 184.745 356.485 185.075 ;
        RECT 356.155 182.435 356.485 182.765 ;
        RECT 356.155 181.585 356.485 181.915 ;
        RECT 356.155 179.275 356.485 179.605 ;
        RECT 356.155 178.425 356.485 178.755 ;
        RECT 356.155 176.115 356.485 176.445 ;
        RECT 356.155 174.535 356.485 174.865 ;
        RECT 356.155 173.685 356.485 174.015 ;
        RECT 356.155 171.375 356.485 171.705 ;
        RECT 356.155 170.525 356.485 170.855 ;
        RECT 356.155 168.215 356.485 168.545 ;
        RECT 356.155 167.365 356.485 167.695 ;
        RECT 356.155 165.055 356.485 165.385 ;
        RECT 356.155 164.205 356.485 164.535 ;
        RECT 356.155 161.895 356.485 162.225 ;
        RECT 356.155 160.315 356.485 160.645 ;
        RECT 356.155 159.465 356.485 159.795 ;
        RECT 356.155 157.155 356.485 157.485 ;
        RECT 356.155 156.305 356.485 156.635 ;
        RECT 356.155 153.995 356.485 154.325 ;
        RECT 356.155 153.145 356.485 153.475 ;
        RECT 356.155 150.835 356.485 151.165 ;
        RECT 356.155 149.985 356.485 150.315 ;
        RECT 356.155 147.675 356.485 148.005 ;
        RECT 356.155 146.095 356.485 146.425 ;
        RECT 356.155 145.245 356.485 145.575 ;
        RECT 356.155 142.935 356.485 143.265 ;
        RECT 356.155 142.085 356.485 142.415 ;
        RECT 356.155 139.775 356.485 140.105 ;
        RECT 356.155 138.925 356.485 139.255 ;
        RECT 356.155 136.615 356.485 136.945 ;
        RECT 356.155 135.765 356.485 136.095 ;
        RECT 356.155 133.455 356.485 133.785 ;
        RECT 356.155 131.875 356.485 132.205 ;
        RECT 356.155 131.025 356.485 131.355 ;
        RECT 356.155 128.715 356.485 129.045 ;
        RECT 356.155 127.865 356.485 128.195 ;
        RECT 356.155 125.555 356.485 125.885 ;
        RECT 356.155 124.705 356.485 125.035 ;
        RECT 356.155 122.395 356.485 122.725 ;
        RECT 356.155 121.545 356.485 121.875 ;
        RECT 356.155 119.235 356.485 119.565 ;
        RECT 356.155 117.655 356.485 117.985 ;
        RECT 356.155 116.805 356.485 117.135 ;
        RECT 356.155 114.495 356.485 114.825 ;
        RECT 356.155 113.645 356.485 113.975 ;
        RECT 356.155 111.335 356.485 111.665 ;
        RECT 356.155 110.485 356.485 110.815 ;
        RECT 356.155 108.175 356.485 108.505 ;
        RECT 356.155 107.325 356.485 107.655 ;
        RECT 356.155 105.015 356.485 105.345 ;
        RECT 356.155 103.435 356.485 103.765 ;
        RECT 356.155 102.585 356.485 102.915 ;
        RECT 356.155 100.275 356.485 100.605 ;
        RECT 356.155 99.425 356.485 99.755 ;
        RECT 356.155 97.115 356.485 97.445 ;
        RECT 356.155 96.265 356.485 96.595 ;
        RECT 356.155 93.955 356.485 94.285 ;
        RECT 356.155 93.105 356.485 93.435 ;
        RECT 356.155 90.795 356.485 91.125 ;
        RECT 356.155 89.215 356.485 89.545 ;
        RECT 356.155 88.365 356.485 88.695 ;
        RECT 356.155 86.055 356.485 86.385 ;
        RECT 356.155 85.205 356.485 85.535 ;
        RECT 356.155 82.895 356.485 83.225 ;
        RECT 356.155 82.045 356.485 82.375 ;
        RECT 356.155 79.735 356.485 80.065 ;
        RECT 356.155 78.885 356.485 79.215 ;
        RECT 356.155 76.575 356.485 76.905 ;
        RECT 356.155 74.995 356.485 75.325 ;
        RECT 356.155 74.145 356.485 74.475 ;
        RECT 356.155 71.835 356.485 72.165 ;
        RECT 356.155 70.985 356.485 71.315 ;
        RECT 356.155 68.675 356.485 69.005 ;
        RECT 356.155 67.825 356.485 68.155 ;
        RECT 356.155 65.515 356.485 65.845 ;
        RECT 356.155 64.665 356.485 64.995 ;
        RECT 356.155 62.355 356.485 62.685 ;
        RECT 356.155 60.775 356.485 61.105 ;
        RECT 356.155 59.925 356.485 60.255 ;
        RECT 356.155 57.615 356.485 57.945 ;
        RECT 356.155 56.765 356.485 57.095 ;
        RECT 356.155 54.455 356.485 54.785 ;
        RECT 356.155 53.605 356.485 53.935 ;
        RECT 356.155 51.295 356.485 51.625 ;
        RECT 356.155 50.445 356.485 50.775 ;
        RECT 356.155 48.135 356.485 48.465 ;
        RECT 356.155 46.555 356.485 46.885 ;
        RECT 356.155 45.705 356.485 46.035 ;
        RECT 356.155 43.395 356.485 43.725 ;
        RECT 356.155 42.545 356.485 42.875 ;
        RECT 356.155 40.235 356.485 40.565 ;
        RECT 356.155 39.385 356.485 39.715 ;
        RECT 356.155 37.075 356.485 37.405 ;
        RECT 356.155 36.225 356.485 36.555 ;
        RECT 356.155 33.915 356.485 34.245 ;
        RECT 356.155 32.335 356.485 32.665 ;
        RECT 356.155 31.485 356.485 31.815 ;
        RECT 356.155 29.175 356.485 29.505 ;
        RECT 356.155 28.325 356.485 28.655 ;
        RECT 356.155 26.015 356.485 26.345 ;
        RECT 356.155 25.165 356.485 25.495 ;
        RECT 356.155 22.855 356.485 23.185 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.995 244.04 314.325 245.17 ;
        RECT 313.995 239.875 314.325 240.205 ;
        RECT 313.995 238.515 314.325 238.845 ;
        RECT 313.995 237.155 314.325 237.485 ;
        RECT 314 237.155 314.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.995 -0.845 314.325 -0.515 ;
        RECT 313.995 -2.205 314.325 -1.875 ;
        RECT 313.995 -3.565 314.325 -3.235 ;
        RECT 314 -3.565 314.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.995 -96.045 314.325 -95.715 ;
        RECT 313.995 -97.405 314.325 -97.075 ;
        RECT 313.995 -98.765 314.325 -98.435 ;
        RECT 313.995 -100.125 314.325 -99.795 ;
        RECT 313.995 -101.485 314.325 -101.155 ;
        RECT 313.995 -102.845 314.325 -102.515 ;
        RECT 313.995 -104.205 314.325 -103.875 ;
        RECT 313.995 -105.565 314.325 -105.235 ;
        RECT 313.995 -106.925 314.325 -106.595 ;
        RECT 313.995 -108.285 314.325 -107.955 ;
        RECT 313.995 -109.645 314.325 -109.315 ;
        RECT 313.995 -111.005 314.325 -110.675 ;
        RECT 313.995 -112.365 314.325 -112.035 ;
        RECT 313.995 -113.725 314.325 -113.395 ;
        RECT 313.995 -115.085 314.325 -114.755 ;
        RECT 313.995 -116.445 314.325 -116.115 ;
        RECT 313.995 -117.805 314.325 -117.475 ;
        RECT 313.995 -119.165 314.325 -118.835 ;
        RECT 313.995 -120.525 314.325 -120.195 ;
        RECT 313.995 -121.885 314.325 -121.555 ;
        RECT 313.995 -123.245 314.325 -122.915 ;
        RECT 313.995 -124.605 314.325 -124.275 ;
        RECT 313.995 -125.965 314.325 -125.635 ;
        RECT 313.995 -127.325 314.325 -126.995 ;
        RECT 313.995 -128.685 314.325 -128.355 ;
        RECT 313.995 -130.045 314.325 -129.715 ;
        RECT 313.995 -131.405 314.325 -131.075 ;
        RECT 313.995 -132.765 314.325 -132.435 ;
        RECT 313.995 -134.125 314.325 -133.795 ;
        RECT 313.995 -135.485 314.325 -135.155 ;
        RECT 313.995 -136.845 314.325 -136.515 ;
        RECT 313.995 -138.205 314.325 -137.875 ;
        RECT 313.995 -139.565 314.325 -139.235 ;
        RECT 313.995 -140.925 314.325 -140.595 ;
        RECT 313.995 -142.285 314.325 -141.955 ;
        RECT 313.995 -143.645 314.325 -143.315 ;
        RECT 313.995 -145.005 314.325 -144.675 ;
        RECT 313.995 -146.365 314.325 -146.035 ;
        RECT 313.995 -147.725 314.325 -147.395 ;
        RECT 313.995 -149.085 314.325 -148.755 ;
        RECT 313.995 -150.445 314.325 -150.115 ;
        RECT 313.995 -151.805 314.325 -151.475 ;
        RECT 313.995 -153.165 314.325 -152.835 ;
        RECT 313.995 -154.525 314.325 -154.195 ;
        RECT 313.995 -155.885 314.325 -155.555 ;
        RECT 313.995 -157.245 314.325 -156.915 ;
        RECT 313.995 -158.605 314.325 -158.275 ;
        RECT 313.995 -159.965 314.325 -159.635 ;
        RECT 313.995 -161.325 314.325 -160.995 ;
        RECT 313.995 -162.685 314.325 -162.355 ;
        RECT 313.995 -164.045 314.325 -163.715 ;
        RECT 313.995 -165.405 314.325 -165.075 ;
        RECT 313.995 -166.765 314.325 -166.435 ;
        RECT 313.995 -168.125 314.325 -167.795 ;
        RECT 313.995 -169.485 314.325 -169.155 ;
        RECT 313.995 -170.845 314.325 -170.515 ;
        RECT 313.995 -172.205 314.325 -171.875 ;
        RECT 313.995 -173.565 314.325 -173.235 ;
        RECT 313.995 -174.925 314.325 -174.595 ;
        RECT 313.995 -176.285 314.325 -175.955 ;
        RECT 313.995 -177.645 314.325 -177.315 ;
        RECT 313.995 -179.005 314.325 -178.675 ;
        RECT 313.995 -184.65 314.325 -183.52 ;
        RECT 314 -184.765 314.32 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.355 244.04 315.685 245.17 ;
        RECT 315.355 239.875 315.685 240.205 ;
        RECT 315.355 238.515 315.685 238.845 ;
        RECT 315.355 237.155 315.685 237.485 ;
        RECT 315.36 237.155 315.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.355 -0.845 315.685 -0.515 ;
        RECT 315.355 -2.205 315.685 -1.875 ;
        RECT 315.355 -3.565 315.685 -3.235 ;
        RECT 315.36 -3.565 315.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 315.355 -96.045 315.685 -95.715 ;
        RECT 315.355 -97.405 315.685 -97.075 ;
        RECT 315.355 -98.765 315.685 -98.435 ;
        RECT 315.355 -100.125 315.685 -99.795 ;
        RECT 315.355 -101.485 315.685 -101.155 ;
        RECT 315.355 -102.845 315.685 -102.515 ;
        RECT 315.355 -104.205 315.685 -103.875 ;
        RECT 315.355 -105.565 315.685 -105.235 ;
        RECT 315.355 -106.925 315.685 -106.595 ;
        RECT 315.355 -108.285 315.685 -107.955 ;
        RECT 315.355 -109.645 315.685 -109.315 ;
        RECT 315.355 -111.005 315.685 -110.675 ;
        RECT 315.355 -112.365 315.685 -112.035 ;
        RECT 315.355 -113.725 315.685 -113.395 ;
        RECT 315.355 -115.085 315.685 -114.755 ;
        RECT 315.355 -116.445 315.685 -116.115 ;
        RECT 315.355 -117.805 315.685 -117.475 ;
        RECT 315.355 -119.165 315.685 -118.835 ;
        RECT 315.355 -120.525 315.685 -120.195 ;
        RECT 315.355 -121.885 315.685 -121.555 ;
        RECT 315.355 -123.245 315.685 -122.915 ;
        RECT 315.355 -124.605 315.685 -124.275 ;
        RECT 315.355 -125.965 315.685 -125.635 ;
        RECT 315.355 -127.325 315.685 -126.995 ;
        RECT 315.355 -128.685 315.685 -128.355 ;
        RECT 315.355 -130.045 315.685 -129.715 ;
        RECT 315.355 -131.405 315.685 -131.075 ;
        RECT 315.355 -132.765 315.685 -132.435 ;
        RECT 315.355 -134.125 315.685 -133.795 ;
        RECT 315.355 -135.485 315.685 -135.155 ;
        RECT 315.355 -136.845 315.685 -136.515 ;
        RECT 315.355 -138.205 315.685 -137.875 ;
        RECT 315.355 -139.565 315.685 -139.235 ;
        RECT 315.355 -140.925 315.685 -140.595 ;
        RECT 315.355 -142.285 315.685 -141.955 ;
        RECT 315.355 -143.645 315.685 -143.315 ;
        RECT 315.355 -145.005 315.685 -144.675 ;
        RECT 315.355 -146.365 315.685 -146.035 ;
        RECT 315.355 -147.725 315.685 -147.395 ;
        RECT 315.355 -149.085 315.685 -148.755 ;
        RECT 315.355 -150.445 315.685 -150.115 ;
        RECT 315.355 -151.805 315.685 -151.475 ;
        RECT 315.355 -153.165 315.685 -152.835 ;
        RECT 315.355 -154.525 315.685 -154.195 ;
        RECT 315.355 -155.885 315.685 -155.555 ;
        RECT 315.355 -157.245 315.685 -156.915 ;
        RECT 315.355 -158.605 315.685 -158.275 ;
        RECT 315.355 -159.965 315.685 -159.635 ;
        RECT 315.355 -161.325 315.685 -160.995 ;
        RECT 315.355 -162.685 315.685 -162.355 ;
        RECT 315.355 -164.045 315.685 -163.715 ;
        RECT 315.355 -165.405 315.685 -165.075 ;
        RECT 315.355 -166.765 315.685 -166.435 ;
        RECT 315.355 -168.125 315.685 -167.795 ;
        RECT 315.355 -169.485 315.685 -169.155 ;
        RECT 315.355 -170.845 315.685 -170.515 ;
        RECT 315.355 -172.205 315.685 -171.875 ;
        RECT 315.355 -173.565 315.685 -173.235 ;
        RECT 315.355 -174.925 315.685 -174.595 ;
        RECT 315.355 -176.285 315.685 -175.955 ;
        RECT 315.355 -177.645 315.685 -177.315 ;
        RECT 315.355 -179.005 315.685 -178.675 ;
        RECT 315.355 -184.65 315.685 -183.52 ;
        RECT 315.36 -184.765 315.68 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.715 244.04 317.045 245.17 ;
        RECT 316.715 239.875 317.045 240.205 ;
        RECT 316.715 238.515 317.045 238.845 ;
        RECT 316.715 237.155 317.045 237.485 ;
        RECT 316.72 237.155 317.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.715 -0.845 317.045 -0.515 ;
        RECT 316.715 -2.205 317.045 -1.875 ;
        RECT 316.715 -3.565 317.045 -3.235 ;
        RECT 316.72 -3.565 317.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.715 -96.045 317.045 -95.715 ;
        RECT 316.715 -97.405 317.045 -97.075 ;
        RECT 316.715 -98.765 317.045 -98.435 ;
        RECT 316.715 -100.125 317.045 -99.795 ;
        RECT 316.715 -101.485 317.045 -101.155 ;
        RECT 316.715 -102.845 317.045 -102.515 ;
        RECT 316.715 -104.205 317.045 -103.875 ;
        RECT 316.715 -105.565 317.045 -105.235 ;
        RECT 316.715 -106.925 317.045 -106.595 ;
        RECT 316.715 -108.285 317.045 -107.955 ;
        RECT 316.715 -109.645 317.045 -109.315 ;
        RECT 316.715 -111.005 317.045 -110.675 ;
        RECT 316.715 -112.365 317.045 -112.035 ;
        RECT 316.715 -113.725 317.045 -113.395 ;
        RECT 316.715 -115.085 317.045 -114.755 ;
        RECT 316.715 -116.445 317.045 -116.115 ;
        RECT 316.715 -117.805 317.045 -117.475 ;
        RECT 316.715 -119.165 317.045 -118.835 ;
        RECT 316.715 -120.525 317.045 -120.195 ;
        RECT 316.715 -121.885 317.045 -121.555 ;
        RECT 316.715 -123.245 317.045 -122.915 ;
        RECT 316.715 -124.605 317.045 -124.275 ;
        RECT 316.715 -125.965 317.045 -125.635 ;
        RECT 316.715 -127.325 317.045 -126.995 ;
        RECT 316.715 -128.685 317.045 -128.355 ;
        RECT 316.715 -130.045 317.045 -129.715 ;
        RECT 316.715 -131.405 317.045 -131.075 ;
        RECT 316.715 -132.765 317.045 -132.435 ;
        RECT 316.715 -134.125 317.045 -133.795 ;
        RECT 316.715 -135.485 317.045 -135.155 ;
        RECT 316.715 -136.845 317.045 -136.515 ;
        RECT 316.715 -138.205 317.045 -137.875 ;
        RECT 316.715 -139.565 317.045 -139.235 ;
        RECT 316.715 -140.925 317.045 -140.595 ;
        RECT 316.715 -142.285 317.045 -141.955 ;
        RECT 316.715 -143.645 317.045 -143.315 ;
        RECT 316.715 -145.005 317.045 -144.675 ;
        RECT 316.715 -146.365 317.045 -146.035 ;
        RECT 316.715 -147.725 317.045 -147.395 ;
        RECT 316.715 -149.085 317.045 -148.755 ;
        RECT 316.715 -150.445 317.045 -150.115 ;
        RECT 316.715 -151.805 317.045 -151.475 ;
        RECT 316.715 -153.165 317.045 -152.835 ;
        RECT 316.715 -154.525 317.045 -154.195 ;
        RECT 316.715 -155.885 317.045 -155.555 ;
        RECT 316.715 -157.245 317.045 -156.915 ;
        RECT 316.715 -158.605 317.045 -158.275 ;
        RECT 316.715 -159.965 317.045 -159.635 ;
        RECT 316.715 -161.325 317.045 -160.995 ;
        RECT 316.715 -162.685 317.045 -162.355 ;
        RECT 316.715 -164.045 317.045 -163.715 ;
        RECT 316.715 -165.405 317.045 -165.075 ;
        RECT 316.715 -166.765 317.045 -166.435 ;
        RECT 316.715 -168.125 317.045 -167.795 ;
        RECT 316.715 -169.485 317.045 -169.155 ;
        RECT 316.715 -170.845 317.045 -170.515 ;
        RECT 316.715 -172.205 317.045 -171.875 ;
        RECT 316.715 -173.565 317.045 -173.235 ;
        RECT 316.715 -174.925 317.045 -174.595 ;
        RECT 316.715 -176.285 317.045 -175.955 ;
        RECT 316.715 -177.645 317.045 -177.315 ;
        RECT 316.715 -179.005 317.045 -178.675 ;
        RECT 316.715 -184.65 317.045 -183.52 ;
        RECT 316.72 -184.765 317.04 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.075 244.04 318.405 245.17 ;
        RECT 318.075 239.875 318.405 240.205 ;
        RECT 318.075 238.515 318.405 238.845 ;
        RECT 318.075 237.155 318.405 237.485 ;
        RECT 318.08 237.155 318.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.075 -0.845 318.405 -0.515 ;
        RECT 318.075 -2.205 318.405 -1.875 ;
        RECT 318.075 -3.565 318.405 -3.235 ;
        RECT 318.08 -3.565 318.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.075 -96.045 318.405 -95.715 ;
        RECT 318.075 -97.405 318.405 -97.075 ;
        RECT 318.075 -98.765 318.405 -98.435 ;
        RECT 318.075 -100.125 318.405 -99.795 ;
        RECT 318.075 -101.485 318.405 -101.155 ;
        RECT 318.075 -102.845 318.405 -102.515 ;
        RECT 318.075 -104.205 318.405 -103.875 ;
        RECT 318.075 -105.565 318.405 -105.235 ;
        RECT 318.075 -106.925 318.405 -106.595 ;
        RECT 318.075 -108.285 318.405 -107.955 ;
        RECT 318.075 -109.645 318.405 -109.315 ;
        RECT 318.075 -111.005 318.405 -110.675 ;
        RECT 318.075 -112.365 318.405 -112.035 ;
        RECT 318.075 -113.725 318.405 -113.395 ;
        RECT 318.075 -115.085 318.405 -114.755 ;
        RECT 318.075 -116.445 318.405 -116.115 ;
        RECT 318.075 -117.805 318.405 -117.475 ;
        RECT 318.075 -119.165 318.405 -118.835 ;
        RECT 318.075 -120.525 318.405 -120.195 ;
        RECT 318.075 -121.885 318.405 -121.555 ;
        RECT 318.075 -123.245 318.405 -122.915 ;
        RECT 318.075 -124.605 318.405 -124.275 ;
        RECT 318.075 -125.965 318.405 -125.635 ;
        RECT 318.075 -127.325 318.405 -126.995 ;
        RECT 318.075 -128.685 318.405 -128.355 ;
        RECT 318.075 -130.045 318.405 -129.715 ;
        RECT 318.075 -131.405 318.405 -131.075 ;
        RECT 318.075 -132.765 318.405 -132.435 ;
        RECT 318.075 -134.125 318.405 -133.795 ;
        RECT 318.075 -135.485 318.405 -135.155 ;
        RECT 318.075 -136.845 318.405 -136.515 ;
        RECT 318.075 -138.205 318.405 -137.875 ;
        RECT 318.075 -139.565 318.405 -139.235 ;
        RECT 318.075 -140.925 318.405 -140.595 ;
        RECT 318.075 -142.285 318.405 -141.955 ;
        RECT 318.075 -143.645 318.405 -143.315 ;
        RECT 318.075 -145.005 318.405 -144.675 ;
        RECT 318.075 -146.365 318.405 -146.035 ;
        RECT 318.075 -147.725 318.405 -147.395 ;
        RECT 318.075 -149.085 318.405 -148.755 ;
        RECT 318.075 -150.445 318.405 -150.115 ;
        RECT 318.075 -151.805 318.405 -151.475 ;
        RECT 318.075 -153.165 318.405 -152.835 ;
        RECT 318.075 -154.525 318.405 -154.195 ;
        RECT 318.075 -155.885 318.405 -155.555 ;
        RECT 318.075 -157.245 318.405 -156.915 ;
        RECT 318.075 -158.605 318.405 -158.275 ;
        RECT 318.075 -159.965 318.405 -159.635 ;
        RECT 318.075 -161.325 318.405 -160.995 ;
        RECT 318.075 -162.685 318.405 -162.355 ;
        RECT 318.075 -164.045 318.405 -163.715 ;
        RECT 318.075 -165.405 318.405 -165.075 ;
        RECT 318.075 -166.765 318.405 -166.435 ;
        RECT 318.075 -168.125 318.405 -167.795 ;
        RECT 318.075 -169.485 318.405 -169.155 ;
        RECT 318.075 -170.845 318.405 -170.515 ;
        RECT 318.075 -172.205 318.405 -171.875 ;
        RECT 318.075 -173.565 318.405 -173.235 ;
        RECT 318.075 -174.925 318.405 -174.595 ;
        RECT 318.075 -176.285 318.405 -175.955 ;
        RECT 318.075 -177.645 318.405 -177.315 ;
        RECT 318.075 -179.005 318.405 -178.675 ;
        RECT 318.075 -184.65 318.405 -183.52 ;
        RECT 318.08 -184.765 318.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.76 -98.075 319.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.435 244.04 319.765 245.17 ;
        RECT 319.435 239.875 319.765 240.205 ;
        RECT 319.435 238.515 319.765 238.845 ;
        RECT 319.435 237.155 319.765 237.485 ;
        RECT 319.44 237.155 319.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.795 244.04 321.125 245.17 ;
        RECT 320.795 239.875 321.125 240.205 ;
        RECT 320.795 238.515 321.125 238.845 ;
        RECT 320.795 237.155 321.125 237.485 ;
        RECT 320.8 237.155 321.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.795 -0.845 321.125 -0.515 ;
        RECT 320.795 -2.205 321.125 -1.875 ;
        RECT 320.795 -3.565 321.125 -3.235 ;
        RECT 320.8 -3.565 321.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.155 244.04 322.485 245.17 ;
        RECT 322.155 239.875 322.485 240.205 ;
        RECT 322.155 238.515 322.485 238.845 ;
        RECT 322.155 237.155 322.485 237.485 ;
        RECT 322.16 237.155 322.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.155 -0.845 322.485 -0.515 ;
        RECT 322.155 -2.205 322.485 -1.875 ;
        RECT 322.155 -3.565 322.485 -3.235 ;
        RECT 322.16 -3.565 322.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.515 244.04 323.845 245.17 ;
        RECT 323.515 239.875 323.845 240.205 ;
        RECT 323.515 238.515 323.845 238.845 ;
        RECT 323.515 237.155 323.845 237.485 ;
        RECT 323.52 237.155 323.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.515 -0.845 323.845 -0.515 ;
        RECT 323.515 -2.205 323.845 -1.875 ;
        RECT 323.515 -3.565 323.845 -3.235 ;
        RECT 323.52 -3.565 323.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 323.515 -96.045 323.845 -95.715 ;
        RECT 323.515 -97.405 323.845 -97.075 ;
        RECT 323.515 -98.765 323.845 -98.435 ;
        RECT 323.515 -100.125 323.845 -99.795 ;
        RECT 323.515 -101.485 323.845 -101.155 ;
        RECT 323.515 -102.845 323.845 -102.515 ;
        RECT 323.515 -104.205 323.845 -103.875 ;
        RECT 323.515 -105.565 323.845 -105.235 ;
        RECT 323.515 -106.925 323.845 -106.595 ;
        RECT 323.515 -108.285 323.845 -107.955 ;
        RECT 323.515 -109.645 323.845 -109.315 ;
        RECT 323.515 -111.005 323.845 -110.675 ;
        RECT 323.515 -112.365 323.845 -112.035 ;
        RECT 323.515 -113.725 323.845 -113.395 ;
        RECT 323.515 -115.085 323.845 -114.755 ;
        RECT 323.515 -116.445 323.845 -116.115 ;
        RECT 323.515 -117.805 323.845 -117.475 ;
        RECT 323.515 -119.165 323.845 -118.835 ;
        RECT 323.515 -120.525 323.845 -120.195 ;
        RECT 323.515 -121.885 323.845 -121.555 ;
        RECT 323.515 -123.245 323.845 -122.915 ;
        RECT 323.515 -124.605 323.845 -124.275 ;
        RECT 323.515 -125.965 323.845 -125.635 ;
        RECT 323.515 -127.325 323.845 -126.995 ;
        RECT 323.515 -128.685 323.845 -128.355 ;
        RECT 323.515 -130.045 323.845 -129.715 ;
        RECT 323.515 -131.405 323.845 -131.075 ;
        RECT 323.515 -132.765 323.845 -132.435 ;
        RECT 323.515 -134.125 323.845 -133.795 ;
        RECT 323.515 -135.485 323.845 -135.155 ;
        RECT 323.515 -136.845 323.845 -136.515 ;
        RECT 323.515 -138.205 323.845 -137.875 ;
        RECT 323.515 -139.565 323.845 -139.235 ;
        RECT 323.515 -140.925 323.845 -140.595 ;
        RECT 323.515 -142.285 323.845 -141.955 ;
        RECT 323.515 -143.645 323.845 -143.315 ;
        RECT 323.515 -145.005 323.845 -144.675 ;
        RECT 323.515 -146.365 323.845 -146.035 ;
        RECT 323.515 -147.725 323.845 -147.395 ;
        RECT 323.515 -149.085 323.845 -148.755 ;
        RECT 323.515 -150.445 323.845 -150.115 ;
        RECT 323.515 -151.805 323.845 -151.475 ;
        RECT 323.515 -153.165 323.845 -152.835 ;
        RECT 323.515 -154.525 323.845 -154.195 ;
        RECT 323.515 -155.885 323.845 -155.555 ;
        RECT 323.515 -157.245 323.845 -156.915 ;
        RECT 323.515 -158.605 323.845 -158.275 ;
        RECT 323.515 -159.965 323.845 -159.635 ;
        RECT 323.515 -161.325 323.845 -160.995 ;
        RECT 323.515 -162.685 323.845 -162.355 ;
        RECT 323.515 -164.045 323.845 -163.715 ;
        RECT 323.515 -165.405 323.845 -165.075 ;
        RECT 323.515 -166.765 323.845 -166.435 ;
        RECT 323.515 -168.125 323.845 -167.795 ;
        RECT 323.515 -169.485 323.845 -169.155 ;
        RECT 323.515 -170.845 323.845 -170.515 ;
        RECT 323.515 -172.205 323.845 -171.875 ;
        RECT 323.515 -173.565 323.845 -173.235 ;
        RECT 323.515 -174.925 323.845 -174.595 ;
        RECT 323.515 -176.285 323.845 -175.955 ;
        RECT 323.515 -177.645 323.845 -177.315 ;
        RECT 323.515 -179.005 323.845 -178.675 ;
        RECT 323.515 -184.65 323.845 -183.52 ;
        RECT 323.52 -184.765 323.84 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.875 244.04 325.205 245.17 ;
        RECT 324.875 239.875 325.205 240.205 ;
        RECT 324.875 238.515 325.205 238.845 ;
        RECT 324.875 237.155 325.205 237.485 ;
        RECT 324.88 237.155 325.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.875 -0.845 325.205 -0.515 ;
        RECT 324.875 -2.205 325.205 -1.875 ;
        RECT 324.875 -3.565 325.205 -3.235 ;
        RECT 324.88 -3.565 325.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.875 -96.045 325.205 -95.715 ;
        RECT 324.875 -97.405 325.205 -97.075 ;
        RECT 324.875 -98.765 325.205 -98.435 ;
        RECT 324.875 -100.125 325.205 -99.795 ;
        RECT 324.875 -101.485 325.205 -101.155 ;
        RECT 324.875 -102.845 325.205 -102.515 ;
        RECT 324.875 -104.205 325.205 -103.875 ;
        RECT 324.875 -105.565 325.205 -105.235 ;
        RECT 324.875 -106.925 325.205 -106.595 ;
        RECT 324.875 -108.285 325.205 -107.955 ;
        RECT 324.875 -109.645 325.205 -109.315 ;
        RECT 324.875 -111.005 325.205 -110.675 ;
        RECT 324.875 -112.365 325.205 -112.035 ;
        RECT 324.875 -113.725 325.205 -113.395 ;
        RECT 324.875 -115.085 325.205 -114.755 ;
        RECT 324.875 -116.445 325.205 -116.115 ;
        RECT 324.875 -117.805 325.205 -117.475 ;
        RECT 324.875 -119.165 325.205 -118.835 ;
        RECT 324.875 -120.525 325.205 -120.195 ;
        RECT 324.875 -121.885 325.205 -121.555 ;
        RECT 324.875 -123.245 325.205 -122.915 ;
        RECT 324.875 -124.605 325.205 -124.275 ;
        RECT 324.875 -125.965 325.205 -125.635 ;
        RECT 324.875 -127.325 325.205 -126.995 ;
        RECT 324.875 -128.685 325.205 -128.355 ;
        RECT 324.875 -130.045 325.205 -129.715 ;
        RECT 324.875 -131.405 325.205 -131.075 ;
        RECT 324.875 -132.765 325.205 -132.435 ;
        RECT 324.875 -134.125 325.205 -133.795 ;
        RECT 324.875 -135.485 325.205 -135.155 ;
        RECT 324.875 -136.845 325.205 -136.515 ;
        RECT 324.875 -138.205 325.205 -137.875 ;
        RECT 324.875 -139.565 325.205 -139.235 ;
        RECT 324.875 -140.925 325.205 -140.595 ;
        RECT 324.875 -142.285 325.205 -141.955 ;
        RECT 324.875 -143.645 325.205 -143.315 ;
        RECT 324.875 -145.005 325.205 -144.675 ;
        RECT 324.875 -146.365 325.205 -146.035 ;
        RECT 324.875 -147.725 325.205 -147.395 ;
        RECT 324.875 -149.085 325.205 -148.755 ;
        RECT 324.875 -150.445 325.205 -150.115 ;
        RECT 324.875 -151.805 325.205 -151.475 ;
        RECT 324.875 -153.165 325.205 -152.835 ;
        RECT 324.875 -154.525 325.205 -154.195 ;
        RECT 324.875 -155.885 325.205 -155.555 ;
        RECT 324.875 -157.245 325.205 -156.915 ;
        RECT 324.875 -158.605 325.205 -158.275 ;
        RECT 324.875 -159.965 325.205 -159.635 ;
        RECT 324.875 -161.325 325.205 -160.995 ;
        RECT 324.875 -162.685 325.205 -162.355 ;
        RECT 324.875 -164.045 325.205 -163.715 ;
        RECT 324.875 -165.405 325.205 -165.075 ;
        RECT 324.875 -166.765 325.205 -166.435 ;
        RECT 324.875 -168.125 325.205 -167.795 ;
        RECT 324.875 -169.485 325.205 -169.155 ;
        RECT 324.875 -170.845 325.205 -170.515 ;
        RECT 324.875 -172.205 325.205 -171.875 ;
        RECT 324.875 -173.565 325.205 -173.235 ;
        RECT 324.875 -174.925 325.205 -174.595 ;
        RECT 324.875 -176.285 325.205 -175.955 ;
        RECT 324.875 -177.645 325.205 -177.315 ;
        RECT 324.875 -179.005 325.205 -178.675 ;
        RECT 324.875 -184.65 325.205 -183.52 ;
        RECT 324.88 -184.765 325.2 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.235 244.04 326.565 245.17 ;
        RECT 326.235 239.875 326.565 240.205 ;
        RECT 326.235 238.515 326.565 238.845 ;
        RECT 326.235 237.155 326.565 237.485 ;
        RECT 326.24 237.155 326.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.235 -0.845 326.565 -0.515 ;
        RECT 326.235 -2.205 326.565 -1.875 ;
        RECT 326.235 -3.565 326.565 -3.235 ;
        RECT 326.24 -3.565 326.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.235 -96.045 326.565 -95.715 ;
        RECT 326.235 -97.405 326.565 -97.075 ;
        RECT 326.235 -98.765 326.565 -98.435 ;
        RECT 326.235 -100.125 326.565 -99.795 ;
        RECT 326.235 -101.485 326.565 -101.155 ;
        RECT 326.235 -102.845 326.565 -102.515 ;
        RECT 326.235 -104.205 326.565 -103.875 ;
        RECT 326.235 -105.565 326.565 -105.235 ;
        RECT 326.235 -106.925 326.565 -106.595 ;
        RECT 326.235 -108.285 326.565 -107.955 ;
        RECT 326.235 -109.645 326.565 -109.315 ;
        RECT 326.235 -111.005 326.565 -110.675 ;
        RECT 326.235 -112.365 326.565 -112.035 ;
        RECT 326.235 -113.725 326.565 -113.395 ;
        RECT 326.235 -115.085 326.565 -114.755 ;
        RECT 326.235 -116.445 326.565 -116.115 ;
        RECT 326.235 -117.805 326.565 -117.475 ;
        RECT 326.235 -119.165 326.565 -118.835 ;
        RECT 326.235 -120.525 326.565 -120.195 ;
        RECT 326.235 -121.885 326.565 -121.555 ;
        RECT 326.235 -123.245 326.565 -122.915 ;
        RECT 326.235 -124.605 326.565 -124.275 ;
        RECT 326.235 -125.965 326.565 -125.635 ;
        RECT 326.235 -127.325 326.565 -126.995 ;
        RECT 326.235 -128.685 326.565 -128.355 ;
        RECT 326.235 -130.045 326.565 -129.715 ;
        RECT 326.235 -131.405 326.565 -131.075 ;
        RECT 326.235 -132.765 326.565 -132.435 ;
        RECT 326.235 -134.125 326.565 -133.795 ;
        RECT 326.235 -135.485 326.565 -135.155 ;
        RECT 326.235 -136.845 326.565 -136.515 ;
        RECT 326.235 -138.205 326.565 -137.875 ;
        RECT 326.235 -139.565 326.565 -139.235 ;
        RECT 326.235 -140.925 326.565 -140.595 ;
        RECT 326.235 -142.285 326.565 -141.955 ;
        RECT 326.235 -143.645 326.565 -143.315 ;
        RECT 326.235 -145.005 326.565 -144.675 ;
        RECT 326.235 -146.365 326.565 -146.035 ;
        RECT 326.235 -147.725 326.565 -147.395 ;
        RECT 326.235 -149.085 326.565 -148.755 ;
        RECT 326.235 -150.445 326.565 -150.115 ;
        RECT 326.235 -151.805 326.565 -151.475 ;
        RECT 326.235 -153.165 326.565 -152.835 ;
        RECT 326.235 -154.525 326.565 -154.195 ;
        RECT 326.235 -155.885 326.565 -155.555 ;
        RECT 326.235 -157.245 326.565 -156.915 ;
        RECT 326.235 -158.605 326.565 -158.275 ;
        RECT 326.235 -159.965 326.565 -159.635 ;
        RECT 326.235 -161.325 326.565 -160.995 ;
        RECT 326.235 -162.685 326.565 -162.355 ;
        RECT 326.235 -164.045 326.565 -163.715 ;
        RECT 326.235 -165.405 326.565 -165.075 ;
        RECT 326.235 -166.765 326.565 -166.435 ;
        RECT 326.235 -168.125 326.565 -167.795 ;
        RECT 326.235 -169.485 326.565 -169.155 ;
        RECT 326.235 -170.845 326.565 -170.515 ;
        RECT 326.235 -172.205 326.565 -171.875 ;
        RECT 326.235 -173.565 326.565 -173.235 ;
        RECT 326.235 -174.925 326.565 -174.595 ;
        RECT 326.235 -176.285 326.565 -175.955 ;
        RECT 326.235 -177.645 326.565 -177.315 ;
        RECT 326.235 -179.005 326.565 -178.675 ;
        RECT 326.235 -184.65 326.565 -183.52 ;
        RECT 326.24 -184.765 326.56 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.595 244.04 327.925 245.17 ;
        RECT 327.595 239.875 327.925 240.205 ;
        RECT 327.595 238.515 327.925 238.845 ;
        RECT 327.595 237.155 327.925 237.485 ;
        RECT 327.6 237.155 327.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.595 -0.845 327.925 -0.515 ;
        RECT 327.595 -2.205 327.925 -1.875 ;
        RECT 327.595 -3.565 327.925 -3.235 ;
        RECT 327.6 -3.565 327.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 327.595 -96.045 327.925 -95.715 ;
        RECT 327.595 -97.405 327.925 -97.075 ;
        RECT 327.595 -98.765 327.925 -98.435 ;
        RECT 327.595 -100.125 327.925 -99.795 ;
        RECT 327.595 -101.485 327.925 -101.155 ;
        RECT 327.595 -102.845 327.925 -102.515 ;
        RECT 327.595 -104.205 327.925 -103.875 ;
        RECT 327.595 -105.565 327.925 -105.235 ;
        RECT 327.595 -106.925 327.925 -106.595 ;
        RECT 327.595 -108.285 327.925 -107.955 ;
        RECT 327.595 -109.645 327.925 -109.315 ;
        RECT 327.595 -111.005 327.925 -110.675 ;
        RECT 327.595 -112.365 327.925 -112.035 ;
        RECT 327.595 -113.725 327.925 -113.395 ;
        RECT 327.595 -115.085 327.925 -114.755 ;
        RECT 327.595 -116.445 327.925 -116.115 ;
        RECT 327.595 -117.805 327.925 -117.475 ;
        RECT 327.595 -119.165 327.925 -118.835 ;
        RECT 327.595 -120.525 327.925 -120.195 ;
        RECT 327.595 -121.885 327.925 -121.555 ;
        RECT 327.595 -123.245 327.925 -122.915 ;
        RECT 327.595 -124.605 327.925 -124.275 ;
        RECT 327.595 -125.965 327.925 -125.635 ;
        RECT 327.595 -127.325 327.925 -126.995 ;
        RECT 327.595 -128.685 327.925 -128.355 ;
        RECT 327.595 -130.045 327.925 -129.715 ;
        RECT 327.595 -131.405 327.925 -131.075 ;
        RECT 327.595 -132.765 327.925 -132.435 ;
        RECT 327.595 -134.125 327.925 -133.795 ;
        RECT 327.595 -135.485 327.925 -135.155 ;
        RECT 327.595 -136.845 327.925 -136.515 ;
        RECT 327.595 -138.205 327.925 -137.875 ;
        RECT 327.595 -139.565 327.925 -139.235 ;
        RECT 327.595 -140.925 327.925 -140.595 ;
        RECT 327.595 -142.285 327.925 -141.955 ;
        RECT 327.595 -143.645 327.925 -143.315 ;
        RECT 327.595 -145.005 327.925 -144.675 ;
        RECT 327.595 -146.365 327.925 -146.035 ;
        RECT 327.595 -147.725 327.925 -147.395 ;
        RECT 327.595 -149.085 327.925 -148.755 ;
        RECT 327.595 -150.445 327.925 -150.115 ;
        RECT 327.595 -151.805 327.925 -151.475 ;
        RECT 327.595 -153.165 327.925 -152.835 ;
        RECT 327.595 -154.525 327.925 -154.195 ;
        RECT 327.595 -155.885 327.925 -155.555 ;
        RECT 327.595 -157.245 327.925 -156.915 ;
        RECT 327.595 -158.605 327.925 -158.275 ;
        RECT 327.595 -159.965 327.925 -159.635 ;
        RECT 327.595 -161.325 327.925 -160.995 ;
        RECT 327.595 -162.685 327.925 -162.355 ;
        RECT 327.595 -164.045 327.925 -163.715 ;
        RECT 327.595 -165.405 327.925 -165.075 ;
        RECT 327.595 -166.765 327.925 -166.435 ;
        RECT 327.595 -168.125 327.925 -167.795 ;
        RECT 327.595 -169.485 327.925 -169.155 ;
        RECT 327.595 -170.845 327.925 -170.515 ;
        RECT 327.595 -172.205 327.925 -171.875 ;
        RECT 327.595 -173.565 327.925 -173.235 ;
        RECT 327.595 -174.925 327.925 -174.595 ;
        RECT 327.595 -176.285 327.925 -175.955 ;
        RECT 327.595 -177.645 327.925 -177.315 ;
        RECT 327.595 -179.005 327.925 -178.675 ;
        RECT 327.595 -184.65 327.925 -183.52 ;
        RECT 327.6 -184.765 327.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.955 244.04 329.285 245.17 ;
        RECT 328.955 239.875 329.285 240.205 ;
        RECT 328.955 238.515 329.285 238.845 ;
        RECT 328.955 237.155 329.285 237.485 ;
        RECT 328.96 237.155 329.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.955 -0.845 329.285 -0.515 ;
        RECT 328.955 -2.205 329.285 -1.875 ;
        RECT 328.955 -3.565 329.285 -3.235 ;
        RECT 328.96 -3.565 329.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.955 -96.045 329.285 -95.715 ;
        RECT 328.955 -97.405 329.285 -97.075 ;
        RECT 328.955 -98.765 329.285 -98.435 ;
        RECT 328.955 -100.125 329.285 -99.795 ;
        RECT 328.955 -101.485 329.285 -101.155 ;
        RECT 328.955 -102.845 329.285 -102.515 ;
        RECT 328.955 -104.205 329.285 -103.875 ;
        RECT 328.955 -105.565 329.285 -105.235 ;
        RECT 328.955 -106.925 329.285 -106.595 ;
        RECT 328.955 -108.285 329.285 -107.955 ;
        RECT 328.955 -109.645 329.285 -109.315 ;
        RECT 328.955 -111.005 329.285 -110.675 ;
        RECT 328.955 -112.365 329.285 -112.035 ;
        RECT 328.955 -113.725 329.285 -113.395 ;
        RECT 328.955 -115.085 329.285 -114.755 ;
        RECT 328.955 -116.445 329.285 -116.115 ;
        RECT 328.955 -117.805 329.285 -117.475 ;
        RECT 328.955 -119.165 329.285 -118.835 ;
        RECT 328.955 -120.525 329.285 -120.195 ;
        RECT 328.955 -121.885 329.285 -121.555 ;
        RECT 328.955 -123.245 329.285 -122.915 ;
        RECT 328.955 -124.605 329.285 -124.275 ;
        RECT 328.955 -125.965 329.285 -125.635 ;
        RECT 328.955 -127.325 329.285 -126.995 ;
        RECT 328.955 -128.685 329.285 -128.355 ;
        RECT 328.955 -130.045 329.285 -129.715 ;
        RECT 328.955 -131.405 329.285 -131.075 ;
        RECT 328.955 -132.765 329.285 -132.435 ;
        RECT 328.955 -134.125 329.285 -133.795 ;
        RECT 328.955 -135.485 329.285 -135.155 ;
        RECT 328.955 -136.845 329.285 -136.515 ;
        RECT 328.955 -138.205 329.285 -137.875 ;
        RECT 328.955 -139.565 329.285 -139.235 ;
        RECT 328.955 -140.925 329.285 -140.595 ;
        RECT 328.955 -142.285 329.285 -141.955 ;
        RECT 328.955 -143.645 329.285 -143.315 ;
        RECT 328.955 -145.005 329.285 -144.675 ;
        RECT 328.955 -146.365 329.285 -146.035 ;
        RECT 328.955 -147.725 329.285 -147.395 ;
        RECT 328.955 -149.085 329.285 -148.755 ;
        RECT 328.955 -150.445 329.285 -150.115 ;
        RECT 328.955 -151.805 329.285 -151.475 ;
        RECT 328.955 -153.165 329.285 -152.835 ;
        RECT 328.955 -154.525 329.285 -154.195 ;
        RECT 328.955 -155.885 329.285 -155.555 ;
        RECT 328.955 -157.245 329.285 -156.915 ;
        RECT 328.955 -158.605 329.285 -158.275 ;
        RECT 328.955 -159.965 329.285 -159.635 ;
        RECT 328.955 -161.325 329.285 -160.995 ;
        RECT 328.955 -162.685 329.285 -162.355 ;
        RECT 328.955 -164.045 329.285 -163.715 ;
        RECT 328.955 -165.405 329.285 -165.075 ;
        RECT 328.955 -166.765 329.285 -166.435 ;
        RECT 328.955 -168.125 329.285 -167.795 ;
        RECT 328.955 -169.485 329.285 -169.155 ;
        RECT 328.955 -170.845 329.285 -170.515 ;
        RECT 328.955 -172.205 329.285 -171.875 ;
        RECT 328.955 -173.565 329.285 -173.235 ;
        RECT 328.955 -174.925 329.285 -174.595 ;
        RECT 328.955 -176.285 329.285 -175.955 ;
        RECT 328.955 -177.645 329.285 -177.315 ;
        RECT 328.955 -179.005 329.285 -178.675 ;
        RECT 328.955 -184.65 329.285 -183.52 ;
        RECT 328.96 -184.765 329.28 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.66 -98.075 329.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.315 244.04 330.645 245.17 ;
        RECT 330.315 239.875 330.645 240.205 ;
        RECT 330.315 238.515 330.645 238.845 ;
        RECT 330.315 237.155 330.645 237.485 ;
        RECT 330.32 237.155 330.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.315 -98.765 330.645 -98.435 ;
        RECT 330.315 -100.125 330.645 -99.795 ;
        RECT 330.315 -101.485 330.645 -101.155 ;
        RECT 330.315 -102.845 330.645 -102.515 ;
        RECT 330.315 -104.205 330.645 -103.875 ;
        RECT 330.315 -105.565 330.645 -105.235 ;
        RECT 330.315 -106.925 330.645 -106.595 ;
        RECT 330.315 -108.285 330.645 -107.955 ;
        RECT 330.315 -109.645 330.645 -109.315 ;
        RECT 330.315 -111.005 330.645 -110.675 ;
        RECT 330.315 -112.365 330.645 -112.035 ;
        RECT 330.315 -113.725 330.645 -113.395 ;
        RECT 330.315 -115.085 330.645 -114.755 ;
        RECT 330.315 -116.445 330.645 -116.115 ;
        RECT 330.315 -117.805 330.645 -117.475 ;
        RECT 330.315 -119.165 330.645 -118.835 ;
        RECT 330.315 -120.525 330.645 -120.195 ;
        RECT 330.315 -121.885 330.645 -121.555 ;
        RECT 330.315 -123.245 330.645 -122.915 ;
        RECT 330.315 -124.605 330.645 -124.275 ;
        RECT 330.315 -125.965 330.645 -125.635 ;
        RECT 330.315 -127.325 330.645 -126.995 ;
        RECT 330.315 -128.685 330.645 -128.355 ;
        RECT 330.315 -130.045 330.645 -129.715 ;
        RECT 330.315 -131.405 330.645 -131.075 ;
        RECT 330.315 -132.765 330.645 -132.435 ;
        RECT 330.315 -134.125 330.645 -133.795 ;
        RECT 330.315 -135.485 330.645 -135.155 ;
        RECT 330.315 -136.845 330.645 -136.515 ;
        RECT 330.315 -138.205 330.645 -137.875 ;
        RECT 330.315 -139.565 330.645 -139.235 ;
        RECT 330.315 -140.925 330.645 -140.595 ;
        RECT 330.315 -142.285 330.645 -141.955 ;
        RECT 330.315 -143.645 330.645 -143.315 ;
        RECT 330.315 -145.005 330.645 -144.675 ;
        RECT 330.315 -146.365 330.645 -146.035 ;
        RECT 330.315 -147.725 330.645 -147.395 ;
        RECT 330.315 -149.085 330.645 -148.755 ;
        RECT 330.315 -150.445 330.645 -150.115 ;
        RECT 330.315 -151.805 330.645 -151.475 ;
        RECT 330.315 -153.165 330.645 -152.835 ;
        RECT 330.315 -154.525 330.645 -154.195 ;
        RECT 330.315 -155.885 330.645 -155.555 ;
        RECT 330.315 -157.245 330.645 -156.915 ;
        RECT 330.315 -158.605 330.645 -158.275 ;
        RECT 330.315 -159.965 330.645 -159.635 ;
        RECT 330.315 -161.325 330.645 -160.995 ;
        RECT 330.315 -162.685 330.645 -162.355 ;
        RECT 330.315 -164.045 330.645 -163.715 ;
        RECT 330.315 -165.405 330.645 -165.075 ;
        RECT 330.315 -166.765 330.645 -166.435 ;
        RECT 330.315 -168.125 330.645 -167.795 ;
        RECT 330.315 -169.485 330.645 -169.155 ;
        RECT 330.315 -170.845 330.645 -170.515 ;
        RECT 330.315 -172.205 330.645 -171.875 ;
        RECT 330.315 -173.565 330.645 -173.235 ;
        RECT 330.315 -174.925 330.645 -174.595 ;
        RECT 330.315 -176.285 330.645 -175.955 ;
        RECT 330.315 -177.645 330.645 -177.315 ;
        RECT 330.315 -179.005 330.645 -178.675 ;
        RECT 330.315 -184.65 330.645 -183.52 ;
        RECT 330.32 -184.765 330.64 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.675 244.04 332.005 245.17 ;
        RECT 331.675 239.875 332.005 240.205 ;
        RECT 331.675 238.515 332.005 238.845 ;
        RECT 331.675 237.155 332.005 237.485 ;
        RECT 331.68 237.155 332 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 331.675 -0.845 332.005 -0.515 ;
        RECT 331.675 -2.205 332.005 -1.875 ;
        RECT 331.675 -3.565 332.005 -3.235 ;
        RECT 331.68 -3.565 332 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.035 244.04 333.365 245.17 ;
        RECT 333.035 239.875 333.365 240.205 ;
        RECT 333.035 238.515 333.365 238.845 ;
        RECT 333.035 237.155 333.365 237.485 ;
        RECT 333.04 237.155 333.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.035 -0.845 333.365 -0.515 ;
        RECT 333.035 -2.205 333.365 -1.875 ;
        RECT 333.035 -3.565 333.365 -3.235 ;
        RECT 333.04 -3.565 333.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.395 244.04 334.725 245.17 ;
        RECT 334.395 239.875 334.725 240.205 ;
        RECT 334.395 238.515 334.725 238.845 ;
        RECT 334.395 237.155 334.725 237.485 ;
        RECT 334.4 237.155 334.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.395 -0.845 334.725 -0.515 ;
        RECT 334.395 -2.205 334.725 -1.875 ;
        RECT 334.395 -3.565 334.725 -3.235 ;
        RECT 334.4 -3.565 334.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 334.395 -96.045 334.725 -95.715 ;
        RECT 334.395 -97.405 334.725 -97.075 ;
        RECT 334.395 -98.765 334.725 -98.435 ;
        RECT 334.395 -100.125 334.725 -99.795 ;
        RECT 334.395 -101.485 334.725 -101.155 ;
        RECT 334.395 -102.845 334.725 -102.515 ;
        RECT 334.395 -104.205 334.725 -103.875 ;
        RECT 334.395 -105.565 334.725 -105.235 ;
        RECT 334.395 -106.925 334.725 -106.595 ;
        RECT 334.395 -108.285 334.725 -107.955 ;
        RECT 334.395 -109.645 334.725 -109.315 ;
        RECT 334.395 -111.005 334.725 -110.675 ;
        RECT 334.395 -112.365 334.725 -112.035 ;
        RECT 334.395 -113.725 334.725 -113.395 ;
        RECT 334.395 -115.085 334.725 -114.755 ;
        RECT 334.395 -116.445 334.725 -116.115 ;
        RECT 334.395 -117.805 334.725 -117.475 ;
        RECT 334.395 -119.165 334.725 -118.835 ;
        RECT 334.395 -120.525 334.725 -120.195 ;
        RECT 334.395 -121.885 334.725 -121.555 ;
        RECT 334.395 -123.245 334.725 -122.915 ;
        RECT 334.395 -124.605 334.725 -124.275 ;
        RECT 334.395 -125.965 334.725 -125.635 ;
        RECT 334.395 -127.325 334.725 -126.995 ;
        RECT 334.395 -128.685 334.725 -128.355 ;
        RECT 334.395 -130.045 334.725 -129.715 ;
        RECT 334.395 -131.405 334.725 -131.075 ;
        RECT 334.395 -132.765 334.725 -132.435 ;
        RECT 334.395 -134.125 334.725 -133.795 ;
        RECT 334.395 -135.485 334.725 -135.155 ;
        RECT 334.395 -136.845 334.725 -136.515 ;
        RECT 334.395 -138.205 334.725 -137.875 ;
        RECT 334.395 -139.565 334.725 -139.235 ;
        RECT 334.395 -140.925 334.725 -140.595 ;
        RECT 334.395 -142.285 334.725 -141.955 ;
        RECT 334.395 -143.645 334.725 -143.315 ;
        RECT 334.395 -145.005 334.725 -144.675 ;
        RECT 334.395 -146.365 334.725 -146.035 ;
        RECT 334.395 -147.725 334.725 -147.395 ;
        RECT 334.395 -149.085 334.725 -148.755 ;
        RECT 334.395 -150.445 334.725 -150.115 ;
        RECT 334.395 -151.805 334.725 -151.475 ;
        RECT 334.395 -153.165 334.725 -152.835 ;
        RECT 334.395 -154.525 334.725 -154.195 ;
        RECT 334.395 -155.885 334.725 -155.555 ;
        RECT 334.395 -157.245 334.725 -156.915 ;
        RECT 334.395 -158.605 334.725 -158.275 ;
        RECT 334.395 -159.965 334.725 -159.635 ;
        RECT 334.395 -161.325 334.725 -160.995 ;
        RECT 334.395 -162.685 334.725 -162.355 ;
        RECT 334.395 -164.045 334.725 -163.715 ;
        RECT 334.395 -165.405 334.725 -165.075 ;
        RECT 334.395 -166.765 334.725 -166.435 ;
        RECT 334.395 -168.125 334.725 -167.795 ;
        RECT 334.395 -169.485 334.725 -169.155 ;
        RECT 334.395 -170.845 334.725 -170.515 ;
        RECT 334.395 -172.205 334.725 -171.875 ;
        RECT 334.395 -173.565 334.725 -173.235 ;
        RECT 334.395 -174.925 334.725 -174.595 ;
        RECT 334.395 -176.285 334.725 -175.955 ;
        RECT 334.395 -177.645 334.725 -177.315 ;
        RECT 334.395 -179.005 334.725 -178.675 ;
        RECT 334.395 -184.65 334.725 -183.52 ;
        RECT 334.4 -184.765 334.72 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.755 244.04 336.085 245.17 ;
        RECT 335.755 239.875 336.085 240.205 ;
        RECT 335.755 238.515 336.085 238.845 ;
        RECT 335.755 237.155 336.085 237.485 ;
        RECT 335.76 237.155 336.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.755 -0.845 336.085 -0.515 ;
        RECT 335.755 -2.205 336.085 -1.875 ;
        RECT 335.755 -3.565 336.085 -3.235 ;
        RECT 335.76 -3.565 336.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.755 -96.045 336.085 -95.715 ;
        RECT 335.755 -97.405 336.085 -97.075 ;
        RECT 335.755 -98.765 336.085 -98.435 ;
        RECT 335.755 -100.125 336.085 -99.795 ;
        RECT 335.755 -101.485 336.085 -101.155 ;
        RECT 335.755 -102.845 336.085 -102.515 ;
        RECT 335.755 -104.205 336.085 -103.875 ;
        RECT 335.755 -105.565 336.085 -105.235 ;
        RECT 335.755 -106.925 336.085 -106.595 ;
        RECT 335.755 -108.285 336.085 -107.955 ;
        RECT 335.755 -109.645 336.085 -109.315 ;
        RECT 335.755 -111.005 336.085 -110.675 ;
        RECT 335.755 -112.365 336.085 -112.035 ;
        RECT 335.755 -113.725 336.085 -113.395 ;
        RECT 335.755 -115.085 336.085 -114.755 ;
        RECT 335.755 -116.445 336.085 -116.115 ;
        RECT 335.755 -117.805 336.085 -117.475 ;
        RECT 335.755 -119.165 336.085 -118.835 ;
        RECT 335.755 -120.525 336.085 -120.195 ;
        RECT 335.755 -121.885 336.085 -121.555 ;
        RECT 335.755 -123.245 336.085 -122.915 ;
        RECT 335.755 -124.605 336.085 -124.275 ;
        RECT 335.755 -125.965 336.085 -125.635 ;
        RECT 335.755 -127.325 336.085 -126.995 ;
        RECT 335.755 -128.685 336.085 -128.355 ;
        RECT 335.755 -130.045 336.085 -129.715 ;
        RECT 335.755 -131.405 336.085 -131.075 ;
        RECT 335.755 -132.765 336.085 -132.435 ;
        RECT 335.755 -134.125 336.085 -133.795 ;
        RECT 335.755 -135.485 336.085 -135.155 ;
        RECT 335.755 -136.845 336.085 -136.515 ;
        RECT 335.755 -138.205 336.085 -137.875 ;
        RECT 335.755 -139.565 336.085 -139.235 ;
        RECT 335.755 -140.925 336.085 -140.595 ;
        RECT 335.755 -142.285 336.085 -141.955 ;
        RECT 335.755 -143.645 336.085 -143.315 ;
        RECT 335.755 -145.005 336.085 -144.675 ;
        RECT 335.755 -146.365 336.085 -146.035 ;
        RECT 335.755 -147.725 336.085 -147.395 ;
        RECT 335.755 -149.085 336.085 -148.755 ;
        RECT 335.755 -150.445 336.085 -150.115 ;
        RECT 335.755 -151.805 336.085 -151.475 ;
        RECT 335.755 -153.165 336.085 -152.835 ;
        RECT 335.755 -154.525 336.085 -154.195 ;
        RECT 335.755 -155.885 336.085 -155.555 ;
        RECT 335.755 -157.245 336.085 -156.915 ;
        RECT 335.755 -158.605 336.085 -158.275 ;
        RECT 335.755 -159.965 336.085 -159.635 ;
        RECT 335.755 -161.325 336.085 -160.995 ;
        RECT 335.755 -162.685 336.085 -162.355 ;
        RECT 335.755 -164.045 336.085 -163.715 ;
        RECT 335.755 -165.405 336.085 -165.075 ;
        RECT 335.755 -166.765 336.085 -166.435 ;
        RECT 335.755 -168.125 336.085 -167.795 ;
        RECT 335.755 -169.485 336.085 -169.155 ;
        RECT 335.755 -170.845 336.085 -170.515 ;
        RECT 335.755 -172.205 336.085 -171.875 ;
        RECT 335.755 -173.565 336.085 -173.235 ;
        RECT 335.755 -174.925 336.085 -174.595 ;
        RECT 335.755 -176.285 336.085 -175.955 ;
        RECT 335.755 -177.645 336.085 -177.315 ;
        RECT 335.755 -179.005 336.085 -178.675 ;
        RECT 335.755 -184.65 336.085 -183.52 ;
        RECT 335.76 -184.765 336.08 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.115 244.04 337.445 245.17 ;
        RECT 337.115 239.875 337.445 240.205 ;
        RECT 337.115 238.515 337.445 238.845 ;
        RECT 337.115 237.155 337.445 237.485 ;
        RECT 337.12 237.155 337.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.115 -0.845 337.445 -0.515 ;
        RECT 337.115 -2.205 337.445 -1.875 ;
        RECT 337.115 -3.565 337.445 -3.235 ;
        RECT 337.12 -3.565 337.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.115 -151.805 337.445 -151.475 ;
        RECT 337.115 -153.165 337.445 -152.835 ;
        RECT 337.115 -154.525 337.445 -154.195 ;
        RECT 337.115 -155.885 337.445 -155.555 ;
        RECT 337.115 -157.245 337.445 -156.915 ;
        RECT 337.115 -158.605 337.445 -158.275 ;
        RECT 337.115 -159.965 337.445 -159.635 ;
        RECT 337.115 -161.325 337.445 -160.995 ;
        RECT 337.115 -162.685 337.445 -162.355 ;
        RECT 337.115 -164.045 337.445 -163.715 ;
        RECT 337.115 -165.405 337.445 -165.075 ;
        RECT 337.115 -166.765 337.445 -166.435 ;
        RECT 337.115 -168.125 337.445 -167.795 ;
        RECT 337.115 -169.485 337.445 -169.155 ;
        RECT 337.115 -170.845 337.445 -170.515 ;
        RECT 337.115 -172.205 337.445 -171.875 ;
        RECT 337.115 -173.565 337.445 -173.235 ;
        RECT 337.115 -174.925 337.445 -174.595 ;
        RECT 337.115 -176.285 337.445 -175.955 ;
        RECT 337.115 -177.645 337.445 -177.315 ;
        RECT 337.115 -179.005 337.445 -178.675 ;
        RECT 337.115 -184.65 337.445 -183.52 ;
        RECT 337.12 -184.765 337.44 -95.04 ;
        RECT 337.115 -96.045 337.445 -95.715 ;
        RECT 337.115 -97.405 337.445 -97.075 ;
        RECT 337.115 -98.765 337.445 -98.435 ;
        RECT 337.115 -100.125 337.445 -99.795 ;
        RECT 337.115 -101.485 337.445 -101.155 ;
        RECT 337.115 -102.845 337.445 -102.515 ;
        RECT 337.115 -104.205 337.445 -103.875 ;
        RECT 337.115 -105.565 337.445 -105.235 ;
        RECT 337.115 -106.925 337.445 -106.595 ;
        RECT 337.115 -108.285 337.445 -107.955 ;
        RECT 337.115 -109.645 337.445 -109.315 ;
        RECT 337.115 -111.005 337.445 -110.675 ;
        RECT 337.115 -112.365 337.445 -112.035 ;
        RECT 337.115 -113.725 337.445 -113.395 ;
        RECT 337.115 -115.085 337.445 -114.755 ;
        RECT 337.115 -116.445 337.445 -116.115 ;
        RECT 337.115 -117.805 337.445 -117.475 ;
        RECT 337.115 -119.165 337.445 -118.835 ;
        RECT 337.115 -120.525 337.445 -120.195 ;
        RECT 337.115 -121.885 337.445 -121.555 ;
        RECT 337.115 -123.245 337.445 -122.915 ;
        RECT 337.115 -124.605 337.445 -124.275 ;
        RECT 337.115 -125.965 337.445 -125.635 ;
        RECT 337.115 -127.325 337.445 -126.995 ;
        RECT 337.115 -128.685 337.445 -128.355 ;
        RECT 337.115 -130.045 337.445 -129.715 ;
        RECT 337.115 -131.405 337.445 -131.075 ;
        RECT 337.115 -132.765 337.445 -132.435 ;
        RECT 337.115 -134.125 337.445 -133.795 ;
        RECT 337.115 -135.485 337.445 -135.155 ;
        RECT 337.115 -136.845 337.445 -136.515 ;
        RECT 337.115 -138.205 337.445 -137.875 ;
        RECT 337.115 -139.565 337.445 -139.235 ;
        RECT 337.115 -140.925 337.445 -140.595 ;
        RECT 337.115 -142.285 337.445 -141.955 ;
        RECT 337.115 -143.645 337.445 -143.315 ;
        RECT 337.115 -145.005 337.445 -144.675 ;
        RECT 337.115 -146.365 337.445 -146.035 ;
        RECT 337.115 -147.725 337.445 -147.395 ;
        RECT 337.115 -149.085 337.445 -148.755 ;
        RECT 337.115 -150.445 337.445 -150.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.435 244.04 285.765 245.17 ;
        RECT 285.435 239.875 285.765 240.205 ;
        RECT 285.435 238.515 285.765 238.845 ;
        RECT 285.435 237.155 285.765 237.485 ;
        RECT 285.44 237.155 285.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 285.435 -98.765 285.765 -98.435 ;
        RECT 285.435 -100.125 285.765 -99.795 ;
        RECT 285.435 -101.485 285.765 -101.155 ;
        RECT 285.435 -102.845 285.765 -102.515 ;
        RECT 285.435 -104.205 285.765 -103.875 ;
        RECT 285.435 -105.565 285.765 -105.235 ;
        RECT 285.435 -106.925 285.765 -106.595 ;
        RECT 285.435 -108.285 285.765 -107.955 ;
        RECT 285.435 -109.645 285.765 -109.315 ;
        RECT 285.435 -111.005 285.765 -110.675 ;
        RECT 285.435 -112.365 285.765 -112.035 ;
        RECT 285.435 -113.725 285.765 -113.395 ;
        RECT 285.435 -115.085 285.765 -114.755 ;
        RECT 285.435 -116.445 285.765 -116.115 ;
        RECT 285.435 -117.805 285.765 -117.475 ;
        RECT 285.435 -119.165 285.765 -118.835 ;
        RECT 285.435 -120.525 285.765 -120.195 ;
        RECT 285.435 -121.885 285.765 -121.555 ;
        RECT 285.435 -123.245 285.765 -122.915 ;
        RECT 285.435 -124.605 285.765 -124.275 ;
        RECT 285.435 -125.965 285.765 -125.635 ;
        RECT 285.435 -127.325 285.765 -126.995 ;
        RECT 285.435 -128.685 285.765 -128.355 ;
        RECT 285.435 -130.045 285.765 -129.715 ;
        RECT 285.435 -131.405 285.765 -131.075 ;
        RECT 285.435 -132.765 285.765 -132.435 ;
        RECT 285.435 -134.125 285.765 -133.795 ;
        RECT 285.435 -135.485 285.765 -135.155 ;
        RECT 285.435 -136.845 285.765 -136.515 ;
        RECT 285.435 -138.205 285.765 -137.875 ;
        RECT 285.435 -139.565 285.765 -139.235 ;
        RECT 285.435 -140.925 285.765 -140.595 ;
        RECT 285.435 -142.285 285.765 -141.955 ;
        RECT 285.435 -143.645 285.765 -143.315 ;
        RECT 285.435 -145.005 285.765 -144.675 ;
        RECT 285.435 -146.365 285.765 -146.035 ;
        RECT 285.435 -147.725 285.765 -147.395 ;
        RECT 285.435 -149.085 285.765 -148.755 ;
        RECT 285.435 -150.445 285.765 -150.115 ;
        RECT 285.435 -151.805 285.765 -151.475 ;
        RECT 285.435 -153.165 285.765 -152.835 ;
        RECT 285.435 -154.525 285.765 -154.195 ;
        RECT 285.435 -155.885 285.765 -155.555 ;
        RECT 285.435 -157.245 285.765 -156.915 ;
        RECT 285.435 -158.605 285.765 -158.275 ;
        RECT 285.435 -159.965 285.765 -159.635 ;
        RECT 285.435 -161.325 285.765 -160.995 ;
        RECT 285.435 -162.685 285.765 -162.355 ;
        RECT 285.435 -164.045 285.765 -163.715 ;
        RECT 285.435 -165.405 285.765 -165.075 ;
        RECT 285.435 -166.765 285.765 -166.435 ;
        RECT 285.435 -168.125 285.765 -167.795 ;
        RECT 285.435 -169.485 285.765 -169.155 ;
        RECT 285.435 -170.845 285.765 -170.515 ;
        RECT 285.435 -172.205 285.765 -171.875 ;
        RECT 285.435 -173.565 285.765 -173.235 ;
        RECT 285.435 -174.925 285.765 -174.595 ;
        RECT 285.435 -176.285 285.765 -175.955 ;
        RECT 285.435 -177.645 285.765 -177.315 ;
        RECT 285.435 -179.005 285.765 -178.675 ;
        RECT 285.435 -184.65 285.765 -183.52 ;
        RECT 285.44 -184.765 285.76 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.06 -98.075 286.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.795 244.04 287.125 245.17 ;
        RECT 286.795 239.875 287.125 240.205 ;
        RECT 286.795 238.515 287.125 238.845 ;
        RECT 286.795 237.155 287.125 237.485 ;
        RECT 286.8 237.155 287.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.155 244.04 288.485 245.17 ;
        RECT 288.155 239.875 288.485 240.205 ;
        RECT 288.155 238.515 288.485 238.845 ;
        RECT 288.155 237.155 288.485 237.485 ;
        RECT 288.16 237.155 288.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.155 -0.845 288.485 -0.515 ;
        RECT 288.155 -2.205 288.485 -1.875 ;
        RECT 288.155 -3.565 288.485 -3.235 ;
        RECT 288.16 -3.565 288.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.155 -96.045 288.485 -95.715 ;
        RECT 288.155 -97.405 288.485 -97.075 ;
        RECT 288.155 -98.765 288.485 -98.435 ;
        RECT 288.155 -100.125 288.485 -99.795 ;
        RECT 288.155 -101.485 288.485 -101.155 ;
        RECT 288.155 -102.845 288.485 -102.515 ;
        RECT 288.155 -104.205 288.485 -103.875 ;
        RECT 288.155 -105.565 288.485 -105.235 ;
        RECT 288.155 -106.925 288.485 -106.595 ;
        RECT 288.155 -108.285 288.485 -107.955 ;
        RECT 288.155 -109.645 288.485 -109.315 ;
        RECT 288.155 -111.005 288.485 -110.675 ;
        RECT 288.155 -112.365 288.485 -112.035 ;
        RECT 288.155 -113.725 288.485 -113.395 ;
        RECT 288.155 -115.085 288.485 -114.755 ;
        RECT 288.155 -116.445 288.485 -116.115 ;
        RECT 288.155 -117.805 288.485 -117.475 ;
        RECT 288.155 -119.165 288.485 -118.835 ;
        RECT 288.155 -120.525 288.485 -120.195 ;
        RECT 288.155 -121.885 288.485 -121.555 ;
        RECT 288.155 -123.245 288.485 -122.915 ;
        RECT 288.155 -124.605 288.485 -124.275 ;
        RECT 288.155 -125.965 288.485 -125.635 ;
        RECT 288.155 -127.325 288.485 -126.995 ;
        RECT 288.155 -128.685 288.485 -128.355 ;
        RECT 288.155 -130.045 288.485 -129.715 ;
        RECT 288.155 -131.405 288.485 -131.075 ;
        RECT 288.155 -132.765 288.485 -132.435 ;
        RECT 288.155 -134.125 288.485 -133.795 ;
        RECT 288.155 -135.485 288.485 -135.155 ;
        RECT 288.155 -136.845 288.485 -136.515 ;
        RECT 288.155 -138.205 288.485 -137.875 ;
        RECT 288.155 -139.565 288.485 -139.235 ;
        RECT 288.155 -140.925 288.485 -140.595 ;
        RECT 288.155 -142.285 288.485 -141.955 ;
        RECT 288.155 -143.645 288.485 -143.315 ;
        RECT 288.155 -145.005 288.485 -144.675 ;
        RECT 288.155 -146.365 288.485 -146.035 ;
        RECT 288.155 -147.725 288.485 -147.395 ;
        RECT 288.155 -149.085 288.485 -148.755 ;
        RECT 288.155 -150.445 288.485 -150.115 ;
        RECT 288.155 -151.805 288.485 -151.475 ;
        RECT 288.155 -153.165 288.485 -152.835 ;
        RECT 288.155 -154.525 288.485 -154.195 ;
        RECT 288.155 -155.885 288.485 -155.555 ;
        RECT 288.155 -157.245 288.485 -156.915 ;
        RECT 288.155 -158.605 288.485 -158.275 ;
        RECT 288.155 -159.965 288.485 -159.635 ;
        RECT 288.155 -161.325 288.485 -160.995 ;
        RECT 288.155 -162.685 288.485 -162.355 ;
        RECT 288.155 -164.045 288.485 -163.715 ;
        RECT 288.155 -165.405 288.485 -165.075 ;
        RECT 288.155 -166.765 288.485 -166.435 ;
        RECT 288.155 -168.125 288.485 -167.795 ;
        RECT 288.155 -169.485 288.485 -169.155 ;
        RECT 288.155 -170.845 288.485 -170.515 ;
        RECT 288.155 -172.205 288.485 -171.875 ;
        RECT 288.155 -173.565 288.485 -173.235 ;
        RECT 288.155 -174.925 288.485 -174.595 ;
        RECT 288.155 -176.285 288.485 -175.955 ;
        RECT 288.155 -177.645 288.485 -177.315 ;
        RECT 288.155 -179.005 288.485 -178.675 ;
        RECT 288.155 -184.65 288.485 -183.52 ;
        RECT 288.16 -184.765 288.48 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.515 244.04 289.845 245.17 ;
        RECT 289.515 239.875 289.845 240.205 ;
        RECT 289.515 238.515 289.845 238.845 ;
        RECT 289.515 237.155 289.845 237.485 ;
        RECT 289.52 237.155 289.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 289.515 -0.845 289.845 -0.515 ;
        RECT 289.515 -2.205 289.845 -1.875 ;
        RECT 289.515 -3.565 289.845 -3.235 ;
        RECT 289.52 -3.565 289.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.875 244.04 291.205 245.17 ;
        RECT 290.875 239.875 291.205 240.205 ;
        RECT 290.875 238.515 291.205 238.845 ;
        RECT 290.875 237.155 291.205 237.485 ;
        RECT 290.88 237.155 291.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.875 -0.845 291.205 -0.515 ;
        RECT 290.875 -2.205 291.205 -1.875 ;
        RECT 290.875 -3.565 291.205 -3.235 ;
        RECT 290.88 -3.565 291.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.875 -96.045 291.205 -95.715 ;
        RECT 290.875 -97.405 291.205 -97.075 ;
        RECT 290.875 -98.765 291.205 -98.435 ;
        RECT 290.875 -100.125 291.205 -99.795 ;
        RECT 290.875 -101.485 291.205 -101.155 ;
        RECT 290.875 -102.845 291.205 -102.515 ;
        RECT 290.875 -104.205 291.205 -103.875 ;
        RECT 290.875 -105.565 291.205 -105.235 ;
        RECT 290.875 -106.925 291.205 -106.595 ;
        RECT 290.875 -108.285 291.205 -107.955 ;
        RECT 290.875 -109.645 291.205 -109.315 ;
        RECT 290.875 -111.005 291.205 -110.675 ;
        RECT 290.875 -112.365 291.205 -112.035 ;
        RECT 290.875 -113.725 291.205 -113.395 ;
        RECT 290.875 -115.085 291.205 -114.755 ;
        RECT 290.875 -116.445 291.205 -116.115 ;
        RECT 290.875 -117.805 291.205 -117.475 ;
        RECT 290.875 -119.165 291.205 -118.835 ;
        RECT 290.875 -120.525 291.205 -120.195 ;
        RECT 290.875 -121.885 291.205 -121.555 ;
        RECT 290.875 -123.245 291.205 -122.915 ;
        RECT 290.875 -124.605 291.205 -124.275 ;
        RECT 290.875 -125.965 291.205 -125.635 ;
        RECT 290.875 -127.325 291.205 -126.995 ;
        RECT 290.875 -128.685 291.205 -128.355 ;
        RECT 290.875 -130.045 291.205 -129.715 ;
        RECT 290.875 -131.405 291.205 -131.075 ;
        RECT 290.875 -132.765 291.205 -132.435 ;
        RECT 290.875 -134.125 291.205 -133.795 ;
        RECT 290.875 -135.485 291.205 -135.155 ;
        RECT 290.875 -136.845 291.205 -136.515 ;
        RECT 290.875 -138.205 291.205 -137.875 ;
        RECT 290.875 -139.565 291.205 -139.235 ;
        RECT 290.875 -140.925 291.205 -140.595 ;
        RECT 290.875 -142.285 291.205 -141.955 ;
        RECT 290.875 -143.645 291.205 -143.315 ;
        RECT 290.875 -145.005 291.205 -144.675 ;
        RECT 290.875 -146.365 291.205 -146.035 ;
        RECT 290.875 -147.725 291.205 -147.395 ;
        RECT 290.875 -149.085 291.205 -148.755 ;
        RECT 290.875 -150.445 291.205 -150.115 ;
        RECT 290.875 -151.805 291.205 -151.475 ;
        RECT 290.875 -153.165 291.205 -152.835 ;
        RECT 290.875 -154.525 291.205 -154.195 ;
        RECT 290.875 -155.885 291.205 -155.555 ;
        RECT 290.875 -157.245 291.205 -156.915 ;
        RECT 290.875 -158.605 291.205 -158.275 ;
        RECT 290.875 -159.965 291.205 -159.635 ;
        RECT 290.875 -161.325 291.205 -160.995 ;
        RECT 290.875 -162.685 291.205 -162.355 ;
        RECT 290.875 -164.045 291.205 -163.715 ;
        RECT 290.875 -165.405 291.205 -165.075 ;
        RECT 290.875 -166.765 291.205 -166.435 ;
        RECT 290.875 -168.125 291.205 -167.795 ;
        RECT 290.875 -169.485 291.205 -169.155 ;
        RECT 290.875 -170.845 291.205 -170.515 ;
        RECT 290.875 -172.205 291.205 -171.875 ;
        RECT 290.875 -173.565 291.205 -173.235 ;
        RECT 290.875 -174.925 291.205 -174.595 ;
        RECT 290.875 -176.285 291.205 -175.955 ;
        RECT 290.875 -177.645 291.205 -177.315 ;
        RECT 290.875 -179.005 291.205 -178.675 ;
        RECT 290.875 -184.65 291.205 -183.52 ;
        RECT 290.88 -184.765 291.2 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.235 244.04 292.565 245.17 ;
        RECT 292.235 239.875 292.565 240.205 ;
        RECT 292.235 238.515 292.565 238.845 ;
        RECT 292.235 237.155 292.565 237.485 ;
        RECT 292.24 237.155 292.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.235 -0.845 292.565 -0.515 ;
        RECT 292.235 -2.205 292.565 -1.875 ;
        RECT 292.235 -3.565 292.565 -3.235 ;
        RECT 292.24 -3.565 292.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.235 -96.045 292.565 -95.715 ;
        RECT 292.235 -97.405 292.565 -97.075 ;
        RECT 292.235 -98.765 292.565 -98.435 ;
        RECT 292.235 -100.125 292.565 -99.795 ;
        RECT 292.235 -101.485 292.565 -101.155 ;
        RECT 292.235 -102.845 292.565 -102.515 ;
        RECT 292.235 -104.205 292.565 -103.875 ;
        RECT 292.235 -105.565 292.565 -105.235 ;
        RECT 292.235 -106.925 292.565 -106.595 ;
        RECT 292.235 -108.285 292.565 -107.955 ;
        RECT 292.235 -109.645 292.565 -109.315 ;
        RECT 292.235 -111.005 292.565 -110.675 ;
        RECT 292.235 -112.365 292.565 -112.035 ;
        RECT 292.235 -113.725 292.565 -113.395 ;
        RECT 292.235 -115.085 292.565 -114.755 ;
        RECT 292.235 -116.445 292.565 -116.115 ;
        RECT 292.235 -117.805 292.565 -117.475 ;
        RECT 292.235 -119.165 292.565 -118.835 ;
        RECT 292.235 -120.525 292.565 -120.195 ;
        RECT 292.235 -121.885 292.565 -121.555 ;
        RECT 292.235 -123.245 292.565 -122.915 ;
        RECT 292.235 -124.605 292.565 -124.275 ;
        RECT 292.235 -125.965 292.565 -125.635 ;
        RECT 292.235 -127.325 292.565 -126.995 ;
        RECT 292.235 -128.685 292.565 -128.355 ;
        RECT 292.235 -130.045 292.565 -129.715 ;
        RECT 292.235 -131.405 292.565 -131.075 ;
        RECT 292.235 -132.765 292.565 -132.435 ;
        RECT 292.235 -134.125 292.565 -133.795 ;
        RECT 292.235 -135.485 292.565 -135.155 ;
        RECT 292.235 -136.845 292.565 -136.515 ;
        RECT 292.235 -138.205 292.565 -137.875 ;
        RECT 292.235 -139.565 292.565 -139.235 ;
        RECT 292.235 -140.925 292.565 -140.595 ;
        RECT 292.235 -142.285 292.565 -141.955 ;
        RECT 292.235 -143.645 292.565 -143.315 ;
        RECT 292.235 -145.005 292.565 -144.675 ;
        RECT 292.235 -146.365 292.565 -146.035 ;
        RECT 292.235 -147.725 292.565 -147.395 ;
        RECT 292.235 -149.085 292.565 -148.755 ;
        RECT 292.235 -150.445 292.565 -150.115 ;
        RECT 292.235 -151.805 292.565 -151.475 ;
        RECT 292.235 -153.165 292.565 -152.835 ;
        RECT 292.235 -154.525 292.565 -154.195 ;
        RECT 292.235 -155.885 292.565 -155.555 ;
        RECT 292.235 -157.245 292.565 -156.915 ;
        RECT 292.235 -158.605 292.565 -158.275 ;
        RECT 292.235 -159.965 292.565 -159.635 ;
        RECT 292.235 -161.325 292.565 -160.995 ;
        RECT 292.235 -162.685 292.565 -162.355 ;
        RECT 292.235 -164.045 292.565 -163.715 ;
        RECT 292.235 -165.405 292.565 -165.075 ;
        RECT 292.235 -166.765 292.565 -166.435 ;
        RECT 292.235 -168.125 292.565 -167.795 ;
        RECT 292.235 -169.485 292.565 -169.155 ;
        RECT 292.235 -170.845 292.565 -170.515 ;
        RECT 292.235 -172.205 292.565 -171.875 ;
        RECT 292.235 -173.565 292.565 -173.235 ;
        RECT 292.235 -174.925 292.565 -174.595 ;
        RECT 292.235 -176.285 292.565 -175.955 ;
        RECT 292.235 -177.645 292.565 -177.315 ;
        RECT 292.235 -179.005 292.565 -178.675 ;
        RECT 292.235 -184.65 292.565 -183.52 ;
        RECT 292.24 -184.765 292.56 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.595 244.04 293.925 245.17 ;
        RECT 293.595 239.875 293.925 240.205 ;
        RECT 293.595 238.515 293.925 238.845 ;
        RECT 293.595 237.155 293.925 237.485 ;
        RECT 293.6 237.155 293.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.595 -0.845 293.925 -0.515 ;
        RECT 293.595 -2.205 293.925 -1.875 ;
        RECT 293.595 -3.565 293.925 -3.235 ;
        RECT 293.6 -3.565 293.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 293.595 -96.045 293.925 -95.715 ;
        RECT 293.595 -97.405 293.925 -97.075 ;
        RECT 293.595 -98.765 293.925 -98.435 ;
        RECT 293.595 -100.125 293.925 -99.795 ;
        RECT 293.595 -101.485 293.925 -101.155 ;
        RECT 293.595 -102.845 293.925 -102.515 ;
        RECT 293.595 -104.205 293.925 -103.875 ;
        RECT 293.595 -105.565 293.925 -105.235 ;
        RECT 293.595 -106.925 293.925 -106.595 ;
        RECT 293.595 -108.285 293.925 -107.955 ;
        RECT 293.595 -109.645 293.925 -109.315 ;
        RECT 293.595 -111.005 293.925 -110.675 ;
        RECT 293.595 -112.365 293.925 -112.035 ;
        RECT 293.595 -113.725 293.925 -113.395 ;
        RECT 293.595 -115.085 293.925 -114.755 ;
        RECT 293.595 -116.445 293.925 -116.115 ;
        RECT 293.595 -117.805 293.925 -117.475 ;
        RECT 293.595 -119.165 293.925 -118.835 ;
        RECT 293.595 -120.525 293.925 -120.195 ;
        RECT 293.595 -121.885 293.925 -121.555 ;
        RECT 293.595 -123.245 293.925 -122.915 ;
        RECT 293.595 -124.605 293.925 -124.275 ;
        RECT 293.595 -125.965 293.925 -125.635 ;
        RECT 293.595 -127.325 293.925 -126.995 ;
        RECT 293.595 -128.685 293.925 -128.355 ;
        RECT 293.595 -130.045 293.925 -129.715 ;
        RECT 293.595 -131.405 293.925 -131.075 ;
        RECT 293.595 -132.765 293.925 -132.435 ;
        RECT 293.595 -134.125 293.925 -133.795 ;
        RECT 293.595 -135.485 293.925 -135.155 ;
        RECT 293.595 -136.845 293.925 -136.515 ;
        RECT 293.595 -138.205 293.925 -137.875 ;
        RECT 293.595 -139.565 293.925 -139.235 ;
        RECT 293.595 -140.925 293.925 -140.595 ;
        RECT 293.595 -142.285 293.925 -141.955 ;
        RECT 293.595 -143.645 293.925 -143.315 ;
        RECT 293.595 -145.005 293.925 -144.675 ;
        RECT 293.595 -146.365 293.925 -146.035 ;
        RECT 293.595 -147.725 293.925 -147.395 ;
        RECT 293.595 -149.085 293.925 -148.755 ;
        RECT 293.595 -150.445 293.925 -150.115 ;
        RECT 293.595 -151.805 293.925 -151.475 ;
        RECT 293.595 -153.165 293.925 -152.835 ;
        RECT 293.595 -154.525 293.925 -154.195 ;
        RECT 293.595 -155.885 293.925 -155.555 ;
        RECT 293.595 -157.245 293.925 -156.915 ;
        RECT 293.595 -158.605 293.925 -158.275 ;
        RECT 293.595 -159.965 293.925 -159.635 ;
        RECT 293.595 -161.325 293.925 -160.995 ;
        RECT 293.595 -162.685 293.925 -162.355 ;
        RECT 293.595 -164.045 293.925 -163.715 ;
        RECT 293.595 -165.405 293.925 -165.075 ;
        RECT 293.595 -166.765 293.925 -166.435 ;
        RECT 293.595 -168.125 293.925 -167.795 ;
        RECT 293.595 -169.485 293.925 -169.155 ;
        RECT 293.595 -170.845 293.925 -170.515 ;
        RECT 293.595 -172.205 293.925 -171.875 ;
        RECT 293.595 -173.565 293.925 -173.235 ;
        RECT 293.595 -174.925 293.925 -174.595 ;
        RECT 293.595 -176.285 293.925 -175.955 ;
        RECT 293.595 -177.645 293.925 -177.315 ;
        RECT 293.595 -179.005 293.925 -178.675 ;
        RECT 293.595 -184.65 293.925 -183.52 ;
        RECT 293.6 -184.765 293.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.955 244.04 295.285 245.17 ;
        RECT 294.955 239.875 295.285 240.205 ;
        RECT 294.955 238.515 295.285 238.845 ;
        RECT 294.955 237.155 295.285 237.485 ;
        RECT 294.96 237.155 295.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.955 -0.845 295.285 -0.515 ;
        RECT 294.955 -2.205 295.285 -1.875 ;
        RECT 294.955 -3.565 295.285 -3.235 ;
        RECT 294.96 -3.565 295.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.955 -96.045 295.285 -95.715 ;
        RECT 294.955 -97.405 295.285 -97.075 ;
        RECT 294.955 -98.765 295.285 -98.435 ;
        RECT 294.955 -100.125 295.285 -99.795 ;
        RECT 294.955 -101.485 295.285 -101.155 ;
        RECT 294.955 -102.845 295.285 -102.515 ;
        RECT 294.955 -104.205 295.285 -103.875 ;
        RECT 294.955 -105.565 295.285 -105.235 ;
        RECT 294.955 -106.925 295.285 -106.595 ;
        RECT 294.955 -108.285 295.285 -107.955 ;
        RECT 294.955 -109.645 295.285 -109.315 ;
        RECT 294.955 -111.005 295.285 -110.675 ;
        RECT 294.955 -112.365 295.285 -112.035 ;
        RECT 294.955 -113.725 295.285 -113.395 ;
        RECT 294.955 -115.085 295.285 -114.755 ;
        RECT 294.955 -116.445 295.285 -116.115 ;
        RECT 294.955 -117.805 295.285 -117.475 ;
        RECT 294.955 -119.165 295.285 -118.835 ;
        RECT 294.955 -120.525 295.285 -120.195 ;
        RECT 294.955 -121.885 295.285 -121.555 ;
        RECT 294.955 -123.245 295.285 -122.915 ;
        RECT 294.955 -124.605 295.285 -124.275 ;
        RECT 294.955 -125.965 295.285 -125.635 ;
        RECT 294.955 -127.325 295.285 -126.995 ;
        RECT 294.955 -128.685 295.285 -128.355 ;
        RECT 294.955 -130.045 295.285 -129.715 ;
        RECT 294.955 -131.405 295.285 -131.075 ;
        RECT 294.955 -132.765 295.285 -132.435 ;
        RECT 294.955 -134.125 295.285 -133.795 ;
        RECT 294.955 -135.485 295.285 -135.155 ;
        RECT 294.955 -136.845 295.285 -136.515 ;
        RECT 294.955 -138.205 295.285 -137.875 ;
        RECT 294.955 -139.565 295.285 -139.235 ;
        RECT 294.955 -140.925 295.285 -140.595 ;
        RECT 294.955 -142.285 295.285 -141.955 ;
        RECT 294.955 -143.645 295.285 -143.315 ;
        RECT 294.955 -145.005 295.285 -144.675 ;
        RECT 294.955 -146.365 295.285 -146.035 ;
        RECT 294.955 -147.725 295.285 -147.395 ;
        RECT 294.955 -149.085 295.285 -148.755 ;
        RECT 294.955 -150.445 295.285 -150.115 ;
        RECT 294.955 -151.805 295.285 -151.475 ;
        RECT 294.955 -153.165 295.285 -152.835 ;
        RECT 294.955 -154.525 295.285 -154.195 ;
        RECT 294.955 -155.885 295.285 -155.555 ;
        RECT 294.955 -157.245 295.285 -156.915 ;
        RECT 294.955 -158.605 295.285 -158.275 ;
        RECT 294.955 -159.965 295.285 -159.635 ;
        RECT 294.955 -161.325 295.285 -160.995 ;
        RECT 294.955 -162.685 295.285 -162.355 ;
        RECT 294.955 -164.045 295.285 -163.715 ;
        RECT 294.955 -165.405 295.285 -165.075 ;
        RECT 294.955 -166.765 295.285 -166.435 ;
        RECT 294.955 -168.125 295.285 -167.795 ;
        RECT 294.955 -169.485 295.285 -169.155 ;
        RECT 294.955 -170.845 295.285 -170.515 ;
        RECT 294.955 -172.205 295.285 -171.875 ;
        RECT 294.955 -173.565 295.285 -173.235 ;
        RECT 294.955 -174.925 295.285 -174.595 ;
        RECT 294.955 -176.285 295.285 -175.955 ;
        RECT 294.955 -177.645 295.285 -177.315 ;
        RECT 294.955 -179.005 295.285 -178.675 ;
        RECT 294.955 -184.65 295.285 -183.52 ;
        RECT 294.96 -184.765 295.28 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.315 244.04 296.645 245.17 ;
        RECT 296.315 239.875 296.645 240.205 ;
        RECT 296.315 238.515 296.645 238.845 ;
        RECT 296.315 237.155 296.645 237.485 ;
        RECT 296.32 237.155 296.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.315 -98.765 296.645 -98.435 ;
        RECT 296.315 -100.125 296.645 -99.795 ;
        RECT 296.315 -101.485 296.645 -101.155 ;
        RECT 296.315 -102.845 296.645 -102.515 ;
        RECT 296.315 -104.205 296.645 -103.875 ;
        RECT 296.315 -105.565 296.645 -105.235 ;
        RECT 296.315 -106.925 296.645 -106.595 ;
        RECT 296.315 -108.285 296.645 -107.955 ;
        RECT 296.315 -109.645 296.645 -109.315 ;
        RECT 296.315 -111.005 296.645 -110.675 ;
        RECT 296.315 -112.365 296.645 -112.035 ;
        RECT 296.315 -113.725 296.645 -113.395 ;
        RECT 296.315 -115.085 296.645 -114.755 ;
        RECT 296.315 -116.445 296.645 -116.115 ;
        RECT 296.315 -117.805 296.645 -117.475 ;
        RECT 296.315 -119.165 296.645 -118.835 ;
        RECT 296.315 -120.525 296.645 -120.195 ;
        RECT 296.315 -121.885 296.645 -121.555 ;
        RECT 296.315 -123.245 296.645 -122.915 ;
        RECT 296.315 -124.605 296.645 -124.275 ;
        RECT 296.315 -125.965 296.645 -125.635 ;
        RECT 296.315 -127.325 296.645 -126.995 ;
        RECT 296.315 -128.685 296.645 -128.355 ;
        RECT 296.315 -130.045 296.645 -129.715 ;
        RECT 296.315 -131.405 296.645 -131.075 ;
        RECT 296.315 -132.765 296.645 -132.435 ;
        RECT 296.315 -134.125 296.645 -133.795 ;
        RECT 296.315 -135.485 296.645 -135.155 ;
        RECT 296.315 -136.845 296.645 -136.515 ;
        RECT 296.315 -138.205 296.645 -137.875 ;
        RECT 296.315 -139.565 296.645 -139.235 ;
        RECT 296.315 -140.925 296.645 -140.595 ;
        RECT 296.315 -142.285 296.645 -141.955 ;
        RECT 296.315 -143.645 296.645 -143.315 ;
        RECT 296.315 -145.005 296.645 -144.675 ;
        RECT 296.315 -146.365 296.645 -146.035 ;
        RECT 296.315 -147.725 296.645 -147.395 ;
        RECT 296.315 -149.085 296.645 -148.755 ;
        RECT 296.315 -150.445 296.645 -150.115 ;
        RECT 296.315 -151.805 296.645 -151.475 ;
        RECT 296.315 -153.165 296.645 -152.835 ;
        RECT 296.315 -154.525 296.645 -154.195 ;
        RECT 296.315 -155.885 296.645 -155.555 ;
        RECT 296.315 -157.245 296.645 -156.915 ;
        RECT 296.315 -158.605 296.645 -158.275 ;
        RECT 296.315 -159.965 296.645 -159.635 ;
        RECT 296.315 -161.325 296.645 -160.995 ;
        RECT 296.315 -162.685 296.645 -162.355 ;
        RECT 296.315 -164.045 296.645 -163.715 ;
        RECT 296.315 -165.405 296.645 -165.075 ;
        RECT 296.315 -166.765 296.645 -166.435 ;
        RECT 296.315 -168.125 296.645 -167.795 ;
        RECT 296.315 -169.485 296.645 -169.155 ;
        RECT 296.315 -170.845 296.645 -170.515 ;
        RECT 296.315 -172.205 296.645 -171.875 ;
        RECT 296.315 -173.565 296.645 -173.235 ;
        RECT 296.315 -174.925 296.645 -174.595 ;
        RECT 296.315 -176.285 296.645 -175.955 ;
        RECT 296.315 -177.645 296.645 -177.315 ;
        RECT 296.315 -179.005 296.645 -178.675 ;
        RECT 296.315 -184.65 296.645 -183.52 ;
        RECT 296.32 -184.765 296.64 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.96 -98.075 297.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.675 244.04 298.005 245.17 ;
        RECT 297.675 239.875 298.005 240.205 ;
        RECT 297.675 238.515 298.005 238.845 ;
        RECT 297.675 237.155 298.005 237.485 ;
        RECT 297.68 237.155 298 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.035 244.04 299.365 245.17 ;
        RECT 299.035 239.875 299.365 240.205 ;
        RECT 299.035 238.515 299.365 238.845 ;
        RECT 299.035 237.155 299.365 237.485 ;
        RECT 299.04 237.155 299.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.035 -0.845 299.365 -0.515 ;
        RECT 299.035 -2.205 299.365 -1.875 ;
        RECT 299.035 -3.565 299.365 -3.235 ;
        RECT 299.04 -3.565 299.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.395 244.04 300.725 245.17 ;
        RECT 300.395 239.875 300.725 240.205 ;
        RECT 300.395 238.515 300.725 238.845 ;
        RECT 300.395 237.155 300.725 237.485 ;
        RECT 300.4 237.155 300.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 300.395 -0.845 300.725 -0.515 ;
        RECT 300.395 -2.205 300.725 -1.875 ;
        RECT 300.395 -3.565 300.725 -3.235 ;
        RECT 300.4 -3.565 300.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.755 244.04 302.085 245.17 ;
        RECT 301.755 239.875 302.085 240.205 ;
        RECT 301.755 238.515 302.085 238.845 ;
        RECT 301.755 237.155 302.085 237.485 ;
        RECT 301.76 237.155 302.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.755 -0.845 302.085 -0.515 ;
        RECT 301.755 -2.205 302.085 -1.875 ;
        RECT 301.755 -3.565 302.085 -3.235 ;
        RECT 301.76 -3.565 302.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.755 -96.045 302.085 -95.715 ;
        RECT 301.755 -97.405 302.085 -97.075 ;
        RECT 301.755 -98.765 302.085 -98.435 ;
        RECT 301.755 -100.125 302.085 -99.795 ;
        RECT 301.755 -101.485 302.085 -101.155 ;
        RECT 301.755 -102.845 302.085 -102.515 ;
        RECT 301.755 -104.205 302.085 -103.875 ;
        RECT 301.755 -105.565 302.085 -105.235 ;
        RECT 301.755 -106.925 302.085 -106.595 ;
        RECT 301.755 -108.285 302.085 -107.955 ;
        RECT 301.755 -109.645 302.085 -109.315 ;
        RECT 301.755 -111.005 302.085 -110.675 ;
        RECT 301.755 -112.365 302.085 -112.035 ;
        RECT 301.755 -113.725 302.085 -113.395 ;
        RECT 301.755 -115.085 302.085 -114.755 ;
        RECT 301.755 -116.445 302.085 -116.115 ;
        RECT 301.755 -117.805 302.085 -117.475 ;
        RECT 301.755 -119.165 302.085 -118.835 ;
        RECT 301.755 -120.525 302.085 -120.195 ;
        RECT 301.755 -121.885 302.085 -121.555 ;
        RECT 301.755 -123.245 302.085 -122.915 ;
        RECT 301.755 -124.605 302.085 -124.275 ;
        RECT 301.755 -125.965 302.085 -125.635 ;
        RECT 301.755 -127.325 302.085 -126.995 ;
        RECT 301.755 -128.685 302.085 -128.355 ;
        RECT 301.755 -130.045 302.085 -129.715 ;
        RECT 301.755 -131.405 302.085 -131.075 ;
        RECT 301.755 -132.765 302.085 -132.435 ;
        RECT 301.755 -134.125 302.085 -133.795 ;
        RECT 301.755 -135.485 302.085 -135.155 ;
        RECT 301.755 -136.845 302.085 -136.515 ;
        RECT 301.755 -138.205 302.085 -137.875 ;
        RECT 301.755 -139.565 302.085 -139.235 ;
        RECT 301.755 -140.925 302.085 -140.595 ;
        RECT 301.755 -142.285 302.085 -141.955 ;
        RECT 301.755 -143.645 302.085 -143.315 ;
        RECT 301.755 -145.005 302.085 -144.675 ;
        RECT 301.755 -146.365 302.085 -146.035 ;
        RECT 301.755 -147.725 302.085 -147.395 ;
        RECT 301.755 -149.085 302.085 -148.755 ;
        RECT 301.755 -150.445 302.085 -150.115 ;
        RECT 301.755 -151.805 302.085 -151.475 ;
        RECT 301.755 -153.165 302.085 -152.835 ;
        RECT 301.755 -154.525 302.085 -154.195 ;
        RECT 301.755 -155.885 302.085 -155.555 ;
        RECT 301.755 -157.245 302.085 -156.915 ;
        RECT 301.755 -158.605 302.085 -158.275 ;
        RECT 301.755 -159.965 302.085 -159.635 ;
        RECT 301.755 -161.325 302.085 -160.995 ;
        RECT 301.755 -162.685 302.085 -162.355 ;
        RECT 301.755 -164.045 302.085 -163.715 ;
        RECT 301.755 -165.405 302.085 -165.075 ;
        RECT 301.755 -166.765 302.085 -166.435 ;
        RECT 301.755 -168.125 302.085 -167.795 ;
        RECT 301.755 -169.485 302.085 -169.155 ;
        RECT 301.755 -170.845 302.085 -170.515 ;
        RECT 301.755 -172.205 302.085 -171.875 ;
        RECT 301.755 -173.565 302.085 -173.235 ;
        RECT 301.755 -174.925 302.085 -174.595 ;
        RECT 301.755 -176.285 302.085 -175.955 ;
        RECT 301.755 -177.645 302.085 -177.315 ;
        RECT 301.755 -179.005 302.085 -178.675 ;
        RECT 301.755 -184.65 302.085 -183.52 ;
        RECT 301.76 -184.765 302.08 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.115 244.04 303.445 245.17 ;
        RECT 303.115 239.875 303.445 240.205 ;
        RECT 303.115 238.515 303.445 238.845 ;
        RECT 303.115 237.155 303.445 237.485 ;
        RECT 303.12 237.155 303.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.115 -0.845 303.445 -0.515 ;
        RECT 303.115 -2.205 303.445 -1.875 ;
        RECT 303.115 -3.565 303.445 -3.235 ;
        RECT 303.12 -3.565 303.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.115 -96.045 303.445 -95.715 ;
        RECT 303.115 -97.405 303.445 -97.075 ;
        RECT 303.115 -98.765 303.445 -98.435 ;
        RECT 303.115 -100.125 303.445 -99.795 ;
        RECT 303.115 -101.485 303.445 -101.155 ;
        RECT 303.115 -102.845 303.445 -102.515 ;
        RECT 303.115 -104.205 303.445 -103.875 ;
        RECT 303.115 -105.565 303.445 -105.235 ;
        RECT 303.115 -106.925 303.445 -106.595 ;
        RECT 303.115 -108.285 303.445 -107.955 ;
        RECT 303.115 -109.645 303.445 -109.315 ;
        RECT 303.115 -111.005 303.445 -110.675 ;
        RECT 303.115 -112.365 303.445 -112.035 ;
        RECT 303.115 -113.725 303.445 -113.395 ;
        RECT 303.115 -115.085 303.445 -114.755 ;
        RECT 303.115 -116.445 303.445 -116.115 ;
        RECT 303.115 -117.805 303.445 -117.475 ;
        RECT 303.115 -119.165 303.445 -118.835 ;
        RECT 303.115 -120.525 303.445 -120.195 ;
        RECT 303.115 -121.885 303.445 -121.555 ;
        RECT 303.115 -123.245 303.445 -122.915 ;
        RECT 303.115 -124.605 303.445 -124.275 ;
        RECT 303.115 -125.965 303.445 -125.635 ;
        RECT 303.115 -127.325 303.445 -126.995 ;
        RECT 303.115 -128.685 303.445 -128.355 ;
        RECT 303.115 -130.045 303.445 -129.715 ;
        RECT 303.115 -131.405 303.445 -131.075 ;
        RECT 303.115 -132.765 303.445 -132.435 ;
        RECT 303.115 -134.125 303.445 -133.795 ;
        RECT 303.115 -135.485 303.445 -135.155 ;
        RECT 303.115 -136.845 303.445 -136.515 ;
        RECT 303.115 -138.205 303.445 -137.875 ;
        RECT 303.115 -139.565 303.445 -139.235 ;
        RECT 303.115 -140.925 303.445 -140.595 ;
        RECT 303.115 -142.285 303.445 -141.955 ;
        RECT 303.115 -143.645 303.445 -143.315 ;
        RECT 303.115 -145.005 303.445 -144.675 ;
        RECT 303.115 -146.365 303.445 -146.035 ;
        RECT 303.115 -147.725 303.445 -147.395 ;
        RECT 303.115 -149.085 303.445 -148.755 ;
        RECT 303.115 -150.445 303.445 -150.115 ;
        RECT 303.115 -151.805 303.445 -151.475 ;
        RECT 303.115 -153.165 303.445 -152.835 ;
        RECT 303.115 -154.525 303.445 -154.195 ;
        RECT 303.115 -155.885 303.445 -155.555 ;
        RECT 303.115 -157.245 303.445 -156.915 ;
        RECT 303.115 -158.605 303.445 -158.275 ;
        RECT 303.115 -159.965 303.445 -159.635 ;
        RECT 303.115 -161.325 303.445 -160.995 ;
        RECT 303.115 -162.685 303.445 -162.355 ;
        RECT 303.115 -164.045 303.445 -163.715 ;
        RECT 303.115 -165.405 303.445 -165.075 ;
        RECT 303.115 -166.765 303.445 -166.435 ;
        RECT 303.115 -168.125 303.445 -167.795 ;
        RECT 303.115 -169.485 303.445 -169.155 ;
        RECT 303.115 -170.845 303.445 -170.515 ;
        RECT 303.115 -172.205 303.445 -171.875 ;
        RECT 303.115 -173.565 303.445 -173.235 ;
        RECT 303.115 -174.925 303.445 -174.595 ;
        RECT 303.115 -176.285 303.445 -175.955 ;
        RECT 303.115 -177.645 303.445 -177.315 ;
        RECT 303.115 -179.005 303.445 -178.675 ;
        RECT 303.115 -184.65 303.445 -183.52 ;
        RECT 303.12 -184.765 303.44 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.475 244.04 304.805 245.17 ;
        RECT 304.475 239.875 304.805 240.205 ;
        RECT 304.475 238.515 304.805 238.845 ;
        RECT 304.475 237.155 304.805 237.485 ;
        RECT 304.48 237.155 304.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.475 -0.845 304.805 -0.515 ;
        RECT 304.475 -2.205 304.805 -1.875 ;
        RECT 304.475 -3.565 304.805 -3.235 ;
        RECT 304.48 -3.565 304.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 304.475 -96.045 304.805 -95.715 ;
        RECT 304.475 -97.405 304.805 -97.075 ;
        RECT 304.475 -98.765 304.805 -98.435 ;
        RECT 304.475 -100.125 304.805 -99.795 ;
        RECT 304.475 -101.485 304.805 -101.155 ;
        RECT 304.475 -102.845 304.805 -102.515 ;
        RECT 304.475 -104.205 304.805 -103.875 ;
        RECT 304.475 -105.565 304.805 -105.235 ;
        RECT 304.475 -106.925 304.805 -106.595 ;
        RECT 304.475 -108.285 304.805 -107.955 ;
        RECT 304.475 -109.645 304.805 -109.315 ;
        RECT 304.475 -111.005 304.805 -110.675 ;
        RECT 304.475 -112.365 304.805 -112.035 ;
        RECT 304.475 -113.725 304.805 -113.395 ;
        RECT 304.475 -115.085 304.805 -114.755 ;
        RECT 304.475 -116.445 304.805 -116.115 ;
        RECT 304.475 -117.805 304.805 -117.475 ;
        RECT 304.475 -119.165 304.805 -118.835 ;
        RECT 304.475 -120.525 304.805 -120.195 ;
        RECT 304.475 -121.885 304.805 -121.555 ;
        RECT 304.475 -123.245 304.805 -122.915 ;
        RECT 304.475 -124.605 304.805 -124.275 ;
        RECT 304.475 -125.965 304.805 -125.635 ;
        RECT 304.475 -127.325 304.805 -126.995 ;
        RECT 304.475 -128.685 304.805 -128.355 ;
        RECT 304.475 -130.045 304.805 -129.715 ;
        RECT 304.475 -131.405 304.805 -131.075 ;
        RECT 304.475 -132.765 304.805 -132.435 ;
        RECT 304.475 -134.125 304.805 -133.795 ;
        RECT 304.475 -135.485 304.805 -135.155 ;
        RECT 304.475 -136.845 304.805 -136.515 ;
        RECT 304.475 -138.205 304.805 -137.875 ;
        RECT 304.475 -139.565 304.805 -139.235 ;
        RECT 304.475 -140.925 304.805 -140.595 ;
        RECT 304.475 -142.285 304.805 -141.955 ;
        RECT 304.475 -143.645 304.805 -143.315 ;
        RECT 304.475 -145.005 304.805 -144.675 ;
        RECT 304.475 -146.365 304.805 -146.035 ;
        RECT 304.475 -147.725 304.805 -147.395 ;
        RECT 304.475 -149.085 304.805 -148.755 ;
        RECT 304.475 -150.445 304.805 -150.115 ;
        RECT 304.475 -151.805 304.805 -151.475 ;
        RECT 304.475 -153.165 304.805 -152.835 ;
        RECT 304.475 -154.525 304.805 -154.195 ;
        RECT 304.475 -155.885 304.805 -155.555 ;
        RECT 304.475 -157.245 304.805 -156.915 ;
        RECT 304.475 -158.605 304.805 -158.275 ;
        RECT 304.475 -159.965 304.805 -159.635 ;
        RECT 304.475 -161.325 304.805 -160.995 ;
        RECT 304.475 -162.685 304.805 -162.355 ;
        RECT 304.475 -164.045 304.805 -163.715 ;
        RECT 304.475 -165.405 304.805 -165.075 ;
        RECT 304.475 -166.765 304.805 -166.435 ;
        RECT 304.475 -168.125 304.805 -167.795 ;
        RECT 304.475 -169.485 304.805 -169.155 ;
        RECT 304.475 -170.845 304.805 -170.515 ;
        RECT 304.475 -172.205 304.805 -171.875 ;
        RECT 304.475 -173.565 304.805 -173.235 ;
        RECT 304.475 -174.925 304.805 -174.595 ;
        RECT 304.475 -176.285 304.805 -175.955 ;
        RECT 304.475 -177.645 304.805 -177.315 ;
        RECT 304.475 -179.005 304.805 -178.675 ;
        RECT 304.475 -184.65 304.805 -183.52 ;
        RECT 304.48 -184.765 304.8 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.835 244.04 306.165 245.17 ;
        RECT 305.835 239.875 306.165 240.205 ;
        RECT 305.835 238.515 306.165 238.845 ;
        RECT 305.835 237.155 306.165 237.485 ;
        RECT 305.84 237.155 306.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.835 -0.845 306.165 -0.515 ;
        RECT 305.835 -2.205 306.165 -1.875 ;
        RECT 305.835 -3.565 306.165 -3.235 ;
        RECT 305.84 -3.565 306.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.835 -96.045 306.165 -95.715 ;
        RECT 305.835 -97.405 306.165 -97.075 ;
        RECT 305.835 -98.765 306.165 -98.435 ;
        RECT 305.835 -100.125 306.165 -99.795 ;
        RECT 305.835 -101.485 306.165 -101.155 ;
        RECT 305.835 -102.845 306.165 -102.515 ;
        RECT 305.835 -104.205 306.165 -103.875 ;
        RECT 305.835 -105.565 306.165 -105.235 ;
        RECT 305.835 -106.925 306.165 -106.595 ;
        RECT 305.835 -108.285 306.165 -107.955 ;
        RECT 305.835 -109.645 306.165 -109.315 ;
        RECT 305.835 -111.005 306.165 -110.675 ;
        RECT 305.835 -112.365 306.165 -112.035 ;
        RECT 305.835 -113.725 306.165 -113.395 ;
        RECT 305.835 -115.085 306.165 -114.755 ;
        RECT 305.835 -116.445 306.165 -116.115 ;
        RECT 305.835 -117.805 306.165 -117.475 ;
        RECT 305.835 -119.165 306.165 -118.835 ;
        RECT 305.835 -120.525 306.165 -120.195 ;
        RECT 305.835 -121.885 306.165 -121.555 ;
        RECT 305.835 -123.245 306.165 -122.915 ;
        RECT 305.835 -124.605 306.165 -124.275 ;
        RECT 305.835 -125.965 306.165 -125.635 ;
        RECT 305.835 -127.325 306.165 -126.995 ;
        RECT 305.835 -128.685 306.165 -128.355 ;
        RECT 305.835 -130.045 306.165 -129.715 ;
        RECT 305.835 -131.405 306.165 -131.075 ;
        RECT 305.835 -132.765 306.165 -132.435 ;
        RECT 305.835 -134.125 306.165 -133.795 ;
        RECT 305.835 -135.485 306.165 -135.155 ;
        RECT 305.835 -136.845 306.165 -136.515 ;
        RECT 305.835 -138.205 306.165 -137.875 ;
        RECT 305.835 -139.565 306.165 -139.235 ;
        RECT 305.835 -140.925 306.165 -140.595 ;
        RECT 305.835 -142.285 306.165 -141.955 ;
        RECT 305.835 -143.645 306.165 -143.315 ;
        RECT 305.835 -145.005 306.165 -144.675 ;
        RECT 305.835 -146.365 306.165 -146.035 ;
        RECT 305.835 -147.725 306.165 -147.395 ;
        RECT 305.835 -149.085 306.165 -148.755 ;
        RECT 305.835 -150.445 306.165 -150.115 ;
        RECT 305.835 -151.805 306.165 -151.475 ;
        RECT 305.835 -153.165 306.165 -152.835 ;
        RECT 305.835 -154.525 306.165 -154.195 ;
        RECT 305.835 -155.885 306.165 -155.555 ;
        RECT 305.835 -157.245 306.165 -156.915 ;
        RECT 305.835 -158.605 306.165 -158.275 ;
        RECT 305.835 -159.965 306.165 -159.635 ;
        RECT 305.835 -161.325 306.165 -160.995 ;
        RECT 305.835 -162.685 306.165 -162.355 ;
        RECT 305.835 -164.045 306.165 -163.715 ;
        RECT 305.835 -165.405 306.165 -165.075 ;
        RECT 305.835 -166.765 306.165 -166.435 ;
        RECT 305.835 -168.125 306.165 -167.795 ;
        RECT 305.835 -169.485 306.165 -169.155 ;
        RECT 305.835 -170.845 306.165 -170.515 ;
        RECT 305.835 -172.205 306.165 -171.875 ;
        RECT 305.835 -173.565 306.165 -173.235 ;
        RECT 305.835 -174.925 306.165 -174.595 ;
        RECT 305.835 -176.285 306.165 -175.955 ;
        RECT 305.835 -177.645 306.165 -177.315 ;
        RECT 305.835 -179.005 306.165 -178.675 ;
        RECT 305.835 -184.65 306.165 -183.52 ;
        RECT 305.84 -184.765 306.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.195 244.04 307.525 245.17 ;
        RECT 307.195 239.875 307.525 240.205 ;
        RECT 307.195 238.515 307.525 238.845 ;
        RECT 307.195 237.155 307.525 237.485 ;
        RECT 307.2 237.155 307.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.195 -98.765 307.525 -98.435 ;
        RECT 307.195 -100.125 307.525 -99.795 ;
        RECT 307.195 -101.485 307.525 -101.155 ;
        RECT 307.195 -102.845 307.525 -102.515 ;
        RECT 307.195 -104.205 307.525 -103.875 ;
        RECT 307.195 -105.565 307.525 -105.235 ;
        RECT 307.195 -106.925 307.525 -106.595 ;
        RECT 307.195 -108.285 307.525 -107.955 ;
        RECT 307.195 -109.645 307.525 -109.315 ;
        RECT 307.195 -111.005 307.525 -110.675 ;
        RECT 307.195 -112.365 307.525 -112.035 ;
        RECT 307.195 -113.725 307.525 -113.395 ;
        RECT 307.195 -115.085 307.525 -114.755 ;
        RECT 307.195 -116.445 307.525 -116.115 ;
        RECT 307.195 -117.805 307.525 -117.475 ;
        RECT 307.195 -119.165 307.525 -118.835 ;
        RECT 307.195 -120.525 307.525 -120.195 ;
        RECT 307.195 -121.885 307.525 -121.555 ;
        RECT 307.195 -123.245 307.525 -122.915 ;
        RECT 307.195 -124.605 307.525 -124.275 ;
        RECT 307.195 -125.965 307.525 -125.635 ;
        RECT 307.195 -127.325 307.525 -126.995 ;
        RECT 307.195 -128.685 307.525 -128.355 ;
        RECT 307.195 -130.045 307.525 -129.715 ;
        RECT 307.195 -131.405 307.525 -131.075 ;
        RECT 307.195 -132.765 307.525 -132.435 ;
        RECT 307.195 -134.125 307.525 -133.795 ;
        RECT 307.195 -135.485 307.525 -135.155 ;
        RECT 307.195 -136.845 307.525 -136.515 ;
        RECT 307.195 -138.205 307.525 -137.875 ;
        RECT 307.195 -139.565 307.525 -139.235 ;
        RECT 307.195 -140.925 307.525 -140.595 ;
        RECT 307.195 -142.285 307.525 -141.955 ;
        RECT 307.195 -143.645 307.525 -143.315 ;
        RECT 307.195 -145.005 307.525 -144.675 ;
        RECT 307.195 -146.365 307.525 -146.035 ;
        RECT 307.195 -147.725 307.525 -147.395 ;
        RECT 307.195 -149.085 307.525 -148.755 ;
        RECT 307.195 -150.445 307.525 -150.115 ;
        RECT 307.195 -151.805 307.525 -151.475 ;
        RECT 307.195 -153.165 307.525 -152.835 ;
        RECT 307.195 -154.525 307.525 -154.195 ;
        RECT 307.195 -155.885 307.525 -155.555 ;
        RECT 307.195 -157.245 307.525 -156.915 ;
        RECT 307.195 -158.605 307.525 -158.275 ;
        RECT 307.195 -159.965 307.525 -159.635 ;
        RECT 307.195 -161.325 307.525 -160.995 ;
        RECT 307.195 -162.685 307.525 -162.355 ;
        RECT 307.195 -164.045 307.525 -163.715 ;
        RECT 307.195 -165.405 307.525 -165.075 ;
        RECT 307.195 -166.765 307.525 -166.435 ;
        RECT 307.195 -168.125 307.525 -167.795 ;
        RECT 307.195 -169.485 307.525 -169.155 ;
        RECT 307.195 -170.845 307.525 -170.515 ;
        RECT 307.195 -172.205 307.525 -171.875 ;
        RECT 307.195 -173.565 307.525 -173.235 ;
        RECT 307.195 -174.925 307.525 -174.595 ;
        RECT 307.195 -176.285 307.525 -175.955 ;
        RECT 307.195 -177.645 307.525 -177.315 ;
        RECT 307.195 -179.005 307.525 -178.675 ;
        RECT 307.195 -184.65 307.525 -183.52 ;
        RECT 307.2 -184.765 307.52 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.86 -98.075 308.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.555 244.04 308.885 245.17 ;
        RECT 308.555 239.875 308.885 240.205 ;
        RECT 308.555 238.515 308.885 238.845 ;
        RECT 308.555 237.155 308.885 237.485 ;
        RECT 308.56 237.155 308.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.915 244.04 310.245 245.17 ;
        RECT 309.915 239.875 310.245 240.205 ;
        RECT 309.915 238.515 310.245 238.845 ;
        RECT 309.915 237.155 310.245 237.485 ;
        RECT 309.92 237.155 310.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.915 -0.845 310.245 -0.515 ;
        RECT 309.915 -2.205 310.245 -1.875 ;
        RECT 309.915 -3.565 310.245 -3.235 ;
        RECT 309.92 -3.565 310.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.275 244.04 311.605 245.17 ;
        RECT 311.275 239.875 311.605 240.205 ;
        RECT 311.275 238.515 311.605 238.845 ;
        RECT 311.275 237.155 311.605 237.485 ;
        RECT 311.28 237.155 311.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.275 -0.845 311.605 -0.515 ;
        RECT 311.275 -2.205 311.605 -1.875 ;
        RECT 311.275 -3.565 311.605 -3.235 ;
        RECT 311.28 -3.565 311.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.635 244.04 312.965 245.17 ;
        RECT 312.635 239.875 312.965 240.205 ;
        RECT 312.635 238.515 312.965 238.845 ;
        RECT 312.635 237.155 312.965 237.485 ;
        RECT 312.64 237.155 312.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.635 -0.845 312.965 -0.515 ;
        RECT 312.635 -2.205 312.965 -1.875 ;
        RECT 312.635 -3.565 312.965 -3.235 ;
        RECT 312.64 -3.565 312.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 312.635 -170.845 312.965 -170.515 ;
        RECT 312.635 -172.205 312.965 -171.875 ;
        RECT 312.635 -173.565 312.965 -173.235 ;
        RECT 312.635 -174.925 312.965 -174.595 ;
        RECT 312.635 -176.285 312.965 -175.955 ;
        RECT 312.635 -177.645 312.965 -177.315 ;
        RECT 312.635 -179.005 312.965 -178.675 ;
        RECT 312.635 -184.65 312.965 -183.52 ;
        RECT 312.64 -184.765 312.96 -95.04 ;
        RECT 312.635 -96.045 312.965 -95.715 ;
        RECT 312.635 -97.405 312.965 -97.075 ;
        RECT 312.635 -98.765 312.965 -98.435 ;
        RECT 312.635 -100.125 312.965 -99.795 ;
        RECT 312.635 -101.485 312.965 -101.155 ;
        RECT 312.635 -102.845 312.965 -102.515 ;
        RECT 312.635 -104.205 312.965 -103.875 ;
        RECT 312.635 -105.565 312.965 -105.235 ;
        RECT 312.635 -106.925 312.965 -106.595 ;
        RECT 312.635 -108.285 312.965 -107.955 ;
        RECT 312.635 -109.645 312.965 -109.315 ;
        RECT 312.635 -111.005 312.965 -110.675 ;
        RECT 312.635 -112.365 312.965 -112.035 ;
        RECT 312.635 -113.725 312.965 -113.395 ;
        RECT 312.635 -115.085 312.965 -114.755 ;
        RECT 312.635 -116.445 312.965 -116.115 ;
        RECT 312.635 -117.805 312.965 -117.475 ;
        RECT 312.635 -119.165 312.965 -118.835 ;
        RECT 312.635 -120.525 312.965 -120.195 ;
        RECT 312.635 -121.885 312.965 -121.555 ;
        RECT 312.635 -123.245 312.965 -122.915 ;
        RECT 312.635 -124.605 312.965 -124.275 ;
        RECT 312.635 -125.965 312.965 -125.635 ;
        RECT 312.635 -127.325 312.965 -126.995 ;
        RECT 312.635 -128.685 312.965 -128.355 ;
        RECT 312.635 -130.045 312.965 -129.715 ;
        RECT 312.635 -131.405 312.965 -131.075 ;
        RECT 312.635 -132.765 312.965 -132.435 ;
        RECT 312.635 -134.125 312.965 -133.795 ;
        RECT 312.635 -135.485 312.965 -135.155 ;
        RECT 312.635 -136.845 312.965 -136.515 ;
        RECT 312.635 -138.205 312.965 -137.875 ;
        RECT 312.635 -139.565 312.965 -139.235 ;
        RECT 312.635 -140.925 312.965 -140.595 ;
        RECT 312.635 -142.285 312.965 -141.955 ;
        RECT 312.635 -143.645 312.965 -143.315 ;
        RECT 312.635 -145.005 312.965 -144.675 ;
        RECT 312.635 -146.365 312.965 -146.035 ;
        RECT 312.635 -147.725 312.965 -147.395 ;
        RECT 312.635 -149.085 312.965 -148.755 ;
        RECT 312.635 -150.445 312.965 -150.115 ;
        RECT 312.635 -151.805 312.965 -151.475 ;
        RECT 312.635 -153.165 312.965 -152.835 ;
        RECT 312.635 -154.525 312.965 -154.195 ;
        RECT 312.635 -155.885 312.965 -155.555 ;
        RECT 312.635 -157.245 312.965 -156.915 ;
        RECT 312.635 -158.605 312.965 -158.275 ;
        RECT 312.635 -159.965 312.965 -159.635 ;
        RECT 312.635 -161.325 312.965 -160.995 ;
        RECT 312.635 -162.685 312.965 -162.355 ;
        RECT 312.635 -164.045 312.965 -163.715 ;
        RECT 312.635 -165.405 312.965 -165.075 ;
        RECT 312.635 -166.765 312.965 -166.435 ;
        RECT 312.635 -168.125 312.965 -167.795 ;
        RECT 312.635 -169.485 312.965 -169.155 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.955 244.04 261.285 245.17 ;
        RECT 260.955 239.875 261.285 240.205 ;
        RECT 260.955 238.515 261.285 238.845 ;
        RECT 260.955 237.155 261.285 237.485 ;
        RECT 260.96 237.155 261.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.955 -0.845 261.285 -0.515 ;
        RECT 260.955 -2.205 261.285 -1.875 ;
        RECT 260.955 -3.565 261.285 -3.235 ;
        RECT 260.96 -3.565 261.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.955 -96.045 261.285 -95.715 ;
        RECT 260.955 -97.405 261.285 -97.075 ;
        RECT 260.955 -98.765 261.285 -98.435 ;
        RECT 260.955 -100.125 261.285 -99.795 ;
        RECT 260.955 -101.485 261.285 -101.155 ;
        RECT 260.955 -102.845 261.285 -102.515 ;
        RECT 260.955 -104.205 261.285 -103.875 ;
        RECT 260.955 -105.565 261.285 -105.235 ;
        RECT 260.955 -106.925 261.285 -106.595 ;
        RECT 260.955 -108.285 261.285 -107.955 ;
        RECT 260.955 -109.645 261.285 -109.315 ;
        RECT 260.955 -111.005 261.285 -110.675 ;
        RECT 260.955 -112.365 261.285 -112.035 ;
        RECT 260.955 -113.725 261.285 -113.395 ;
        RECT 260.955 -115.085 261.285 -114.755 ;
        RECT 260.955 -116.445 261.285 -116.115 ;
        RECT 260.955 -117.805 261.285 -117.475 ;
        RECT 260.955 -119.165 261.285 -118.835 ;
        RECT 260.955 -120.525 261.285 -120.195 ;
        RECT 260.955 -121.885 261.285 -121.555 ;
        RECT 260.955 -123.245 261.285 -122.915 ;
        RECT 260.955 -124.605 261.285 -124.275 ;
        RECT 260.955 -125.965 261.285 -125.635 ;
        RECT 260.955 -127.325 261.285 -126.995 ;
        RECT 260.955 -128.685 261.285 -128.355 ;
        RECT 260.955 -130.045 261.285 -129.715 ;
        RECT 260.955 -131.405 261.285 -131.075 ;
        RECT 260.955 -132.765 261.285 -132.435 ;
        RECT 260.955 -134.125 261.285 -133.795 ;
        RECT 260.955 -135.485 261.285 -135.155 ;
        RECT 260.955 -136.845 261.285 -136.515 ;
        RECT 260.955 -138.205 261.285 -137.875 ;
        RECT 260.955 -139.565 261.285 -139.235 ;
        RECT 260.955 -140.925 261.285 -140.595 ;
        RECT 260.955 -142.285 261.285 -141.955 ;
        RECT 260.955 -143.645 261.285 -143.315 ;
        RECT 260.955 -145.005 261.285 -144.675 ;
        RECT 260.955 -146.365 261.285 -146.035 ;
        RECT 260.955 -147.725 261.285 -147.395 ;
        RECT 260.955 -149.085 261.285 -148.755 ;
        RECT 260.955 -150.445 261.285 -150.115 ;
        RECT 260.955 -151.805 261.285 -151.475 ;
        RECT 260.955 -153.165 261.285 -152.835 ;
        RECT 260.955 -154.525 261.285 -154.195 ;
        RECT 260.955 -155.885 261.285 -155.555 ;
        RECT 260.955 -157.245 261.285 -156.915 ;
        RECT 260.955 -158.605 261.285 -158.275 ;
        RECT 260.955 -159.965 261.285 -159.635 ;
        RECT 260.955 -161.325 261.285 -160.995 ;
        RECT 260.955 -162.685 261.285 -162.355 ;
        RECT 260.955 -164.045 261.285 -163.715 ;
        RECT 260.955 -165.405 261.285 -165.075 ;
        RECT 260.955 -166.765 261.285 -166.435 ;
        RECT 260.955 -168.125 261.285 -167.795 ;
        RECT 260.955 -169.485 261.285 -169.155 ;
        RECT 260.955 -170.845 261.285 -170.515 ;
        RECT 260.955 -172.205 261.285 -171.875 ;
        RECT 260.955 -173.565 261.285 -173.235 ;
        RECT 260.955 -174.925 261.285 -174.595 ;
        RECT 260.955 -176.285 261.285 -175.955 ;
        RECT 260.955 -177.645 261.285 -177.315 ;
        RECT 260.955 -179.005 261.285 -178.675 ;
        RECT 260.955 -184.65 261.285 -183.52 ;
        RECT 260.96 -184.765 261.28 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.315 244.04 262.645 245.17 ;
        RECT 262.315 239.875 262.645 240.205 ;
        RECT 262.315 238.515 262.645 238.845 ;
        RECT 262.315 237.155 262.645 237.485 ;
        RECT 262.32 237.155 262.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.315 -0.845 262.645 -0.515 ;
        RECT 262.315 -2.205 262.645 -1.875 ;
        RECT 262.315 -3.565 262.645 -3.235 ;
        RECT 262.32 -3.565 262.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.315 -96.045 262.645 -95.715 ;
        RECT 262.315 -97.405 262.645 -97.075 ;
        RECT 262.315 -98.765 262.645 -98.435 ;
        RECT 262.315 -100.125 262.645 -99.795 ;
        RECT 262.315 -101.485 262.645 -101.155 ;
        RECT 262.315 -102.845 262.645 -102.515 ;
        RECT 262.315 -104.205 262.645 -103.875 ;
        RECT 262.315 -105.565 262.645 -105.235 ;
        RECT 262.315 -106.925 262.645 -106.595 ;
        RECT 262.315 -108.285 262.645 -107.955 ;
        RECT 262.315 -109.645 262.645 -109.315 ;
        RECT 262.315 -111.005 262.645 -110.675 ;
        RECT 262.315 -112.365 262.645 -112.035 ;
        RECT 262.315 -113.725 262.645 -113.395 ;
        RECT 262.315 -115.085 262.645 -114.755 ;
        RECT 262.315 -116.445 262.645 -116.115 ;
        RECT 262.315 -117.805 262.645 -117.475 ;
        RECT 262.315 -119.165 262.645 -118.835 ;
        RECT 262.315 -120.525 262.645 -120.195 ;
        RECT 262.315 -121.885 262.645 -121.555 ;
        RECT 262.315 -123.245 262.645 -122.915 ;
        RECT 262.315 -124.605 262.645 -124.275 ;
        RECT 262.315 -125.965 262.645 -125.635 ;
        RECT 262.315 -127.325 262.645 -126.995 ;
        RECT 262.315 -128.685 262.645 -128.355 ;
        RECT 262.315 -130.045 262.645 -129.715 ;
        RECT 262.315 -131.405 262.645 -131.075 ;
        RECT 262.315 -132.765 262.645 -132.435 ;
        RECT 262.315 -134.125 262.645 -133.795 ;
        RECT 262.315 -135.485 262.645 -135.155 ;
        RECT 262.315 -136.845 262.645 -136.515 ;
        RECT 262.315 -138.205 262.645 -137.875 ;
        RECT 262.315 -139.565 262.645 -139.235 ;
        RECT 262.315 -140.925 262.645 -140.595 ;
        RECT 262.315 -142.285 262.645 -141.955 ;
        RECT 262.315 -143.645 262.645 -143.315 ;
        RECT 262.315 -145.005 262.645 -144.675 ;
        RECT 262.315 -146.365 262.645 -146.035 ;
        RECT 262.315 -147.725 262.645 -147.395 ;
        RECT 262.315 -149.085 262.645 -148.755 ;
        RECT 262.315 -150.445 262.645 -150.115 ;
        RECT 262.315 -151.805 262.645 -151.475 ;
        RECT 262.315 -153.165 262.645 -152.835 ;
        RECT 262.315 -154.525 262.645 -154.195 ;
        RECT 262.315 -155.885 262.645 -155.555 ;
        RECT 262.315 -157.245 262.645 -156.915 ;
        RECT 262.315 -158.605 262.645 -158.275 ;
        RECT 262.315 -159.965 262.645 -159.635 ;
        RECT 262.315 -161.325 262.645 -160.995 ;
        RECT 262.315 -162.685 262.645 -162.355 ;
        RECT 262.315 -164.045 262.645 -163.715 ;
        RECT 262.315 -165.405 262.645 -165.075 ;
        RECT 262.315 -166.765 262.645 -166.435 ;
        RECT 262.315 -168.125 262.645 -167.795 ;
        RECT 262.315 -169.485 262.645 -169.155 ;
        RECT 262.315 -170.845 262.645 -170.515 ;
        RECT 262.315 -172.205 262.645 -171.875 ;
        RECT 262.315 -173.565 262.645 -173.235 ;
        RECT 262.315 -174.925 262.645 -174.595 ;
        RECT 262.315 -176.285 262.645 -175.955 ;
        RECT 262.315 -177.645 262.645 -177.315 ;
        RECT 262.315 -179.005 262.645 -178.675 ;
        RECT 262.315 -184.65 262.645 -183.52 ;
        RECT 262.32 -184.765 262.64 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.675 244.04 264.005 245.17 ;
        RECT 263.675 239.875 264.005 240.205 ;
        RECT 263.675 238.515 264.005 238.845 ;
        RECT 263.675 237.155 264.005 237.485 ;
        RECT 263.68 237.155 264 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 263.675 -98.765 264.005 -98.435 ;
        RECT 263.675 -100.125 264.005 -99.795 ;
        RECT 263.675 -101.485 264.005 -101.155 ;
        RECT 263.675 -102.845 264.005 -102.515 ;
        RECT 263.675 -104.205 264.005 -103.875 ;
        RECT 263.675 -105.565 264.005 -105.235 ;
        RECT 263.675 -106.925 264.005 -106.595 ;
        RECT 263.675 -108.285 264.005 -107.955 ;
        RECT 263.675 -109.645 264.005 -109.315 ;
        RECT 263.675 -111.005 264.005 -110.675 ;
        RECT 263.675 -112.365 264.005 -112.035 ;
        RECT 263.675 -113.725 264.005 -113.395 ;
        RECT 263.675 -115.085 264.005 -114.755 ;
        RECT 263.675 -116.445 264.005 -116.115 ;
        RECT 263.675 -117.805 264.005 -117.475 ;
        RECT 263.675 -119.165 264.005 -118.835 ;
        RECT 263.675 -120.525 264.005 -120.195 ;
        RECT 263.675 -121.885 264.005 -121.555 ;
        RECT 263.675 -123.245 264.005 -122.915 ;
        RECT 263.675 -124.605 264.005 -124.275 ;
        RECT 263.675 -125.965 264.005 -125.635 ;
        RECT 263.675 -127.325 264.005 -126.995 ;
        RECT 263.675 -128.685 264.005 -128.355 ;
        RECT 263.675 -130.045 264.005 -129.715 ;
        RECT 263.675 -131.405 264.005 -131.075 ;
        RECT 263.675 -132.765 264.005 -132.435 ;
        RECT 263.675 -134.125 264.005 -133.795 ;
        RECT 263.675 -135.485 264.005 -135.155 ;
        RECT 263.675 -136.845 264.005 -136.515 ;
        RECT 263.675 -138.205 264.005 -137.875 ;
        RECT 263.675 -139.565 264.005 -139.235 ;
        RECT 263.675 -140.925 264.005 -140.595 ;
        RECT 263.675 -142.285 264.005 -141.955 ;
        RECT 263.675 -143.645 264.005 -143.315 ;
        RECT 263.675 -145.005 264.005 -144.675 ;
        RECT 263.675 -146.365 264.005 -146.035 ;
        RECT 263.675 -147.725 264.005 -147.395 ;
        RECT 263.675 -149.085 264.005 -148.755 ;
        RECT 263.675 -150.445 264.005 -150.115 ;
        RECT 263.675 -151.805 264.005 -151.475 ;
        RECT 263.675 -153.165 264.005 -152.835 ;
        RECT 263.675 -154.525 264.005 -154.195 ;
        RECT 263.675 -155.885 264.005 -155.555 ;
        RECT 263.675 -157.245 264.005 -156.915 ;
        RECT 263.675 -158.605 264.005 -158.275 ;
        RECT 263.675 -159.965 264.005 -159.635 ;
        RECT 263.675 -161.325 264.005 -160.995 ;
        RECT 263.675 -162.685 264.005 -162.355 ;
        RECT 263.675 -164.045 264.005 -163.715 ;
        RECT 263.675 -165.405 264.005 -165.075 ;
        RECT 263.675 -166.765 264.005 -166.435 ;
        RECT 263.675 -168.125 264.005 -167.795 ;
        RECT 263.675 -169.485 264.005 -169.155 ;
        RECT 263.675 -170.845 264.005 -170.515 ;
        RECT 263.675 -172.205 264.005 -171.875 ;
        RECT 263.675 -173.565 264.005 -173.235 ;
        RECT 263.675 -174.925 264.005 -174.595 ;
        RECT 263.675 -176.285 264.005 -175.955 ;
        RECT 263.675 -177.645 264.005 -177.315 ;
        RECT 263.675 -179.005 264.005 -178.675 ;
        RECT 263.675 -184.65 264.005 -183.52 ;
        RECT 263.68 -184.765 264 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.26 -98.075 264.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.035 244.04 265.365 245.17 ;
        RECT 265.035 239.875 265.365 240.205 ;
        RECT 265.035 238.515 265.365 238.845 ;
        RECT 265.035 237.155 265.365 237.485 ;
        RECT 265.04 237.155 265.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.395 244.04 266.725 245.17 ;
        RECT 266.395 239.875 266.725 240.205 ;
        RECT 266.395 238.515 266.725 238.845 ;
        RECT 266.395 237.155 266.725 237.485 ;
        RECT 266.4 237.155 266.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.395 -0.845 266.725 -0.515 ;
        RECT 266.395 -2.205 266.725 -1.875 ;
        RECT 266.395 -3.565 266.725 -3.235 ;
        RECT 266.4 -3.565 266.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 266.395 -96.045 266.725 -95.715 ;
        RECT 266.395 -97.405 266.725 -97.075 ;
        RECT 266.395 -98.765 266.725 -98.435 ;
        RECT 266.395 -100.125 266.725 -99.795 ;
        RECT 266.395 -101.485 266.725 -101.155 ;
        RECT 266.395 -102.845 266.725 -102.515 ;
        RECT 266.395 -104.205 266.725 -103.875 ;
        RECT 266.395 -105.565 266.725 -105.235 ;
        RECT 266.395 -106.925 266.725 -106.595 ;
        RECT 266.395 -108.285 266.725 -107.955 ;
        RECT 266.395 -109.645 266.725 -109.315 ;
        RECT 266.395 -111.005 266.725 -110.675 ;
        RECT 266.395 -112.365 266.725 -112.035 ;
        RECT 266.395 -113.725 266.725 -113.395 ;
        RECT 266.395 -115.085 266.725 -114.755 ;
        RECT 266.395 -116.445 266.725 -116.115 ;
        RECT 266.395 -117.805 266.725 -117.475 ;
        RECT 266.395 -119.165 266.725 -118.835 ;
        RECT 266.395 -120.525 266.725 -120.195 ;
        RECT 266.395 -121.885 266.725 -121.555 ;
        RECT 266.395 -123.245 266.725 -122.915 ;
        RECT 266.395 -124.605 266.725 -124.275 ;
        RECT 266.395 -125.965 266.725 -125.635 ;
        RECT 266.395 -127.325 266.725 -126.995 ;
        RECT 266.395 -128.685 266.725 -128.355 ;
        RECT 266.395 -130.045 266.725 -129.715 ;
        RECT 266.395 -131.405 266.725 -131.075 ;
        RECT 266.395 -132.765 266.725 -132.435 ;
        RECT 266.395 -134.125 266.725 -133.795 ;
        RECT 266.395 -135.485 266.725 -135.155 ;
        RECT 266.395 -136.845 266.725 -136.515 ;
        RECT 266.395 -138.205 266.725 -137.875 ;
        RECT 266.395 -139.565 266.725 -139.235 ;
        RECT 266.395 -140.925 266.725 -140.595 ;
        RECT 266.395 -142.285 266.725 -141.955 ;
        RECT 266.395 -143.645 266.725 -143.315 ;
        RECT 266.395 -145.005 266.725 -144.675 ;
        RECT 266.395 -146.365 266.725 -146.035 ;
        RECT 266.395 -147.725 266.725 -147.395 ;
        RECT 266.395 -149.085 266.725 -148.755 ;
        RECT 266.395 -150.445 266.725 -150.115 ;
        RECT 266.395 -151.805 266.725 -151.475 ;
        RECT 266.395 -153.165 266.725 -152.835 ;
        RECT 266.395 -154.525 266.725 -154.195 ;
        RECT 266.395 -155.885 266.725 -155.555 ;
        RECT 266.395 -157.245 266.725 -156.915 ;
        RECT 266.395 -158.605 266.725 -158.275 ;
        RECT 266.395 -159.965 266.725 -159.635 ;
        RECT 266.395 -161.325 266.725 -160.995 ;
        RECT 266.395 -162.685 266.725 -162.355 ;
        RECT 266.395 -164.045 266.725 -163.715 ;
        RECT 266.395 -165.405 266.725 -165.075 ;
        RECT 266.395 -166.765 266.725 -166.435 ;
        RECT 266.395 -168.125 266.725 -167.795 ;
        RECT 266.395 -169.485 266.725 -169.155 ;
        RECT 266.395 -170.845 266.725 -170.515 ;
        RECT 266.395 -172.205 266.725 -171.875 ;
        RECT 266.395 -173.565 266.725 -173.235 ;
        RECT 266.395 -174.925 266.725 -174.595 ;
        RECT 266.395 -176.285 266.725 -175.955 ;
        RECT 266.395 -177.645 266.725 -177.315 ;
        RECT 266.395 -179.005 266.725 -178.675 ;
        RECT 266.395 -184.65 266.725 -183.52 ;
        RECT 266.4 -184.765 266.72 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.755 244.04 268.085 245.17 ;
        RECT 267.755 239.875 268.085 240.205 ;
        RECT 267.755 238.515 268.085 238.845 ;
        RECT 267.755 237.155 268.085 237.485 ;
        RECT 267.76 237.155 268.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.755 -0.845 268.085 -0.515 ;
        RECT 267.755 -2.205 268.085 -1.875 ;
        RECT 267.755 -3.565 268.085 -3.235 ;
        RECT 267.76 -3.565 268.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.115 244.04 269.445 245.17 ;
        RECT 269.115 239.875 269.445 240.205 ;
        RECT 269.115 238.515 269.445 238.845 ;
        RECT 269.115 237.155 269.445 237.485 ;
        RECT 269.12 237.155 269.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.115 -0.845 269.445 -0.515 ;
        RECT 269.115 -2.205 269.445 -1.875 ;
        RECT 269.115 -3.565 269.445 -3.235 ;
        RECT 269.12 -3.565 269.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.115 -96.045 269.445 -95.715 ;
        RECT 269.115 -97.405 269.445 -97.075 ;
        RECT 269.115 -98.765 269.445 -98.435 ;
        RECT 269.115 -100.125 269.445 -99.795 ;
        RECT 269.115 -101.485 269.445 -101.155 ;
        RECT 269.115 -102.845 269.445 -102.515 ;
        RECT 269.115 -104.205 269.445 -103.875 ;
        RECT 269.115 -105.565 269.445 -105.235 ;
        RECT 269.115 -106.925 269.445 -106.595 ;
        RECT 269.115 -108.285 269.445 -107.955 ;
        RECT 269.115 -109.645 269.445 -109.315 ;
        RECT 269.115 -111.005 269.445 -110.675 ;
        RECT 269.115 -112.365 269.445 -112.035 ;
        RECT 269.115 -113.725 269.445 -113.395 ;
        RECT 269.115 -115.085 269.445 -114.755 ;
        RECT 269.115 -116.445 269.445 -116.115 ;
        RECT 269.115 -117.805 269.445 -117.475 ;
        RECT 269.115 -119.165 269.445 -118.835 ;
        RECT 269.115 -120.525 269.445 -120.195 ;
        RECT 269.115 -121.885 269.445 -121.555 ;
        RECT 269.115 -123.245 269.445 -122.915 ;
        RECT 269.115 -124.605 269.445 -124.275 ;
        RECT 269.115 -125.965 269.445 -125.635 ;
        RECT 269.115 -127.325 269.445 -126.995 ;
        RECT 269.115 -128.685 269.445 -128.355 ;
        RECT 269.115 -130.045 269.445 -129.715 ;
        RECT 269.115 -131.405 269.445 -131.075 ;
        RECT 269.115 -132.765 269.445 -132.435 ;
        RECT 269.115 -134.125 269.445 -133.795 ;
        RECT 269.115 -135.485 269.445 -135.155 ;
        RECT 269.115 -136.845 269.445 -136.515 ;
        RECT 269.115 -138.205 269.445 -137.875 ;
        RECT 269.115 -139.565 269.445 -139.235 ;
        RECT 269.115 -140.925 269.445 -140.595 ;
        RECT 269.115 -142.285 269.445 -141.955 ;
        RECT 269.115 -143.645 269.445 -143.315 ;
        RECT 269.115 -145.005 269.445 -144.675 ;
        RECT 269.115 -146.365 269.445 -146.035 ;
        RECT 269.115 -147.725 269.445 -147.395 ;
        RECT 269.115 -149.085 269.445 -148.755 ;
        RECT 269.115 -150.445 269.445 -150.115 ;
        RECT 269.115 -151.805 269.445 -151.475 ;
        RECT 269.115 -153.165 269.445 -152.835 ;
        RECT 269.115 -154.525 269.445 -154.195 ;
        RECT 269.115 -155.885 269.445 -155.555 ;
        RECT 269.115 -157.245 269.445 -156.915 ;
        RECT 269.115 -158.605 269.445 -158.275 ;
        RECT 269.115 -159.965 269.445 -159.635 ;
        RECT 269.115 -161.325 269.445 -160.995 ;
        RECT 269.115 -162.685 269.445 -162.355 ;
        RECT 269.115 -164.045 269.445 -163.715 ;
        RECT 269.115 -165.405 269.445 -165.075 ;
        RECT 269.115 -166.765 269.445 -166.435 ;
        RECT 269.115 -168.125 269.445 -167.795 ;
        RECT 269.115 -169.485 269.445 -169.155 ;
        RECT 269.115 -170.845 269.445 -170.515 ;
        RECT 269.115 -172.205 269.445 -171.875 ;
        RECT 269.115 -173.565 269.445 -173.235 ;
        RECT 269.115 -174.925 269.445 -174.595 ;
        RECT 269.115 -176.285 269.445 -175.955 ;
        RECT 269.115 -177.645 269.445 -177.315 ;
        RECT 269.115 -179.005 269.445 -178.675 ;
        RECT 269.115 -184.65 269.445 -183.52 ;
        RECT 269.12 -184.765 269.44 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.475 244.04 270.805 245.17 ;
        RECT 270.475 239.875 270.805 240.205 ;
        RECT 270.475 238.515 270.805 238.845 ;
        RECT 270.475 237.155 270.805 237.485 ;
        RECT 270.48 237.155 270.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.475 -0.845 270.805 -0.515 ;
        RECT 270.475 -2.205 270.805 -1.875 ;
        RECT 270.475 -3.565 270.805 -3.235 ;
        RECT 270.48 -3.565 270.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 270.475 -96.045 270.805 -95.715 ;
        RECT 270.475 -97.405 270.805 -97.075 ;
        RECT 270.475 -98.765 270.805 -98.435 ;
        RECT 270.475 -100.125 270.805 -99.795 ;
        RECT 270.475 -101.485 270.805 -101.155 ;
        RECT 270.475 -102.845 270.805 -102.515 ;
        RECT 270.475 -104.205 270.805 -103.875 ;
        RECT 270.475 -105.565 270.805 -105.235 ;
        RECT 270.475 -106.925 270.805 -106.595 ;
        RECT 270.475 -108.285 270.805 -107.955 ;
        RECT 270.475 -109.645 270.805 -109.315 ;
        RECT 270.475 -111.005 270.805 -110.675 ;
        RECT 270.475 -112.365 270.805 -112.035 ;
        RECT 270.475 -113.725 270.805 -113.395 ;
        RECT 270.475 -115.085 270.805 -114.755 ;
        RECT 270.475 -116.445 270.805 -116.115 ;
        RECT 270.475 -117.805 270.805 -117.475 ;
        RECT 270.475 -119.165 270.805 -118.835 ;
        RECT 270.475 -120.525 270.805 -120.195 ;
        RECT 270.475 -121.885 270.805 -121.555 ;
        RECT 270.475 -123.245 270.805 -122.915 ;
        RECT 270.475 -124.605 270.805 -124.275 ;
        RECT 270.475 -125.965 270.805 -125.635 ;
        RECT 270.475 -127.325 270.805 -126.995 ;
        RECT 270.475 -128.685 270.805 -128.355 ;
        RECT 270.475 -130.045 270.805 -129.715 ;
        RECT 270.475 -131.405 270.805 -131.075 ;
        RECT 270.475 -132.765 270.805 -132.435 ;
        RECT 270.475 -134.125 270.805 -133.795 ;
        RECT 270.475 -135.485 270.805 -135.155 ;
        RECT 270.475 -136.845 270.805 -136.515 ;
        RECT 270.475 -138.205 270.805 -137.875 ;
        RECT 270.475 -139.565 270.805 -139.235 ;
        RECT 270.475 -140.925 270.805 -140.595 ;
        RECT 270.475 -142.285 270.805 -141.955 ;
        RECT 270.475 -143.645 270.805 -143.315 ;
        RECT 270.475 -145.005 270.805 -144.675 ;
        RECT 270.475 -146.365 270.805 -146.035 ;
        RECT 270.475 -147.725 270.805 -147.395 ;
        RECT 270.475 -149.085 270.805 -148.755 ;
        RECT 270.475 -150.445 270.805 -150.115 ;
        RECT 270.475 -151.805 270.805 -151.475 ;
        RECT 270.475 -153.165 270.805 -152.835 ;
        RECT 270.475 -154.525 270.805 -154.195 ;
        RECT 270.475 -155.885 270.805 -155.555 ;
        RECT 270.475 -157.245 270.805 -156.915 ;
        RECT 270.475 -158.605 270.805 -158.275 ;
        RECT 270.475 -159.965 270.805 -159.635 ;
        RECT 270.475 -161.325 270.805 -160.995 ;
        RECT 270.475 -162.685 270.805 -162.355 ;
        RECT 270.475 -164.045 270.805 -163.715 ;
        RECT 270.475 -165.405 270.805 -165.075 ;
        RECT 270.475 -166.765 270.805 -166.435 ;
        RECT 270.475 -168.125 270.805 -167.795 ;
        RECT 270.475 -169.485 270.805 -169.155 ;
        RECT 270.475 -170.845 270.805 -170.515 ;
        RECT 270.475 -172.205 270.805 -171.875 ;
        RECT 270.475 -173.565 270.805 -173.235 ;
        RECT 270.475 -174.925 270.805 -174.595 ;
        RECT 270.475 -176.285 270.805 -175.955 ;
        RECT 270.475 -177.645 270.805 -177.315 ;
        RECT 270.475 -179.005 270.805 -178.675 ;
        RECT 270.475 -184.65 270.805 -183.52 ;
        RECT 270.48 -184.765 270.8 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.835 244.04 272.165 245.17 ;
        RECT 271.835 239.875 272.165 240.205 ;
        RECT 271.835 238.515 272.165 238.845 ;
        RECT 271.835 237.155 272.165 237.485 ;
        RECT 271.84 237.155 272.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.835 -0.845 272.165 -0.515 ;
        RECT 271.835 -2.205 272.165 -1.875 ;
        RECT 271.835 -3.565 272.165 -3.235 ;
        RECT 271.84 -3.565 272.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.835 -96.045 272.165 -95.715 ;
        RECT 271.835 -97.405 272.165 -97.075 ;
        RECT 271.835 -98.765 272.165 -98.435 ;
        RECT 271.835 -100.125 272.165 -99.795 ;
        RECT 271.835 -101.485 272.165 -101.155 ;
        RECT 271.835 -102.845 272.165 -102.515 ;
        RECT 271.835 -104.205 272.165 -103.875 ;
        RECT 271.835 -105.565 272.165 -105.235 ;
        RECT 271.835 -106.925 272.165 -106.595 ;
        RECT 271.835 -108.285 272.165 -107.955 ;
        RECT 271.835 -109.645 272.165 -109.315 ;
        RECT 271.835 -111.005 272.165 -110.675 ;
        RECT 271.835 -112.365 272.165 -112.035 ;
        RECT 271.835 -113.725 272.165 -113.395 ;
        RECT 271.835 -115.085 272.165 -114.755 ;
        RECT 271.835 -116.445 272.165 -116.115 ;
        RECT 271.835 -117.805 272.165 -117.475 ;
        RECT 271.835 -119.165 272.165 -118.835 ;
        RECT 271.835 -120.525 272.165 -120.195 ;
        RECT 271.835 -121.885 272.165 -121.555 ;
        RECT 271.835 -123.245 272.165 -122.915 ;
        RECT 271.835 -124.605 272.165 -124.275 ;
        RECT 271.835 -125.965 272.165 -125.635 ;
        RECT 271.835 -127.325 272.165 -126.995 ;
        RECT 271.835 -128.685 272.165 -128.355 ;
        RECT 271.835 -130.045 272.165 -129.715 ;
        RECT 271.835 -131.405 272.165 -131.075 ;
        RECT 271.835 -132.765 272.165 -132.435 ;
        RECT 271.835 -134.125 272.165 -133.795 ;
        RECT 271.835 -135.485 272.165 -135.155 ;
        RECT 271.835 -136.845 272.165 -136.515 ;
        RECT 271.835 -138.205 272.165 -137.875 ;
        RECT 271.835 -139.565 272.165 -139.235 ;
        RECT 271.835 -140.925 272.165 -140.595 ;
        RECT 271.835 -142.285 272.165 -141.955 ;
        RECT 271.835 -143.645 272.165 -143.315 ;
        RECT 271.835 -145.005 272.165 -144.675 ;
        RECT 271.835 -146.365 272.165 -146.035 ;
        RECT 271.835 -147.725 272.165 -147.395 ;
        RECT 271.835 -149.085 272.165 -148.755 ;
        RECT 271.835 -150.445 272.165 -150.115 ;
        RECT 271.835 -151.805 272.165 -151.475 ;
        RECT 271.835 -153.165 272.165 -152.835 ;
        RECT 271.835 -154.525 272.165 -154.195 ;
        RECT 271.835 -155.885 272.165 -155.555 ;
        RECT 271.835 -157.245 272.165 -156.915 ;
        RECT 271.835 -158.605 272.165 -158.275 ;
        RECT 271.835 -159.965 272.165 -159.635 ;
        RECT 271.835 -161.325 272.165 -160.995 ;
        RECT 271.835 -162.685 272.165 -162.355 ;
        RECT 271.835 -164.045 272.165 -163.715 ;
        RECT 271.835 -165.405 272.165 -165.075 ;
        RECT 271.835 -166.765 272.165 -166.435 ;
        RECT 271.835 -168.125 272.165 -167.795 ;
        RECT 271.835 -169.485 272.165 -169.155 ;
        RECT 271.835 -170.845 272.165 -170.515 ;
        RECT 271.835 -172.205 272.165 -171.875 ;
        RECT 271.835 -173.565 272.165 -173.235 ;
        RECT 271.835 -174.925 272.165 -174.595 ;
        RECT 271.835 -176.285 272.165 -175.955 ;
        RECT 271.835 -177.645 272.165 -177.315 ;
        RECT 271.835 -179.005 272.165 -178.675 ;
        RECT 271.835 -184.65 272.165 -183.52 ;
        RECT 271.84 -184.765 272.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.195 244.04 273.525 245.17 ;
        RECT 273.195 239.875 273.525 240.205 ;
        RECT 273.195 238.515 273.525 238.845 ;
        RECT 273.195 237.155 273.525 237.485 ;
        RECT 273.2 237.155 273.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.195 -0.845 273.525 -0.515 ;
        RECT 273.195 -2.205 273.525 -1.875 ;
        RECT 273.195 -3.565 273.525 -3.235 ;
        RECT 273.2 -3.565 273.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.195 -96.045 273.525 -95.715 ;
        RECT 273.195 -97.405 273.525 -97.075 ;
        RECT 273.195 -98.765 273.525 -98.435 ;
        RECT 273.195 -100.125 273.525 -99.795 ;
        RECT 273.195 -101.485 273.525 -101.155 ;
        RECT 273.195 -102.845 273.525 -102.515 ;
        RECT 273.195 -104.205 273.525 -103.875 ;
        RECT 273.195 -105.565 273.525 -105.235 ;
        RECT 273.195 -106.925 273.525 -106.595 ;
        RECT 273.195 -108.285 273.525 -107.955 ;
        RECT 273.195 -109.645 273.525 -109.315 ;
        RECT 273.195 -111.005 273.525 -110.675 ;
        RECT 273.195 -112.365 273.525 -112.035 ;
        RECT 273.195 -113.725 273.525 -113.395 ;
        RECT 273.195 -115.085 273.525 -114.755 ;
        RECT 273.195 -116.445 273.525 -116.115 ;
        RECT 273.195 -117.805 273.525 -117.475 ;
        RECT 273.195 -119.165 273.525 -118.835 ;
        RECT 273.195 -120.525 273.525 -120.195 ;
        RECT 273.195 -121.885 273.525 -121.555 ;
        RECT 273.195 -123.245 273.525 -122.915 ;
        RECT 273.195 -124.605 273.525 -124.275 ;
        RECT 273.195 -125.965 273.525 -125.635 ;
        RECT 273.195 -127.325 273.525 -126.995 ;
        RECT 273.195 -128.685 273.525 -128.355 ;
        RECT 273.195 -130.045 273.525 -129.715 ;
        RECT 273.195 -131.405 273.525 -131.075 ;
        RECT 273.195 -132.765 273.525 -132.435 ;
        RECT 273.195 -134.125 273.525 -133.795 ;
        RECT 273.195 -135.485 273.525 -135.155 ;
        RECT 273.195 -136.845 273.525 -136.515 ;
        RECT 273.195 -138.205 273.525 -137.875 ;
        RECT 273.195 -139.565 273.525 -139.235 ;
        RECT 273.195 -140.925 273.525 -140.595 ;
        RECT 273.195 -142.285 273.525 -141.955 ;
        RECT 273.195 -143.645 273.525 -143.315 ;
        RECT 273.195 -145.005 273.525 -144.675 ;
        RECT 273.195 -146.365 273.525 -146.035 ;
        RECT 273.195 -147.725 273.525 -147.395 ;
        RECT 273.195 -149.085 273.525 -148.755 ;
        RECT 273.195 -150.445 273.525 -150.115 ;
        RECT 273.195 -151.805 273.525 -151.475 ;
        RECT 273.195 -153.165 273.525 -152.835 ;
        RECT 273.195 -154.525 273.525 -154.195 ;
        RECT 273.195 -155.885 273.525 -155.555 ;
        RECT 273.195 -157.245 273.525 -156.915 ;
        RECT 273.195 -158.605 273.525 -158.275 ;
        RECT 273.195 -159.965 273.525 -159.635 ;
        RECT 273.195 -161.325 273.525 -160.995 ;
        RECT 273.195 -162.685 273.525 -162.355 ;
        RECT 273.195 -164.045 273.525 -163.715 ;
        RECT 273.195 -165.405 273.525 -165.075 ;
        RECT 273.195 -166.765 273.525 -166.435 ;
        RECT 273.195 -168.125 273.525 -167.795 ;
        RECT 273.195 -169.485 273.525 -169.155 ;
        RECT 273.195 -170.845 273.525 -170.515 ;
        RECT 273.195 -172.205 273.525 -171.875 ;
        RECT 273.195 -173.565 273.525 -173.235 ;
        RECT 273.195 -174.925 273.525 -174.595 ;
        RECT 273.195 -176.285 273.525 -175.955 ;
        RECT 273.195 -177.645 273.525 -177.315 ;
        RECT 273.195 -179.005 273.525 -178.675 ;
        RECT 273.195 -184.65 273.525 -183.52 ;
        RECT 273.2 -184.765 273.52 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.555 244.04 274.885 245.17 ;
        RECT 274.555 239.875 274.885 240.205 ;
        RECT 274.555 238.515 274.885 238.845 ;
        RECT 274.555 237.155 274.885 237.485 ;
        RECT 274.56 237.155 274.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 274.555 -98.765 274.885 -98.435 ;
        RECT 274.555 -100.125 274.885 -99.795 ;
        RECT 274.555 -101.485 274.885 -101.155 ;
        RECT 274.555 -102.845 274.885 -102.515 ;
        RECT 274.555 -104.205 274.885 -103.875 ;
        RECT 274.555 -105.565 274.885 -105.235 ;
        RECT 274.555 -106.925 274.885 -106.595 ;
        RECT 274.555 -108.285 274.885 -107.955 ;
        RECT 274.555 -109.645 274.885 -109.315 ;
        RECT 274.555 -111.005 274.885 -110.675 ;
        RECT 274.555 -112.365 274.885 -112.035 ;
        RECT 274.555 -113.725 274.885 -113.395 ;
        RECT 274.555 -115.085 274.885 -114.755 ;
        RECT 274.555 -116.445 274.885 -116.115 ;
        RECT 274.555 -117.805 274.885 -117.475 ;
        RECT 274.555 -119.165 274.885 -118.835 ;
        RECT 274.555 -120.525 274.885 -120.195 ;
        RECT 274.555 -121.885 274.885 -121.555 ;
        RECT 274.555 -123.245 274.885 -122.915 ;
        RECT 274.555 -124.605 274.885 -124.275 ;
        RECT 274.555 -125.965 274.885 -125.635 ;
        RECT 274.555 -127.325 274.885 -126.995 ;
        RECT 274.555 -128.685 274.885 -128.355 ;
        RECT 274.555 -130.045 274.885 -129.715 ;
        RECT 274.555 -131.405 274.885 -131.075 ;
        RECT 274.555 -132.765 274.885 -132.435 ;
        RECT 274.555 -134.125 274.885 -133.795 ;
        RECT 274.555 -135.485 274.885 -135.155 ;
        RECT 274.555 -136.845 274.885 -136.515 ;
        RECT 274.555 -138.205 274.885 -137.875 ;
        RECT 274.555 -139.565 274.885 -139.235 ;
        RECT 274.555 -140.925 274.885 -140.595 ;
        RECT 274.555 -142.285 274.885 -141.955 ;
        RECT 274.555 -143.645 274.885 -143.315 ;
        RECT 274.555 -145.005 274.885 -144.675 ;
        RECT 274.555 -146.365 274.885 -146.035 ;
        RECT 274.555 -147.725 274.885 -147.395 ;
        RECT 274.555 -149.085 274.885 -148.755 ;
        RECT 274.555 -150.445 274.885 -150.115 ;
        RECT 274.555 -151.805 274.885 -151.475 ;
        RECT 274.555 -153.165 274.885 -152.835 ;
        RECT 274.555 -154.525 274.885 -154.195 ;
        RECT 274.555 -155.885 274.885 -155.555 ;
        RECT 274.555 -157.245 274.885 -156.915 ;
        RECT 274.555 -158.605 274.885 -158.275 ;
        RECT 274.555 -159.965 274.885 -159.635 ;
        RECT 274.555 -161.325 274.885 -160.995 ;
        RECT 274.555 -162.685 274.885 -162.355 ;
        RECT 274.555 -164.045 274.885 -163.715 ;
        RECT 274.555 -165.405 274.885 -165.075 ;
        RECT 274.555 -166.765 274.885 -166.435 ;
        RECT 274.555 -168.125 274.885 -167.795 ;
        RECT 274.555 -169.485 274.885 -169.155 ;
        RECT 274.555 -170.845 274.885 -170.515 ;
        RECT 274.555 -172.205 274.885 -171.875 ;
        RECT 274.555 -173.565 274.885 -173.235 ;
        RECT 274.555 -174.925 274.885 -174.595 ;
        RECT 274.555 -176.285 274.885 -175.955 ;
        RECT 274.555 -177.645 274.885 -177.315 ;
        RECT 274.555 -179.005 274.885 -178.675 ;
        RECT 274.555 -184.65 274.885 -183.52 ;
        RECT 274.56 -184.765 274.88 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.16 -98.075 275.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.915 244.04 276.245 245.17 ;
        RECT 275.915 239.875 276.245 240.205 ;
        RECT 275.915 238.515 276.245 238.845 ;
        RECT 275.915 237.155 276.245 237.485 ;
        RECT 275.92 237.155 276.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.275 244.04 277.605 245.17 ;
        RECT 277.275 239.875 277.605 240.205 ;
        RECT 277.275 238.515 277.605 238.845 ;
        RECT 277.275 237.155 277.605 237.485 ;
        RECT 277.28 237.155 277.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.275 -0.845 277.605 -0.515 ;
        RECT 277.275 -2.205 277.605 -1.875 ;
        RECT 277.275 -3.565 277.605 -3.235 ;
        RECT 277.28 -3.565 277.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.275 -96.045 277.605 -95.715 ;
        RECT 277.275 -97.405 277.605 -97.075 ;
        RECT 277.275 -98.765 277.605 -98.435 ;
        RECT 277.275 -100.125 277.605 -99.795 ;
        RECT 277.275 -101.485 277.605 -101.155 ;
        RECT 277.275 -102.845 277.605 -102.515 ;
        RECT 277.275 -104.205 277.605 -103.875 ;
        RECT 277.275 -105.565 277.605 -105.235 ;
        RECT 277.275 -106.925 277.605 -106.595 ;
        RECT 277.275 -108.285 277.605 -107.955 ;
        RECT 277.275 -109.645 277.605 -109.315 ;
        RECT 277.275 -111.005 277.605 -110.675 ;
        RECT 277.275 -112.365 277.605 -112.035 ;
        RECT 277.275 -113.725 277.605 -113.395 ;
        RECT 277.275 -115.085 277.605 -114.755 ;
        RECT 277.275 -116.445 277.605 -116.115 ;
        RECT 277.275 -117.805 277.605 -117.475 ;
        RECT 277.275 -119.165 277.605 -118.835 ;
        RECT 277.275 -120.525 277.605 -120.195 ;
        RECT 277.275 -121.885 277.605 -121.555 ;
        RECT 277.275 -123.245 277.605 -122.915 ;
        RECT 277.275 -124.605 277.605 -124.275 ;
        RECT 277.275 -125.965 277.605 -125.635 ;
        RECT 277.275 -127.325 277.605 -126.995 ;
        RECT 277.275 -128.685 277.605 -128.355 ;
        RECT 277.275 -130.045 277.605 -129.715 ;
        RECT 277.275 -131.405 277.605 -131.075 ;
        RECT 277.275 -132.765 277.605 -132.435 ;
        RECT 277.275 -134.125 277.605 -133.795 ;
        RECT 277.275 -135.485 277.605 -135.155 ;
        RECT 277.275 -136.845 277.605 -136.515 ;
        RECT 277.275 -138.205 277.605 -137.875 ;
        RECT 277.275 -139.565 277.605 -139.235 ;
        RECT 277.275 -140.925 277.605 -140.595 ;
        RECT 277.275 -142.285 277.605 -141.955 ;
        RECT 277.275 -143.645 277.605 -143.315 ;
        RECT 277.275 -145.005 277.605 -144.675 ;
        RECT 277.275 -146.365 277.605 -146.035 ;
        RECT 277.275 -147.725 277.605 -147.395 ;
        RECT 277.275 -149.085 277.605 -148.755 ;
        RECT 277.275 -150.445 277.605 -150.115 ;
        RECT 277.275 -151.805 277.605 -151.475 ;
        RECT 277.275 -153.165 277.605 -152.835 ;
        RECT 277.275 -154.525 277.605 -154.195 ;
        RECT 277.275 -155.885 277.605 -155.555 ;
        RECT 277.275 -157.245 277.605 -156.915 ;
        RECT 277.275 -158.605 277.605 -158.275 ;
        RECT 277.275 -159.965 277.605 -159.635 ;
        RECT 277.275 -161.325 277.605 -160.995 ;
        RECT 277.275 -162.685 277.605 -162.355 ;
        RECT 277.275 -164.045 277.605 -163.715 ;
        RECT 277.275 -165.405 277.605 -165.075 ;
        RECT 277.275 -166.765 277.605 -166.435 ;
        RECT 277.275 -168.125 277.605 -167.795 ;
        RECT 277.275 -169.485 277.605 -169.155 ;
        RECT 277.275 -170.845 277.605 -170.515 ;
        RECT 277.275 -172.205 277.605 -171.875 ;
        RECT 277.275 -173.565 277.605 -173.235 ;
        RECT 277.275 -174.925 277.605 -174.595 ;
        RECT 277.275 -176.285 277.605 -175.955 ;
        RECT 277.275 -177.645 277.605 -177.315 ;
        RECT 277.275 -179.005 277.605 -178.675 ;
        RECT 277.275 -184.65 277.605 -183.52 ;
        RECT 277.28 -184.765 277.6 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.635 244.04 278.965 245.17 ;
        RECT 278.635 239.875 278.965 240.205 ;
        RECT 278.635 238.515 278.965 238.845 ;
        RECT 278.635 237.155 278.965 237.485 ;
        RECT 278.64 237.155 278.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 278.635 -0.845 278.965 -0.515 ;
        RECT 278.635 -2.205 278.965 -1.875 ;
        RECT 278.635 -3.565 278.965 -3.235 ;
        RECT 278.64 -3.565 278.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.995 244.04 280.325 245.17 ;
        RECT 279.995 239.875 280.325 240.205 ;
        RECT 279.995 238.515 280.325 238.845 ;
        RECT 279.995 237.155 280.325 237.485 ;
        RECT 280 237.155 280.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.995 -0.845 280.325 -0.515 ;
        RECT 279.995 -2.205 280.325 -1.875 ;
        RECT 279.995 -3.565 280.325 -3.235 ;
        RECT 280 -3.565 280.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.995 -96.045 280.325 -95.715 ;
        RECT 279.995 -97.405 280.325 -97.075 ;
        RECT 279.995 -98.765 280.325 -98.435 ;
        RECT 279.995 -100.125 280.325 -99.795 ;
        RECT 279.995 -101.485 280.325 -101.155 ;
        RECT 279.995 -102.845 280.325 -102.515 ;
        RECT 279.995 -104.205 280.325 -103.875 ;
        RECT 279.995 -105.565 280.325 -105.235 ;
        RECT 279.995 -106.925 280.325 -106.595 ;
        RECT 279.995 -108.285 280.325 -107.955 ;
        RECT 279.995 -109.645 280.325 -109.315 ;
        RECT 279.995 -111.005 280.325 -110.675 ;
        RECT 279.995 -112.365 280.325 -112.035 ;
        RECT 279.995 -113.725 280.325 -113.395 ;
        RECT 279.995 -115.085 280.325 -114.755 ;
        RECT 279.995 -116.445 280.325 -116.115 ;
        RECT 279.995 -117.805 280.325 -117.475 ;
        RECT 279.995 -119.165 280.325 -118.835 ;
        RECT 279.995 -120.525 280.325 -120.195 ;
        RECT 279.995 -121.885 280.325 -121.555 ;
        RECT 279.995 -123.245 280.325 -122.915 ;
        RECT 279.995 -124.605 280.325 -124.275 ;
        RECT 279.995 -125.965 280.325 -125.635 ;
        RECT 279.995 -127.325 280.325 -126.995 ;
        RECT 279.995 -128.685 280.325 -128.355 ;
        RECT 279.995 -130.045 280.325 -129.715 ;
        RECT 279.995 -131.405 280.325 -131.075 ;
        RECT 279.995 -132.765 280.325 -132.435 ;
        RECT 279.995 -134.125 280.325 -133.795 ;
        RECT 279.995 -135.485 280.325 -135.155 ;
        RECT 279.995 -136.845 280.325 -136.515 ;
        RECT 279.995 -138.205 280.325 -137.875 ;
        RECT 279.995 -139.565 280.325 -139.235 ;
        RECT 279.995 -140.925 280.325 -140.595 ;
        RECT 279.995 -142.285 280.325 -141.955 ;
        RECT 279.995 -143.645 280.325 -143.315 ;
        RECT 279.995 -145.005 280.325 -144.675 ;
        RECT 279.995 -146.365 280.325 -146.035 ;
        RECT 279.995 -147.725 280.325 -147.395 ;
        RECT 279.995 -149.085 280.325 -148.755 ;
        RECT 279.995 -150.445 280.325 -150.115 ;
        RECT 279.995 -151.805 280.325 -151.475 ;
        RECT 279.995 -153.165 280.325 -152.835 ;
        RECT 279.995 -154.525 280.325 -154.195 ;
        RECT 279.995 -155.885 280.325 -155.555 ;
        RECT 279.995 -157.245 280.325 -156.915 ;
        RECT 279.995 -158.605 280.325 -158.275 ;
        RECT 279.995 -159.965 280.325 -159.635 ;
        RECT 279.995 -161.325 280.325 -160.995 ;
        RECT 279.995 -162.685 280.325 -162.355 ;
        RECT 279.995 -164.045 280.325 -163.715 ;
        RECT 279.995 -165.405 280.325 -165.075 ;
        RECT 279.995 -166.765 280.325 -166.435 ;
        RECT 279.995 -168.125 280.325 -167.795 ;
        RECT 279.995 -169.485 280.325 -169.155 ;
        RECT 279.995 -170.845 280.325 -170.515 ;
        RECT 279.995 -172.205 280.325 -171.875 ;
        RECT 279.995 -173.565 280.325 -173.235 ;
        RECT 279.995 -174.925 280.325 -174.595 ;
        RECT 279.995 -176.285 280.325 -175.955 ;
        RECT 279.995 -177.645 280.325 -177.315 ;
        RECT 279.995 -179.005 280.325 -178.675 ;
        RECT 279.995 -184.65 280.325 -183.52 ;
        RECT 280 -184.765 280.32 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.355 244.04 281.685 245.17 ;
        RECT 281.355 239.875 281.685 240.205 ;
        RECT 281.355 238.515 281.685 238.845 ;
        RECT 281.355 237.155 281.685 237.485 ;
        RECT 281.36 237.155 281.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.355 -0.845 281.685 -0.515 ;
        RECT 281.355 -2.205 281.685 -1.875 ;
        RECT 281.355 -3.565 281.685 -3.235 ;
        RECT 281.36 -3.565 281.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 281.355 -96.045 281.685 -95.715 ;
        RECT 281.355 -97.405 281.685 -97.075 ;
        RECT 281.355 -98.765 281.685 -98.435 ;
        RECT 281.355 -100.125 281.685 -99.795 ;
        RECT 281.355 -101.485 281.685 -101.155 ;
        RECT 281.355 -102.845 281.685 -102.515 ;
        RECT 281.355 -104.205 281.685 -103.875 ;
        RECT 281.355 -105.565 281.685 -105.235 ;
        RECT 281.355 -106.925 281.685 -106.595 ;
        RECT 281.355 -108.285 281.685 -107.955 ;
        RECT 281.355 -109.645 281.685 -109.315 ;
        RECT 281.355 -111.005 281.685 -110.675 ;
        RECT 281.355 -112.365 281.685 -112.035 ;
        RECT 281.355 -113.725 281.685 -113.395 ;
        RECT 281.355 -115.085 281.685 -114.755 ;
        RECT 281.355 -116.445 281.685 -116.115 ;
        RECT 281.355 -117.805 281.685 -117.475 ;
        RECT 281.355 -119.165 281.685 -118.835 ;
        RECT 281.355 -120.525 281.685 -120.195 ;
        RECT 281.355 -121.885 281.685 -121.555 ;
        RECT 281.355 -123.245 281.685 -122.915 ;
        RECT 281.355 -124.605 281.685 -124.275 ;
        RECT 281.355 -125.965 281.685 -125.635 ;
        RECT 281.355 -127.325 281.685 -126.995 ;
        RECT 281.355 -128.685 281.685 -128.355 ;
        RECT 281.355 -130.045 281.685 -129.715 ;
        RECT 281.355 -131.405 281.685 -131.075 ;
        RECT 281.355 -132.765 281.685 -132.435 ;
        RECT 281.355 -134.125 281.685 -133.795 ;
        RECT 281.355 -135.485 281.685 -135.155 ;
        RECT 281.355 -136.845 281.685 -136.515 ;
        RECT 281.355 -138.205 281.685 -137.875 ;
        RECT 281.355 -139.565 281.685 -139.235 ;
        RECT 281.355 -140.925 281.685 -140.595 ;
        RECT 281.355 -142.285 281.685 -141.955 ;
        RECT 281.355 -143.645 281.685 -143.315 ;
        RECT 281.355 -145.005 281.685 -144.675 ;
        RECT 281.355 -146.365 281.685 -146.035 ;
        RECT 281.355 -147.725 281.685 -147.395 ;
        RECT 281.355 -149.085 281.685 -148.755 ;
        RECT 281.355 -150.445 281.685 -150.115 ;
        RECT 281.355 -151.805 281.685 -151.475 ;
        RECT 281.355 -153.165 281.685 -152.835 ;
        RECT 281.355 -154.525 281.685 -154.195 ;
        RECT 281.355 -155.885 281.685 -155.555 ;
        RECT 281.355 -157.245 281.685 -156.915 ;
        RECT 281.355 -158.605 281.685 -158.275 ;
        RECT 281.355 -159.965 281.685 -159.635 ;
        RECT 281.355 -161.325 281.685 -160.995 ;
        RECT 281.355 -162.685 281.685 -162.355 ;
        RECT 281.355 -164.045 281.685 -163.715 ;
        RECT 281.355 -165.405 281.685 -165.075 ;
        RECT 281.355 -166.765 281.685 -166.435 ;
        RECT 281.355 -168.125 281.685 -167.795 ;
        RECT 281.355 -169.485 281.685 -169.155 ;
        RECT 281.355 -170.845 281.685 -170.515 ;
        RECT 281.355 -172.205 281.685 -171.875 ;
        RECT 281.355 -173.565 281.685 -173.235 ;
        RECT 281.355 -174.925 281.685 -174.595 ;
        RECT 281.355 -176.285 281.685 -175.955 ;
        RECT 281.355 -177.645 281.685 -177.315 ;
        RECT 281.355 -179.005 281.685 -178.675 ;
        RECT 281.355 -184.65 281.685 -183.52 ;
        RECT 281.36 -184.765 281.68 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.715 244.04 283.045 245.17 ;
        RECT 282.715 239.875 283.045 240.205 ;
        RECT 282.715 238.515 283.045 238.845 ;
        RECT 282.715 237.155 283.045 237.485 ;
        RECT 282.72 237.155 283.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.715 -0.845 283.045 -0.515 ;
        RECT 282.715 -2.205 283.045 -1.875 ;
        RECT 282.715 -3.565 283.045 -3.235 ;
        RECT 282.72 -3.565 283.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.715 -96.045 283.045 -95.715 ;
        RECT 282.715 -97.405 283.045 -97.075 ;
        RECT 282.715 -98.765 283.045 -98.435 ;
        RECT 282.715 -100.125 283.045 -99.795 ;
        RECT 282.715 -101.485 283.045 -101.155 ;
        RECT 282.715 -102.845 283.045 -102.515 ;
        RECT 282.715 -104.205 283.045 -103.875 ;
        RECT 282.715 -105.565 283.045 -105.235 ;
        RECT 282.715 -106.925 283.045 -106.595 ;
        RECT 282.715 -108.285 283.045 -107.955 ;
        RECT 282.715 -109.645 283.045 -109.315 ;
        RECT 282.715 -111.005 283.045 -110.675 ;
        RECT 282.715 -112.365 283.045 -112.035 ;
        RECT 282.715 -113.725 283.045 -113.395 ;
        RECT 282.715 -115.085 283.045 -114.755 ;
        RECT 282.715 -116.445 283.045 -116.115 ;
        RECT 282.715 -117.805 283.045 -117.475 ;
        RECT 282.715 -119.165 283.045 -118.835 ;
        RECT 282.715 -120.525 283.045 -120.195 ;
        RECT 282.715 -121.885 283.045 -121.555 ;
        RECT 282.715 -123.245 283.045 -122.915 ;
        RECT 282.715 -124.605 283.045 -124.275 ;
        RECT 282.715 -125.965 283.045 -125.635 ;
        RECT 282.715 -127.325 283.045 -126.995 ;
        RECT 282.715 -128.685 283.045 -128.355 ;
        RECT 282.715 -130.045 283.045 -129.715 ;
        RECT 282.715 -131.405 283.045 -131.075 ;
        RECT 282.715 -132.765 283.045 -132.435 ;
        RECT 282.715 -134.125 283.045 -133.795 ;
        RECT 282.715 -135.485 283.045 -135.155 ;
        RECT 282.715 -136.845 283.045 -136.515 ;
        RECT 282.715 -138.205 283.045 -137.875 ;
        RECT 282.715 -139.565 283.045 -139.235 ;
        RECT 282.715 -140.925 283.045 -140.595 ;
        RECT 282.715 -142.285 283.045 -141.955 ;
        RECT 282.715 -143.645 283.045 -143.315 ;
        RECT 282.715 -145.005 283.045 -144.675 ;
        RECT 282.715 -146.365 283.045 -146.035 ;
        RECT 282.715 -147.725 283.045 -147.395 ;
        RECT 282.715 -149.085 283.045 -148.755 ;
        RECT 282.715 -150.445 283.045 -150.115 ;
        RECT 282.715 -151.805 283.045 -151.475 ;
        RECT 282.715 -153.165 283.045 -152.835 ;
        RECT 282.715 -154.525 283.045 -154.195 ;
        RECT 282.715 -155.885 283.045 -155.555 ;
        RECT 282.715 -157.245 283.045 -156.915 ;
        RECT 282.715 -158.605 283.045 -158.275 ;
        RECT 282.715 -159.965 283.045 -159.635 ;
        RECT 282.715 -161.325 283.045 -160.995 ;
        RECT 282.715 -162.685 283.045 -162.355 ;
        RECT 282.715 -164.045 283.045 -163.715 ;
        RECT 282.715 -165.405 283.045 -165.075 ;
        RECT 282.715 -166.765 283.045 -166.435 ;
        RECT 282.715 -168.125 283.045 -167.795 ;
        RECT 282.715 -169.485 283.045 -169.155 ;
        RECT 282.715 -170.845 283.045 -170.515 ;
        RECT 282.715 -172.205 283.045 -171.875 ;
        RECT 282.715 -173.565 283.045 -173.235 ;
        RECT 282.715 -174.925 283.045 -174.595 ;
        RECT 282.715 -176.285 283.045 -175.955 ;
        RECT 282.715 -177.645 283.045 -177.315 ;
        RECT 282.715 -179.005 283.045 -178.675 ;
        RECT 282.715 -184.65 283.045 -183.52 ;
        RECT 282.72 -184.765 283.04 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.075 244.04 284.405 245.17 ;
        RECT 284.075 239.875 284.405 240.205 ;
        RECT 284.075 238.515 284.405 238.845 ;
        RECT 284.075 237.155 284.405 237.485 ;
        RECT 284.08 237.155 284.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.075 -0.845 284.405 -0.515 ;
        RECT 284.075 -2.205 284.405 -1.875 ;
        RECT 284.075 -3.565 284.405 -3.235 ;
        RECT 284.08 -3.565 284.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.075 -179.005 284.405 -178.675 ;
        RECT 284.075 -184.65 284.405 -183.52 ;
        RECT 284.08 -184.765 284.4 -95.04 ;
        RECT 284.075 -96.045 284.405 -95.715 ;
        RECT 284.075 -97.405 284.405 -97.075 ;
        RECT 284.075 -98.765 284.405 -98.435 ;
        RECT 284.075 -100.125 284.405 -99.795 ;
        RECT 284.075 -101.485 284.405 -101.155 ;
        RECT 284.075 -102.845 284.405 -102.515 ;
        RECT 284.075 -104.205 284.405 -103.875 ;
        RECT 284.075 -105.565 284.405 -105.235 ;
        RECT 284.075 -106.925 284.405 -106.595 ;
        RECT 284.075 -108.285 284.405 -107.955 ;
        RECT 284.075 -109.645 284.405 -109.315 ;
        RECT 284.075 -111.005 284.405 -110.675 ;
        RECT 284.075 -112.365 284.405 -112.035 ;
        RECT 284.075 -113.725 284.405 -113.395 ;
        RECT 284.075 -115.085 284.405 -114.755 ;
        RECT 284.075 -116.445 284.405 -116.115 ;
        RECT 284.075 -117.805 284.405 -117.475 ;
        RECT 284.075 -119.165 284.405 -118.835 ;
        RECT 284.075 -120.525 284.405 -120.195 ;
        RECT 284.075 -121.885 284.405 -121.555 ;
        RECT 284.075 -123.245 284.405 -122.915 ;
        RECT 284.075 -124.605 284.405 -124.275 ;
        RECT 284.075 -125.965 284.405 -125.635 ;
        RECT 284.075 -127.325 284.405 -126.995 ;
        RECT 284.075 -128.685 284.405 -128.355 ;
        RECT 284.075 -130.045 284.405 -129.715 ;
        RECT 284.075 -131.405 284.405 -131.075 ;
        RECT 284.075 -132.765 284.405 -132.435 ;
        RECT 284.075 -134.125 284.405 -133.795 ;
        RECT 284.075 -135.485 284.405 -135.155 ;
        RECT 284.075 -136.845 284.405 -136.515 ;
        RECT 284.075 -138.205 284.405 -137.875 ;
        RECT 284.075 -139.565 284.405 -139.235 ;
        RECT 284.075 -140.925 284.405 -140.595 ;
        RECT 284.075 -142.285 284.405 -141.955 ;
        RECT 284.075 -143.645 284.405 -143.315 ;
        RECT 284.075 -145.005 284.405 -144.675 ;
        RECT 284.075 -146.365 284.405 -146.035 ;
        RECT 284.075 -147.725 284.405 -147.395 ;
        RECT 284.075 -149.085 284.405 -148.755 ;
        RECT 284.075 -150.445 284.405 -150.115 ;
        RECT 284.075 -151.805 284.405 -151.475 ;
        RECT 284.075 -153.165 284.405 -152.835 ;
        RECT 284.075 -154.525 284.405 -154.195 ;
        RECT 284.075 -155.885 284.405 -155.555 ;
        RECT 284.075 -157.245 284.405 -156.915 ;
        RECT 284.075 -158.605 284.405 -158.275 ;
        RECT 284.075 -159.965 284.405 -159.635 ;
        RECT 284.075 -161.325 284.405 -160.995 ;
        RECT 284.075 -162.685 284.405 -162.355 ;
        RECT 284.075 -164.045 284.405 -163.715 ;
        RECT 284.075 -165.405 284.405 -165.075 ;
        RECT 284.075 -166.765 284.405 -166.435 ;
        RECT 284.075 -168.125 284.405 -167.795 ;
        RECT 284.075 -169.485 284.405 -169.155 ;
        RECT 284.075 -170.845 284.405 -170.515 ;
        RECT 284.075 -172.205 284.405 -171.875 ;
        RECT 284.075 -173.565 284.405 -173.235 ;
        RECT 284.075 -174.925 284.405 -174.595 ;
        RECT 284.075 -176.285 284.405 -175.955 ;
        RECT 284.075 -177.645 284.405 -177.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.835 244.04 238.165 245.17 ;
        RECT 237.835 239.875 238.165 240.205 ;
        RECT 237.835 238.515 238.165 238.845 ;
        RECT 237.835 237.155 238.165 237.485 ;
        RECT 237.84 237.155 238.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.835 -0.845 238.165 -0.515 ;
        RECT 237.835 -2.205 238.165 -1.875 ;
        RECT 237.835 -3.565 238.165 -3.235 ;
        RECT 237.84 -3.565 238.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.835 -96.045 238.165 -95.715 ;
        RECT 237.835 -97.405 238.165 -97.075 ;
        RECT 237.835 -98.765 238.165 -98.435 ;
        RECT 237.835 -100.125 238.165 -99.795 ;
        RECT 237.835 -101.485 238.165 -101.155 ;
        RECT 237.835 -102.845 238.165 -102.515 ;
        RECT 237.835 -104.205 238.165 -103.875 ;
        RECT 237.835 -105.565 238.165 -105.235 ;
        RECT 237.835 -106.925 238.165 -106.595 ;
        RECT 237.835 -108.285 238.165 -107.955 ;
        RECT 237.835 -109.645 238.165 -109.315 ;
        RECT 237.835 -111.005 238.165 -110.675 ;
        RECT 237.835 -112.365 238.165 -112.035 ;
        RECT 237.835 -113.725 238.165 -113.395 ;
        RECT 237.835 -115.085 238.165 -114.755 ;
        RECT 237.835 -116.445 238.165 -116.115 ;
        RECT 237.835 -117.805 238.165 -117.475 ;
        RECT 237.835 -119.165 238.165 -118.835 ;
        RECT 237.835 -120.525 238.165 -120.195 ;
        RECT 237.835 -121.885 238.165 -121.555 ;
        RECT 237.835 -123.245 238.165 -122.915 ;
        RECT 237.835 -124.605 238.165 -124.275 ;
        RECT 237.835 -125.965 238.165 -125.635 ;
        RECT 237.835 -127.325 238.165 -126.995 ;
        RECT 237.835 -128.685 238.165 -128.355 ;
        RECT 237.835 -130.045 238.165 -129.715 ;
        RECT 237.835 -131.405 238.165 -131.075 ;
        RECT 237.835 -132.765 238.165 -132.435 ;
        RECT 237.835 -134.125 238.165 -133.795 ;
        RECT 237.835 -135.485 238.165 -135.155 ;
        RECT 237.835 -136.845 238.165 -136.515 ;
        RECT 237.835 -138.205 238.165 -137.875 ;
        RECT 237.835 -139.565 238.165 -139.235 ;
        RECT 237.835 -140.925 238.165 -140.595 ;
        RECT 237.835 -142.285 238.165 -141.955 ;
        RECT 237.835 -143.645 238.165 -143.315 ;
        RECT 237.835 -145.005 238.165 -144.675 ;
        RECT 237.835 -146.365 238.165 -146.035 ;
        RECT 237.835 -147.725 238.165 -147.395 ;
        RECT 237.835 -149.085 238.165 -148.755 ;
        RECT 237.835 -150.445 238.165 -150.115 ;
        RECT 237.835 -151.805 238.165 -151.475 ;
        RECT 237.835 -153.165 238.165 -152.835 ;
        RECT 237.835 -154.525 238.165 -154.195 ;
        RECT 237.835 -155.885 238.165 -155.555 ;
        RECT 237.835 -157.245 238.165 -156.915 ;
        RECT 237.835 -158.605 238.165 -158.275 ;
        RECT 237.835 -159.965 238.165 -159.635 ;
        RECT 237.835 -161.325 238.165 -160.995 ;
        RECT 237.835 -162.685 238.165 -162.355 ;
        RECT 237.835 -164.045 238.165 -163.715 ;
        RECT 237.835 -165.405 238.165 -165.075 ;
        RECT 237.835 -166.765 238.165 -166.435 ;
        RECT 237.835 -168.125 238.165 -167.795 ;
        RECT 237.835 -169.485 238.165 -169.155 ;
        RECT 237.835 -170.845 238.165 -170.515 ;
        RECT 237.835 -172.205 238.165 -171.875 ;
        RECT 237.835 -173.565 238.165 -173.235 ;
        RECT 237.835 -174.925 238.165 -174.595 ;
        RECT 237.835 -176.285 238.165 -175.955 ;
        RECT 237.835 -177.645 238.165 -177.315 ;
        RECT 237.835 -179.005 238.165 -178.675 ;
        RECT 237.835 -184.65 238.165 -183.52 ;
        RECT 237.84 -184.765 238.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.195 244.04 239.525 245.17 ;
        RECT 239.195 239.875 239.525 240.205 ;
        RECT 239.195 238.515 239.525 238.845 ;
        RECT 239.195 237.155 239.525 237.485 ;
        RECT 239.2 237.155 239.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.195 -0.845 239.525 -0.515 ;
        RECT 239.195 -2.205 239.525 -1.875 ;
        RECT 239.195 -3.565 239.525 -3.235 ;
        RECT 239.2 -3.565 239.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.195 -96.045 239.525 -95.715 ;
        RECT 239.195 -97.405 239.525 -97.075 ;
        RECT 239.195 -98.765 239.525 -98.435 ;
        RECT 239.195 -100.125 239.525 -99.795 ;
        RECT 239.195 -101.485 239.525 -101.155 ;
        RECT 239.195 -102.845 239.525 -102.515 ;
        RECT 239.195 -104.205 239.525 -103.875 ;
        RECT 239.195 -105.565 239.525 -105.235 ;
        RECT 239.195 -106.925 239.525 -106.595 ;
        RECT 239.195 -108.285 239.525 -107.955 ;
        RECT 239.195 -109.645 239.525 -109.315 ;
        RECT 239.195 -111.005 239.525 -110.675 ;
        RECT 239.195 -112.365 239.525 -112.035 ;
        RECT 239.195 -113.725 239.525 -113.395 ;
        RECT 239.195 -115.085 239.525 -114.755 ;
        RECT 239.195 -116.445 239.525 -116.115 ;
        RECT 239.195 -117.805 239.525 -117.475 ;
        RECT 239.195 -119.165 239.525 -118.835 ;
        RECT 239.195 -120.525 239.525 -120.195 ;
        RECT 239.195 -121.885 239.525 -121.555 ;
        RECT 239.195 -123.245 239.525 -122.915 ;
        RECT 239.195 -124.605 239.525 -124.275 ;
        RECT 239.195 -125.965 239.525 -125.635 ;
        RECT 239.195 -127.325 239.525 -126.995 ;
        RECT 239.195 -128.685 239.525 -128.355 ;
        RECT 239.195 -130.045 239.525 -129.715 ;
        RECT 239.195 -131.405 239.525 -131.075 ;
        RECT 239.195 -132.765 239.525 -132.435 ;
        RECT 239.195 -134.125 239.525 -133.795 ;
        RECT 239.195 -135.485 239.525 -135.155 ;
        RECT 239.195 -136.845 239.525 -136.515 ;
        RECT 239.195 -138.205 239.525 -137.875 ;
        RECT 239.195 -139.565 239.525 -139.235 ;
        RECT 239.195 -140.925 239.525 -140.595 ;
        RECT 239.195 -142.285 239.525 -141.955 ;
        RECT 239.195 -143.645 239.525 -143.315 ;
        RECT 239.195 -145.005 239.525 -144.675 ;
        RECT 239.195 -146.365 239.525 -146.035 ;
        RECT 239.195 -147.725 239.525 -147.395 ;
        RECT 239.195 -149.085 239.525 -148.755 ;
        RECT 239.195 -150.445 239.525 -150.115 ;
        RECT 239.195 -151.805 239.525 -151.475 ;
        RECT 239.195 -153.165 239.525 -152.835 ;
        RECT 239.195 -154.525 239.525 -154.195 ;
        RECT 239.195 -155.885 239.525 -155.555 ;
        RECT 239.195 -157.245 239.525 -156.915 ;
        RECT 239.195 -158.605 239.525 -158.275 ;
        RECT 239.195 -159.965 239.525 -159.635 ;
        RECT 239.195 -161.325 239.525 -160.995 ;
        RECT 239.195 -162.685 239.525 -162.355 ;
        RECT 239.195 -164.045 239.525 -163.715 ;
        RECT 239.195 -165.405 239.525 -165.075 ;
        RECT 239.195 -166.765 239.525 -166.435 ;
        RECT 239.195 -168.125 239.525 -167.795 ;
        RECT 239.195 -169.485 239.525 -169.155 ;
        RECT 239.195 -170.845 239.525 -170.515 ;
        RECT 239.195 -172.205 239.525 -171.875 ;
        RECT 239.195 -173.565 239.525 -173.235 ;
        RECT 239.195 -174.925 239.525 -174.595 ;
        RECT 239.195 -176.285 239.525 -175.955 ;
        RECT 239.195 -177.645 239.525 -177.315 ;
        RECT 239.195 -179.005 239.525 -178.675 ;
        RECT 239.195 -184.65 239.525 -183.52 ;
        RECT 239.2 -184.765 239.52 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.555 244.04 240.885 245.17 ;
        RECT 240.555 239.875 240.885 240.205 ;
        RECT 240.555 238.515 240.885 238.845 ;
        RECT 240.555 237.155 240.885 237.485 ;
        RECT 240.56 237.155 240.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.555 -0.845 240.885 -0.515 ;
        RECT 240.555 -2.205 240.885 -1.875 ;
        RECT 240.555 -3.565 240.885 -3.235 ;
        RECT 240.56 -3.565 240.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 240.555 -96.045 240.885 -95.715 ;
        RECT 240.555 -97.405 240.885 -97.075 ;
        RECT 240.555 -98.765 240.885 -98.435 ;
        RECT 240.555 -100.125 240.885 -99.795 ;
        RECT 240.555 -101.485 240.885 -101.155 ;
        RECT 240.555 -102.845 240.885 -102.515 ;
        RECT 240.555 -104.205 240.885 -103.875 ;
        RECT 240.555 -105.565 240.885 -105.235 ;
        RECT 240.555 -106.925 240.885 -106.595 ;
        RECT 240.555 -108.285 240.885 -107.955 ;
        RECT 240.555 -109.645 240.885 -109.315 ;
        RECT 240.555 -111.005 240.885 -110.675 ;
        RECT 240.555 -112.365 240.885 -112.035 ;
        RECT 240.555 -113.725 240.885 -113.395 ;
        RECT 240.555 -115.085 240.885 -114.755 ;
        RECT 240.555 -116.445 240.885 -116.115 ;
        RECT 240.555 -117.805 240.885 -117.475 ;
        RECT 240.555 -119.165 240.885 -118.835 ;
        RECT 240.555 -120.525 240.885 -120.195 ;
        RECT 240.555 -121.885 240.885 -121.555 ;
        RECT 240.555 -123.245 240.885 -122.915 ;
        RECT 240.555 -124.605 240.885 -124.275 ;
        RECT 240.555 -125.965 240.885 -125.635 ;
        RECT 240.555 -127.325 240.885 -126.995 ;
        RECT 240.555 -128.685 240.885 -128.355 ;
        RECT 240.555 -130.045 240.885 -129.715 ;
        RECT 240.555 -131.405 240.885 -131.075 ;
        RECT 240.555 -132.765 240.885 -132.435 ;
        RECT 240.555 -134.125 240.885 -133.795 ;
        RECT 240.555 -135.485 240.885 -135.155 ;
        RECT 240.555 -136.845 240.885 -136.515 ;
        RECT 240.555 -138.205 240.885 -137.875 ;
        RECT 240.555 -139.565 240.885 -139.235 ;
        RECT 240.555 -140.925 240.885 -140.595 ;
        RECT 240.555 -142.285 240.885 -141.955 ;
        RECT 240.555 -143.645 240.885 -143.315 ;
        RECT 240.555 -145.005 240.885 -144.675 ;
        RECT 240.555 -146.365 240.885 -146.035 ;
        RECT 240.555 -147.725 240.885 -147.395 ;
        RECT 240.555 -149.085 240.885 -148.755 ;
        RECT 240.555 -150.445 240.885 -150.115 ;
        RECT 240.555 -151.805 240.885 -151.475 ;
        RECT 240.555 -153.165 240.885 -152.835 ;
        RECT 240.555 -154.525 240.885 -154.195 ;
        RECT 240.555 -155.885 240.885 -155.555 ;
        RECT 240.555 -157.245 240.885 -156.915 ;
        RECT 240.555 -158.605 240.885 -158.275 ;
        RECT 240.555 -159.965 240.885 -159.635 ;
        RECT 240.555 -161.325 240.885 -160.995 ;
        RECT 240.555 -162.685 240.885 -162.355 ;
        RECT 240.555 -164.045 240.885 -163.715 ;
        RECT 240.555 -165.405 240.885 -165.075 ;
        RECT 240.555 -166.765 240.885 -166.435 ;
        RECT 240.555 -168.125 240.885 -167.795 ;
        RECT 240.555 -169.485 240.885 -169.155 ;
        RECT 240.555 -170.845 240.885 -170.515 ;
        RECT 240.555 -172.205 240.885 -171.875 ;
        RECT 240.555 -173.565 240.885 -173.235 ;
        RECT 240.555 -174.925 240.885 -174.595 ;
        RECT 240.555 -176.285 240.885 -175.955 ;
        RECT 240.555 -177.645 240.885 -177.315 ;
        RECT 240.555 -179.005 240.885 -178.675 ;
        RECT 240.555 -184.65 240.885 -183.52 ;
        RECT 240.56 -184.765 240.88 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.915 244.04 242.245 245.17 ;
        RECT 241.915 239.875 242.245 240.205 ;
        RECT 241.915 238.515 242.245 238.845 ;
        RECT 241.915 237.155 242.245 237.485 ;
        RECT 241.92 237.155 242.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.915 -98.765 242.245 -98.435 ;
        RECT 241.915 -100.125 242.245 -99.795 ;
        RECT 241.915 -101.485 242.245 -101.155 ;
        RECT 241.915 -102.845 242.245 -102.515 ;
        RECT 241.915 -104.205 242.245 -103.875 ;
        RECT 241.915 -105.565 242.245 -105.235 ;
        RECT 241.915 -106.925 242.245 -106.595 ;
        RECT 241.915 -108.285 242.245 -107.955 ;
        RECT 241.915 -109.645 242.245 -109.315 ;
        RECT 241.915 -111.005 242.245 -110.675 ;
        RECT 241.915 -112.365 242.245 -112.035 ;
        RECT 241.915 -113.725 242.245 -113.395 ;
        RECT 241.915 -115.085 242.245 -114.755 ;
        RECT 241.915 -116.445 242.245 -116.115 ;
        RECT 241.915 -117.805 242.245 -117.475 ;
        RECT 241.915 -119.165 242.245 -118.835 ;
        RECT 241.915 -120.525 242.245 -120.195 ;
        RECT 241.915 -121.885 242.245 -121.555 ;
        RECT 241.915 -123.245 242.245 -122.915 ;
        RECT 241.915 -124.605 242.245 -124.275 ;
        RECT 241.915 -125.965 242.245 -125.635 ;
        RECT 241.915 -127.325 242.245 -126.995 ;
        RECT 241.915 -128.685 242.245 -128.355 ;
        RECT 241.915 -130.045 242.245 -129.715 ;
        RECT 241.915 -131.405 242.245 -131.075 ;
        RECT 241.915 -132.765 242.245 -132.435 ;
        RECT 241.915 -134.125 242.245 -133.795 ;
        RECT 241.915 -135.485 242.245 -135.155 ;
        RECT 241.915 -136.845 242.245 -136.515 ;
        RECT 241.915 -138.205 242.245 -137.875 ;
        RECT 241.915 -139.565 242.245 -139.235 ;
        RECT 241.915 -140.925 242.245 -140.595 ;
        RECT 241.915 -142.285 242.245 -141.955 ;
        RECT 241.915 -143.645 242.245 -143.315 ;
        RECT 241.915 -145.005 242.245 -144.675 ;
        RECT 241.915 -146.365 242.245 -146.035 ;
        RECT 241.915 -147.725 242.245 -147.395 ;
        RECT 241.915 -149.085 242.245 -148.755 ;
        RECT 241.915 -150.445 242.245 -150.115 ;
        RECT 241.915 -151.805 242.245 -151.475 ;
        RECT 241.915 -153.165 242.245 -152.835 ;
        RECT 241.915 -154.525 242.245 -154.195 ;
        RECT 241.915 -155.885 242.245 -155.555 ;
        RECT 241.915 -157.245 242.245 -156.915 ;
        RECT 241.915 -158.605 242.245 -158.275 ;
        RECT 241.915 -159.965 242.245 -159.635 ;
        RECT 241.915 -161.325 242.245 -160.995 ;
        RECT 241.915 -162.685 242.245 -162.355 ;
        RECT 241.915 -164.045 242.245 -163.715 ;
        RECT 241.915 -165.405 242.245 -165.075 ;
        RECT 241.915 -166.765 242.245 -166.435 ;
        RECT 241.915 -168.125 242.245 -167.795 ;
        RECT 241.915 -169.485 242.245 -169.155 ;
        RECT 241.915 -170.845 242.245 -170.515 ;
        RECT 241.915 -172.205 242.245 -171.875 ;
        RECT 241.915 -173.565 242.245 -173.235 ;
        RECT 241.915 -174.925 242.245 -174.595 ;
        RECT 241.915 -176.285 242.245 -175.955 ;
        RECT 241.915 -177.645 242.245 -177.315 ;
        RECT 241.915 -179.005 242.245 -178.675 ;
        RECT 241.915 -184.65 242.245 -183.52 ;
        RECT 241.92 -184.765 242.24 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.46 -98.075 242.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.275 244.04 243.605 245.17 ;
        RECT 243.275 239.875 243.605 240.205 ;
        RECT 243.275 238.515 243.605 238.845 ;
        RECT 243.275 237.155 243.605 237.485 ;
        RECT 243.28 237.155 243.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.635 244.04 244.965 245.17 ;
        RECT 244.635 239.875 244.965 240.205 ;
        RECT 244.635 238.515 244.965 238.845 ;
        RECT 244.635 237.155 244.965 237.485 ;
        RECT 244.64 237.155 244.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.635 -0.845 244.965 -0.515 ;
        RECT 244.635 -2.205 244.965 -1.875 ;
        RECT 244.635 -3.565 244.965 -3.235 ;
        RECT 244.64 -3.565 244.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 244.635 -96.045 244.965 -95.715 ;
        RECT 244.635 -97.405 244.965 -97.075 ;
        RECT 244.635 -98.765 244.965 -98.435 ;
        RECT 244.635 -100.125 244.965 -99.795 ;
        RECT 244.635 -101.485 244.965 -101.155 ;
        RECT 244.635 -102.845 244.965 -102.515 ;
        RECT 244.635 -104.205 244.965 -103.875 ;
        RECT 244.635 -105.565 244.965 -105.235 ;
        RECT 244.635 -106.925 244.965 -106.595 ;
        RECT 244.635 -108.285 244.965 -107.955 ;
        RECT 244.635 -109.645 244.965 -109.315 ;
        RECT 244.635 -111.005 244.965 -110.675 ;
        RECT 244.635 -112.365 244.965 -112.035 ;
        RECT 244.635 -113.725 244.965 -113.395 ;
        RECT 244.635 -115.085 244.965 -114.755 ;
        RECT 244.635 -116.445 244.965 -116.115 ;
        RECT 244.635 -117.805 244.965 -117.475 ;
        RECT 244.635 -119.165 244.965 -118.835 ;
        RECT 244.635 -120.525 244.965 -120.195 ;
        RECT 244.635 -121.885 244.965 -121.555 ;
        RECT 244.635 -123.245 244.965 -122.915 ;
        RECT 244.635 -124.605 244.965 -124.275 ;
        RECT 244.635 -125.965 244.965 -125.635 ;
        RECT 244.635 -127.325 244.965 -126.995 ;
        RECT 244.635 -128.685 244.965 -128.355 ;
        RECT 244.635 -130.045 244.965 -129.715 ;
        RECT 244.635 -131.405 244.965 -131.075 ;
        RECT 244.635 -132.765 244.965 -132.435 ;
        RECT 244.635 -134.125 244.965 -133.795 ;
        RECT 244.635 -135.485 244.965 -135.155 ;
        RECT 244.635 -136.845 244.965 -136.515 ;
        RECT 244.635 -138.205 244.965 -137.875 ;
        RECT 244.635 -139.565 244.965 -139.235 ;
        RECT 244.635 -140.925 244.965 -140.595 ;
        RECT 244.635 -142.285 244.965 -141.955 ;
        RECT 244.635 -143.645 244.965 -143.315 ;
        RECT 244.635 -145.005 244.965 -144.675 ;
        RECT 244.635 -146.365 244.965 -146.035 ;
        RECT 244.635 -147.725 244.965 -147.395 ;
        RECT 244.635 -149.085 244.965 -148.755 ;
        RECT 244.635 -150.445 244.965 -150.115 ;
        RECT 244.635 -151.805 244.965 -151.475 ;
        RECT 244.635 -153.165 244.965 -152.835 ;
        RECT 244.635 -154.525 244.965 -154.195 ;
        RECT 244.635 -155.885 244.965 -155.555 ;
        RECT 244.635 -157.245 244.965 -156.915 ;
        RECT 244.635 -158.605 244.965 -158.275 ;
        RECT 244.635 -159.965 244.965 -159.635 ;
        RECT 244.635 -161.325 244.965 -160.995 ;
        RECT 244.635 -162.685 244.965 -162.355 ;
        RECT 244.635 -164.045 244.965 -163.715 ;
        RECT 244.635 -165.405 244.965 -165.075 ;
        RECT 244.635 -166.765 244.965 -166.435 ;
        RECT 244.635 -168.125 244.965 -167.795 ;
        RECT 244.635 -169.485 244.965 -169.155 ;
        RECT 244.635 -170.845 244.965 -170.515 ;
        RECT 244.635 -172.205 244.965 -171.875 ;
        RECT 244.635 -173.565 244.965 -173.235 ;
        RECT 244.635 -174.925 244.965 -174.595 ;
        RECT 244.635 -176.285 244.965 -175.955 ;
        RECT 244.635 -177.645 244.965 -177.315 ;
        RECT 244.635 -179.005 244.965 -178.675 ;
        RECT 244.635 -184.65 244.965 -183.52 ;
        RECT 244.64 -184.765 244.96 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.995 244.04 246.325 245.17 ;
        RECT 245.995 239.875 246.325 240.205 ;
        RECT 245.995 238.515 246.325 238.845 ;
        RECT 245.995 237.155 246.325 237.485 ;
        RECT 246 237.155 246.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.995 -0.845 246.325 -0.515 ;
        RECT 245.995 -2.205 246.325 -1.875 ;
        RECT 245.995 -3.565 246.325 -3.235 ;
        RECT 246 -3.565 246.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.355 244.04 247.685 245.17 ;
        RECT 247.355 239.875 247.685 240.205 ;
        RECT 247.355 238.515 247.685 238.845 ;
        RECT 247.355 237.155 247.685 237.485 ;
        RECT 247.36 237.155 247.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.355 -0.845 247.685 -0.515 ;
        RECT 247.355 -2.205 247.685 -1.875 ;
        RECT 247.355 -3.565 247.685 -3.235 ;
        RECT 247.36 -3.565 247.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 247.355 -96.045 247.685 -95.715 ;
        RECT 247.355 -97.405 247.685 -97.075 ;
        RECT 247.355 -98.765 247.685 -98.435 ;
        RECT 247.355 -100.125 247.685 -99.795 ;
        RECT 247.355 -101.485 247.685 -101.155 ;
        RECT 247.355 -102.845 247.685 -102.515 ;
        RECT 247.355 -104.205 247.685 -103.875 ;
        RECT 247.355 -105.565 247.685 -105.235 ;
        RECT 247.355 -106.925 247.685 -106.595 ;
        RECT 247.355 -108.285 247.685 -107.955 ;
        RECT 247.355 -109.645 247.685 -109.315 ;
        RECT 247.355 -111.005 247.685 -110.675 ;
        RECT 247.355 -112.365 247.685 -112.035 ;
        RECT 247.355 -113.725 247.685 -113.395 ;
        RECT 247.355 -115.085 247.685 -114.755 ;
        RECT 247.355 -116.445 247.685 -116.115 ;
        RECT 247.355 -117.805 247.685 -117.475 ;
        RECT 247.355 -119.165 247.685 -118.835 ;
        RECT 247.355 -120.525 247.685 -120.195 ;
        RECT 247.355 -121.885 247.685 -121.555 ;
        RECT 247.355 -123.245 247.685 -122.915 ;
        RECT 247.355 -124.605 247.685 -124.275 ;
        RECT 247.355 -125.965 247.685 -125.635 ;
        RECT 247.355 -127.325 247.685 -126.995 ;
        RECT 247.355 -128.685 247.685 -128.355 ;
        RECT 247.355 -130.045 247.685 -129.715 ;
        RECT 247.355 -131.405 247.685 -131.075 ;
        RECT 247.355 -132.765 247.685 -132.435 ;
        RECT 247.355 -134.125 247.685 -133.795 ;
        RECT 247.355 -135.485 247.685 -135.155 ;
        RECT 247.355 -136.845 247.685 -136.515 ;
        RECT 247.355 -138.205 247.685 -137.875 ;
        RECT 247.355 -139.565 247.685 -139.235 ;
        RECT 247.355 -140.925 247.685 -140.595 ;
        RECT 247.355 -142.285 247.685 -141.955 ;
        RECT 247.355 -143.645 247.685 -143.315 ;
        RECT 247.355 -145.005 247.685 -144.675 ;
        RECT 247.355 -146.365 247.685 -146.035 ;
        RECT 247.355 -147.725 247.685 -147.395 ;
        RECT 247.355 -149.085 247.685 -148.755 ;
        RECT 247.355 -150.445 247.685 -150.115 ;
        RECT 247.355 -151.805 247.685 -151.475 ;
        RECT 247.355 -153.165 247.685 -152.835 ;
        RECT 247.355 -154.525 247.685 -154.195 ;
        RECT 247.355 -155.885 247.685 -155.555 ;
        RECT 247.355 -157.245 247.685 -156.915 ;
        RECT 247.355 -158.605 247.685 -158.275 ;
        RECT 247.355 -159.965 247.685 -159.635 ;
        RECT 247.355 -161.325 247.685 -160.995 ;
        RECT 247.355 -162.685 247.685 -162.355 ;
        RECT 247.355 -164.045 247.685 -163.715 ;
        RECT 247.355 -165.405 247.685 -165.075 ;
        RECT 247.355 -166.765 247.685 -166.435 ;
        RECT 247.355 -168.125 247.685 -167.795 ;
        RECT 247.355 -169.485 247.685 -169.155 ;
        RECT 247.355 -170.845 247.685 -170.515 ;
        RECT 247.355 -172.205 247.685 -171.875 ;
        RECT 247.355 -173.565 247.685 -173.235 ;
        RECT 247.355 -174.925 247.685 -174.595 ;
        RECT 247.355 -176.285 247.685 -175.955 ;
        RECT 247.355 -177.645 247.685 -177.315 ;
        RECT 247.355 -179.005 247.685 -178.675 ;
        RECT 247.355 -184.65 247.685 -183.52 ;
        RECT 247.36 -184.765 247.68 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.715 244.04 249.045 245.17 ;
        RECT 248.715 239.875 249.045 240.205 ;
        RECT 248.715 238.515 249.045 238.845 ;
        RECT 248.715 237.155 249.045 237.485 ;
        RECT 248.72 237.155 249.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.715 -0.845 249.045 -0.515 ;
        RECT 248.715 -2.205 249.045 -1.875 ;
        RECT 248.715 -3.565 249.045 -3.235 ;
        RECT 248.72 -3.565 249.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.715 -96.045 249.045 -95.715 ;
        RECT 248.715 -97.405 249.045 -97.075 ;
        RECT 248.715 -98.765 249.045 -98.435 ;
        RECT 248.715 -100.125 249.045 -99.795 ;
        RECT 248.715 -101.485 249.045 -101.155 ;
        RECT 248.715 -102.845 249.045 -102.515 ;
        RECT 248.715 -104.205 249.045 -103.875 ;
        RECT 248.715 -105.565 249.045 -105.235 ;
        RECT 248.715 -106.925 249.045 -106.595 ;
        RECT 248.715 -108.285 249.045 -107.955 ;
        RECT 248.715 -109.645 249.045 -109.315 ;
        RECT 248.715 -111.005 249.045 -110.675 ;
        RECT 248.715 -112.365 249.045 -112.035 ;
        RECT 248.715 -113.725 249.045 -113.395 ;
        RECT 248.715 -115.085 249.045 -114.755 ;
        RECT 248.715 -116.445 249.045 -116.115 ;
        RECT 248.715 -117.805 249.045 -117.475 ;
        RECT 248.715 -119.165 249.045 -118.835 ;
        RECT 248.715 -120.525 249.045 -120.195 ;
        RECT 248.715 -121.885 249.045 -121.555 ;
        RECT 248.715 -123.245 249.045 -122.915 ;
        RECT 248.715 -124.605 249.045 -124.275 ;
        RECT 248.715 -125.965 249.045 -125.635 ;
        RECT 248.715 -127.325 249.045 -126.995 ;
        RECT 248.715 -128.685 249.045 -128.355 ;
        RECT 248.715 -130.045 249.045 -129.715 ;
        RECT 248.715 -131.405 249.045 -131.075 ;
        RECT 248.715 -132.765 249.045 -132.435 ;
        RECT 248.715 -134.125 249.045 -133.795 ;
        RECT 248.715 -135.485 249.045 -135.155 ;
        RECT 248.715 -136.845 249.045 -136.515 ;
        RECT 248.715 -138.205 249.045 -137.875 ;
        RECT 248.715 -139.565 249.045 -139.235 ;
        RECT 248.715 -140.925 249.045 -140.595 ;
        RECT 248.715 -142.285 249.045 -141.955 ;
        RECT 248.715 -143.645 249.045 -143.315 ;
        RECT 248.715 -145.005 249.045 -144.675 ;
        RECT 248.715 -146.365 249.045 -146.035 ;
        RECT 248.715 -147.725 249.045 -147.395 ;
        RECT 248.715 -149.085 249.045 -148.755 ;
        RECT 248.715 -150.445 249.045 -150.115 ;
        RECT 248.715 -151.805 249.045 -151.475 ;
        RECT 248.715 -153.165 249.045 -152.835 ;
        RECT 248.715 -154.525 249.045 -154.195 ;
        RECT 248.715 -155.885 249.045 -155.555 ;
        RECT 248.715 -157.245 249.045 -156.915 ;
        RECT 248.715 -158.605 249.045 -158.275 ;
        RECT 248.715 -159.965 249.045 -159.635 ;
        RECT 248.715 -161.325 249.045 -160.995 ;
        RECT 248.715 -162.685 249.045 -162.355 ;
        RECT 248.715 -164.045 249.045 -163.715 ;
        RECT 248.715 -165.405 249.045 -165.075 ;
        RECT 248.715 -166.765 249.045 -166.435 ;
        RECT 248.715 -168.125 249.045 -167.795 ;
        RECT 248.715 -169.485 249.045 -169.155 ;
        RECT 248.715 -170.845 249.045 -170.515 ;
        RECT 248.715 -172.205 249.045 -171.875 ;
        RECT 248.715 -173.565 249.045 -173.235 ;
        RECT 248.715 -174.925 249.045 -174.595 ;
        RECT 248.715 -176.285 249.045 -175.955 ;
        RECT 248.715 -177.645 249.045 -177.315 ;
        RECT 248.715 -179.005 249.045 -178.675 ;
        RECT 248.715 -184.65 249.045 -183.52 ;
        RECT 248.72 -184.765 249.04 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.075 244.04 250.405 245.17 ;
        RECT 250.075 239.875 250.405 240.205 ;
        RECT 250.075 238.515 250.405 238.845 ;
        RECT 250.075 237.155 250.405 237.485 ;
        RECT 250.08 237.155 250.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.075 -0.845 250.405 -0.515 ;
        RECT 250.075 -2.205 250.405 -1.875 ;
        RECT 250.075 -3.565 250.405 -3.235 ;
        RECT 250.08 -3.565 250.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.075 -96.045 250.405 -95.715 ;
        RECT 250.075 -97.405 250.405 -97.075 ;
        RECT 250.075 -98.765 250.405 -98.435 ;
        RECT 250.075 -100.125 250.405 -99.795 ;
        RECT 250.075 -101.485 250.405 -101.155 ;
        RECT 250.075 -102.845 250.405 -102.515 ;
        RECT 250.075 -104.205 250.405 -103.875 ;
        RECT 250.075 -105.565 250.405 -105.235 ;
        RECT 250.075 -106.925 250.405 -106.595 ;
        RECT 250.075 -108.285 250.405 -107.955 ;
        RECT 250.075 -109.645 250.405 -109.315 ;
        RECT 250.075 -111.005 250.405 -110.675 ;
        RECT 250.075 -112.365 250.405 -112.035 ;
        RECT 250.075 -113.725 250.405 -113.395 ;
        RECT 250.075 -115.085 250.405 -114.755 ;
        RECT 250.075 -116.445 250.405 -116.115 ;
        RECT 250.075 -117.805 250.405 -117.475 ;
        RECT 250.075 -119.165 250.405 -118.835 ;
        RECT 250.075 -120.525 250.405 -120.195 ;
        RECT 250.075 -121.885 250.405 -121.555 ;
        RECT 250.075 -123.245 250.405 -122.915 ;
        RECT 250.075 -124.605 250.405 -124.275 ;
        RECT 250.075 -125.965 250.405 -125.635 ;
        RECT 250.075 -127.325 250.405 -126.995 ;
        RECT 250.075 -128.685 250.405 -128.355 ;
        RECT 250.075 -130.045 250.405 -129.715 ;
        RECT 250.075 -131.405 250.405 -131.075 ;
        RECT 250.075 -132.765 250.405 -132.435 ;
        RECT 250.075 -134.125 250.405 -133.795 ;
        RECT 250.075 -135.485 250.405 -135.155 ;
        RECT 250.075 -136.845 250.405 -136.515 ;
        RECT 250.075 -138.205 250.405 -137.875 ;
        RECT 250.075 -139.565 250.405 -139.235 ;
        RECT 250.075 -140.925 250.405 -140.595 ;
        RECT 250.075 -142.285 250.405 -141.955 ;
        RECT 250.075 -143.645 250.405 -143.315 ;
        RECT 250.075 -145.005 250.405 -144.675 ;
        RECT 250.075 -146.365 250.405 -146.035 ;
        RECT 250.075 -147.725 250.405 -147.395 ;
        RECT 250.075 -149.085 250.405 -148.755 ;
        RECT 250.075 -150.445 250.405 -150.115 ;
        RECT 250.075 -151.805 250.405 -151.475 ;
        RECT 250.075 -153.165 250.405 -152.835 ;
        RECT 250.075 -154.525 250.405 -154.195 ;
        RECT 250.075 -155.885 250.405 -155.555 ;
        RECT 250.075 -157.245 250.405 -156.915 ;
        RECT 250.075 -158.605 250.405 -158.275 ;
        RECT 250.075 -159.965 250.405 -159.635 ;
        RECT 250.075 -161.325 250.405 -160.995 ;
        RECT 250.075 -162.685 250.405 -162.355 ;
        RECT 250.075 -164.045 250.405 -163.715 ;
        RECT 250.075 -165.405 250.405 -165.075 ;
        RECT 250.075 -166.765 250.405 -166.435 ;
        RECT 250.075 -168.125 250.405 -167.795 ;
        RECT 250.075 -169.485 250.405 -169.155 ;
        RECT 250.075 -170.845 250.405 -170.515 ;
        RECT 250.075 -172.205 250.405 -171.875 ;
        RECT 250.075 -173.565 250.405 -173.235 ;
        RECT 250.075 -174.925 250.405 -174.595 ;
        RECT 250.075 -176.285 250.405 -175.955 ;
        RECT 250.075 -177.645 250.405 -177.315 ;
        RECT 250.075 -179.005 250.405 -178.675 ;
        RECT 250.075 -184.65 250.405 -183.52 ;
        RECT 250.08 -184.765 250.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.435 244.04 251.765 245.17 ;
        RECT 251.435 239.875 251.765 240.205 ;
        RECT 251.435 238.515 251.765 238.845 ;
        RECT 251.435 237.155 251.765 237.485 ;
        RECT 251.44 237.155 251.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.435 -0.845 251.765 -0.515 ;
        RECT 251.435 -2.205 251.765 -1.875 ;
        RECT 251.435 -3.565 251.765 -3.235 ;
        RECT 251.44 -3.565 251.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 251.435 -96.045 251.765 -95.715 ;
        RECT 251.435 -97.405 251.765 -97.075 ;
        RECT 251.435 -98.765 251.765 -98.435 ;
        RECT 251.435 -100.125 251.765 -99.795 ;
        RECT 251.435 -101.485 251.765 -101.155 ;
        RECT 251.435 -102.845 251.765 -102.515 ;
        RECT 251.435 -104.205 251.765 -103.875 ;
        RECT 251.435 -105.565 251.765 -105.235 ;
        RECT 251.435 -106.925 251.765 -106.595 ;
        RECT 251.435 -108.285 251.765 -107.955 ;
        RECT 251.435 -109.645 251.765 -109.315 ;
        RECT 251.435 -111.005 251.765 -110.675 ;
        RECT 251.435 -112.365 251.765 -112.035 ;
        RECT 251.435 -113.725 251.765 -113.395 ;
        RECT 251.435 -115.085 251.765 -114.755 ;
        RECT 251.435 -116.445 251.765 -116.115 ;
        RECT 251.435 -117.805 251.765 -117.475 ;
        RECT 251.435 -119.165 251.765 -118.835 ;
        RECT 251.435 -120.525 251.765 -120.195 ;
        RECT 251.435 -121.885 251.765 -121.555 ;
        RECT 251.435 -123.245 251.765 -122.915 ;
        RECT 251.435 -124.605 251.765 -124.275 ;
        RECT 251.435 -125.965 251.765 -125.635 ;
        RECT 251.435 -127.325 251.765 -126.995 ;
        RECT 251.435 -128.685 251.765 -128.355 ;
        RECT 251.435 -130.045 251.765 -129.715 ;
        RECT 251.435 -131.405 251.765 -131.075 ;
        RECT 251.435 -132.765 251.765 -132.435 ;
        RECT 251.435 -134.125 251.765 -133.795 ;
        RECT 251.435 -135.485 251.765 -135.155 ;
        RECT 251.435 -136.845 251.765 -136.515 ;
        RECT 251.435 -138.205 251.765 -137.875 ;
        RECT 251.435 -139.565 251.765 -139.235 ;
        RECT 251.435 -140.925 251.765 -140.595 ;
        RECT 251.435 -142.285 251.765 -141.955 ;
        RECT 251.435 -143.645 251.765 -143.315 ;
        RECT 251.435 -145.005 251.765 -144.675 ;
        RECT 251.435 -146.365 251.765 -146.035 ;
        RECT 251.435 -147.725 251.765 -147.395 ;
        RECT 251.435 -149.085 251.765 -148.755 ;
        RECT 251.435 -150.445 251.765 -150.115 ;
        RECT 251.435 -151.805 251.765 -151.475 ;
        RECT 251.435 -153.165 251.765 -152.835 ;
        RECT 251.435 -154.525 251.765 -154.195 ;
        RECT 251.435 -155.885 251.765 -155.555 ;
        RECT 251.435 -157.245 251.765 -156.915 ;
        RECT 251.435 -158.605 251.765 -158.275 ;
        RECT 251.435 -159.965 251.765 -159.635 ;
        RECT 251.435 -161.325 251.765 -160.995 ;
        RECT 251.435 -162.685 251.765 -162.355 ;
        RECT 251.435 -164.045 251.765 -163.715 ;
        RECT 251.435 -165.405 251.765 -165.075 ;
        RECT 251.435 -166.765 251.765 -166.435 ;
        RECT 251.435 -168.125 251.765 -167.795 ;
        RECT 251.435 -169.485 251.765 -169.155 ;
        RECT 251.435 -170.845 251.765 -170.515 ;
        RECT 251.435 -172.205 251.765 -171.875 ;
        RECT 251.435 -173.565 251.765 -173.235 ;
        RECT 251.435 -174.925 251.765 -174.595 ;
        RECT 251.435 -176.285 251.765 -175.955 ;
        RECT 251.435 -177.645 251.765 -177.315 ;
        RECT 251.435 -179.005 251.765 -178.675 ;
        RECT 251.435 -184.65 251.765 -183.52 ;
        RECT 251.44 -184.765 251.76 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.795 244.04 253.125 245.17 ;
        RECT 252.795 239.875 253.125 240.205 ;
        RECT 252.795 238.515 253.125 238.845 ;
        RECT 252.795 237.155 253.125 237.485 ;
        RECT 252.8 237.155 253.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.795 -98.765 253.125 -98.435 ;
        RECT 252.795 -100.125 253.125 -99.795 ;
        RECT 252.795 -101.485 253.125 -101.155 ;
        RECT 252.795 -102.845 253.125 -102.515 ;
        RECT 252.795 -104.205 253.125 -103.875 ;
        RECT 252.795 -105.565 253.125 -105.235 ;
        RECT 252.795 -106.925 253.125 -106.595 ;
        RECT 252.795 -108.285 253.125 -107.955 ;
        RECT 252.795 -109.645 253.125 -109.315 ;
        RECT 252.795 -111.005 253.125 -110.675 ;
        RECT 252.795 -112.365 253.125 -112.035 ;
        RECT 252.795 -113.725 253.125 -113.395 ;
        RECT 252.795 -115.085 253.125 -114.755 ;
        RECT 252.795 -116.445 253.125 -116.115 ;
        RECT 252.795 -117.805 253.125 -117.475 ;
        RECT 252.795 -119.165 253.125 -118.835 ;
        RECT 252.795 -120.525 253.125 -120.195 ;
        RECT 252.795 -121.885 253.125 -121.555 ;
        RECT 252.795 -123.245 253.125 -122.915 ;
        RECT 252.795 -124.605 253.125 -124.275 ;
        RECT 252.795 -125.965 253.125 -125.635 ;
        RECT 252.795 -127.325 253.125 -126.995 ;
        RECT 252.795 -128.685 253.125 -128.355 ;
        RECT 252.795 -130.045 253.125 -129.715 ;
        RECT 252.795 -131.405 253.125 -131.075 ;
        RECT 252.795 -132.765 253.125 -132.435 ;
        RECT 252.795 -134.125 253.125 -133.795 ;
        RECT 252.795 -135.485 253.125 -135.155 ;
        RECT 252.795 -136.845 253.125 -136.515 ;
        RECT 252.795 -138.205 253.125 -137.875 ;
        RECT 252.795 -139.565 253.125 -139.235 ;
        RECT 252.795 -140.925 253.125 -140.595 ;
        RECT 252.795 -142.285 253.125 -141.955 ;
        RECT 252.795 -143.645 253.125 -143.315 ;
        RECT 252.795 -145.005 253.125 -144.675 ;
        RECT 252.795 -146.365 253.125 -146.035 ;
        RECT 252.795 -147.725 253.125 -147.395 ;
        RECT 252.795 -149.085 253.125 -148.755 ;
        RECT 252.795 -150.445 253.125 -150.115 ;
        RECT 252.795 -151.805 253.125 -151.475 ;
        RECT 252.795 -153.165 253.125 -152.835 ;
        RECT 252.795 -154.525 253.125 -154.195 ;
        RECT 252.795 -155.885 253.125 -155.555 ;
        RECT 252.795 -157.245 253.125 -156.915 ;
        RECT 252.795 -158.605 253.125 -158.275 ;
        RECT 252.795 -159.965 253.125 -159.635 ;
        RECT 252.795 -161.325 253.125 -160.995 ;
        RECT 252.795 -162.685 253.125 -162.355 ;
        RECT 252.795 -164.045 253.125 -163.715 ;
        RECT 252.795 -165.405 253.125 -165.075 ;
        RECT 252.795 -166.765 253.125 -166.435 ;
        RECT 252.795 -168.125 253.125 -167.795 ;
        RECT 252.795 -169.485 253.125 -169.155 ;
        RECT 252.795 -170.845 253.125 -170.515 ;
        RECT 252.795 -172.205 253.125 -171.875 ;
        RECT 252.795 -173.565 253.125 -173.235 ;
        RECT 252.795 -174.925 253.125 -174.595 ;
        RECT 252.795 -176.285 253.125 -175.955 ;
        RECT 252.795 -177.645 253.125 -177.315 ;
        RECT 252.795 -179.005 253.125 -178.675 ;
        RECT 252.795 -184.65 253.125 -183.52 ;
        RECT 252.8 -184.765 253.12 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.36 -98.075 253.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.155 244.04 254.485 245.17 ;
        RECT 254.155 239.875 254.485 240.205 ;
        RECT 254.155 238.515 254.485 238.845 ;
        RECT 254.155 237.155 254.485 237.485 ;
        RECT 254.16 237.155 254.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.515 244.04 255.845 245.17 ;
        RECT 255.515 239.875 255.845 240.205 ;
        RECT 255.515 238.515 255.845 238.845 ;
        RECT 255.515 237.155 255.845 237.485 ;
        RECT 255.52 237.155 255.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.515 -0.845 255.845 -0.515 ;
        RECT 255.515 -2.205 255.845 -1.875 ;
        RECT 255.515 -3.565 255.845 -3.235 ;
        RECT 255.52 -3.565 255.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 255.515 -96.045 255.845 -95.715 ;
        RECT 255.515 -97.405 255.845 -97.075 ;
        RECT 255.515 -98.765 255.845 -98.435 ;
        RECT 255.515 -100.125 255.845 -99.795 ;
        RECT 255.515 -101.485 255.845 -101.155 ;
        RECT 255.515 -102.845 255.845 -102.515 ;
        RECT 255.515 -104.205 255.845 -103.875 ;
        RECT 255.515 -105.565 255.845 -105.235 ;
        RECT 255.515 -106.925 255.845 -106.595 ;
        RECT 255.515 -108.285 255.845 -107.955 ;
        RECT 255.515 -109.645 255.845 -109.315 ;
        RECT 255.515 -111.005 255.845 -110.675 ;
        RECT 255.515 -112.365 255.845 -112.035 ;
        RECT 255.515 -113.725 255.845 -113.395 ;
        RECT 255.515 -115.085 255.845 -114.755 ;
        RECT 255.515 -116.445 255.845 -116.115 ;
        RECT 255.515 -117.805 255.845 -117.475 ;
        RECT 255.515 -119.165 255.845 -118.835 ;
        RECT 255.515 -120.525 255.845 -120.195 ;
        RECT 255.515 -121.885 255.845 -121.555 ;
        RECT 255.515 -123.245 255.845 -122.915 ;
        RECT 255.515 -124.605 255.845 -124.275 ;
        RECT 255.515 -125.965 255.845 -125.635 ;
        RECT 255.515 -127.325 255.845 -126.995 ;
        RECT 255.515 -128.685 255.845 -128.355 ;
        RECT 255.515 -130.045 255.845 -129.715 ;
        RECT 255.515 -131.405 255.845 -131.075 ;
        RECT 255.515 -132.765 255.845 -132.435 ;
        RECT 255.515 -134.125 255.845 -133.795 ;
        RECT 255.515 -135.485 255.845 -135.155 ;
        RECT 255.515 -136.845 255.845 -136.515 ;
        RECT 255.515 -138.205 255.845 -137.875 ;
        RECT 255.515 -139.565 255.845 -139.235 ;
        RECT 255.515 -140.925 255.845 -140.595 ;
        RECT 255.515 -142.285 255.845 -141.955 ;
        RECT 255.515 -143.645 255.845 -143.315 ;
        RECT 255.515 -145.005 255.845 -144.675 ;
        RECT 255.515 -146.365 255.845 -146.035 ;
        RECT 255.515 -147.725 255.845 -147.395 ;
        RECT 255.515 -149.085 255.845 -148.755 ;
        RECT 255.515 -150.445 255.845 -150.115 ;
        RECT 255.515 -151.805 255.845 -151.475 ;
        RECT 255.515 -153.165 255.845 -152.835 ;
        RECT 255.515 -154.525 255.845 -154.195 ;
        RECT 255.515 -155.885 255.845 -155.555 ;
        RECT 255.515 -157.245 255.845 -156.915 ;
        RECT 255.515 -158.605 255.845 -158.275 ;
        RECT 255.515 -159.965 255.845 -159.635 ;
        RECT 255.515 -161.325 255.845 -160.995 ;
        RECT 255.515 -162.685 255.845 -162.355 ;
        RECT 255.515 -164.045 255.845 -163.715 ;
        RECT 255.515 -165.405 255.845 -165.075 ;
        RECT 255.515 -166.765 255.845 -166.435 ;
        RECT 255.515 -168.125 255.845 -167.795 ;
        RECT 255.515 -169.485 255.845 -169.155 ;
        RECT 255.515 -170.845 255.845 -170.515 ;
        RECT 255.515 -172.205 255.845 -171.875 ;
        RECT 255.515 -173.565 255.845 -173.235 ;
        RECT 255.515 -174.925 255.845 -174.595 ;
        RECT 255.515 -176.285 255.845 -175.955 ;
        RECT 255.515 -177.645 255.845 -177.315 ;
        RECT 255.515 -179.005 255.845 -178.675 ;
        RECT 255.515 -184.65 255.845 -183.52 ;
        RECT 255.52 -184.765 255.84 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.875 244.04 257.205 245.17 ;
        RECT 256.875 239.875 257.205 240.205 ;
        RECT 256.875 238.515 257.205 238.845 ;
        RECT 256.875 237.155 257.205 237.485 ;
        RECT 256.88 237.155 257.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.875 -0.845 257.205 -0.515 ;
        RECT 256.875 -2.205 257.205 -1.875 ;
        RECT 256.875 -3.565 257.205 -3.235 ;
        RECT 256.88 -3.565 257.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.235 244.04 258.565 245.17 ;
        RECT 258.235 239.875 258.565 240.205 ;
        RECT 258.235 238.515 258.565 238.845 ;
        RECT 258.235 237.155 258.565 237.485 ;
        RECT 258.24 237.155 258.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.235 -0.845 258.565 -0.515 ;
        RECT 258.235 -2.205 258.565 -1.875 ;
        RECT 258.235 -3.565 258.565 -3.235 ;
        RECT 258.24 -3.565 258.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.235 -96.045 258.565 -95.715 ;
        RECT 258.235 -97.405 258.565 -97.075 ;
        RECT 258.235 -98.765 258.565 -98.435 ;
        RECT 258.235 -100.125 258.565 -99.795 ;
        RECT 258.235 -101.485 258.565 -101.155 ;
        RECT 258.235 -102.845 258.565 -102.515 ;
        RECT 258.235 -104.205 258.565 -103.875 ;
        RECT 258.235 -105.565 258.565 -105.235 ;
        RECT 258.235 -106.925 258.565 -106.595 ;
        RECT 258.235 -108.285 258.565 -107.955 ;
        RECT 258.235 -109.645 258.565 -109.315 ;
        RECT 258.235 -111.005 258.565 -110.675 ;
        RECT 258.235 -112.365 258.565 -112.035 ;
        RECT 258.235 -113.725 258.565 -113.395 ;
        RECT 258.235 -115.085 258.565 -114.755 ;
        RECT 258.235 -116.445 258.565 -116.115 ;
        RECT 258.235 -117.805 258.565 -117.475 ;
        RECT 258.235 -119.165 258.565 -118.835 ;
        RECT 258.235 -120.525 258.565 -120.195 ;
        RECT 258.235 -121.885 258.565 -121.555 ;
        RECT 258.235 -123.245 258.565 -122.915 ;
        RECT 258.235 -124.605 258.565 -124.275 ;
        RECT 258.235 -125.965 258.565 -125.635 ;
        RECT 258.235 -127.325 258.565 -126.995 ;
        RECT 258.235 -128.685 258.565 -128.355 ;
        RECT 258.235 -130.045 258.565 -129.715 ;
        RECT 258.235 -131.405 258.565 -131.075 ;
        RECT 258.235 -132.765 258.565 -132.435 ;
        RECT 258.235 -134.125 258.565 -133.795 ;
        RECT 258.235 -135.485 258.565 -135.155 ;
        RECT 258.235 -136.845 258.565 -136.515 ;
        RECT 258.235 -138.205 258.565 -137.875 ;
        RECT 258.235 -139.565 258.565 -139.235 ;
        RECT 258.235 -140.925 258.565 -140.595 ;
        RECT 258.235 -142.285 258.565 -141.955 ;
        RECT 258.235 -143.645 258.565 -143.315 ;
        RECT 258.235 -145.005 258.565 -144.675 ;
        RECT 258.235 -146.365 258.565 -146.035 ;
        RECT 258.235 -147.725 258.565 -147.395 ;
        RECT 258.235 -149.085 258.565 -148.755 ;
        RECT 258.235 -150.445 258.565 -150.115 ;
        RECT 258.235 -151.805 258.565 -151.475 ;
        RECT 258.235 -153.165 258.565 -152.835 ;
        RECT 258.235 -154.525 258.565 -154.195 ;
        RECT 258.235 -155.885 258.565 -155.555 ;
        RECT 258.235 -157.245 258.565 -156.915 ;
        RECT 258.235 -158.605 258.565 -158.275 ;
        RECT 258.235 -159.965 258.565 -159.635 ;
        RECT 258.235 -161.325 258.565 -160.995 ;
        RECT 258.235 -162.685 258.565 -162.355 ;
        RECT 258.235 -164.045 258.565 -163.715 ;
        RECT 258.235 -165.405 258.565 -165.075 ;
        RECT 258.235 -166.765 258.565 -166.435 ;
        RECT 258.235 -168.125 258.565 -167.795 ;
        RECT 258.235 -169.485 258.565 -169.155 ;
        RECT 258.235 -170.845 258.565 -170.515 ;
        RECT 258.235 -172.205 258.565 -171.875 ;
        RECT 258.235 -173.565 258.565 -173.235 ;
        RECT 258.235 -174.925 258.565 -174.595 ;
        RECT 258.235 -176.285 258.565 -175.955 ;
        RECT 258.235 -177.645 258.565 -177.315 ;
        RECT 258.235 -179.005 258.565 -178.675 ;
        RECT 258.235 -184.65 258.565 -183.52 ;
        RECT 258.24 -184.765 258.56 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.595 244.04 259.925 245.17 ;
        RECT 259.595 239.875 259.925 240.205 ;
        RECT 259.595 238.515 259.925 238.845 ;
        RECT 259.595 237.155 259.925 237.485 ;
        RECT 259.6 237.155 259.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.595 -0.845 259.925 -0.515 ;
        RECT 259.595 -2.205 259.925 -1.875 ;
        RECT 259.595 -3.565 259.925 -3.235 ;
        RECT 259.6 -3.565 259.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 259.595 -124.605 259.925 -124.275 ;
        RECT 259.595 -125.965 259.925 -125.635 ;
        RECT 259.595 -127.325 259.925 -126.995 ;
        RECT 259.595 -128.685 259.925 -128.355 ;
        RECT 259.595 -130.045 259.925 -129.715 ;
        RECT 259.595 -131.405 259.925 -131.075 ;
        RECT 259.595 -132.765 259.925 -132.435 ;
        RECT 259.595 -134.125 259.925 -133.795 ;
        RECT 259.595 -135.485 259.925 -135.155 ;
        RECT 259.595 -136.845 259.925 -136.515 ;
        RECT 259.595 -138.205 259.925 -137.875 ;
        RECT 259.595 -139.565 259.925 -139.235 ;
        RECT 259.595 -140.925 259.925 -140.595 ;
        RECT 259.595 -142.285 259.925 -141.955 ;
        RECT 259.595 -143.645 259.925 -143.315 ;
        RECT 259.595 -145.005 259.925 -144.675 ;
        RECT 259.595 -146.365 259.925 -146.035 ;
        RECT 259.595 -147.725 259.925 -147.395 ;
        RECT 259.595 -149.085 259.925 -148.755 ;
        RECT 259.595 -150.445 259.925 -150.115 ;
        RECT 259.595 -151.805 259.925 -151.475 ;
        RECT 259.595 -153.165 259.925 -152.835 ;
        RECT 259.595 -154.525 259.925 -154.195 ;
        RECT 259.595 -155.885 259.925 -155.555 ;
        RECT 259.595 -157.245 259.925 -156.915 ;
        RECT 259.595 -158.605 259.925 -158.275 ;
        RECT 259.595 -159.965 259.925 -159.635 ;
        RECT 259.595 -161.325 259.925 -160.995 ;
        RECT 259.595 -162.685 259.925 -162.355 ;
        RECT 259.595 -164.045 259.925 -163.715 ;
        RECT 259.595 -165.405 259.925 -165.075 ;
        RECT 259.595 -166.765 259.925 -166.435 ;
        RECT 259.595 -168.125 259.925 -167.795 ;
        RECT 259.595 -169.485 259.925 -169.155 ;
        RECT 259.595 -170.845 259.925 -170.515 ;
        RECT 259.595 -172.205 259.925 -171.875 ;
        RECT 259.595 -173.565 259.925 -173.235 ;
        RECT 259.595 -174.925 259.925 -174.595 ;
        RECT 259.595 -176.285 259.925 -175.955 ;
        RECT 259.595 -177.645 259.925 -177.315 ;
        RECT 259.595 -179.005 259.925 -178.675 ;
        RECT 259.595 -184.65 259.925 -183.52 ;
        RECT 259.6 -184.765 259.92 -95.04 ;
        RECT 259.595 -96.045 259.925 -95.715 ;
        RECT 259.595 -97.405 259.925 -97.075 ;
        RECT 259.595 -98.765 259.925 -98.435 ;
        RECT 259.595 -100.125 259.925 -99.795 ;
        RECT 259.595 -101.485 259.925 -101.155 ;
        RECT 259.595 -102.845 259.925 -102.515 ;
        RECT 259.595 -104.205 259.925 -103.875 ;
        RECT 259.595 -105.565 259.925 -105.235 ;
        RECT 259.595 -106.925 259.925 -106.595 ;
        RECT 259.595 -108.285 259.925 -107.955 ;
        RECT 259.595 -109.645 259.925 -109.315 ;
        RECT 259.595 -111.005 259.925 -110.675 ;
        RECT 259.595 -112.365 259.925 -112.035 ;
        RECT 259.595 -113.725 259.925 -113.395 ;
        RECT 259.595 -115.085 259.925 -114.755 ;
        RECT 259.595 -116.445 259.925 -116.115 ;
        RECT 259.595 -117.805 259.925 -117.475 ;
        RECT 259.595 -119.165 259.925 -118.835 ;
        RECT 259.595 -120.525 259.925 -120.195 ;
        RECT 259.595 -121.885 259.925 -121.555 ;
        RECT 259.595 -123.245 259.925 -122.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.635 244.04 210.965 245.17 ;
        RECT 210.635 239.875 210.965 240.205 ;
        RECT 210.635 238.515 210.965 238.845 ;
        RECT 210.635 237.155 210.965 237.485 ;
        RECT 210.64 237.155 210.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.995 244.04 212.325 245.17 ;
        RECT 211.995 239.875 212.325 240.205 ;
        RECT 211.995 238.515 212.325 238.845 ;
        RECT 211.995 237.155 212.325 237.485 ;
        RECT 212 237.155 212.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.995 -0.845 212.325 -0.515 ;
        RECT 211.995 -2.205 212.325 -1.875 ;
        RECT 211.995 -3.565 212.325 -3.235 ;
        RECT 212 -3.565 212.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.995 -96.045 212.325 -95.715 ;
        RECT 211.995 -97.405 212.325 -97.075 ;
        RECT 211.995 -98.765 212.325 -98.435 ;
        RECT 211.995 -100.125 212.325 -99.795 ;
        RECT 211.995 -101.485 212.325 -101.155 ;
        RECT 211.995 -102.845 212.325 -102.515 ;
        RECT 211.995 -104.205 212.325 -103.875 ;
        RECT 211.995 -105.565 212.325 -105.235 ;
        RECT 211.995 -106.925 212.325 -106.595 ;
        RECT 211.995 -108.285 212.325 -107.955 ;
        RECT 211.995 -109.645 212.325 -109.315 ;
        RECT 211.995 -111.005 212.325 -110.675 ;
        RECT 211.995 -112.365 212.325 -112.035 ;
        RECT 211.995 -113.725 212.325 -113.395 ;
        RECT 211.995 -115.085 212.325 -114.755 ;
        RECT 211.995 -116.445 212.325 -116.115 ;
        RECT 211.995 -117.805 212.325 -117.475 ;
        RECT 211.995 -119.165 212.325 -118.835 ;
        RECT 211.995 -120.525 212.325 -120.195 ;
        RECT 211.995 -121.885 212.325 -121.555 ;
        RECT 211.995 -123.245 212.325 -122.915 ;
        RECT 211.995 -124.605 212.325 -124.275 ;
        RECT 211.995 -125.965 212.325 -125.635 ;
        RECT 211.995 -127.325 212.325 -126.995 ;
        RECT 211.995 -128.685 212.325 -128.355 ;
        RECT 211.995 -130.045 212.325 -129.715 ;
        RECT 211.995 -131.405 212.325 -131.075 ;
        RECT 211.995 -132.765 212.325 -132.435 ;
        RECT 211.995 -134.125 212.325 -133.795 ;
        RECT 211.995 -135.485 212.325 -135.155 ;
        RECT 211.995 -136.845 212.325 -136.515 ;
        RECT 211.995 -138.205 212.325 -137.875 ;
        RECT 211.995 -139.565 212.325 -139.235 ;
        RECT 211.995 -140.925 212.325 -140.595 ;
        RECT 211.995 -142.285 212.325 -141.955 ;
        RECT 211.995 -143.645 212.325 -143.315 ;
        RECT 211.995 -145.005 212.325 -144.675 ;
        RECT 211.995 -146.365 212.325 -146.035 ;
        RECT 211.995 -147.725 212.325 -147.395 ;
        RECT 211.995 -149.085 212.325 -148.755 ;
        RECT 211.995 -150.445 212.325 -150.115 ;
        RECT 211.995 -151.805 212.325 -151.475 ;
        RECT 211.995 -153.165 212.325 -152.835 ;
        RECT 211.995 -154.525 212.325 -154.195 ;
        RECT 211.995 -155.885 212.325 -155.555 ;
        RECT 211.995 -157.245 212.325 -156.915 ;
        RECT 211.995 -158.605 212.325 -158.275 ;
        RECT 211.995 -159.965 212.325 -159.635 ;
        RECT 211.995 -161.325 212.325 -160.995 ;
        RECT 211.995 -162.685 212.325 -162.355 ;
        RECT 211.995 -164.045 212.325 -163.715 ;
        RECT 211.995 -165.405 212.325 -165.075 ;
        RECT 211.995 -166.765 212.325 -166.435 ;
        RECT 211.995 -168.125 212.325 -167.795 ;
        RECT 211.995 -169.485 212.325 -169.155 ;
        RECT 211.995 -170.845 212.325 -170.515 ;
        RECT 211.995 -172.205 212.325 -171.875 ;
        RECT 211.995 -173.565 212.325 -173.235 ;
        RECT 211.995 -174.925 212.325 -174.595 ;
        RECT 211.995 -176.285 212.325 -175.955 ;
        RECT 211.995 -177.645 212.325 -177.315 ;
        RECT 211.995 -179.005 212.325 -178.675 ;
        RECT 211.995 -184.65 212.325 -183.52 ;
        RECT 212 -184.765 212.32 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.355 244.04 213.685 245.17 ;
        RECT 213.355 239.875 213.685 240.205 ;
        RECT 213.355 238.515 213.685 238.845 ;
        RECT 213.355 237.155 213.685 237.485 ;
        RECT 213.36 237.155 213.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 213.355 -0.845 213.685 -0.515 ;
        RECT 213.355 -2.205 213.685 -1.875 ;
        RECT 213.355 -3.565 213.685 -3.235 ;
        RECT 213.36 -3.565 213.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.715 244.04 215.045 245.17 ;
        RECT 214.715 239.875 215.045 240.205 ;
        RECT 214.715 238.515 215.045 238.845 ;
        RECT 214.715 237.155 215.045 237.485 ;
        RECT 214.72 237.155 215.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.715 -0.845 215.045 -0.515 ;
        RECT 214.715 -2.205 215.045 -1.875 ;
        RECT 214.715 -3.565 215.045 -3.235 ;
        RECT 214.72 -3.565 215.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.715 -96.045 215.045 -95.715 ;
        RECT 214.715 -97.405 215.045 -97.075 ;
        RECT 214.715 -98.765 215.045 -98.435 ;
        RECT 214.715 -100.125 215.045 -99.795 ;
        RECT 214.715 -101.485 215.045 -101.155 ;
        RECT 214.715 -102.845 215.045 -102.515 ;
        RECT 214.715 -104.205 215.045 -103.875 ;
        RECT 214.715 -105.565 215.045 -105.235 ;
        RECT 214.715 -106.925 215.045 -106.595 ;
        RECT 214.715 -108.285 215.045 -107.955 ;
        RECT 214.715 -109.645 215.045 -109.315 ;
        RECT 214.715 -111.005 215.045 -110.675 ;
        RECT 214.715 -112.365 215.045 -112.035 ;
        RECT 214.715 -113.725 215.045 -113.395 ;
        RECT 214.715 -115.085 215.045 -114.755 ;
        RECT 214.715 -116.445 215.045 -116.115 ;
        RECT 214.715 -117.805 215.045 -117.475 ;
        RECT 214.715 -119.165 215.045 -118.835 ;
        RECT 214.715 -120.525 215.045 -120.195 ;
        RECT 214.715 -121.885 215.045 -121.555 ;
        RECT 214.715 -123.245 215.045 -122.915 ;
        RECT 214.715 -124.605 215.045 -124.275 ;
        RECT 214.715 -125.965 215.045 -125.635 ;
        RECT 214.715 -127.325 215.045 -126.995 ;
        RECT 214.715 -128.685 215.045 -128.355 ;
        RECT 214.715 -130.045 215.045 -129.715 ;
        RECT 214.715 -131.405 215.045 -131.075 ;
        RECT 214.715 -132.765 215.045 -132.435 ;
        RECT 214.715 -134.125 215.045 -133.795 ;
        RECT 214.715 -135.485 215.045 -135.155 ;
        RECT 214.715 -136.845 215.045 -136.515 ;
        RECT 214.715 -138.205 215.045 -137.875 ;
        RECT 214.715 -139.565 215.045 -139.235 ;
        RECT 214.715 -140.925 215.045 -140.595 ;
        RECT 214.715 -142.285 215.045 -141.955 ;
        RECT 214.715 -143.645 215.045 -143.315 ;
        RECT 214.715 -145.005 215.045 -144.675 ;
        RECT 214.715 -146.365 215.045 -146.035 ;
        RECT 214.715 -147.725 215.045 -147.395 ;
        RECT 214.715 -149.085 215.045 -148.755 ;
        RECT 214.715 -150.445 215.045 -150.115 ;
        RECT 214.715 -151.805 215.045 -151.475 ;
        RECT 214.715 -153.165 215.045 -152.835 ;
        RECT 214.715 -154.525 215.045 -154.195 ;
        RECT 214.715 -155.885 215.045 -155.555 ;
        RECT 214.715 -157.245 215.045 -156.915 ;
        RECT 214.715 -158.605 215.045 -158.275 ;
        RECT 214.715 -159.965 215.045 -159.635 ;
        RECT 214.715 -161.325 215.045 -160.995 ;
        RECT 214.715 -162.685 215.045 -162.355 ;
        RECT 214.715 -164.045 215.045 -163.715 ;
        RECT 214.715 -165.405 215.045 -165.075 ;
        RECT 214.715 -166.765 215.045 -166.435 ;
        RECT 214.715 -168.125 215.045 -167.795 ;
        RECT 214.715 -169.485 215.045 -169.155 ;
        RECT 214.715 -170.845 215.045 -170.515 ;
        RECT 214.715 -172.205 215.045 -171.875 ;
        RECT 214.715 -173.565 215.045 -173.235 ;
        RECT 214.715 -174.925 215.045 -174.595 ;
        RECT 214.715 -176.285 215.045 -175.955 ;
        RECT 214.715 -177.645 215.045 -177.315 ;
        RECT 214.715 -179.005 215.045 -178.675 ;
        RECT 214.715 -184.65 215.045 -183.52 ;
        RECT 214.72 -184.765 215.04 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.075 244.04 216.405 245.17 ;
        RECT 216.075 239.875 216.405 240.205 ;
        RECT 216.075 238.515 216.405 238.845 ;
        RECT 216.075 237.155 216.405 237.485 ;
        RECT 216.08 237.155 216.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.075 -0.845 216.405 -0.515 ;
        RECT 216.075 -2.205 216.405 -1.875 ;
        RECT 216.075 -3.565 216.405 -3.235 ;
        RECT 216.08 -3.565 216.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.075 -96.045 216.405 -95.715 ;
        RECT 216.075 -97.405 216.405 -97.075 ;
        RECT 216.075 -98.765 216.405 -98.435 ;
        RECT 216.075 -100.125 216.405 -99.795 ;
        RECT 216.075 -101.485 216.405 -101.155 ;
        RECT 216.075 -102.845 216.405 -102.515 ;
        RECT 216.075 -104.205 216.405 -103.875 ;
        RECT 216.075 -105.565 216.405 -105.235 ;
        RECT 216.075 -106.925 216.405 -106.595 ;
        RECT 216.075 -108.285 216.405 -107.955 ;
        RECT 216.075 -109.645 216.405 -109.315 ;
        RECT 216.075 -111.005 216.405 -110.675 ;
        RECT 216.075 -112.365 216.405 -112.035 ;
        RECT 216.075 -113.725 216.405 -113.395 ;
        RECT 216.075 -115.085 216.405 -114.755 ;
        RECT 216.075 -116.445 216.405 -116.115 ;
        RECT 216.075 -117.805 216.405 -117.475 ;
        RECT 216.075 -119.165 216.405 -118.835 ;
        RECT 216.075 -120.525 216.405 -120.195 ;
        RECT 216.075 -121.885 216.405 -121.555 ;
        RECT 216.075 -123.245 216.405 -122.915 ;
        RECT 216.075 -124.605 216.405 -124.275 ;
        RECT 216.075 -125.965 216.405 -125.635 ;
        RECT 216.075 -127.325 216.405 -126.995 ;
        RECT 216.075 -128.685 216.405 -128.355 ;
        RECT 216.075 -130.045 216.405 -129.715 ;
        RECT 216.075 -131.405 216.405 -131.075 ;
        RECT 216.075 -132.765 216.405 -132.435 ;
        RECT 216.075 -134.125 216.405 -133.795 ;
        RECT 216.075 -135.485 216.405 -135.155 ;
        RECT 216.075 -136.845 216.405 -136.515 ;
        RECT 216.075 -138.205 216.405 -137.875 ;
        RECT 216.075 -139.565 216.405 -139.235 ;
        RECT 216.075 -140.925 216.405 -140.595 ;
        RECT 216.075 -142.285 216.405 -141.955 ;
        RECT 216.075 -143.645 216.405 -143.315 ;
        RECT 216.075 -145.005 216.405 -144.675 ;
        RECT 216.075 -146.365 216.405 -146.035 ;
        RECT 216.075 -147.725 216.405 -147.395 ;
        RECT 216.075 -149.085 216.405 -148.755 ;
        RECT 216.075 -150.445 216.405 -150.115 ;
        RECT 216.075 -151.805 216.405 -151.475 ;
        RECT 216.075 -153.165 216.405 -152.835 ;
        RECT 216.075 -154.525 216.405 -154.195 ;
        RECT 216.075 -155.885 216.405 -155.555 ;
        RECT 216.075 -157.245 216.405 -156.915 ;
        RECT 216.075 -158.605 216.405 -158.275 ;
        RECT 216.075 -159.965 216.405 -159.635 ;
        RECT 216.075 -161.325 216.405 -160.995 ;
        RECT 216.075 -162.685 216.405 -162.355 ;
        RECT 216.075 -164.045 216.405 -163.715 ;
        RECT 216.075 -165.405 216.405 -165.075 ;
        RECT 216.075 -166.765 216.405 -166.435 ;
        RECT 216.075 -168.125 216.405 -167.795 ;
        RECT 216.075 -169.485 216.405 -169.155 ;
        RECT 216.075 -170.845 216.405 -170.515 ;
        RECT 216.075 -172.205 216.405 -171.875 ;
        RECT 216.075 -173.565 216.405 -173.235 ;
        RECT 216.075 -174.925 216.405 -174.595 ;
        RECT 216.075 -176.285 216.405 -175.955 ;
        RECT 216.075 -177.645 216.405 -177.315 ;
        RECT 216.075 -179.005 216.405 -178.675 ;
        RECT 216.075 -184.65 216.405 -183.52 ;
        RECT 216.08 -184.765 216.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.435 244.04 217.765 245.17 ;
        RECT 217.435 239.875 217.765 240.205 ;
        RECT 217.435 238.515 217.765 238.845 ;
        RECT 217.435 237.155 217.765 237.485 ;
        RECT 217.44 237.155 217.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.435 -0.845 217.765 -0.515 ;
        RECT 217.435 -2.205 217.765 -1.875 ;
        RECT 217.435 -3.565 217.765 -3.235 ;
        RECT 217.44 -3.565 217.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 217.435 -96.045 217.765 -95.715 ;
        RECT 217.435 -97.405 217.765 -97.075 ;
        RECT 217.435 -98.765 217.765 -98.435 ;
        RECT 217.435 -100.125 217.765 -99.795 ;
        RECT 217.435 -101.485 217.765 -101.155 ;
        RECT 217.435 -102.845 217.765 -102.515 ;
        RECT 217.435 -104.205 217.765 -103.875 ;
        RECT 217.435 -105.565 217.765 -105.235 ;
        RECT 217.435 -106.925 217.765 -106.595 ;
        RECT 217.435 -108.285 217.765 -107.955 ;
        RECT 217.435 -109.645 217.765 -109.315 ;
        RECT 217.435 -111.005 217.765 -110.675 ;
        RECT 217.435 -112.365 217.765 -112.035 ;
        RECT 217.435 -113.725 217.765 -113.395 ;
        RECT 217.435 -115.085 217.765 -114.755 ;
        RECT 217.435 -116.445 217.765 -116.115 ;
        RECT 217.435 -117.805 217.765 -117.475 ;
        RECT 217.435 -119.165 217.765 -118.835 ;
        RECT 217.435 -120.525 217.765 -120.195 ;
        RECT 217.435 -121.885 217.765 -121.555 ;
        RECT 217.435 -123.245 217.765 -122.915 ;
        RECT 217.435 -124.605 217.765 -124.275 ;
        RECT 217.435 -125.965 217.765 -125.635 ;
        RECT 217.435 -127.325 217.765 -126.995 ;
        RECT 217.435 -128.685 217.765 -128.355 ;
        RECT 217.435 -130.045 217.765 -129.715 ;
        RECT 217.435 -131.405 217.765 -131.075 ;
        RECT 217.435 -132.765 217.765 -132.435 ;
        RECT 217.435 -134.125 217.765 -133.795 ;
        RECT 217.435 -135.485 217.765 -135.155 ;
        RECT 217.435 -136.845 217.765 -136.515 ;
        RECT 217.435 -138.205 217.765 -137.875 ;
        RECT 217.435 -139.565 217.765 -139.235 ;
        RECT 217.435 -140.925 217.765 -140.595 ;
        RECT 217.435 -142.285 217.765 -141.955 ;
        RECT 217.435 -143.645 217.765 -143.315 ;
        RECT 217.435 -145.005 217.765 -144.675 ;
        RECT 217.435 -146.365 217.765 -146.035 ;
        RECT 217.435 -147.725 217.765 -147.395 ;
        RECT 217.435 -149.085 217.765 -148.755 ;
        RECT 217.435 -150.445 217.765 -150.115 ;
        RECT 217.435 -151.805 217.765 -151.475 ;
        RECT 217.435 -153.165 217.765 -152.835 ;
        RECT 217.435 -154.525 217.765 -154.195 ;
        RECT 217.435 -155.885 217.765 -155.555 ;
        RECT 217.435 -157.245 217.765 -156.915 ;
        RECT 217.435 -158.605 217.765 -158.275 ;
        RECT 217.435 -159.965 217.765 -159.635 ;
        RECT 217.435 -161.325 217.765 -160.995 ;
        RECT 217.435 -162.685 217.765 -162.355 ;
        RECT 217.435 -164.045 217.765 -163.715 ;
        RECT 217.435 -165.405 217.765 -165.075 ;
        RECT 217.435 -166.765 217.765 -166.435 ;
        RECT 217.435 -168.125 217.765 -167.795 ;
        RECT 217.435 -169.485 217.765 -169.155 ;
        RECT 217.435 -170.845 217.765 -170.515 ;
        RECT 217.435 -172.205 217.765 -171.875 ;
        RECT 217.435 -173.565 217.765 -173.235 ;
        RECT 217.435 -174.925 217.765 -174.595 ;
        RECT 217.435 -176.285 217.765 -175.955 ;
        RECT 217.435 -177.645 217.765 -177.315 ;
        RECT 217.435 -179.005 217.765 -178.675 ;
        RECT 217.435 -184.65 217.765 -183.52 ;
        RECT 217.44 -184.765 217.76 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.795 244.04 219.125 245.17 ;
        RECT 218.795 239.875 219.125 240.205 ;
        RECT 218.795 238.515 219.125 238.845 ;
        RECT 218.795 237.155 219.125 237.485 ;
        RECT 218.8 237.155 219.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.795 -0.845 219.125 -0.515 ;
        RECT 218.795 -2.205 219.125 -1.875 ;
        RECT 218.795 -3.565 219.125 -3.235 ;
        RECT 218.8 -3.565 219.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.795 -96.045 219.125 -95.715 ;
        RECT 218.795 -97.405 219.125 -97.075 ;
        RECT 218.795 -98.765 219.125 -98.435 ;
        RECT 218.795 -100.125 219.125 -99.795 ;
        RECT 218.795 -101.485 219.125 -101.155 ;
        RECT 218.795 -102.845 219.125 -102.515 ;
        RECT 218.795 -104.205 219.125 -103.875 ;
        RECT 218.795 -105.565 219.125 -105.235 ;
        RECT 218.795 -106.925 219.125 -106.595 ;
        RECT 218.795 -108.285 219.125 -107.955 ;
        RECT 218.795 -109.645 219.125 -109.315 ;
        RECT 218.795 -111.005 219.125 -110.675 ;
        RECT 218.795 -112.365 219.125 -112.035 ;
        RECT 218.795 -113.725 219.125 -113.395 ;
        RECT 218.795 -115.085 219.125 -114.755 ;
        RECT 218.795 -116.445 219.125 -116.115 ;
        RECT 218.795 -117.805 219.125 -117.475 ;
        RECT 218.795 -119.165 219.125 -118.835 ;
        RECT 218.795 -120.525 219.125 -120.195 ;
        RECT 218.795 -121.885 219.125 -121.555 ;
        RECT 218.795 -123.245 219.125 -122.915 ;
        RECT 218.795 -124.605 219.125 -124.275 ;
        RECT 218.795 -125.965 219.125 -125.635 ;
        RECT 218.795 -127.325 219.125 -126.995 ;
        RECT 218.795 -128.685 219.125 -128.355 ;
        RECT 218.795 -130.045 219.125 -129.715 ;
        RECT 218.795 -131.405 219.125 -131.075 ;
        RECT 218.795 -132.765 219.125 -132.435 ;
        RECT 218.795 -134.125 219.125 -133.795 ;
        RECT 218.795 -135.485 219.125 -135.155 ;
        RECT 218.795 -136.845 219.125 -136.515 ;
        RECT 218.795 -138.205 219.125 -137.875 ;
        RECT 218.795 -139.565 219.125 -139.235 ;
        RECT 218.795 -140.925 219.125 -140.595 ;
        RECT 218.795 -142.285 219.125 -141.955 ;
        RECT 218.795 -143.645 219.125 -143.315 ;
        RECT 218.795 -145.005 219.125 -144.675 ;
        RECT 218.795 -146.365 219.125 -146.035 ;
        RECT 218.795 -147.725 219.125 -147.395 ;
        RECT 218.795 -149.085 219.125 -148.755 ;
        RECT 218.795 -150.445 219.125 -150.115 ;
        RECT 218.795 -151.805 219.125 -151.475 ;
        RECT 218.795 -153.165 219.125 -152.835 ;
        RECT 218.795 -154.525 219.125 -154.195 ;
        RECT 218.795 -155.885 219.125 -155.555 ;
        RECT 218.795 -157.245 219.125 -156.915 ;
        RECT 218.795 -158.605 219.125 -158.275 ;
        RECT 218.795 -159.965 219.125 -159.635 ;
        RECT 218.795 -161.325 219.125 -160.995 ;
        RECT 218.795 -162.685 219.125 -162.355 ;
        RECT 218.795 -164.045 219.125 -163.715 ;
        RECT 218.795 -165.405 219.125 -165.075 ;
        RECT 218.795 -166.765 219.125 -166.435 ;
        RECT 218.795 -168.125 219.125 -167.795 ;
        RECT 218.795 -169.485 219.125 -169.155 ;
        RECT 218.795 -170.845 219.125 -170.515 ;
        RECT 218.795 -172.205 219.125 -171.875 ;
        RECT 218.795 -173.565 219.125 -173.235 ;
        RECT 218.795 -174.925 219.125 -174.595 ;
        RECT 218.795 -176.285 219.125 -175.955 ;
        RECT 218.795 -177.645 219.125 -177.315 ;
        RECT 218.795 -179.005 219.125 -178.675 ;
        RECT 218.795 -184.65 219.125 -183.52 ;
        RECT 218.8 -184.765 219.12 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.155 244.04 220.485 245.17 ;
        RECT 220.155 239.875 220.485 240.205 ;
        RECT 220.155 238.515 220.485 238.845 ;
        RECT 220.155 237.155 220.485 237.485 ;
        RECT 220.16 237.155 220.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.155 -98.765 220.485 -98.435 ;
        RECT 220.155 -100.125 220.485 -99.795 ;
        RECT 220.155 -101.485 220.485 -101.155 ;
        RECT 220.155 -102.845 220.485 -102.515 ;
        RECT 220.155 -104.205 220.485 -103.875 ;
        RECT 220.155 -105.565 220.485 -105.235 ;
        RECT 220.155 -106.925 220.485 -106.595 ;
        RECT 220.155 -108.285 220.485 -107.955 ;
        RECT 220.155 -109.645 220.485 -109.315 ;
        RECT 220.155 -111.005 220.485 -110.675 ;
        RECT 220.155 -112.365 220.485 -112.035 ;
        RECT 220.155 -113.725 220.485 -113.395 ;
        RECT 220.155 -115.085 220.485 -114.755 ;
        RECT 220.155 -116.445 220.485 -116.115 ;
        RECT 220.155 -117.805 220.485 -117.475 ;
        RECT 220.155 -119.165 220.485 -118.835 ;
        RECT 220.155 -120.525 220.485 -120.195 ;
        RECT 220.155 -121.885 220.485 -121.555 ;
        RECT 220.155 -123.245 220.485 -122.915 ;
        RECT 220.155 -124.605 220.485 -124.275 ;
        RECT 220.155 -125.965 220.485 -125.635 ;
        RECT 220.155 -127.325 220.485 -126.995 ;
        RECT 220.155 -128.685 220.485 -128.355 ;
        RECT 220.155 -130.045 220.485 -129.715 ;
        RECT 220.155 -131.405 220.485 -131.075 ;
        RECT 220.155 -132.765 220.485 -132.435 ;
        RECT 220.155 -134.125 220.485 -133.795 ;
        RECT 220.155 -135.485 220.485 -135.155 ;
        RECT 220.155 -136.845 220.485 -136.515 ;
        RECT 220.155 -138.205 220.485 -137.875 ;
        RECT 220.155 -139.565 220.485 -139.235 ;
        RECT 220.155 -140.925 220.485 -140.595 ;
        RECT 220.155 -142.285 220.485 -141.955 ;
        RECT 220.155 -143.645 220.485 -143.315 ;
        RECT 220.155 -145.005 220.485 -144.675 ;
        RECT 220.155 -146.365 220.485 -146.035 ;
        RECT 220.155 -147.725 220.485 -147.395 ;
        RECT 220.155 -149.085 220.485 -148.755 ;
        RECT 220.155 -150.445 220.485 -150.115 ;
        RECT 220.155 -151.805 220.485 -151.475 ;
        RECT 220.155 -153.165 220.485 -152.835 ;
        RECT 220.155 -154.525 220.485 -154.195 ;
        RECT 220.155 -155.885 220.485 -155.555 ;
        RECT 220.155 -157.245 220.485 -156.915 ;
        RECT 220.155 -158.605 220.485 -158.275 ;
        RECT 220.155 -159.965 220.485 -159.635 ;
        RECT 220.155 -161.325 220.485 -160.995 ;
        RECT 220.155 -162.685 220.485 -162.355 ;
        RECT 220.155 -164.045 220.485 -163.715 ;
        RECT 220.155 -165.405 220.485 -165.075 ;
        RECT 220.155 -166.765 220.485 -166.435 ;
        RECT 220.155 -168.125 220.485 -167.795 ;
        RECT 220.155 -169.485 220.485 -169.155 ;
        RECT 220.155 -170.845 220.485 -170.515 ;
        RECT 220.155 -172.205 220.485 -171.875 ;
        RECT 220.155 -173.565 220.485 -173.235 ;
        RECT 220.155 -174.925 220.485 -174.595 ;
        RECT 220.155 -176.285 220.485 -175.955 ;
        RECT 220.155 -177.645 220.485 -177.315 ;
        RECT 220.155 -179.005 220.485 -178.675 ;
        RECT 220.155 -184.65 220.485 -183.52 ;
        RECT 220.16 -184.765 220.48 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.66 -98.075 220.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.515 244.04 221.845 245.17 ;
        RECT 221.515 239.875 221.845 240.205 ;
        RECT 221.515 238.515 221.845 238.845 ;
        RECT 221.515 237.155 221.845 237.485 ;
        RECT 221.52 237.155 221.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.875 244.04 223.205 245.17 ;
        RECT 222.875 239.875 223.205 240.205 ;
        RECT 222.875 238.515 223.205 238.845 ;
        RECT 222.875 237.155 223.205 237.485 ;
        RECT 222.88 237.155 223.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.875 -0.845 223.205 -0.515 ;
        RECT 222.875 -2.205 223.205 -1.875 ;
        RECT 222.875 -3.565 223.205 -3.235 ;
        RECT 222.88 -3.565 223.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.875 -96.045 223.205 -95.715 ;
        RECT 222.875 -97.405 223.205 -97.075 ;
        RECT 222.875 -98.765 223.205 -98.435 ;
        RECT 222.875 -100.125 223.205 -99.795 ;
        RECT 222.875 -101.485 223.205 -101.155 ;
        RECT 222.875 -102.845 223.205 -102.515 ;
        RECT 222.875 -104.205 223.205 -103.875 ;
        RECT 222.875 -105.565 223.205 -105.235 ;
        RECT 222.875 -106.925 223.205 -106.595 ;
        RECT 222.875 -108.285 223.205 -107.955 ;
        RECT 222.875 -109.645 223.205 -109.315 ;
        RECT 222.875 -111.005 223.205 -110.675 ;
        RECT 222.875 -112.365 223.205 -112.035 ;
        RECT 222.875 -113.725 223.205 -113.395 ;
        RECT 222.875 -115.085 223.205 -114.755 ;
        RECT 222.875 -116.445 223.205 -116.115 ;
        RECT 222.875 -117.805 223.205 -117.475 ;
        RECT 222.875 -119.165 223.205 -118.835 ;
        RECT 222.875 -120.525 223.205 -120.195 ;
        RECT 222.875 -121.885 223.205 -121.555 ;
        RECT 222.875 -123.245 223.205 -122.915 ;
        RECT 222.875 -124.605 223.205 -124.275 ;
        RECT 222.875 -125.965 223.205 -125.635 ;
        RECT 222.875 -127.325 223.205 -126.995 ;
        RECT 222.875 -128.685 223.205 -128.355 ;
        RECT 222.875 -130.045 223.205 -129.715 ;
        RECT 222.875 -131.405 223.205 -131.075 ;
        RECT 222.875 -132.765 223.205 -132.435 ;
        RECT 222.875 -134.125 223.205 -133.795 ;
        RECT 222.875 -135.485 223.205 -135.155 ;
        RECT 222.875 -136.845 223.205 -136.515 ;
        RECT 222.875 -138.205 223.205 -137.875 ;
        RECT 222.875 -139.565 223.205 -139.235 ;
        RECT 222.875 -140.925 223.205 -140.595 ;
        RECT 222.875 -142.285 223.205 -141.955 ;
        RECT 222.875 -143.645 223.205 -143.315 ;
        RECT 222.875 -145.005 223.205 -144.675 ;
        RECT 222.875 -146.365 223.205 -146.035 ;
        RECT 222.875 -147.725 223.205 -147.395 ;
        RECT 222.875 -149.085 223.205 -148.755 ;
        RECT 222.875 -150.445 223.205 -150.115 ;
        RECT 222.875 -151.805 223.205 -151.475 ;
        RECT 222.875 -153.165 223.205 -152.835 ;
        RECT 222.875 -154.525 223.205 -154.195 ;
        RECT 222.875 -155.885 223.205 -155.555 ;
        RECT 222.875 -157.245 223.205 -156.915 ;
        RECT 222.875 -158.605 223.205 -158.275 ;
        RECT 222.875 -159.965 223.205 -159.635 ;
        RECT 222.875 -161.325 223.205 -160.995 ;
        RECT 222.875 -162.685 223.205 -162.355 ;
        RECT 222.875 -164.045 223.205 -163.715 ;
        RECT 222.875 -165.405 223.205 -165.075 ;
        RECT 222.875 -166.765 223.205 -166.435 ;
        RECT 222.875 -168.125 223.205 -167.795 ;
        RECT 222.875 -169.485 223.205 -169.155 ;
        RECT 222.875 -170.845 223.205 -170.515 ;
        RECT 222.875 -172.205 223.205 -171.875 ;
        RECT 222.875 -173.565 223.205 -173.235 ;
        RECT 222.875 -174.925 223.205 -174.595 ;
        RECT 222.875 -176.285 223.205 -175.955 ;
        RECT 222.875 -177.645 223.205 -177.315 ;
        RECT 222.875 -179.005 223.205 -178.675 ;
        RECT 222.875 -184.65 223.205 -183.52 ;
        RECT 222.88 -184.765 223.2 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.235 244.04 224.565 245.17 ;
        RECT 224.235 239.875 224.565 240.205 ;
        RECT 224.235 238.515 224.565 238.845 ;
        RECT 224.235 237.155 224.565 237.485 ;
        RECT 224.24 237.155 224.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.235 -0.845 224.565 -0.515 ;
        RECT 224.235 -2.205 224.565 -1.875 ;
        RECT 224.235 -3.565 224.565 -3.235 ;
        RECT 224.24 -3.565 224.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.595 244.04 225.925 245.17 ;
        RECT 225.595 239.875 225.925 240.205 ;
        RECT 225.595 238.515 225.925 238.845 ;
        RECT 225.595 237.155 225.925 237.485 ;
        RECT 225.6 237.155 225.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.595 -0.845 225.925 -0.515 ;
        RECT 225.595 -2.205 225.925 -1.875 ;
        RECT 225.595 -3.565 225.925 -3.235 ;
        RECT 225.6 -3.565 225.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 225.595 -96.045 225.925 -95.715 ;
        RECT 225.595 -97.405 225.925 -97.075 ;
        RECT 225.595 -98.765 225.925 -98.435 ;
        RECT 225.595 -100.125 225.925 -99.795 ;
        RECT 225.595 -101.485 225.925 -101.155 ;
        RECT 225.595 -102.845 225.925 -102.515 ;
        RECT 225.595 -104.205 225.925 -103.875 ;
        RECT 225.595 -105.565 225.925 -105.235 ;
        RECT 225.595 -106.925 225.925 -106.595 ;
        RECT 225.595 -108.285 225.925 -107.955 ;
        RECT 225.595 -109.645 225.925 -109.315 ;
        RECT 225.595 -111.005 225.925 -110.675 ;
        RECT 225.595 -112.365 225.925 -112.035 ;
        RECT 225.595 -113.725 225.925 -113.395 ;
        RECT 225.595 -115.085 225.925 -114.755 ;
        RECT 225.595 -116.445 225.925 -116.115 ;
        RECT 225.595 -117.805 225.925 -117.475 ;
        RECT 225.595 -119.165 225.925 -118.835 ;
        RECT 225.595 -120.525 225.925 -120.195 ;
        RECT 225.595 -121.885 225.925 -121.555 ;
        RECT 225.595 -123.245 225.925 -122.915 ;
        RECT 225.595 -124.605 225.925 -124.275 ;
        RECT 225.595 -125.965 225.925 -125.635 ;
        RECT 225.595 -127.325 225.925 -126.995 ;
        RECT 225.595 -128.685 225.925 -128.355 ;
        RECT 225.595 -130.045 225.925 -129.715 ;
        RECT 225.595 -131.405 225.925 -131.075 ;
        RECT 225.595 -132.765 225.925 -132.435 ;
        RECT 225.595 -134.125 225.925 -133.795 ;
        RECT 225.595 -135.485 225.925 -135.155 ;
        RECT 225.595 -136.845 225.925 -136.515 ;
        RECT 225.595 -138.205 225.925 -137.875 ;
        RECT 225.595 -139.565 225.925 -139.235 ;
        RECT 225.595 -140.925 225.925 -140.595 ;
        RECT 225.595 -142.285 225.925 -141.955 ;
        RECT 225.595 -143.645 225.925 -143.315 ;
        RECT 225.595 -145.005 225.925 -144.675 ;
        RECT 225.595 -146.365 225.925 -146.035 ;
        RECT 225.595 -147.725 225.925 -147.395 ;
        RECT 225.595 -149.085 225.925 -148.755 ;
        RECT 225.595 -150.445 225.925 -150.115 ;
        RECT 225.595 -151.805 225.925 -151.475 ;
        RECT 225.595 -153.165 225.925 -152.835 ;
        RECT 225.595 -154.525 225.925 -154.195 ;
        RECT 225.595 -155.885 225.925 -155.555 ;
        RECT 225.595 -157.245 225.925 -156.915 ;
        RECT 225.595 -158.605 225.925 -158.275 ;
        RECT 225.595 -159.965 225.925 -159.635 ;
        RECT 225.595 -161.325 225.925 -160.995 ;
        RECT 225.595 -162.685 225.925 -162.355 ;
        RECT 225.595 -164.045 225.925 -163.715 ;
        RECT 225.595 -165.405 225.925 -165.075 ;
        RECT 225.595 -166.765 225.925 -166.435 ;
        RECT 225.595 -168.125 225.925 -167.795 ;
        RECT 225.595 -169.485 225.925 -169.155 ;
        RECT 225.595 -170.845 225.925 -170.515 ;
        RECT 225.595 -172.205 225.925 -171.875 ;
        RECT 225.595 -173.565 225.925 -173.235 ;
        RECT 225.595 -174.925 225.925 -174.595 ;
        RECT 225.595 -176.285 225.925 -175.955 ;
        RECT 225.595 -177.645 225.925 -177.315 ;
        RECT 225.595 -179.005 225.925 -178.675 ;
        RECT 225.595 -184.65 225.925 -183.52 ;
        RECT 225.6 -184.765 225.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.955 244.04 227.285 245.17 ;
        RECT 226.955 239.875 227.285 240.205 ;
        RECT 226.955 238.515 227.285 238.845 ;
        RECT 226.955 237.155 227.285 237.485 ;
        RECT 226.96 237.155 227.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.955 -0.845 227.285 -0.515 ;
        RECT 226.955 -2.205 227.285 -1.875 ;
        RECT 226.955 -3.565 227.285 -3.235 ;
        RECT 226.96 -3.565 227.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.955 -96.045 227.285 -95.715 ;
        RECT 226.955 -97.405 227.285 -97.075 ;
        RECT 226.955 -98.765 227.285 -98.435 ;
        RECT 226.955 -100.125 227.285 -99.795 ;
        RECT 226.955 -101.485 227.285 -101.155 ;
        RECT 226.955 -102.845 227.285 -102.515 ;
        RECT 226.955 -104.205 227.285 -103.875 ;
        RECT 226.955 -105.565 227.285 -105.235 ;
        RECT 226.955 -106.925 227.285 -106.595 ;
        RECT 226.955 -108.285 227.285 -107.955 ;
        RECT 226.955 -109.645 227.285 -109.315 ;
        RECT 226.955 -111.005 227.285 -110.675 ;
        RECT 226.955 -112.365 227.285 -112.035 ;
        RECT 226.955 -113.725 227.285 -113.395 ;
        RECT 226.955 -115.085 227.285 -114.755 ;
        RECT 226.955 -116.445 227.285 -116.115 ;
        RECT 226.955 -117.805 227.285 -117.475 ;
        RECT 226.955 -119.165 227.285 -118.835 ;
        RECT 226.955 -120.525 227.285 -120.195 ;
        RECT 226.955 -121.885 227.285 -121.555 ;
        RECT 226.955 -123.245 227.285 -122.915 ;
        RECT 226.955 -124.605 227.285 -124.275 ;
        RECT 226.955 -125.965 227.285 -125.635 ;
        RECT 226.955 -127.325 227.285 -126.995 ;
        RECT 226.955 -128.685 227.285 -128.355 ;
        RECT 226.955 -130.045 227.285 -129.715 ;
        RECT 226.955 -131.405 227.285 -131.075 ;
        RECT 226.955 -132.765 227.285 -132.435 ;
        RECT 226.955 -134.125 227.285 -133.795 ;
        RECT 226.955 -135.485 227.285 -135.155 ;
        RECT 226.955 -136.845 227.285 -136.515 ;
        RECT 226.955 -138.205 227.285 -137.875 ;
        RECT 226.955 -139.565 227.285 -139.235 ;
        RECT 226.955 -140.925 227.285 -140.595 ;
        RECT 226.955 -142.285 227.285 -141.955 ;
        RECT 226.955 -143.645 227.285 -143.315 ;
        RECT 226.955 -145.005 227.285 -144.675 ;
        RECT 226.955 -146.365 227.285 -146.035 ;
        RECT 226.955 -147.725 227.285 -147.395 ;
        RECT 226.955 -149.085 227.285 -148.755 ;
        RECT 226.955 -150.445 227.285 -150.115 ;
        RECT 226.955 -151.805 227.285 -151.475 ;
        RECT 226.955 -153.165 227.285 -152.835 ;
        RECT 226.955 -154.525 227.285 -154.195 ;
        RECT 226.955 -155.885 227.285 -155.555 ;
        RECT 226.955 -157.245 227.285 -156.915 ;
        RECT 226.955 -158.605 227.285 -158.275 ;
        RECT 226.955 -159.965 227.285 -159.635 ;
        RECT 226.955 -161.325 227.285 -160.995 ;
        RECT 226.955 -162.685 227.285 -162.355 ;
        RECT 226.955 -164.045 227.285 -163.715 ;
        RECT 226.955 -165.405 227.285 -165.075 ;
        RECT 226.955 -166.765 227.285 -166.435 ;
        RECT 226.955 -168.125 227.285 -167.795 ;
        RECT 226.955 -169.485 227.285 -169.155 ;
        RECT 226.955 -170.845 227.285 -170.515 ;
        RECT 226.955 -172.205 227.285 -171.875 ;
        RECT 226.955 -173.565 227.285 -173.235 ;
        RECT 226.955 -174.925 227.285 -174.595 ;
        RECT 226.955 -176.285 227.285 -175.955 ;
        RECT 226.955 -177.645 227.285 -177.315 ;
        RECT 226.955 -179.005 227.285 -178.675 ;
        RECT 226.955 -184.65 227.285 -183.52 ;
        RECT 226.96 -184.765 227.28 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.315 244.04 228.645 245.17 ;
        RECT 228.315 239.875 228.645 240.205 ;
        RECT 228.315 238.515 228.645 238.845 ;
        RECT 228.315 237.155 228.645 237.485 ;
        RECT 228.32 237.155 228.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.315 -0.845 228.645 -0.515 ;
        RECT 228.315 -2.205 228.645 -1.875 ;
        RECT 228.315 -3.565 228.645 -3.235 ;
        RECT 228.32 -3.565 228.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.315 -96.045 228.645 -95.715 ;
        RECT 228.315 -97.405 228.645 -97.075 ;
        RECT 228.315 -98.765 228.645 -98.435 ;
        RECT 228.315 -100.125 228.645 -99.795 ;
        RECT 228.315 -101.485 228.645 -101.155 ;
        RECT 228.315 -102.845 228.645 -102.515 ;
        RECT 228.315 -104.205 228.645 -103.875 ;
        RECT 228.315 -105.565 228.645 -105.235 ;
        RECT 228.315 -106.925 228.645 -106.595 ;
        RECT 228.315 -108.285 228.645 -107.955 ;
        RECT 228.315 -109.645 228.645 -109.315 ;
        RECT 228.315 -111.005 228.645 -110.675 ;
        RECT 228.315 -112.365 228.645 -112.035 ;
        RECT 228.315 -113.725 228.645 -113.395 ;
        RECT 228.315 -115.085 228.645 -114.755 ;
        RECT 228.315 -116.445 228.645 -116.115 ;
        RECT 228.315 -117.805 228.645 -117.475 ;
        RECT 228.315 -119.165 228.645 -118.835 ;
        RECT 228.315 -120.525 228.645 -120.195 ;
        RECT 228.315 -121.885 228.645 -121.555 ;
        RECT 228.315 -123.245 228.645 -122.915 ;
        RECT 228.315 -124.605 228.645 -124.275 ;
        RECT 228.315 -125.965 228.645 -125.635 ;
        RECT 228.315 -127.325 228.645 -126.995 ;
        RECT 228.315 -128.685 228.645 -128.355 ;
        RECT 228.315 -130.045 228.645 -129.715 ;
        RECT 228.315 -131.405 228.645 -131.075 ;
        RECT 228.315 -132.765 228.645 -132.435 ;
        RECT 228.315 -134.125 228.645 -133.795 ;
        RECT 228.315 -135.485 228.645 -135.155 ;
        RECT 228.315 -136.845 228.645 -136.515 ;
        RECT 228.315 -138.205 228.645 -137.875 ;
        RECT 228.315 -139.565 228.645 -139.235 ;
        RECT 228.315 -140.925 228.645 -140.595 ;
        RECT 228.315 -142.285 228.645 -141.955 ;
        RECT 228.315 -143.645 228.645 -143.315 ;
        RECT 228.315 -145.005 228.645 -144.675 ;
        RECT 228.315 -146.365 228.645 -146.035 ;
        RECT 228.315 -147.725 228.645 -147.395 ;
        RECT 228.315 -149.085 228.645 -148.755 ;
        RECT 228.315 -150.445 228.645 -150.115 ;
        RECT 228.315 -151.805 228.645 -151.475 ;
        RECT 228.315 -153.165 228.645 -152.835 ;
        RECT 228.315 -154.525 228.645 -154.195 ;
        RECT 228.315 -155.885 228.645 -155.555 ;
        RECT 228.315 -157.245 228.645 -156.915 ;
        RECT 228.315 -158.605 228.645 -158.275 ;
        RECT 228.315 -159.965 228.645 -159.635 ;
        RECT 228.315 -161.325 228.645 -160.995 ;
        RECT 228.315 -162.685 228.645 -162.355 ;
        RECT 228.315 -164.045 228.645 -163.715 ;
        RECT 228.315 -165.405 228.645 -165.075 ;
        RECT 228.315 -166.765 228.645 -166.435 ;
        RECT 228.315 -168.125 228.645 -167.795 ;
        RECT 228.315 -169.485 228.645 -169.155 ;
        RECT 228.315 -170.845 228.645 -170.515 ;
        RECT 228.315 -172.205 228.645 -171.875 ;
        RECT 228.315 -173.565 228.645 -173.235 ;
        RECT 228.315 -174.925 228.645 -174.595 ;
        RECT 228.315 -176.285 228.645 -175.955 ;
        RECT 228.315 -177.645 228.645 -177.315 ;
        RECT 228.315 -179.005 228.645 -178.675 ;
        RECT 228.315 -184.65 228.645 -183.52 ;
        RECT 228.32 -184.765 228.64 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.675 244.04 230.005 245.17 ;
        RECT 229.675 239.875 230.005 240.205 ;
        RECT 229.675 238.515 230.005 238.845 ;
        RECT 229.675 237.155 230.005 237.485 ;
        RECT 229.68 237.155 230 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.675 -0.845 230.005 -0.515 ;
        RECT 229.675 -2.205 230.005 -1.875 ;
        RECT 229.675 -3.565 230.005 -3.235 ;
        RECT 229.68 -3.565 230 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 229.675 -96.045 230.005 -95.715 ;
        RECT 229.675 -97.405 230.005 -97.075 ;
        RECT 229.675 -98.765 230.005 -98.435 ;
        RECT 229.675 -100.125 230.005 -99.795 ;
        RECT 229.675 -101.485 230.005 -101.155 ;
        RECT 229.675 -102.845 230.005 -102.515 ;
        RECT 229.675 -104.205 230.005 -103.875 ;
        RECT 229.675 -105.565 230.005 -105.235 ;
        RECT 229.675 -106.925 230.005 -106.595 ;
        RECT 229.675 -108.285 230.005 -107.955 ;
        RECT 229.675 -109.645 230.005 -109.315 ;
        RECT 229.675 -111.005 230.005 -110.675 ;
        RECT 229.675 -112.365 230.005 -112.035 ;
        RECT 229.675 -113.725 230.005 -113.395 ;
        RECT 229.675 -115.085 230.005 -114.755 ;
        RECT 229.675 -116.445 230.005 -116.115 ;
        RECT 229.675 -117.805 230.005 -117.475 ;
        RECT 229.675 -119.165 230.005 -118.835 ;
        RECT 229.675 -120.525 230.005 -120.195 ;
        RECT 229.675 -121.885 230.005 -121.555 ;
        RECT 229.675 -123.245 230.005 -122.915 ;
        RECT 229.675 -124.605 230.005 -124.275 ;
        RECT 229.675 -125.965 230.005 -125.635 ;
        RECT 229.675 -127.325 230.005 -126.995 ;
        RECT 229.675 -128.685 230.005 -128.355 ;
        RECT 229.675 -130.045 230.005 -129.715 ;
        RECT 229.675 -131.405 230.005 -131.075 ;
        RECT 229.675 -132.765 230.005 -132.435 ;
        RECT 229.675 -134.125 230.005 -133.795 ;
        RECT 229.675 -135.485 230.005 -135.155 ;
        RECT 229.675 -136.845 230.005 -136.515 ;
        RECT 229.675 -138.205 230.005 -137.875 ;
        RECT 229.675 -139.565 230.005 -139.235 ;
        RECT 229.675 -140.925 230.005 -140.595 ;
        RECT 229.675 -142.285 230.005 -141.955 ;
        RECT 229.675 -143.645 230.005 -143.315 ;
        RECT 229.675 -145.005 230.005 -144.675 ;
        RECT 229.675 -146.365 230.005 -146.035 ;
        RECT 229.675 -147.725 230.005 -147.395 ;
        RECT 229.675 -149.085 230.005 -148.755 ;
        RECT 229.675 -150.445 230.005 -150.115 ;
        RECT 229.675 -151.805 230.005 -151.475 ;
        RECT 229.675 -153.165 230.005 -152.835 ;
        RECT 229.675 -154.525 230.005 -154.195 ;
        RECT 229.675 -155.885 230.005 -155.555 ;
        RECT 229.675 -157.245 230.005 -156.915 ;
        RECT 229.675 -158.605 230.005 -158.275 ;
        RECT 229.675 -159.965 230.005 -159.635 ;
        RECT 229.675 -161.325 230.005 -160.995 ;
        RECT 229.675 -162.685 230.005 -162.355 ;
        RECT 229.675 -164.045 230.005 -163.715 ;
        RECT 229.675 -165.405 230.005 -165.075 ;
        RECT 229.675 -166.765 230.005 -166.435 ;
        RECT 229.675 -168.125 230.005 -167.795 ;
        RECT 229.675 -169.485 230.005 -169.155 ;
        RECT 229.675 -170.845 230.005 -170.515 ;
        RECT 229.675 -172.205 230.005 -171.875 ;
        RECT 229.675 -173.565 230.005 -173.235 ;
        RECT 229.675 -174.925 230.005 -174.595 ;
        RECT 229.675 -176.285 230.005 -175.955 ;
        RECT 229.675 -177.645 230.005 -177.315 ;
        RECT 229.675 -179.005 230.005 -178.675 ;
        RECT 229.675 -184.65 230.005 -183.52 ;
        RECT 229.68 -184.765 230 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.035 244.04 231.365 245.17 ;
        RECT 231.035 239.875 231.365 240.205 ;
        RECT 231.035 238.515 231.365 238.845 ;
        RECT 231.035 237.155 231.365 237.485 ;
        RECT 231.04 237.155 231.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.035 -98.765 231.365 -98.435 ;
        RECT 231.035 -100.125 231.365 -99.795 ;
        RECT 231.035 -101.485 231.365 -101.155 ;
        RECT 231.035 -102.845 231.365 -102.515 ;
        RECT 231.035 -104.205 231.365 -103.875 ;
        RECT 231.035 -105.565 231.365 -105.235 ;
        RECT 231.035 -106.925 231.365 -106.595 ;
        RECT 231.035 -108.285 231.365 -107.955 ;
        RECT 231.035 -109.645 231.365 -109.315 ;
        RECT 231.035 -111.005 231.365 -110.675 ;
        RECT 231.035 -112.365 231.365 -112.035 ;
        RECT 231.035 -113.725 231.365 -113.395 ;
        RECT 231.035 -115.085 231.365 -114.755 ;
        RECT 231.035 -116.445 231.365 -116.115 ;
        RECT 231.035 -117.805 231.365 -117.475 ;
        RECT 231.035 -119.165 231.365 -118.835 ;
        RECT 231.035 -120.525 231.365 -120.195 ;
        RECT 231.035 -121.885 231.365 -121.555 ;
        RECT 231.035 -123.245 231.365 -122.915 ;
        RECT 231.035 -124.605 231.365 -124.275 ;
        RECT 231.035 -125.965 231.365 -125.635 ;
        RECT 231.035 -127.325 231.365 -126.995 ;
        RECT 231.035 -128.685 231.365 -128.355 ;
        RECT 231.035 -130.045 231.365 -129.715 ;
        RECT 231.035 -131.405 231.365 -131.075 ;
        RECT 231.035 -132.765 231.365 -132.435 ;
        RECT 231.035 -134.125 231.365 -133.795 ;
        RECT 231.035 -135.485 231.365 -135.155 ;
        RECT 231.035 -136.845 231.365 -136.515 ;
        RECT 231.035 -138.205 231.365 -137.875 ;
        RECT 231.035 -139.565 231.365 -139.235 ;
        RECT 231.035 -140.925 231.365 -140.595 ;
        RECT 231.035 -142.285 231.365 -141.955 ;
        RECT 231.035 -143.645 231.365 -143.315 ;
        RECT 231.035 -145.005 231.365 -144.675 ;
        RECT 231.035 -146.365 231.365 -146.035 ;
        RECT 231.035 -147.725 231.365 -147.395 ;
        RECT 231.035 -149.085 231.365 -148.755 ;
        RECT 231.035 -150.445 231.365 -150.115 ;
        RECT 231.035 -151.805 231.365 -151.475 ;
        RECT 231.035 -153.165 231.365 -152.835 ;
        RECT 231.035 -154.525 231.365 -154.195 ;
        RECT 231.035 -155.885 231.365 -155.555 ;
        RECT 231.035 -157.245 231.365 -156.915 ;
        RECT 231.035 -158.605 231.365 -158.275 ;
        RECT 231.035 -159.965 231.365 -159.635 ;
        RECT 231.035 -161.325 231.365 -160.995 ;
        RECT 231.035 -162.685 231.365 -162.355 ;
        RECT 231.035 -164.045 231.365 -163.715 ;
        RECT 231.035 -165.405 231.365 -165.075 ;
        RECT 231.035 -166.765 231.365 -166.435 ;
        RECT 231.035 -168.125 231.365 -167.795 ;
        RECT 231.035 -169.485 231.365 -169.155 ;
        RECT 231.035 -170.845 231.365 -170.515 ;
        RECT 231.035 -172.205 231.365 -171.875 ;
        RECT 231.035 -173.565 231.365 -173.235 ;
        RECT 231.035 -174.925 231.365 -174.595 ;
        RECT 231.035 -176.285 231.365 -175.955 ;
        RECT 231.035 -177.645 231.365 -177.315 ;
        RECT 231.035 -179.005 231.365 -178.675 ;
        RECT 231.035 -184.65 231.365 -183.52 ;
        RECT 231.04 -184.765 231.36 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.56 -98.075 231.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.395 244.04 232.725 245.17 ;
        RECT 232.395 239.875 232.725 240.205 ;
        RECT 232.395 238.515 232.725 238.845 ;
        RECT 232.395 237.155 232.725 237.485 ;
        RECT 232.4 237.155 232.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.755 244.04 234.085 245.17 ;
        RECT 233.755 239.875 234.085 240.205 ;
        RECT 233.755 238.515 234.085 238.845 ;
        RECT 233.755 237.155 234.085 237.485 ;
        RECT 233.76 237.155 234.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.755 -0.845 234.085 -0.515 ;
        RECT 233.755 -2.205 234.085 -1.875 ;
        RECT 233.755 -3.565 234.085 -3.235 ;
        RECT 233.76 -3.565 234.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.755 -96.045 234.085 -95.715 ;
        RECT 233.755 -97.405 234.085 -97.075 ;
        RECT 233.755 -98.765 234.085 -98.435 ;
        RECT 233.755 -100.125 234.085 -99.795 ;
        RECT 233.755 -101.485 234.085 -101.155 ;
        RECT 233.755 -102.845 234.085 -102.515 ;
        RECT 233.755 -104.205 234.085 -103.875 ;
        RECT 233.755 -105.565 234.085 -105.235 ;
        RECT 233.755 -106.925 234.085 -106.595 ;
        RECT 233.755 -108.285 234.085 -107.955 ;
        RECT 233.755 -109.645 234.085 -109.315 ;
        RECT 233.755 -111.005 234.085 -110.675 ;
        RECT 233.755 -112.365 234.085 -112.035 ;
        RECT 233.755 -113.725 234.085 -113.395 ;
        RECT 233.755 -115.085 234.085 -114.755 ;
        RECT 233.755 -116.445 234.085 -116.115 ;
        RECT 233.755 -117.805 234.085 -117.475 ;
        RECT 233.755 -119.165 234.085 -118.835 ;
        RECT 233.755 -120.525 234.085 -120.195 ;
        RECT 233.755 -121.885 234.085 -121.555 ;
        RECT 233.755 -123.245 234.085 -122.915 ;
        RECT 233.755 -124.605 234.085 -124.275 ;
        RECT 233.755 -125.965 234.085 -125.635 ;
        RECT 233.755 -127.325 234.085 -126.995 ;
        RECT 233.755 -128.685 234.085 -128.355 ;
        RECT 233.755 -130.045 234.085 -129.715 ;
        RECT 233.755 -131.405 234.085 -131.075 ;
        RECT 233.755 -132.765 234.085 -132.435 ;
        RECT 233.755 -134.125 234.085 -133.795 ;
        RECT 233.755 -135.485 234.085 -135.155 ;
        RECT 233.755 -136.845 234.085 -136.515 ;
        RECT 233.755 -138.205 234.085 -137.875 ;
        RECT 233.755 -139.565 234.085 -139.235 ;
        RECT 233.755 -140.925 234.085 -140.595 ;
        RECT 233.755 -142.285 234.085 -141.955 ;
        RECT 233.755 -143.645 234.085 -143.315 ;
        RECT 233.755 -145.005 234.085 -144.675 ;
        RECT 233.755 -146.365 234.085 -146.035 ;
        RECT 233.755 -147.725 234.085 -147.395 ;
        RECT 233.755 -149.085 234.085 -148.755 ;
        RECT 233.755 -150.445 234.085 -150.115 ;
        RECT 233.755 -151.805 234.085 -151.475 ;
        RECT 233.755 -153.165 234.085 -152.835 ;
        RECT 233.755 -154.525 234.085 -154.195 ;
        RECT 233.755 -155.885 234.085 -155.555 ;
        RECT 233.755 -157.245 234.085 -156.915 ;
        RECT 233.755 -158.605 234.085 -158.275 ;
        RECT 233.755 -159.965 234.085 -159.635 ;
        RECT 233.755 -161.325 234.085 -160.995 ;
        RECT 233.755 -162.685 234.085 -162.355 ;
        RECT 233.755 -164.045 234.085 -163.715 ;
        RECT 233.755 -165.405 234.085 -165.075 ;
        RECT 233.755 -166.765 234.085 -166.435 ;
        RECT 233.755 -168.125 234.085 -167.795 ;
        RECT 233.755 -169.485 234.085 -169.155 ;
        RECT 233.755 -170.845 234.085 -170.515 ;
        RECT 233.755 -172.205 234.085 -171.875 ;
        RECT 233.755 -173.565 234.085 -173.235 ;
        RECT 233.755 -174.925 234.085 -174.595 ;
        RECT 233.755 -176.285 234.085 -175.955 ;
        RECT 233.755 -177.645 234.085 -177.315 ;
        RECT 233.755 -179.005 234.085 -178.675 ;
        RECT 233.755 -184.65 234.085 -183.52 ;
        RECT 233.76 -184.765 234.08 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.115 244.04 235.445 245.17 ;
        RECT 235.115 239.875 235.445 240.205 ;
        RECT 235.115 238.515 235.445 238.845 ;
        RECT 235.115 237.155 235.445 237.485 ;
        RECT 235.12 237.155 235.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.115 -0.845 235.445 -0.515 ;
        RECT 235.115 -2.205 235.445 -1.875 ;
        RECT 235.115 -3.565 235.445 -3.235 ;
        RECT 235.12 -3.565 235.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.475 244.04 236.805 245.17 ;
        RECT 236.475 239.875 236.805 240.205 ;
        RECT 236.475 238.515 236.805 238.845 ;
        RECT 236.475 237.155 236.805 237.485 ;
        RECT 236.48 237.155 236.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.475 -0.845 236.805 -0.515 ;
        RECT 236.475 -2.205 236.805 -1.875 ;
        RECT 236.475 -3.565 236.805 -3.235 ;
        RECT 236.48 -3.565 236.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 236.475 -169.485 236.805 -169.155 ;
        RECT 236.475 -170.845 236.805 -170.515 ;
        RECT 236.475 -172.205 236.805 -171.875 ;
        RECT 236.475 -173.565 236.805 -173.235 ;
        RECT 236.475 -174.925 236.805 -174.595 ;
        RECT 236.475 -176.285 236.805 -175.955 ;
        RECT 236.475 -177.645 236.805 -177.315 ;
        RECT 236.475 -179.005 236.805 -178.675 ;
        RECT 236.475 -184.65 236.805 -183.52 ;
        RECT 236.48 -184.765 236.8 -95.04 ;
        RECT 236.475 -96.045 236.805 -95.715 ;
        RECT 236.475 -97.405 236.805 -97.075 ;
        RECT 236.475 -98.765 236.805 -98.435 ;
        RECT 236.475 -100.125 236.805 -99.795 ;
        RECT 236.475 -101.485 236.805 -101.155 ;
        RECT 236.475 -102.845 236.805 -102.515 ;
        RECT 236.475 -104.205 236.805 -103.875 ;
        RECT 236.475 -105.565 236.805 -105.235 ;
        RECT 236.475 -106.925 236.805 -106.595 ;
        RECT 236.475 -108.285 236.805 -107.955 ;
        RECT 236.475 -109.645 236.805 -109.315 ;
        RECT 236.475 -111.005 236.805 -110.675 ;
        RECT 236.475 -112.365 236.805 -112.035 ;
        RECT 236.475 -113.725 236.805 -113.395 ;
        RECT 236.475 -115.085 236.805 -114.755 ;
        RECT 236.475 -116.445 236.805 -116.115 ;
        RECT 236.475 -117.805 236.805 -117.475 ;
        RECT 236.475 -119.165 236.805 -118.835 ;
        RECT 236.475 -120.525 236.805 -120.195 ;
        RECT 236.475 -121.885 236.805 -121.555 ;
        RECT 236.475 -123.245 236.805 -122.915 ;
        RECT 236.475 -124.605 236.805 -124.275 ;
        RECT 236.475 -125.965 236.805 -125.635 ;
        RECT 236.475 -127.325 236.805 -126.995 ;
        RECT 236.475 -128.685 236.805 -128.355 ;
        RECT 236.475 -130.045 236.805 -129.715 ;
        RECT 236.475 -131.405 236.805 -131.075 ;
        RECT 236.475 -132.765 236.805 -132.435 ;
        RECT 236.475 -134.125 236.805 -133.795 ;
        RECT 236.475 -135.485 236.805 -135.155 ;
        RECT 236.475 -136.845 236.805 -136.515 ;
        RECT 236.475 -138.205 236.805 -137.875 ;
        RECT 236.475 -139.565 236.805 -139.235 ;
        RECT 236.475 -140.925 236.805 -140.595 ;
        RECT 236.475 -142.285 236.805 -141.955 ;
        RECT 236.475 -143.645 236.805 -143.315 ;
        RECT 236.475 -145.005 236.805 -144.675 ;
        RECT 236.475 -146.365 236.805 -146.035 ;
        RECT 236.475 -147.725 236.805 -147.395 ;
        RECT 236.475 -149.085 236.805 -148.755 ;
        RECT 236.475 -150.445 236.805 -150.115 ;
        RECT 236.475 -151.805 236.805 -151.475 ;
        RECT 236.475 -153.165 236.805 -152.835 ;
        RECT 236.475 -154.525 236.805 -154.195 ;
        RECT 236.475 -155.885 236.805 -155.555 ;
        RECT 236.475 -157.245 236.805 -156.915 ;
        RECT 236.475 -158.605 236.805 -158.275 ;
        RECT 236.475 -159.965 236.805 -159.635 ;
        RECT 236.475 -161.325 236.805 -160.995 ;
        RECT 236.475 -162.685 236.805 -162.355 ;
        RECT 236.475 -164.045 236.805 -163.715 ;
        RECT 236.475 -165.405 236.805 -165.075 ;
        RECT 236.475 -166.765 236.805 -166.435 ;
        RECT 236.475 -168.125 236.805 -167.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 244.04 186.485 245.17 ;
        RECT 186.155 239.875 186.485 240.205 ;
        RECT 186.155 238.515 186.485 238.845 ;
        RECT 186.155 237.155 186.485 237.485 ;
        RECT 186.16 237.155 186.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 -0.845 186.485 -0.515 ;
        RECT 186.155 -2.205 186.485 -1.875 ;
        RECT 186.155 -3.565 186.485 -3.235 ;
        RECT 186.16 -3.565 186.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.155 -96.045 186.485 -95.715 ;
        RECT 186.155 -97.405 186.485 -97.075 ;
        RECT 186.155 -98.765 186.485 -98.435 ;
        RECT 186.155 -100.125 186.485 -99.795 ;
        RECT 186.155 -101.485 186.485 -101.155 ;
        RECT 186.155 -102.845 186.485 -102.515 ;
        RECT 186.155 -104.205 186.485 -103.875 ;
        RECT 186.155 -105.565 186.485 -105.235 ;
        RECT 186.155 -106.925 186.485 -106.595 ;
        RECT 186.155 -108.285 186.485 -107.955 ;
        RECT 186.155 -109.645 186.485 -109.315 ;
        RECT 186.155 -111.005 186.485 -110.675 ;
        RECT 186.155 -112.365 186.485 -112.035 ;
        RECT 186.155 -113.725 186.485 -113.395 ;
        RECT 186.155 -115.085 186.485 -114.755 ;
        RECT 186.155 -116.445 186.485 -116.115 ;
        RECT 186.155 -117.805 186.485 -117.475 ;
        RECT 186.155 -119.165 186.485 -118.835 ;
        RECT 186.155 -120.525 186.485 -120.195 ;
        RECT 186.155 -121.885 186.485 -121.555 ;
        RECT 186.155 -123.245 186.485 -122.915 ;
        RECT 186.155 -124.605 186.485 -124.275 ;
        RECT 186.155 -125.965 186.485 -125.635 ;
        RECT 186.155 -127.325 186.485 -126.995 ;
        RECT 186.155 -128.685 186.485 -128.355 ;
        RECT 186.155 -130.045 186.485 -129.715 ;
        RECT 186.155 -131.405 186.485 -131.075 ;
        RECT 186.155 -132.765 186.485 -132.435 ;
        RECT 186.155 -134.125 186.485 -133.795 ;
        RECT 186.155 -135.485 186.485 -135.155 ;
        RECT 186.155 -136.845 186.485 -136.515 ;
        RECT 186.155 -138.205 186.485 -137.875 ;
        RECT 186.155 -139.565 186.485 -139.235 ;
        RECT 186.155 -140.925 186.485 -140.595 ;
        RECT 186.155 -142.285 186.485 -141.955 ;
        RECT 186.155 -143.645 186.485 -143.315 ;
        RECT 186.155 -145.005 186.485 -144.675 ;
        RECT 186.155 -146.365 186.485 -146.035 ;
        RECT 186.155 -147.725 186.485 -147.395 ;
        RECT 186.155 -149.085 186.485 -148.755 ;
        RECT 186.155 -150.445 186.485 -150.115 ;
        RECT 186.155 -151.805 186.485 -151.475 ;
        RECT 186.155 -153.165 186.485 -152.835 ;
        RECT 186.155 -154.525 186.485 -154.195 ;
        RECT 186.155 -155.885 186.485 -155.555 ;
        RECT 186.155 -157.245 186.485 -156.915 ;
        RECT 186.155 -158.605 186.485 -158.275 ;
        RECT 186.155 -159.965 186.485 -159.635 ;
        RECT 186.155 -161.325 186.485 -160.995 ;
        RECT 186.155 -162.685 186.485 -162.355 ;
        RECT 186.155 -164.045 186.485 -163.715 ;
        RECT 186.155 -165.405 186.485 -165.075 ;
        RECT 186.155 -166.765 186.485 -166.435 ;
        RECT 186.155 -168.125 186.485 -167.795 ;
        RECT 186.155 -169.485 186.485 -169.155 ;
        RECT 186.155 -170.845 186.485 -170.515 ;
        RECT 186.155 -172.205 186.485 -171.875 ;
        RECT 186.155 -173.565 186.485 -173.235 ;
        RECT 186.155 -174.925 186.485 -174.595 ;
        RECT 186.155 -176.285 186.485 -175.955 ;
        RECT 186.155 -177.645 186.485 -177.315 ;
        RECT 186.155 -179.005 186.485 -178.675 ;
        RECT 186.155 -184.65 186.485 -183.52 ;
        RECT 186.16 -184.765 186.48 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 244.04 187.845 245.17 ;
        RECT 187.515 239.875 187.845 240.205 ;
        RECT 187.515 238.515 187.845 238.845 ;
        RECT 187.515 237.155 187.845 237.485 ;
        RECT 187.52 237.155 187.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.515 -98.765 187.845 -98.435 ;
        RECT 187.515 -100.125 187.845 -99.795 ;
        RECT 187.515 -101.485 187.845 -101.155 ;
        RECT 187.515 -102.845 187.845 -102.515 ;
        RECT 187.515 -104.205 187.845 -103.875 ;
        RECT 187.515 -105.565 187.845 -105.235 ;
        RECT 187.515 -106.925 187.845 -106.595 ;
        RECT 187.515 -108.285 187.845 -107.955 ;
        RECT 187.515 -109.645 187.845 -109.315 ;
        RECT 187.515 -111.005 187.845 -110.675 ;
        RECT 187.515 -112.365 187.845 -112.035 ;
        RECT 187.515 -113.725 187.845 -113.395 ;
        RECT 187.515 -115.085 187.845 -114.755 ;
        RECT 187.515 -116.445 187.845 -116.115 ;
        RECT 187.515 -117.805 187.845 -117.475 ;
        RECT 187.515 -119.165 187.845 -118.835 ;
        RECT 187.515 -120.525 187.845 -120.195 ;
        RECT 187.515 -121.885 187.845 -121.555 ;
        RECT 187.515 -123.245 187.845 -122.915 ;
        RECT 187.515 -124.605 187.845 -124.275 ;
        RECT 187.515 -125.965 187.845 -125.635 ;
        RECT 187.515 -127.325 187.845 -126.995 ;
        RECT 187.515 -128.685 187.845 -128.355 ;
        RECT 187.515 -130.045 187.845 -129.715 ;
        RECT 187.515 -131.405 187.845 -131.075 ;
        RECT 187.515 -132.765 187.845 -132.435 ;
        RECT 187.515 -134.125 187.845 -133.795 ;
        RECT 187.515 -135.485 187.845 -135.155 ;
        RECT 187.515 -136.845 187.845 -136.515 ;
        RECT 187.515 -138.205 187.845 -137.875 ;
        RECT 187.515 -139.565 187.845 -139.235 ;
        RECT 187.515 -140.925 187.845 -140.595 ;
        RECT 187.515 -142.285 187.845 -141.955 ;
        RECT 187.515 -143.645 187.845 -143.315 ;
        RECT 187.515 -145.005 187.845 -144.675 ;
        RECT 187.515 -146.365 187.845 -146.035 ;
        RECT 187.515 -147.725 187.845 -147.395 ;
        RECT 187.515 -149.085 187.845 -148.755 ;
        RECT 187.515 -150.445 187.845 -150.115 ;
        RECT 187.515 -151.805 187.845 -151.475 ;
        RECT 187.515 -153.165 187.845 -152.835 ;
        RECT 187.515 -154.525 187.845 -154.195 ;
        RECT 187.515 -155.885 187.845 -155.555 ;
        RECT 187.515 -157.245 187.845 -156.915 ;
        RECT 187.515 -158.605 187.845 -158.275 ;
        RECT 187.515 -159.965 187.845 -159.635 ;
        RECT 187.515 -161.325 187.845 -160.995 ;
        RECT 187.515 -162.685 187.845 -162.355 ;
        RECT 187.515 -164.045 187.845 -163.715 ;
        RECT 187.515 -165.405 187.845 -165.075 ;
        RECT 187.515 -166.765 187.845 -166.435 ;
        RECT 187.515 -168.125 187.845 -167.795 ;
        RECT 187.515 -169.485 187.845 -169.155 ;
        RECT 187.515 -170.845 187.845 -170.515 ;
        RECT 187.515 -172.205 187.845 -171.875 ;
        RECT 187.515 -173.565 187.845 -173.235 ;
        RECT 187.515 -174.925 187.845 -174.595 ;
        RECT 187.515 -176.285 187.845 -175.955 ;
        RECT 187.515 -177.645 187.845 -177.315 ;
        RECT 187.515 -179.005 187.845 -178.675 ;
        RECT 187.515 -184.65 187.845 -183.52 ;
        RECT 187.52 -184.765 187.84 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 187.96 -98.075 188.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.875 244.04 189.205 245.17 ;
        RECT 188.875 239.875 189.205 240.205 ;
        RECT 188.875 238.515 189.205 238.845 ;
        RECT 188.875 237.155 189.205 237.485 ;
        RECT 188.88 237.155 189.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 244.04 190.565 245.17 ;
        RECT 190.235 239.875 190.565 240.205 ;
        RECT 190.235 238.515 190.565 238.845 ;
        RECT 190.235 237.155 190.565 237.485 ;
        RECT 190.24 237.155 190.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.235 -0.845 190.565 -0.515 ;
        RECT 190.235 -2.205 190.565 -1.875 ;
        RECT 190.235 -3.565 190.565 -3.235 ;
        RECT 190.24 -3.565 190.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 244.04 191.925 245.17 ;
        RECT 191.595 239.875 191.925 240.205 ;
        RECT 191.595 238.515 191.925 238.845 ;
        RECT 191.595 237.155 191.925 237.485 ;
        RECT 191.6 237.155 191.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 191.595 -0.845 191.925 -0.515 ;
        RECT 191.595 -2.205 191.925 -1.875 ;
        RECT 191.595 -3.565 191.925 -3.235 ;
        RECT 191.6 -3.565 191.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.955 244.04 193.285 245.17 ;
        RECT 192.955 239.875 193.285 240.205 ;
        RECT 192.955 238.515 193.285 238.845 ;
        RECT 192.955 237.155 193.285 237.485 ;
        RECT 192.96 237.155 193.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.955 -0.845 193.285 -0.515 ;
        RECT 192.955 -2.205 193.285 -1.875 ;
        RECT 192.955 -3.565 193.285 -3.235 ;
        RECT 192.96 -3.565 193.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.955 -96.045 193.285 -95.715 ;
        RECT 192.955 -97.405 193.285 -97.075 ;
        RECT 192.955 -98.765 193.285 -98.435 ;
        RECT 192.955 -100.125 193.285 -99.795 ;
        RECT 192.955 -101.485 193.285 -101.155 ;
        RECT 192.955 -102.845 193.285 -102.515 ;
        RECT 192.955 -104.205 193.285 -103.875 ;
        RECT 192.955 -105.565 193.285 -105.235 ;
        RECT 192.955 -106.925 193.285 -106.595 ;
        RECT 192.955 -108.285 193.285 -107.955 ;
        RECT 192.955 -109.645 193.285 -109.315 ;
        RECT 192.955 -111.005 193.285 -110.675 ;
        RECT 192.955 -112.365 193.285 -112.035 ;
        RECT 192.955 -113.725 193.285 -113.395 ;
        RECT 192.955 -115.085 193.285 -114.755 ;
        RECT 192.955 -116.445 193.285 -116.115 ;
        RECT 192.955 -117.805 193.285 -117.475 ;
        RECT 192.955 -119.165 193.285 -118.835 ;
        RECT 192.955 -120.525 193.285 -120.195 ;
        RECT 192.955 -121.885 193.285 -121.555 ;
        RECT 192.955 -123.245 193.285 -122.915 ;
        RECT 192.955 -124.605 193.285 -124.275 ;
        RECT 192.955 -125.965 193.285 -125.635 ;
        RECT 192.955 -127.325 193.285 -126.995 ;
        RECT 192.955 -128.685 193.285 -128.355 ;
        RECT 192.955 -130.045 193.285 -129.715 ;
        RECT 192.955 -131.405 193.285 -131.075 ;
        RECT 192.955 -132.765 193.285 -132.435 ;
        RECT 192.955 -134.125 193.285 -133.795 ;
        RECT 192.955 -135.485 193.285 -135.155 ;
        RECT 192.955 -136.845 193.285 -136.515 ;
        RECT 192.955 -138.205 193.285 -137.875 ;
        RECT 192.955 -139.565 193.285 -139.235 ;
        RECT 192.955 -140.925 193.285 -140.595 ;
        RECT 192.955 -142.285 193.285 -141.955 ;
        RECT 192.955 -143.645 193.285 -143.315 ;
        RECT 192.955 -145.005 193.285 -144.675 ;
        RECT 192.955 -146.365 193.285 -146.035 ;
        RECT 192.955 -147.725 193.285 -147.395 ;
        RECT 192.955 -149.085 193.285 -148.755 ;
        RECT 192.955 -150.445 193.285 -150.115 ;
        RECT 192.955 -151.805 193.285 -151.475 ;
        RECT 192.955 -153.165 193.285 -152.835 ;
        RECT 192.955 -154.525 193.285 -154.195 ;
        RECT 192.955 -155.885 193.285 -155.555 ;
        RECT 192.955 -157.245 193.285 -156.915 ;
        RECT 192.955 -158.605 193.285 -158.275 ;
        RECT 192.955 -159.965 193.285 -159.635 ;
        RECT 192.955 -161.325 193.285 -160.995 ;
        RECT 192.955 -162.685 193.285 -162.355 ;
        RECT 192.955 -164.045 193.285 -163.715 ;
        RECT 192.955 -165.405 193.285 -165.075 ;
        RECT 192.955 -166.765 193.285 -166.435 ;
        RECT 192.955 -168.125 193.285 -167.795 ;
        RECT 192.955 -169.485 193.285 -169.155 ;
        RECT 192.955 -170.845 193.285 -170.515 ;
        RECT 192.955 -172.205 193.285 -171.875 ;
        RECT 192.955 -173.565 193.285 -173.235 ;
        RECT 192.955 -174.925 193.285 -174.595 ;
        RECT 192.955 -176.285 193.285 -175.955 ;
        RECT 192.955 -177.645 193.285 -177.315 ;
        RECT 192.955 -179.005 193.285 -178.675 ;
        RECT 192.955 -184.65 193.285 -183.52 ;
        RECT 192.96 -184.765 193.28 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 244.04 194.645 245.17 ;
        RECT 194.315 239.875 194.645 240.205 ;
        RECT 194.315 238.515 194.645 238.845 ;
        RECT 194.315 237.155 194.645 237.485 ;
        RECT 194.32 237.155 194.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 -0.845 194.645 -0.515 ;
        RECT 194.315 -2.205 194.645 -1.875 ;
        RECT 194.315 -3.565 194.645 -3.235 ;
        RECT 194.32 -3.565 194.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.315 -96.045 194.645 -95.715 ;
        RECT 194.315 -97.405 194.645 -97.075 ;
        RECT 194.315 -98.765 194.645 -98.435 ;
        RECT 194.315 -100.125 194.645 -99.795 ;
        RECT 194.315 -101.485 194.645 -101.155 ;
        RECT 194.315 -102.845 194.645 -102.515 ;
        RECT 194.315 -104.205 194.645 -103.875 ;
        RECT 194.315 -105.565 194.645 -105.235 ;
        RECT 194.315 -106.925 194.645 -106.595 ;
        RECT 194.315 -108.285 194.645 -107.955 ;
        RECT 194.315 -109.645 194.645 -109.315 ;
        RECT 194.315 -111.005 194.645 -110.675 ;
        RECT 194.315 -112.365 194.645 -112.035 ;
        RECT 194.315 -113.725 194.645 -113.395 ;
        RECT 194.315 -115.085 194.645 -114.755 ;
        RECT 194.315 -116.445 194.645 -116.115 ;
        RECT 194.315 -117.805 194.645 -117.475 ;
        RECT 194.315 -119.165 194.645 -118.835 ;
        RECT 194.315 -120.525 194.645 -120.195 ;
        RECT 194.315 -121.885 194.645 -121.555 ;
        RECT 194.315 -123.245 194.645 -122.915 ;
        RECT 194.315 -124.605 194.645 -124.275 ;
        RECT 194.315 -125.965 194.645 -125.635 ;
        RECT 194.315 -127.325 194.645 -126.995 ;
        RECT 194.315 -128.685 194.645 -128.355 ;
        RECT 194.315 -130.045 194.645 -129.715 ;
        RECT 194.315 -131.405 194.645 -131.075 ;
        RECT 194.315 -132.765 194.645 -132.435 ;
        RECT 194.315 -134.125 194.645 -133.795 ;
        RECT 194.315 -135.485 194.645 -135.155 ;
        RECT 194.315 -136.845 194.645 -136.515 ;
        RECT 194.315 -138.205 194.645 -137.875 ;
        RECT 194.315 -139.565 194.645 -139.235 ;
        RECT 194.315 -140.925 194.645 -140.595 ;
        RECT 194.315 -142.285 194.645 -141.955 ;
        RECT 194.315 -143.645 194.645 -143.315 ;
        RECT 194.315 -145.005 194.645 -144.675 ;
        RECT 194.315 -146.365 194.645 -146.035 ;
        RECT 194.315 -147.725 194.645 -147.395 ;
        RECT 194.315 -149.085 194.645 -148.755 ;
        RECT 194.315 -150.445 194.645 -150.115 ;
        RECT 194.315 -151.805 194.645 -151.475 ;
        RECT 194.315 -153.165 194.645 -152.835 ;
        RECT 194.315 -154.525 194.645 -154.195 ;
        RECT 194.315 -155.885 194.645 -155.555 ;
        RECT 194.315 -157.245 194.645 -156.915 ;
        RECT 194.315 -158.605 194.645 -158.275 ;
        RECT 194.315 -159.965 194.645 -159.635 ;
        RECT 194.315 -161.325 194.645 -160.995 ;
        RECT 194.315 -162.685 194.645 -162.355 ;
        RECT 194.315 -164.045 194.645 -163.715 ;
        RECT 194.315 -165.405 194.645 -165.075 ;
        RECT 194.315 -166.765 194.645 -166.435 ;
        RECT 194.315 -168.125 194.645 -167.795 ;
        RECT 194.315 -169.485 194.645 -169.155 ;
        RECT 194.315 -170.845 194.645 -170.515 ;
        RECT 194.315 -172.205 194.645 -171.875 ;
        RECT 194.315 -173.565 194.645 -173.235 ;
        RECT 194.315 -174.925 194.645 -174.595 ;
        RECT 194.315 -176.285 194.645 -175.955 ;
        RECT 194.315 -177.645 194.645 -177.315 ;
        RECT 194.315 -179.005 194.645 -178.675 ;
        RECT 194.315 -184.65 194.645 -183.52 ;
        RECT 194.32 -184.765 194.64 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 244.04 196.005 245.17 ;
        RECT 195.675 239.875 196.005 240.205 ;
        RECT 195.675 238.515 196.005 238.845 ;
        RECT 195.675 237.155 196.005 237.485 ;
        RECT 195.68 237.155 196 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 -0.845 196.005 -0.515 ;
        RECT 195.675 -2.205 196.005 -1.875 ;
        RECT 195.675 -3.565 196.005 -3.235 ;
        RECT 195.68 -3.565 196 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 195.675 -96.045 196.005 -95.715 ;
        RECT 195.675 -97.405 196.005 -97.075 ;
        RECT 195.675 -98.765 196.005 -98.435 ;
        RECT 195.675 -100.125 196.005 -99.795 ;
        RECT 195.675 -101.485 196.005 -101.155 ;
        RECT 195.675 -102.845 196.005 -102.515 ;
        RECT 195.675 -104.205 196.005 -103.875 ;
        RECT 195.675 -105.565 196.005 -105.235 ;
        RECT 195.675 -106.925 196.005 -106.595 ;
        RECT 195.675 -108.285 196.005 -107.955 ;
        RECT 195.675 -109.645 196.005 -109.315 ;
        RECT 195.675 -111.005 196.005 -110.675 ;
        RECT 195.675 -112.365 196.005 -112.035 ;
        RECT 195.675 -113.725 196.005 -113.395 ;
        RECT 195.675 -115.085 196.005 -114.755 ;
        RECT 195.675 -116.445 196.005 -116.115 ;
        RECT 195.675 -117.805 196.005 -117.475 ;
        RECT 195.675 -119.165 196.005 -118.835 ;
        RECT 195.675 -120.525 196.005 -120.195 ;
        RECT 195.675 -121.885 196.005 -121.555 ;
        RECT 195.675 -123.245 196.005 -122.915 ;
        RECT 195.675 -124.605 196.005 -124.275 ;
        RECT 195.675 -125.965 196.005 -125.635 ;
        RECT 195.675 -127.325 196.005 -126.995 ;
        RECT 195.675 -128.685 196.005 -128.355 ;
        RECT 195.675 -130.045 196.005 -129.715 ;
        RECT 195.675 -131.405 196.005 -131.075 ;
        RECT 195.675 -132.765 196.005 -132.435 ;
        RECT 195.675 -134.125 196.005 -133.795 ;
        RECT 195.675 -135.485 196.005 -135.155 ;
        RECT 195.675 -136.845 196.005 -136.515 ;
        RECT 195.675 -138.205 196.005 -137.875 ;
        RECT 195.675 -139.565 196.005 -139.235 ;
        RECT 195.675 -140.925 196.005 -140.595 ;
        RECT 195.675 -142.285 196.005 -141.955 ;
        RECT 195.675 -143.645 196.005 -143.315 ;
        RECT 195.675 -145.005 196.005 -144.675 ;
        RECT 195.675 -146.365 196.005 -146.035 ;
        RECT 195.675 -147.725 196.005 -147.395 ;
        RECT 195.675 -149.085 196.005 -148.755 ;
        RECT 195.675 -150.445 196.005 -150.115 ;
        RECT 195.675 -151.805 196.005 -151.475 ;
        RECT 195.675 -153.165 196.005 -152.835 ;
        RECT 195.675 -154.525 196.005 -154.195 ;
        RECT 195.675 -155.885 196.005 -155.555 ;
        RECT 195.675 -157.245 196.005 -156.915 ;
        RECT 195.675 -158.605 196.005 -158.275 ;
        RECT 195.675 -159.965 196.005 -159.635 ;
        RECT 195.675 -161.325 196.005 -160.995 ;
        RECT 195.675 -162.685 196.005 -162.355 ;
        RECT 195.675 -164.045 196.005 -163.715 ;
        RECT 195.675 -165.405 196.005 -165.075 ;
        RECT 195.675 -166.765 196.005 -166.435 ;
        RECT 195.675 -168.125 196.005 -167.795 ;
        RECT 195.675 -169.485 196.005 -169.155 ;
        RECT 195.675 -170.845 196.005 -170.515 ;
        RECT 195.675 -172.205 196.005 -171.875 ;
        RECT 195.675 -173.565 196.005 -173.235 ;
        RECT 195.675 -174.925 196.005 -174.595 ;
        RECT 195.675 -176.285 196.005 -175.955 ;
        RECT 195.675 -177.645 196.005 -177.315 ;
        RECT 195.675 -179.005 196.005 -178.675 ;
        RECT 195.675 -184.65 196.005 -183.52 ;
        RECT 195.68 -184.765 196 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 244.04 197.365 245.17 ;
        RECT 197.035 239.875 197.365 240.205 ;
        RECT 197.035 238.515 197.365 238.845 ;
        RECT 197.035 237.155 197.365 237.485 ;
        RECT 197.04 237.155 197.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 -0.845 197.365 -0.515 ;
        RECT 197.035 -2.205 197.365 -1.875 ;
        RECT 197.035 -3.565 197.365 -3.235 ;
        RECT 197.04 -3.565 197.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.035 -96.045 197.365 -95.715 ;
        RECT 197.035 -97.405 197.365 -97.075 ;
        RECT 197.035 -98.765 197.365 -98.435 ;
        RECT 197.035 -100.125 197.365 -99.795 ;
        RECT 197.035 -101.485 197.365 -101.155 ;
        RECT 197.035 -102.845 197.365 -102.515 ;
        RECT 197.035 -104.205 197.365 -103.875 ;
        RECT 197.035 -105.565 197.365 -105.235 ;
        RECT 197.035 -106.925 197.365 -106.595 ;
        RECT 197.035 -108.285 197.365 -107.955 ;
        RECT 197.035 -109.645 197.365 -109.315 ;
        RECT 197.035 -111.005 197.365 -110.675 ;
        RECT 197.035 -112.365 197.365 -112.035 ;
        RECT 197.035 -113.725 197.365 -113.395 ;
        RECT 197.035 -115.085 197.365 -114.755 ;
        RECT 197.035 -116.445 197.365 -116.115 ;
        RECT 197.035 -117.805 197.365 -117.475 ;
        RECT 197.035 -119.165 197.365 -118.835 ;
        RECT 197.035 -120.525 197.365 -120.195 ;
        RECT 197.035 -121.885 197.365 -121.555 ;
        RECT 197.035 -123.245 197.365 -122.915 ;
        RECT 197.035 -124.605 197.365 -124.275 ;
        RECT 197.035 -125.965 197.365 -125.635 ;
        RECT 197.035 -127.325 197.365 -126.995 ;
        RECT 197.035 -128.685 197.365 -128.355 ;
        RECT 197.035 -130.045 197.365 -129.715 ;
        RECT 197.035 -131.405 197.365 -131.075 ;
        RECT 197.035 -132.765 197.365 -132.435 ;
        RECT 197.035 -134.125 197.365 -133.795 ;
        RECT 197.035 -135.485 197.365 -135.155 ;
        RECT 197.035 -136.845 197.365 -136.515 ;
        RECT 197.035 -138.205 197.365 -137.875 ;
        RECT 197.035 -139.565 197.365 -139.235 ;
        RECT 197.035 -140.925 197.365 -140.595 ;
        RECT 197.035 -142.285 197.365 -141.955 ;
        RECT 197.035 -143.645 197.365 -143.315 ;
        RECT 197.035 -145.005 197.365 -144.675 ;
        RECT 197.035 -146.365 197.365 -146.035 ;
        RECT 197.035 -147.725 197.365 -147.395 ;
        RECT 197.035 -149.085 197.365 -148.755 ;
        RECT 197.035 -150.445 197.365 -150.115 ;
        RECT 197.035 -151.805 197.365 -151.475 ;
        RECT 197.035 -153.165 197.365 -152.835 ;
        RECT 197.035 -154.525 197.365 -154.195 ;
        RECT 197.035 -155.885 197.365 -155.555 ;
        RECT 197.035 -157.245 197.365 -156.915 ;
        RECT 197.035 -158.605 197.365 -158.275 ;
        RECT 197.035 -159.965 197.365 -159.635 ;
        RECT 197.035 -161.325 197.365 -160.995 ;
        RECT 197.035 -162.685 197.365 -162.355 ;
        RECT 197.035 -164.045 197.365 -163.715 ;
        RECT 197.035 -165.405 197.365 -165.075 ;
        RECT 197.035 -166.765 197.365 -166.435 ;
        RECT 197.035 -168.125 197.365 -167.795 ;
        RECT 197.035 -169.485 197.365 -169.155 ;
        RECT 197.035 -170.845 197.365 -170.515 ;
        RECT 197.035 -172.205 197.365 -171.875 ;
        RECT 197.035 -173.565 197.365 -173.235 ;
        RECT 197.035 -174.925 197.365 -174.595 ;
        RECT 197.035 -176.285 197.365 -175.955 ;
        RECT 197.035 -177.645 197.365 -177.315 ;
        RECT 197.035 -179.005 197.365 -178.675 ;
        RECT 197.035 -184.65 197.365 -183.52 ;
        RECT 197.04 -184.765 197.36 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 244.04 198.725 245.17 ;
        RECT 198.395 239.875 198.725 240.205 ;
        RECT 198.395 238.515 198.725 238.845 ;
        RECT 198.395 237.155 198.725 237.485 ;
        RECT 198.4 237.155 198.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.395 -98.765 198.725 -98.435 ;
        RECT 198.395 -100.125 198.725 -99.795 ;
        RECT 198.395 -101.485 198.725 -101.155 ;
        RECT 198.395 -102.845 198.725 -102.515 ;
        RECT 198.395 -104.205 198.725 -103.875 ;
        RECT 198.395 -105.565 198.725 -105.235 ;
        RECT 198.395 -106.925 198.725 -106.595 ;
        RECT 198.395 -108.285 198.725 -107.955 ;
        RECT 198.395 -109.645 198.725 -109.315 ;
        RECT 198.395 -111.005 198.725 -110.675 ;
        RECT 198.395 -112.365 198.725 -112.035 ;
        RECT 198.395 -113.725 198.725 -113.395 ;
        RECT 198.395 -115.085 198.725 -114.755 ;
        RECT 198.395 -116.445 198.725 -116.115 ;
        RECT 198.395 -117.805 198.725 -117.475 ;
        RECT 198.395 -119.165 198.725 -118.835 ;
        RECT 198.395 -120.525 198.725 -120.195 ;
        RECT 198.395 -121.885 198.725 -121.555 ;
        RECT 198.395 -123.245 198.725 -122.915 ;
        RECT 198.395 -124.605 198.725 -124.275 ;
        RECT 198.395 -125.965 198.725 -125.635 ;
        RECT 198.395 -127.325 198.725 -126.995 ;
        RECT 198.395 -128.685 198.725 -128.355 ;
        RECT 198.395 -130.045 198.725 -129.715 ;
        RECT 198.395 -131.405 198.725 -131.075 ;
        RECT 198.395 -132.765 198.725 -132.435 ;
        RECT 198.395 -134.125 198.725 -133.795 ;
        RECT 198.395 -135.485 198.725 -135.155 ;
        RECT 198.395 -136.845 198.725 -136.515 ;
        RECT 198.395 -138.205 198.725 -137.875 ;
        RECT 198.395 -139.565 198.725 -139.235 ;
        RECT 198.395 -140.925 198.725 -140.595 ;
        RECT 198.395 -142.285 198.725 -141.955 ;
        RECT 198.395 -143.645 198.725 -143.315 ;
        RECT 198.395 -145.005 198.725 -144.675 ;
        RECT 198.395 -146.365 198.725 -146.035 ;
        RECT 198.395 -147.725 198.725 -147.395 ;
        RECT 198.395 -149.085 198.725 -148.755 ;
        RECT 198.395 -150.445 198.725 -150.115 ;
        RECT 198.395 -151.805 198.725 -151.475 ;
        RECT 198.395 -153.165 198.725 -152.835 ;
        RECT 198.395 -154.525 198.725 -154.195 ;
        RECT 198.395 -155.885 198.725 -155.555 ;
        RECT 198.395 -157.245 198.725 -156.915 ;
        RECT 198.395 -158.605 198.725 -158.275 ;
        RECT 198.395 -159.965 198.725 -159.635 ;
        RECT 198.395 -161.325 198.725 -160.995 ;
        RECT 198.395 -162.685 198.725 -162.355 ;
        RECT 198.395 -164.045 198.725 -163.715 ;
        RECT 198.395 -165.405 198.725 -165.075 ;
        RECT 198.395 -166.765 198.725 -166.435 ;
        RECT 198.395 -168.125 198.725 -167.795 ;
        RECT 198.395 -169.485 198.725 -169.155 ;
        RECT 198.395 -170.845 198.725 -170.515 ;
        RECT 198.395 -172.205 198.725 -171.875 ;
        RECT 198.395 -173.565 198.725 -173.235 ;
        RECT 198.395 -174.925 198.725 -174.595 ;
        RECT 198.395 -176.285 198.725 -175.955 ;
        RECT 198.395 -177.645 198.725 -177.315 ;
        RECT 198.395 -179.005 198.725 -178.675 ;
        RECT 198.395 -184.65 198.725 -183.52 ;
        RECT 198.4 -184.765 198.72 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 198.86 -98.075 199.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.755 244.04 200.085 245.17 ;
        RECT 199.755 239.875 200.085 240.205 ;
        RECT 199.755 238.515 200.085 238.845 ;
        RECT 199.755 237.155 200.085 237.485 ;
        RECT 199.76 237.155 200.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 244.04 201.445 245.17 ;
        RECT 201.115 239.875 201.445 240.205 ;
        RECT 201.115 238.515 201.445 238.845 ;
        RECT 201.115 237.155 201.445 237.485 ;
        RECT 201.12 237.155 201.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 -0.845 201.445 -0.515 ;
        RECT 201.115 -2.205 201.445 -1.875 ;
        RECT 201.115 -3.565 201.445 -3.235 ;
        RECT 201.12 -3.565 201.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.115 -96.045 201.445 -95.715 ;
        RECT 201.115 -97.405 201.445 -97.075 ;
        RECT 201.115 -98.765 201.445 -98.435 ;
        RECT 201.115 -100.125 201.445 -99.795 ;
        RECT 201.115 -101.485 201.445 -101.155 ;
        RECT 201.115 -102.845 201.445 -102.515 ;
        RECT 201.115 -104.205 201.445 -103.875 ;
        RECT 201.115 -105.565 201.445 -105.235 ;
        RECT 201.115 -106.925 201.445 -106.595 ;
        RECT 201.115 -108.285 201.445 -107.955 ;
        RECT 201.115 -109.645 201.445 -109.315 ;
        RECT 201.115 -111.005 201.445 -110.675 ;
        RECT 201.115 -112.365 201.445 -112.035 ;
        RECT 201.115 -113.725 201.445 -113.395 ;
        RECT 201.115 -115.085 201.445 -114.755 ;
        RECT 201.115 -116.445 201.445 -116.115 ;
        RECT 201.115 -117.805 201.445 -117.475 ;
        RECT 201.115 -119.165 201.445 -118.835 ;
        RECT 201.115 -120.525 201.445 -120.195 ;
        RECT 201.115 -121.885 201.445 -121.555 ;
        RECT 201.115 -123.245 201.445 -122.915 ;
        RECT 201.115 -124.605 201.445 -124.275 ;
        RECT 201.115 -125.965 201.445 -125.635 ;
        RECT 201.115 -127.325 201.445 -126.995 ;
        RECT 201.115 -128.685 201.445 -128.355 ;
        RECT 201.115 -130.045 201.445 -129.715 ;
        RECT 201.115 -131.405 201.445 -131.075 ;
        RECT 201.115 -132.765 201.445 -132.435 ;
        RECT 201.115 -134.125 201.445 -133.795 ;
        RECT 201.115 -135.485 201.445 -135.155 ;
        RECT 201.115 -136.845 201.445 -136.515 ;
        RECT 201.115 -138.205 201.445 -137.875 ;
        RECT 201.115 -139.565 201.445 -139.235 ;
        RECT 201.115 -140.925 201.445 -140.595 ;
        RECT 201.115 -142.285 201.445 -141.955 ;
        RECT 201.115 -143.645 201.445 -143.315 ;
        RECT 201.115 -145.005 201.445 -144.675 ;
        RECT 201.115 -146.365 201.445 -146.035 ;
        RECT 201.115 -147.725 201.445 -147.395 ;
        RECT 201.115 -149.085 201.445 -148.755 ;
        RECT 201.115 -150.445 201.445 -150.115 ;
        RECT 201.115 -151.805 201.445 -151.475 ;
        RECT 201.115 -153.165 201.445 -152.835 ;
        RECT 201.115 -154.525 201.445 -154.195 ;
        RECT 201.115 -155.885 201.445 -155.555 ;
        RECT 201.115 -157.245 201.445 -156.915 ;
        RECT 201.115 -158.605 201.445 -158.275 ;
        RECT 201.115 -159.965 201.445 -159.635 ;
        RECT 201.115 -161.325 201.445 -160.995 ;
        RECT 201.115 -162.685 201.445 -162.355 ;
        RECT 201.115 -164.045 201.445 -163.715 ;
        RECT 201.115 -165.405 201.445 -165.075 ;
        RECT 201.115 -166.765 201.445 -166.435 ;
        RECT 201.115 -168.125 201.445 -167.795 ;
        RECT 201.115 -169.485 201.445 -169.155 ;
        RECT 201.115 -170.845 201.445 -170.515 ;
        RECT 201.115 -172.205 201.445 -171.875 ;
        RECT 201.115 -173.565 201.445 -173.235 ;
        RECT 201.115 -174.925 201.445 -174.595 ;
        RECT 201.115 -176.285 201.445 -175.955 ;
        RECT 201.115 -177.645 201.445 -177.315 ;
        RECT 201.115 -179.005 201.445 -178.675 ;
        RECT 201.115 -184.65 201.445 -183.52 ;
        RECT 201.12 -184.765 201.44 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.475 244.04 202.805 245.17 ;
        RECT 202.475 239.875 202.805 240.205 ;
        RECT 202.475 238.515 202.805 238.845 ;
        RECT 202.475 237.155 202.805 237.485 ;
        RECT 202.48 237.155 202.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 202.475 -0.845 202.805 -0.515 ;
        RECT 202.475 -2.205 202.805 -1.875 ;
        RECT 202.475 -3.565 202.805 -3.235 ;
        RECT 202.48 -3.565 202.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 244.04 204.165 245.17 ;
        RECT 203.835 239.875 204.165 240.205 ;
        RECT 203.835 238.515 204.165 238.845 ;
        RECT 203.835 237.155 204.165 237.485 ;
        RECT 203.84 237.155 204.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 -0.845 204.165 -0.515 ;
        RECT 203.835 -2.205 204.165 -1.875 ;
        RECT 203.835 -3.565 204.165 -3.235 ;
        RECT 203.84 -3.565 204.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.835 -96.045 204.165 -95.715 ;
        RECT 203.835 -97.405 204.165 -97.075 ;
        RECT 203.835 -98.765 204.165 -98.435 ;
        RECT 203.835 -100.125 204.165 -99.795 ;
        RECT 203.835 -101.485 204.165 -101.155 ;
        RECT 203.835 -102.845 204.165 -102.515 ;
        RECT 203.835 -104.205 204.165 -103.875 ;
        RECT 203.835 -105.565 204.165 -105.235 ;
        RECT 203.835 -106.925 204.165 -106.595 ;
        RECT 203.835 -108.285 204.165 -107.955 ;
        RECT 203.835 -109.645 204.165 -109.315 ;
        RECT 203.835 -111.005 204.165 -110.675 ;
        RECT 203.835 -112.365 204.165 -112.035 ;
        RECT 203.835 -113.725 204.165 -113.395 ;
        RECT 203.835 -115.085 204.165 -114.755 ;
        RECT 203.835 -116.445 204.165 -116.115 ;
        RECT 203.835 -117.805 204.165 -117.475 ;
        RECT 203.835 -119.165 204.165 -118.835 ;
        RECT 203.835 -120.525 204.165 -120.195 ;
        RECT 203.835 -121.885 204.165 -121.555 ;
        RECT 203.835 -123.245 204.165 -122.915 ;
        RECT 203.835 -124.605 204.165 -124.275 ;
        RECT 203.835 -125.965 204.165 -125.635 ;
        RECT 203.835 -127.325 204.165 -126.995 ;
        RECT 203.835 -128.685 204.165 -128.355 ;
        RECT 203.835 -130.045 204.165 -129.715 ;
        RECT 203.835 -131.405 204.165 -131.075 ;
        RECT 203.835 -132.765 204.165 -132.435 ;
        RECT 203.835 -134.125 204.165 -133.795 ;
        RECT 203.835 -135.485 204.165 -135.155 ;
        RECT 203.835 -136.845 204.165 -136.515 ;
        RECT 203.835 -138.205 204.165 -137.875 ;
        RECT 203.835 -139.565 204.165 -139.235 ;
        RECT 203.835 -140.925 204.165 -140.595 ;
        RECT 203.835 -142.285 204.165 -141.955 ;
        RECT 203.835 -143.645 204.165 -143.315 ;
        RECT 203.835 -145.005 204.165 -144.675 ;
        RECT 203.835 -146.365 204.165 -146.035 ;
        RECT 203.835 -147.725 204.165 -147.395 ;
        RECT 203.835 -149.085 204.165 -148.755 ;
        RECT 203.835 -150.445 204.165 -150.115 ;
        RECT 203.835 -151.805 204.165 -151.475 ;
        RECT 203.835 -153.165 204.165 -152.835 ;
        RECT 203.835 -154.525 204.165 -154.195 ;
        RECT 203.835 -155.885 204.165 -155.555 ;
        RECT 203.835 -157.245 204.165 -156.915 ;
        RECT 203.835 -158.605 204.165 -158.275 ;
        RECT 203.835 -159.965 204.165 -159.635 ;
        RECT 203.835 -161.325 204.165 -160.995 ;
        RECT 203.835 -162.685 204.165 -162.355 ;
        RECT 203.835 -164.045 204.165 -163.715 ;
        RECT 203.835 -165.405 204.165 -165.075 ;
        RECT 203.835 -166.765 204.165 -166.435 ;
        RECT 203.835 -168.125 204.165 -167.795 ;
        RECT 203.835 -169.485 204.165 -169.155 ;
        RECT 203.835 -170.845 204.165 -170.515 ;
        RECT 203.835 -172.205 204.165 -171.875 ;
        RECT 203.835 -173.565 204.165 -173.235 ;
        RECT 203.835 -174.925 204.165 -174.595 ;
        RECT 203.835 -176.285 204.165 -175.955 ;
        RECT 203.835 -177.645 204.165 -177.315 ;
        RECT 203.835 -179.005 204.165 -178.675 ;
        RECT 203.835 -184.65 204.165 -183.52 ;
        RECT 203.84 -184.765 204.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.195 244.04 205.525 245.17 ;
        RECT 205.195 239.875 205.525 240.205 ;
        RECT 205.195 238.515 205.525 238.845 ;
        RECT 205.195 237.155 205.525 237.485 ;
        RECT 205.2 237.155 205.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.195 -0.845 205.525 -0.515 ;
        RECT 205.195 -2.205 205.525 -1.875 ;
        RECT 205.195 -3.565 205.525 -3.235 ;
        RECT 205.2 -3.565 205.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.195 -96.045 205.525 -95.715 ;
        RECT 205.195 -97.405 205.525 -97.075 ;
        RECT 205.195 -98.765 205.525 -98.435 ;
        RECT 205.195 -100.125 205.525 -99.795 ;
        RECT 205.195 -101.485 205.525 -101.155 ;
        RECT 205.195 -102.845 205.525 -102.515 ;
        RECT 205.195 -104.205 205.525 -103.875 ;
        RECT 205.195 -105.565 205.525 -105.235 ;
        RECT 205.195 -106.925 205.525 -106.595 ;
        RECT 205.195 -108.285 205.525 -107.955 ;
        RECT 205.195 -109.645 205.525 -109.315 ;
        RECT 205.195 -111.005 205.525 -110.675 ;
        RECT 205.195 -112.365 205.525 -112.035 ;
        RECT 205.195 -113.725 205.525 -113.395 ;
        RECT 205.195 -115.085 205.525 -114.755 ;
        RECT 205.195 -116.445 205.525 -116.115 ;
        RECT 205.195 -117.805 205.525 -117.475 ;
        RECT 205.195 -119.165 205.525 -118.835 ;
        RECT 205.195 -120.525 205.525 -120.195 ;
        RECT 205.195 -121.885 205.525 -121.555 ;
        RECT 205.195 -123.245 205.525 -122.915 ;
        RECT 205.195 -124.605 205.525 -124.275 ;
        RECT 205.195 -125.965 205.525 -125.635 ;
        RECT 205.195 -127.325 205.525 -126.995 ;
        RECT 205.195 -128.685 205.525 -128.355 ;
        RECT 205.195 -130.045 205.525 -129.715 ;
        RECT 205.195 -131.405 205.525 -131.075 ;
        RECT 205.195 -132.765 205.525 -132.435 ;
        RECT 205.195 -134.125 205.525 -133.795 ;
        RECT 205.195 -135.485 205.525 -135.155 ;
        RECT 205.195 -136.845 205.525 -136.515 ;
        RECT 205.195 -138.205 205.525 -137.875 ;
        RECT 205.195 -139.565 205.525 -139.235 ;
        RECT 205.195 -140.925 205.525 -140.595 ;
        RECT 205.195 -142.285 205.525 -141.955 ;
        RECT 205.195 -143.645 205.525 -143.315 ;
        RECT 205.195 -145.005 205.525 -144.675 ;
        RECT 205.195 -146.365 205.525 -146.035 ;
        RECT 205.195 -147.725 205.525 -147.395 ;
        RECT 205.195 -149.085 205.525 -148.755 ;
        RECT 205.195 -150.445 205.525 -150.115 ;
        RECT 205.195 -151.805 205.525 -151.475 ;
        RECT 205.195 -153.165 205.525 -152.835 ;
        RECT 205.195 -154.525 205.525 -154.195 ;
        RECT 205.195 -155.885 205.525 -155.555 ;
        RECT 205.195 -157.245 205.525 -156.915 ;
        RECT 205.195 -158.605 205.525 -158.275 ;
        RECT 205.195 -159.965 205.525 -159.635 ;
        RECT 205.195 -161.325 205.525 -160.995 ;
        RECT 205.195 -162.685 205.525 -162.355 ;
        RECT 205.195 -164.045 205.525 -163.715 ;
        RECT 205.195 -165.405 205.525 -165.075 ;
        RECT 205.195 -166.765 205.525 -166.435 ;
        RECT 205.195 -168.125 205.525 -167.795 ;
        RECT 205.195 -169.485 205.525 -169.155 ;
        RECT 205.195 -170.845 205.525 -170.515 ;
        RECT 205.195 -172.205 205.525 -171.875 ;
        RECT 205.195 -173.565 205.525 -173.235 ;
        RECT 205.195 -174.925 205.525 -174.595 ;
        RECT 205.195 -176.285 205.525 -175.955 ;
        RECT 205.195 -177.645 205.525 -177.315 ;
        RECT 205.195 -179.005 205.525 -178.675 ;
        RECT 205.195 -184.65 205.525 -183.52 ;
        RECT 205.2 -184.765 205.52 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.555 244.04 206.885 245.17 ;
        RECT 206.555 239.875 206.885 240.205 ;
        RECT 206.555 238.515 206.885 238.845 ;
        RECT 206.555 237.155 206.885 237.485 ;
        RECT 206.56 237.155 206.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.555 -0.845 206.885 -0.515 ;
        RECT 206.555 -2.205 206.885 -1.875 ;
        RECT 206.555 -3.565 206.885 -3.235 ;
        RECT 206.56 -3.565 206.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 206.555 -96.045 206.885 -95.715 ;
        RECT 206.555 -97.405 206.885 -97.075 ;
        RECT 206.555 -98.765 206.885 -98.435 ;
        RECT 206.555 -100.125 206.885 -99.795 ;
        RECT 206.555 -101.485 206.885 -101.155 ;
        RECT 206.555 -102.845 206.885 -102.515 ;
        RECT 206.555 -104.205 206.885 -103.875 ;
        RECT 206.555 -105.565 206.885 -105.235 ;
        RECT 206.555 -106.925 206.885 -106.595 ;
        RECT 206.555 -108.285 206.885 -107.955 ;
        RECT 206.555 -109.645 206.885 -109.315 ;
        RECT 206.555 -111.005 206.885 -110.675 ;
        RECT 206.555 -112.365 206.885 -112.035 ;
        RECT 206.555 -113.725 206.885 -113.395 ;
        RECT 206.555 -115.085 206.885 -114.755 ;
        RECT 206.555 -116.445 206.885 -116.115 ;
        RECT 206.555 -117.805 206.885 -117.475 ;
        RECT 206.555 -119.165 206.885 -118.835 ;
        RECT 206.555 -120.525 206.885 -120.195 ;
        RECT 206.555 -121.885 206.885 -121.555 ;
        RECT 206.555 -123.245 206.885 -122.915 ;
        RECT 206.555 -124.605 206.885 -124.275 ;
        RECT 206.555 -125.965 206.885 -125.635 ;
        RECT 206.555 -127.325 206.885 -126.995 ;
        RECT 206.555 -128.685 206.885 -128.355 ;
        RECT 206.555 -130.045 206.885 -129.715 ;
        RECT 206.555 -131.405 206.885 -131.075 ;
        RECT 206.555 -132.765 206.885 -132.435 ;
        RECT 206.555 -134.125 206.885 -133.795 ;
        RECT 206.555 -135.485 206.885 -135.155 ;
        RECT 206.555 -136.845 206.885 -136.515 ;
        RECT 206.555 -138.205 206.885 -137.875 ;
        RECT 206.555 -139.565 206.885 -139.235 ;
        RECT 206.555 -140.925 206.885 -140.595 ;
        RECT 206.555 -142.285 206.885 -141.955 ;
        RECT 206.555 -143.645 206.885 -143.315 ;
        RECT 206.555 -145.005 206.885 -144.675 ;
        RECT 206.555 -146.365 206.885 -146.035 ;
        RECT 206.555 -147.725 206.885 -147.395 ;
        RECT 206.555 -149.085 206.885 -148.755 ;
        RECT 206.555 -150.445 206.885 -150.115 ;
        RECT 206.555 -151.805 206.885 -151.475 ;
        RECT 206.555 -153.165 206.885 -152.835 ;
        RECT 206.555 -154.525 206.885 -154.195 ;
        RECT 206.555 -155.885 206.885 -155.555 ;
        RECT 206.555 -157.245 206.885 -156.915 ;
        RECT 206.555 -158.605 206.885 -158.275 ;
        RECT 206.555 -159.965 206.885 -159.635 ;
        RECT 206.555 -161.325 206.885 -160.995 ;
        RECT 206.555 -162.685 206.885 -162.355 ;
        RECT 206.555 -164.045 206.885 -163.715 ;
        RECT 206.555 -165.405 206.885 -165.075 ;
        RECT 206.555 -166.765 206.885 -166.435 ;
        RECT 206.555 -168.125 206.885 -167.795 ;
        RECT 206.555 -169.485 206.885 -169.155 ;
        RECT 206.555 -170.845 206.885 -170.515 ;
        RECT 206.555 -172.205 206.885 -171.875 ;
        RECT 206.555 -173.565 206.885 -173.235 ;
        RECT 206.555 -174.925 206.885 -174.595 ;
        RECT 206.555 -176.285 206.885 -175.955 ;
        RECT 206.555 -177.645 206.885 -177.315 ;
        RECT 206.555 -179.005 206.885 -178.675 ;
        RECT 206.555 -184.65 206.885 -183.52 ;
        RECT 206.56 -184.765 206.88 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 244.04 208.245 245.17 ;
        RECT 207.915 239.875 208.245 240.205 ;
        RECT 207.915 238.515 208.245 238.845 ;
        RECT 207.915 237.155 208.245 237.485 ;
        RECT 207.92 237.155 208.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 -0.845 208.245 -0.515 ;
        RECT 207.915 -2.205 208.245 -1.875 ;
        RECT 207.915 -3.565 208.245 -3.235 ;
        RECT 207.92 -3.565 208.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.915 -96.045 208.245 -95.715 ;
        RECT 207.915 -97.405 208.245 -97.075 ;
        RECT 207.915 -98.765 208.245 -98.435 ;
        RECT 207.915 -100.125 208.245 -99.795 ;
        RECT 207.915 -101.485 208.245 -101.155 ;
        RECT 207.915 -102.845 208.245 -102.515 ;
        RECT 207.915 -104.205 208.245 -103.875 ;
        RECT 207.915 -105.565 208.245 -105.235 ;
        RECT 207.915 -106.925 208.245 -106.595 ;
        RECT 207.915 -108.285 208.245 -107.955 ;
        RECT 207.915 -109.645 208.245 -109.315 ;
        RECT 207.915 -111.005 208.245 -110.675 ;
        RECT 207.915 -112.365 208.245 -112.035 ;
        RECT 207.915 -113.725 208.245 -113.395 ;
        RECT 207.915 -115.085 208.245 -114.755 ;
        RECT 207.915 -116.445 208.245 -116.115 ;
        RECT 207.915 -117.805 208.245 -117.475 ;
        RECT 207.915 -119.165 208.245 -118.835 ;
        RECT 207.915 -120.525 208.245 -120.195 ;
        RECT 207.915 -121.885 208.245 -121.555 ;
        RECT 207.915 -123.245 208.245 -122.915 ;
        RECT 207.915 -124.605 208.245 -124.275 ;
        RECT 207.915 -125.965 208.245 -125.635 ;
        RECT 207.915 -127.325 208.245 -126.995 ;
        RECT 207.915 -128.685 208.245 -128.355 ;
        RECT 207.915 -130.045 208.245 -129.715 ;
        RECT 207.915 -131.405 208.245 -131.075 ;
        RECT 207.915 -132.765 208.245 -132.435 ;
        RECT 207.915 -134.125 208.245 -133.795 ;
        RECT 207.915 -135.485 208.245 -135.155 ;
        RECT 207.915 -136.845 208.245 -136.515 ;
        RECT 207.915 -138.205 208.245 -137.875 ;
        RECT 207.915 -139.565 208.245 -139.235 ;
        RECT 207.915 -140.925 208.245 -140.595 ;
        RECT 207.915 -142.285 208.245 -141.955 ;
        RECT 207.915 -143.645 208.245 -143.315 ;
        RECT 207.915 -145.005 208.245 -144.675 ;
        RECT 207.915 -146.365 208.245 -146.035 ;
        RECT 207.915 -147.725 208.245 -147.395 ;
        RECT 207.915 -149.085 208.245 -148.755 ;
        RECT 207.915 -150.445 208.245 -150.115 ;
        RECT 207.915 -151.805 208.245 -151.475 ;
        RECT 207.915 -153.165 208.245 -152.835 ;
        RECT 207.915 -154.525 208.245 -154.195 ;
        RECT 207.915 -155.885 208.245 -155.555 ;
        RECT 207.915 -157.245 208.245 -156.915 ;
        RECT 207.915 -158.605 208.245 -158.275 ;
        RECT 207.915 -159.965 208.245 -159.635 ;
        RECT 207.915 -161.325 208.245 -160.995 ;
        RECT 207.915 -162.685 208.245 -162.355 ;
        RECT 207.915 -164.045 208.245 -163.715 ;
        RECT 207.915 -165.405 208.245 -165.075 ;
        RECT 207.915 -166.765 208.245 -166.435 ;
        RECT 207.915 -168.125 208.245 -167.795 ;
        RECT 207.915 -169.485 208.245 -169.155 ;
        RECT 207.915 -170.845 208.245 -170.515 ;
        RECT 207.915 -172.205 208.245 -171.875 ;
        RECT 207.915 -173.565 208.245 -173.235 ;
        RECT 207.915 -174.925 208.245 -174.595 ;
        RECT 207.915 -176.285 208.245 -175.955 ;
        RECT 207.915 -177.645 208.245 -177.315 ;
        RECT 207.915 -179.005 208.245 -178.675 ;
        RECT 207.915 -184.65 208.245 -183.52 ;
        RECT 207.92 -184.765 208.24 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.275 244.04 209.605 245.17 ;
        RECT 209.275 239.875 209.605 240.205 ;
        RECT 209.275 238.515 209.605 238.845 ;
        RECT 209.275 237.155 209.605 237.485 ;
        RECT 209.28 237.155 209.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.275 -98.765 209.605 -98.435 ;
        RECT 209.275 -100.125 209.605 -99.795 ;
        RECT 209.275 -101.485 209.605 -101.155 ;
        RECT 209.275 -102.845 209.605 -102.515 ;
        RECT 209.275 -104.205 209.605 -103.875 ;
        RECT 209.275 -105.565 209.605 -105.235 ;
        RECT 209.275 -106.925 209.605 -106.595 ;
        RECT 209.275 -108.285 209.605 -107.955 ;
        RECT 209.275 -109.645 209.605 -109.315 ;
        RECT 209.275 -111.005 209.605 -110.675 ;
        RECT 209.275 -112.365 209.605 -112.035 ;
        RECT 209.275 -113.725 209.605 -113.395 ;
        RECT 209.275 -115.085 209.605 -114.755 ;
        RECT 209.275 -116.445 209.605 -116.115 ;
        RECT 209.275 -117.805 209.605 -117.475 ;
        RECT 209.275 -119.165 209.605 -118.835 ;
        RECT 209.275 -120.525 209.605 -120.195 ;
        RECT 209.275 -121.885 209.605 -121.555 ;
        RECT 209.275 -123.245 209.605 -122.915 ;
        RECT 209.275 -124.605 209.605 -124.275 ;
        RECT 209.275 -125.965 209.605 -125.635 ;
        RECT 209.275 -127.325 209.605 -126.995 ;
        RECT 209.275 -128.685 209.605 -128.355 ;
        RECT 209.275 -130.045 209.605 -129.715 ;
        RECT 209.275 -131.405 209.605 -131.075 ;
        RECT 209.275 -132.765 209.605 -132.435 ;
        RECT 209.275 -134.125 209.605 -133.795 ;
        RECT 209.275 -135.485 209.605 -135.155 ;
        RECT 209.275 -136.845 209.605 -136.515 ;
        RECT 209.275 -138.205 209.605 -137.875 ;
        RECT 209.275 -139.565 209.605 -139.235 ;
        RECT 209.275 -140.925 209.605 -140.595 ;
        RECT 209.275 -142.285 209.605 -141.955 ;
        RECT 209.275 -143.645 209.605 -143.315 ;
        RECT 209.275 -145.005 209.605 -144.675 ;
        RECT 209.275 -146.365 209.605 -146.035 ;
        RECT 209.275 -147.725 209.605 -147.395 ;
        RECT 209.275 -149.085 209.605 -148.755 ;
        RECT 209.275 -150.445 209.605 -150.115 ;
        RECT 209.275 -151.805 209.605 -151.475 ;
        RECT 209.275 -153.165 209.605 -152.835 ;
        RECT 209.275 -154.525 209.605 -154.195 ;
        RECT 209.275 -155.885 209.605 -155.555 ;
        RECT 209.275 -157.245 209.605 -156.915 ;
        RECT 209.275 -158.605 209.605 -158.275 ;
        RECT 209.275 -159.965 209.605 -159.635 ;
        RECT 209.275 -161.325 209.605 -160.995 ;
        RECT 209.275 -162.685 209.605 -162.355 ;
        RECT 209.275 -164.045 209.605 -163.715 ;
        RECT 209.275 -165.405 209.605 -165.075 ;
        RECT 209.275 -166.765 209.605 -166.435 ;
        RECT 209.275 -168.125 209.605 -167.795 ;
        RECT 209.275 -169.485 209.605 -169.155 ;
        RECT 209.275 -170.845 209.605 -170.515 ;
        RECT 209.275 -172.205 209.605 -171.875 ;
        RECT 209.275 -173.565 209.605 -173.235 ;
        RECT 209.275 -174.925 209.605 -174.595 ;
        RECT 209.275 -176.285 209.605 -175.955 ;
        RECT 209.275 -177.645 209.605 -177.315 ;
        RECT 209.275 -179.005 209.605 -178.675 ;
        RECT 209.275 -184.65 209.605 -183.52 ;
        RECT 209.28 -184.765 209.6 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.76 -98.075 210.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 244.04 160.645 245.17 ;
        RECT 160.315 239.875 160.645 240.205 ;
        RECT 160.315 238.515 160.645 238.845 ;
        RECT 160.315 237.155 160.645 237.485 ;
        RECT 160.32 237.155 160.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 -0.845 160.645 -0.515 ;
        RECT 160.315 -2.205 160.645 -1.875 ;
        RECT 160.315 -3.565 160.645 -3.235 ;
        RECT 160.32 -3.565 160.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.315 -96.045 160.645 -95.715 ;
        RECT 160.315 -97.405 160.645 -97.075 ;
        RECT 160.315 -98.765 160.645 -98.435 ;
        RECT 160.315 -100.125 160.645 -99.795 ;
        RECT 160.315 -101.485 160.645 -101.155 ;
        RECT 160.315 -102.845 160.645 -102.515 ;
        RECT 160.315 -104.205 160.645 -103.875 ;
        RECT 160.315 -105.565 160.645 -105.235 ;
        RECT 160.315 -106.925 160.645 -106.595 ;
        RECT 160.315 -108.285 160.645 -107.955 ;
        RECT 160.315 -109.645 160.645 -109.315 ;
        RECT 160.315 -111.005 160.645 -110.675 ;
        RECT 160.315 -112.365 160.645 -112.035 ;
        RECT 160.315 -113.725 160.645 -113.395 ;
        RECT 160.315 -115.085 160.645 -114.755 ;
        RECT 160.315 -116.445 160.645 -116.115 ;
        RECT 160.315 -117.805 160.645 -117.475 ;
        RECT 160.315 -119.165 160.645 -118.835 ;
        RECT 160.315 -120.525 160.645 -120.195 ;
        RECT 160.315 -121.885 160.645 -121.555 ;
        RECT 160.315 -123.245 160.645 -122.915 ;
        RECT 160.315 -124.605 160.645 -124.275 ;
        RECT 160.315 -125.965 160.645 -125.635 ;
        RECT 160.315 -127.325 160.645 -126.995 ;
        RECT 160.315 -128.685 160.645 -128.355 ;
        RECT 160.315 -130.045 160.645 -129.715 ;
        RECT 160.315 -131.405 160.645 -131.075 ;
        RECT 160.315 -132.765 160.645 -132.435 ;
        RECT 160.315 -134.125 160.645 -133.795 ;
        RECT 160.315 -135.485 160.645 -135.155 ;
        RECT 160.315 -136.845 160.645 -136.515 ;
        RECT 160.315 -138.205 160.645 -137.875 ;
        RECT 160.315 -139.565 160.645 -139.235 ;
        RECT 160.315 -140.925 160.645 -140.595 ;
        RECT 160.315 -142.285 160.645 -141.955 ;
        RECT 160.315 -143.645 160.645 -143.315 ;
        RECT 160.315 -145.005 160.645 -144.675 ;
        RECT 160.315 -146.365 160.645 -146.035 ;
        RECT 160.315 -147.725 160.645 -147.395 ;
        RECT 160.315 -149.085 160.645 -148.755 ;
        RECT 160.315 -150.445 160.645 -150.115 ;
        RECT 160.315 -151.805 160.645 -151.475 ;
        RECT 160.315 -153.165 160.645 -152.835 ;
        RECT 160.315 -154.525 160.645 -154.195 ;
        RECT 160.315 -155.885 160.645 -155.555 ;
        RECT 160.315 -157.245 160.645 -156.915 ;
        RECT 160.315 -158.605 160.645 -158.275 ;
        RECT 160.315 -159.965 160.645 -159.635 ;
        RECT 160.315 -161.325 160.645 -160.995 ;
        RECT 160.315 -162.685 160.645 -162.355 ;
        RECT 160.315 -164.045 160.645 -163.715 ;
        RECT 160.315 -165.405 160.645 -165.075 ;
        RECT 160.315 -166.765 160.645 -166.435 ;
        RECT 160.315 -168.125 160.645 -167.795 ;
        RECT 160.315 -169.485 160.645 -169.155 ;
        RECT 160.315 -170.845 160.645 -170.515 ;
        RECT 160.315 -172.205 160.645 -171.875 ;
        RECT 160.315 -173.565 160.645 -173.235 ;
        RECT 160.315 -174.925 160.645 -174.595 ;
        RECT 160.315 -176.285 160.645 -175.955 ;
        RECT 160.315 -177.645 160.645 -177.315 ;
        RECT 160.315 -179.005 160.645 -178.675 ;
        RECT 160.315 -184.65 160.645 -183.52 ;
        RECT 160.32 -184.765 160.64 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 244.04 162.005 245.17 ;
        RECT 161.675 239.875 162.005 240.205 ;
        RECT 161.675 238.515 162.005 238.845 ;
        RECT 161.675 237.155 162.005 237.485 ;
        RECT 161.68 237.155 162 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 -0.845 162.005 -0.515 ;
        RECT 161.675 -2.205 162.005 -1.875 ;
        RECT 161.675 -3.565 162.005 -3.235 ;
        RECT 161.68 -3.565 162 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 161.675 -96.045 162.005 -95.715 ;
        RECT 161.675 -97.405 162.005 -97.075 ;
        RECT 161.675 -98.765 162.005 -98.435 ;
        RECT 161.675 -100.125 162.005 -99.795 ;
        RECT 161.675 -101.485 162.005 -101.155 ;
        RECT 161.675 -102.845 162.005 -102.515 ;
        RECT 161.675 -104.205 162.005 -103.875 ;
        RECT 161.675 -105.565 162.005 -105.235 ;
        RECT 161.675 -106.925 162.005 -106.595 ;
        RECT 161.675 -108.285 162.005 -107.955 ;
        RECT 161.675 -109.645 162.005 -109.315 ;
        RECT 161.675 -111.005 162.005 -110.675 ;
        RECT 161.675 -112.365 162.005 -112.035 ;
        RECT 161.675 -113.725 162.005 -113.395 ;
        RECT 161.675 -115.085 162.005 -114.755 ;
        RECT 161.675 -116.445 162.005 -116.115 ;
        RECT 161.675 -117.805 162.005 -117.475 ;
        RECT 161.675 -119.165 162.005 -118.835 ;
        RECT 161.675 -120.525 162.005 -120.195 ;
        RECT 161.675 -121.885 162.005 -121.555 ;
        RECT 161.675 -123.245 162.005 -122.915 ;
        RECT 161.675 -124.605 162.005 -124.275 ;
        RECT 161.675 -125.965 162.005 -125.635 ;
        RECT 161.675 -127.325 162.005 -126.995 ;
        RECT 161.675 -128.685 162.005 -128.355 ;
        RECT 161.675 -130.045 162.005 -129.715 ;
        RECT 161.675 -131.405 162.005 -131.075 ;
        RECT 161.675 -132.765 162.005 -132.435 ;
        RECT 161.675 -134.125 162.005 -133.795 ;
        RECT 161.675 -135.485 162.005 -135.155 ;
        RECT 161.675 -136.845 162.005 -136.515 ;
        RECT 161.675 -138.205 162.005 -137.875 ;
        RECT 161.675 -139.565 162.005 -139.235 ;
        RECT 161.675 -140.925 162.005 -140.595 ;
        RECT 161.675 -142.285 162.005 -141.955 ;
        RECT 161.675 -143.645 162.005 -143.315 ;
        RECT 161.675 -145.005 162.005 -144.675 ;
        RECT 161.675 -146.365 162.005 -146.035 ;
        RECT 161.675 -147.725 162.005 -147.395 ;
        RECT 161.675 -149.085 162.005 -148.755 ;
        RECT 161.675 -150.445 162.005 -150.115 ;
        RECT 161.675 -151.805 162.005 -151.475 ;
        RECT 161.675 -153.165 162.005 -152.835 ;
        RECT 161.675 -154.525 162.005 -154.195 ;
        RECT 161.675 -155.885 162.005 -155.555 ;
        RECT 161.675 -157.245 162.005 -156.915 ;
        RECT 161.675 -158.605 162.005 -158.275 ;
        RECT 161.675 -159.965 162.005 -159.635 ;
        RECT 161.675 -161.325 162.005 -160.995 ;
        RECT 161.675 -162.685 162.005 -162.355 ;
        RECT 161.675 -164.045 162.005 -163.715 ;
        RECT 161.675 -165.405 162.005 -165.075 ;
        RECT 161.675 -166.765 162.005 -166.435 ;
        RECT 161.675 -168.125 162.005 -167.795 ;
        RECT 161.675 -169.485 162.005 -169.155 ;
        RECT 161.675 -170.845 162.005 -170.515 ;
        RECT 161.675 -172.205 162.005 -171.875 ;
        RECT 161.675 -173.565 162.005 -173.235 ;
        RECT 161.675 -174.925 162.005 -174.595 ;
        RECT 161.675 -176.285 162.005 -175.955 ;
        RECT 161.675 -177.645 162.005 -177.315 ;
        RECT 161.675 -179.005 162.005 -178.675 ;
        RECT 161.675 -184.65 162.005 -183.52 ;
        RECT 161.68 -184.765 162 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 244.04 163.365 245.17 ;
        RECT 163.035 239.875 163.365 240.205 ;
        RECT 163.035 238.515 163.365 238.845 ;
        RECT 163.035 237.155 163.365 237.485 ;
        RECT 163.04 237.155 163.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 -0.845 163.365 -0.515 ;
        RECT 163.035 -2.205 163.365 -1.875 ;
        RECT 163.035 -3.565 163.365 -3.235 ;
        RECT 163.04 -3.565 163.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.035 -96.045 163.365 -95.715 ;
        RECT 163.035 -97.405 163.365 -97.075 ;
        RECT 163.035 -98.765 163.365 -98.435 ;
        RECT 163.035 -100.125 163.365 -99.795 ;
        RECT 163.035 -101.485 163.365 -101.155 ;
        RECT 163.035 -102.845 163.365 -102.515 ;
        RECT 163.035 -104.205 163.365 -103.875 ;
        RECT 163.035 -105.565 163.365 -105.235 ;
        RECT 163.035 -106.925 163.365 -106.595 ;
        RECT 163.035 -108.285 163.365 -107.955 ;
        RECT 163.035 -109.645 163.365 -109.315 ;
        RECT 163.035 -111.005 163.365 -110.675 ;
        RECT 163.035 -112.365 163.365 -112.035 ;
        RECT 163.035 -113.725 163.365 -113.395 ;
        RECT 163.035 -115.085 163.365 -114.755 ;
        RECT 163.035 -116.445 163.365 -116.115 ;
        RECT 163.035 -117.805 163.365 -117.475 ;
        RECT 163.035 -119.165 163.365 -118.835 ;
        RECT 163.035 -120.525 163.365 -120.195 ;
        RECT 163.035 -121.885 163.365 -121.555 ;
        RECT 163.035 -123.245 163.365 -122.915 ;
        RECT 163.035 -124.605 163.365 -124.275 ;
        RECT 163.035 -125.965 163.365 -125.635 ;
        RECT 163.035 -127.325 163.365 -126.995 ;
        RECT 163.035 -128.685 163.365 -128.355 ;
        RECT 163.035 -130.045 163.365 -129.715 ;
        RECT 163.035 -131.405 163.365 -131.075 ;
        RECT 163.035 -132.765 163.365 -132.435 ;
        RECT 163.035 -134.125 163.365 -133.795 ;
        RECT 163.035 -135.485 163.365 -135.155 ;
        RECT 163.035 -136.845 163.365 -136.515 ;
        RECT 163.035 -138.205 163.365 -137.875 ;
        RECT 163.035 -139.565 163.365 -139.235 ;
        RECT 163.035 -140.925 163.365 -140.595 ;
        RECT 163.035 -142.285 163.365 -141.955 ;
        RECT 163.035 -143.645 163.365 -143.315 ;
        RECT 163.035 -145.005 163.365 -144.675 ;
        RECT 163.035 -146.365 163.365 -146.035 ;
        RECT 163.035 -147.725 163.365 -147.395 ;
        RECT 163.035 -149.085 163.365 -148.755 ;
        RECT 163.035 -150.445 163.365 -150.115 ;
        RECT 163.035 -151.805 163.365 -151.475 ;
        RECT 163.035 -153.165 163.365 -152.835 ;
        RECT 163.035 -154.525 163.365 -154.195 ;
        RECT 163.035 -155.885 163.365 -155.555 ;
        RECT 163.035 -157.245 163.365 -156.915 ;
        RECT 163.035 -158.605 163.365 -158.275 ;
        RECT 163.035 -159.965 163.365 -159.635 ;
        RECT 163.035 -161.325 163.365 -160.995 ;
        RECT 163.035 -162.685 163.365 -162.355 ;
        RECT 163.035 -164.045 163.365 -163.715 ;
        RECT 163.035 -165.405 163.365 -165.075 ;
        RECT 163.035 -166.765 163.365 -166.435 ;
        RECT 163.035 -168.125 163.365 -167.795 ;
        RECT 163.035 -169.485 163.365 -169.155 ;
        RECT 163.035 -170.845 163.365 -170.515 ;
        RECT 163.035 -172.205 163.365 -171.875 ;
        RECT 163.035 -173.565 163.365 -173.235 ;
        RECT 163.035 -174.925 163.365 -174.595 ;
        RECT 163.035 -176.285 163.365 -175.955 ;
        RECT 163.035 -177.645 163.365 -177.315 ;
        RECT 163.035 -179.005 163.365 -178.675 ;
        RECT 163.035 -184.65 163.365 -183.52 ;
        RECT 163.04 -184.765 163.36 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 244.04 164.725 245.17 ;
        RECT 164.395 239.875 164.725 240.205 ;
        RECT 164.395 238.515 164.725 238.845 ;
        RECT 164.395 237.155 164.725 237.485 ;
        RECT 164.4 237.155 164.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 -0.845 164.725 -0.515 ;
        RECT 164.395 -2.205 164.725 -1.875 ;
        RECT 164.395 -3.565 164.725 -3.235 ;
        RECT 164.4 -3.565 164.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 164.395 -96.045 164.725 -95.715 ;
        RECT 164.395 -97.405 164.725 -97.075 ;
        RECT 164.395 -98.765 164.725 -98.435 ;
        RECT 164.395 -100.125 164.725 -99.795 ;
        RECT 164.395 -101.485 164.725 -101.155 ;
        RECT 164.395 -102.845 164.725 -102.515 ;
        RECT 164.395 -104.205 164.725 -103.875 ;
        RECT 164.395 -105.565 164.725 -105.235 ;
        RECT 164.395 -106.925 164.725 -106.595 ;
        RECT 164.395 -108.285 164.725 -107.955 ;
        RECT 164.395 -109.645 164.725 -109.315 ;
        RECT 164.395 -111.005 164.725 -110.675 ;
        RECT 164.395 -112.365 164.725 -112.035 ;
        RECT 164.395 -113.725 164.725 -113.395 ;
        RECT 164.395 -115.085 164.725 -114.755 ;
        RECT 164.395 -116.445 164.725 -116.115 ;
        RECT 164.395 -117.805 164.725 -117.475 ;
        RECT 164.395 -119.165 164.725 -118.835 ;
        RECT 164.395 -120.525 164.725 -120.195 ;
        RECT 164.395 -121.885 164.725 -121.555 ;
        RECT 164.395 -123.245 164.725 -122.915 ;
        RECT 164.395 -124.605 164.725 -124.275 ;
        RECT 164.395 -125.965 164.725 -125.635 ;
        RECT 164.395 -127.325 164.725 -126.995 ;
        RECT 164.395 -128.685 164.725 -128.355 ;
        RECT 164.395 -130.045 164.725 -129.715 ;
        RECT 164.395 -131.405 164.725 -131.075 ;
        RECT 164.395 -132.765 164.725 -132.435 ;
        RECT 164.395 -134.125 164.725 -133.795 ;
        RECT 164.395 -135.485 164.725 -135.155 ;
        RECT 164.395 -136.845 164.725 -136.515 ;
        RECT 164.395 -138.205 164.725 -137.875 ;
        RECT 164.395 -139.565 164.725 -139.235 ;
        RECT 164.395 -140.925 164.725 -140.595 ;
        RECT 164.395 -142.285 164.725 -141.955 ;
        RECT 164.395 -143.645 164.725 -143.315 ;
        RECT 164.395 -145.005 164.725 -144.675 ;
        RECT 164.395 -146.365 164.725 -146.035 ;
        RECT 164.395 -147.725 164.725 -147.395 ;
        RECT 164.395 -149.085 164.725 -148.755 ;
        RECT 164.395 -150.445 164.725 -150.115 ;
        RECT 164.395 -151.805 164.725 -151.475 ;
        RECT 164.395 -153.165 164.725 -152.835 ;
        RECT 164.395 -154.525 164.725 -154.195 ;
        RECT 164.395 -155.885 164.725 -155.555 ;
        RECT 164.395 -157.245 164.725 -156.915 ;
        RECT 164.395 -158.605 164.725 -158.275 ;
        RECT 164.395 -159.965 164.725 -159.635 ;
        RECT 164.395 -161.325 164.725 -160.995 ;
        RECT 164.395 -162.685 164.725 -162.355 ;
        RECT 164.395 -164.045 164.725 -163.715 ;
        RECT 164.395 -165.405 164.725 -165.075 ;
        RECT 164.395 -166.765 164.725 -166.435 ;
        RECT 164.395 -168.125 164.725 -167.795 ;
        RECT 164.395 -169.485 164.725 -169.155 ;
        RECT 164.395 -170.845 164.725 -170.515 ;
        RECT 164.395 -172.205 164.725 -171.875 ;
        RECT 164.395 -173.565 164.725 -173.235 ;
        RECT 164.395 -174.925 164.725 -174.595 ;
        RECT 164.395 -176.285 164.725 -175.955 ;
        RECT 164.395 -177.645 164.725 -177.315 ;
        RECT 164.395 -179.005 164.725 -178.675 ;
        RECT 164.395 -184.65 164.725 -183.52 ;
        RECT 164.4 -184.765 164.72 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 244.04 166.085 245.17 ;
        RECT 165.755 239.875 166.085 240.205 ;
        RECT 165.755 238.515 166.085 238.845 ;
        RECT 165.755 237.155 166.085 237.485 ;
        RECT 165.76 237.155 166.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.755 -98.765 166.085 -98.435 ;
        RECT 165.755 -100.125 166.085 -99.795 ;
        RECT 165.755 -101.485 166.085 -101.155 ;
        RECT 165.755 -102.845 166.085 -102.515 ;
        RECT 165.755 -104.205 166.085 -103.875 ;
        RECT 165.755 -105.565 166.085 -105.235 ;
        RECT 165.755 -106.925 166.085 -106.595 ;
        RECT 165.755 -108.285 166.085 -107.955 ;
        RECT 165.755 -109.645 166.085 -109.315 ;
        RECT 165.755 -111.005 166.085 -110.675 ;
        RECT 165.755 -112.365 166.085 -112.035 ;
        RECT 165.755 -113.725 166.085 -113.395 ;
        RECT 165.755 -115.085 166.085 -114.755 ;
        RECT 165.755 -116.445 166.085 -116.115 ;
        RECT 165.755 -117.805 166.085 -117.475 ;
        RECT 165.755 -119.165 166.085 -118.835 ;
        RECT 165.755 -120.525 166.085 -120.195 ;
        RECT 165.755 -121.885 166.085 -121.555 ;
        RECT 165.755 -123.245 166.085 -122.915 ;
        RECT 165.755 -124.605 166.085 -124.275 ;
        RECT 165.755 -125.965 166.085 -125.635 ;
        RECT 165.755 -127.325 166.085 -126.995 ;
        RECT 165.755 -128.685 166.085 -128.355 ;
        RECT 165.755 -130.045 166.085 -129.715 ;
        RECT 165.755 -131.405 166.085 -131.075 ;
        RECT 165.755 -132.765 166.085 -132.435 ;
        RECT 165.755 -134.125 166.085 -133.795 ;
        RECT 165.755 -135.485 166.085 -135.155 ;
        RECT 165.755 -136.845 166.085 -136.515 ;
        RECT 165.755 -138.205 166.085 -137.875 ;
        RECT 165.755 -139.565 166.085 -139.235 ;
        RECT 165.755 -140.925 166.085 -140.595 ;
        RECT 165.755 -142.285 166.085 -141.955 ;
        RECT 165.755 -143.645 166.085 -143.315 ;
        RECT 165.755 -145.005 166.085 -144.675 ;
        RECT 165.755 -146.365 166.085 -146.035 ;
        RECT 165.755 -147.725 166.085 -147.395 ;
        RECT 165.755 -149.085 166.085 -148.755 ;
        RECT 165.755 -150.445 166.085 -150.115 ;
        RECT 165.755 -151.805 166.085 -151.475 ;
        RECT 165.755 -153.165 166.085 -152.835 ;
        RECT 165.755 -154.525 166.085 -154.195 ;
        RECT 165.755 -155.885 166.085 -155.555 ;
        RECT 165.755 -157.245 166.085 -156.915 ;
        RECT 165.755 -158.605 166.085 -158.275 ;
        RECT 165.755 -159.965 166.085 -159.635 ;
        RECT 165.755 -161.325 166.085 -160.995 ;
        RECT 165.755 -162.685 166.085 -162.355 ;
        RECT 165.755 -164.045 166.085 -163.715 ;
        RECT 165.755 -165.405 166.085 -165.075 ;
        RECT 165.755 -166.765 166.085 -166.435 ;
        RECT 165.755 -168.125 166.085 -167.795 ;
        RECT 165.755 -169.485 166.085 -169.155 ;
        RECT 165.755 -170.845 166.085 -170.515 ;
        RECT 165.755 -172.205 166.085 -171.875 ;
        RECT 165.755 -173.565 166.085 -173.235 ;
        RECT 165.755 -174.925 166.085 -174.595 ;
        RECT 165.755 -176.285 166.085 -175.955 ;
        RECT 165.755 -177.645 166.085 -177.315 ;
        RECT 165.755 -179.005 166.085 -178.675 ;
        RECT 165.755 -184.65 166.085 -183.52 ;
        RECT 165.76 -184.765 166.08 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.16 -98.075 166.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.115 244.04 167.445 245.17 ;
        RECT 167.115 239.875 167.445 240.205 ;
        RECT 167.115 238.515 167.445 238.845 ;
        RECT 167.115 237.155 167.445 237.485 ;
        RECT 167.12 237.155 167.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.475 244.04 168.805 245.17 ;
        RECT 168.475 239.875 168.805 240.205 ;
        RECT 168.475 238.515 168.805 238.845 ;
        RECT 168.475 237.155 168.805 237.485 ;
        RECT 168.48 237.155 168.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 168.475 -0.845 168.805 -0.515 ;
        RECT 168.475 -2.205 168.805 -1.875 ;
        RECT 168.475 -3.565 168.805 -3.235 ;
        RECT 168.48 -3.565 168.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 244.04 170.165 245.17 ;
        RECT 169.835 239.875 170.165 240.205 ;
        RECT 169.835 238.515 170.165 238.845 ;
        RECT 169.835 237.155 170.165 237.485 ;
        RECT 169.84 237.155 170.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.835 -0.845 170.165 -0.515 ;
        RECT 169.835 -2.205 170.165 -1.875 ;
        RECT 169.835 -3.565 170.165 -3.235 ;
        RECT 169.84 -3.565 170.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 244.04 171.525 245.17 ;
        RECT 171.195 239.875 171.525 240.205 ;
        RECT 171.195 238.515 171.525 238.845 ;
        RECT 171.195 237.155 171.525 237.485 ;
        RECT 171.2 237.155 171.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 -0.845 171.525 -0.515 ;
        RECT 171.195 -2.205 171.525 -1.875 ;
        RECT 171.195 -3.565 171.525 -3.235 ;
        RECT 171.2 -3.565 171.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.195 -96.045 171.525 -95.715 ;
        RECT 171.195 -97.405 171.525 -97.075 ;
        RECT 171.195 -98.765 171.525 -98.435 ;
        RECT 171.195 -100.125 171.525 -99.795 ;
        RECT 171.195 -101.485 171.525 -101.155 ;
        RECT 171.195 -102.845 171.525 -102.515 ;
        RECT 171.195 -104.205 171.525 -103.875 ;
        RECT 171.195 -105.565 171.525 -105.235 ;
        RECT 171.195 -106.925 171.525 -106.595 ;
        RECT 171.195 -108.285 171.525 -107.955 ;
        RECT 171.195 -109.645 171.525 -109.315 ;
        RECT 171.195 -111.005 171.525 -110.675 ;
        RECT 171.195 -112.365 171.525 -112.035 ;
        RECT 171.195 -113.725 171.525 -113.395 ;
        RECT 171.195 -115.085 171.525 -114.755 ;
        RECT 171.195 -116.445 171.525 -116.115 ;
        RECT 171.195 -117.805 171.525 -117.475 ;
        RECT 171.195 -119.165 171.525 -118.835 ;
        RECT 171.195 -120.525 171.525 -120.195 ;
        RECT 171.195 -121.885 171.525 -121.555 ;
        RECT 171.195 -123.245 171.525 -122.915 ;
        RECT 171.195 -124.605 171.525 -124.275 ;
        RECT 171.195 -125.965 171.525 -125.635 ;
        RECT 171.195 -127.325 171.525 -126.995 ;
        RECT 171.195 -128.685 171.525 -128.355 ;
        RECT 171.195 -130.045 171.525 -129.715 ;
        RECT 171.195 -131.405 171.525 -131.075 ;
        RECT 171.195 -132.765 171.525 -132.435 ;
        RECT 171.195 -134.125 171.525 -133.795 ;
        RECT 171.195 -135.485 171.525 -135.155 ;
        RECT 171.195 -136.845 171.525 -136.515 ;
        RECT 171.195 -138.205 171.525 -137.875 ;
        RECT 171.195 -139.565 171.525 -139.235 ;
        RECT 171.195 -140.925 171.525 -140.595 ;
        RECT 171.195 -142.285 171.525 -141.955 ;
        RECT 171.195 -143.645 171.525 -143.315 ;
        RECT 171.195 -145.005 171.525 -144.675 ;
        RECT 171.195 -146.365 171.525 -146.035 ;
        RECT 171.195 -147.725 171.525 -147.395 ;
        RECT 171.195 -149.085 171.525 -148.755 ;
        RECT 171.195 -150.445 171.525 -150.115 ;
        RECT 171.195 -151.805 171.525 -151.475 ;
        RECT 171.195 -153.165 171.525 -152.835 ;
        RECT 171.195 -154.525 171.525 -154.195 ;
        RECT 171.195 -155.885 171.525 -155.555 ;
        RECT 171.195 -157.245 171.525 -156.915 ;
        RECT 171.195 -158.605 171.525 -158.275 ;
        RECT 171.195 -159.965 171.525 -159.635 ;
        RECT 171.195 -161.325 171.525 -160.995 ;
        RECT 171.195 -162.685 171.525 -162.355 ;
        RECT 171.195 -164.045 171.525 -163.715 ;
        RECT 171.195 -165.405 171.525 -165.075 ;
        RECT 171.195 -166.765 171.525 -166.435 ;
        RECT 171.195 -168.125 171.525 -167.795 ;
        RECT 171.195 -169.485 171.525 -169.155 ;
        RECT 171.195 -170.845 171.525 -170.515 ;
        RECT 171.195 -172.205 171.525 -171.875 ;
        RECT 171.195 -173.565 171.525 -173.235 ;
        RECT 171.195 -174.925 171.525 -174.595 ;
        RECT 171.195 -176.285 171.525 -175.955 ;
        RECT 171.195 -177.645 171.525 -177.315 ;
        RECT 171.195 -179.005 171.525 -178.675 ;
        RECT 171.195 -184.65 171.525 -183.52 ;
        RECT 171.2 -184.765 171.52 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 244.04 172.885 245.17 ;
        RECT 172.555 239.875 172.885 240.205 ;
        RECT 172.555 238.515 172.885 238.845 ;
        RECT 172.555 237.155 172.885 237.485 ;
        RECT 172.56 237.155 172.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 -0.845 172.885 -0.515 ;
        RECT 172.555 -2.205 172.885 -1.875 ;
        RECT 172.555 -3.565 172.885 -3.235 ;
        RECT 172.56 -3.565 172.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 172.555 -96.045 172.885 -95.715 ;
        RECT 172.555 -97.405 172.885 -97.075 ;
        RECT 172.555 -98.765 172.885 -98.435 ;
        RECT 172.555 -100.125 172.885 -99.795 ;
        RECT 172.555 -101.485 172.885 -101.155 ;
        RECT 172.555 -102.845 172.885 -102.515 ;
        RECT 172.555 -104.205 172.885 -103.875 ;
        RECT 172.555 -105.565 172.885 -105.235 ;
        RECT 172.555 -106.925 172.885 -106.595 ;
        RECT 172.555 -108.285 172.885 -107.955 ;
        RECT 172.555 -109.645 172.885 -109.315 ;
        RECT 172.555 -111.005 172.885 -110.675 ;
        RECT 172.555 -112.365 172.885 -112.035 ;
        RECT 172.555 -113.725 172.885 -113.395 ;
        RECT 172.555 -115.085 172.885 -114.755 ;
        RECT 172.555 -116.445 172.885 -116.115 ;
        RECT 172.555 -117.805 172.885 -117.475 ;
        RECT 172.555 -119.165 172.885 -118.835 ;
        RECT 172.555 -120.525 172.885 -120.195 ;
        RECT 172.555 -121.885 172.885 -121.555 ;
        RECT 172.555 -123.245 172.885 -122.915 ;
        RECT 172.555 -124.605 172.885 -124.275 ;
        RECT 172.555 -125.965 172.885 -125.635 ;
        RECT 172.555 -127.325 172.885 -126.995 ;
        RECT 172.555 -128.685 172.885 -128.355 ;
        RECT 172.555 -130.045 172.885 -129.715 ;
        RECT 172.555 -131.405 172.885 -131.075 ;
        RECT 172.555 -132.765 172.885 -132.435 ;
        RECT 172.555 -134.125 172.885 -133.795 ;
        RECT 172.555 -135.485 172.885 -135.155 ;
        RECT 172.555 -136.845 172.885 -136.515 ;
        RECT 172.555 -138.205 172.885 -137.875 ;
        RECT 172.555 -139.565 172.885 -139.235 ;
        RECT 172.555 -140.925 172.885 -140.595 ;
        RECT 172.555 -142.285 172.885 -141.955 ;
        RECT 172.555 -143.645 172.885 -143.315 ;
        RECT 172.555 -145.005 172.885 -144.675 ;
        RECT 172.555 -146.365 172.885 -146.035 ;
        RECT 172.555 -147.725 172.885 -147.395 ;
        RECT 172.555 -149.085 172.885 -148.755 ;
        RECT 172.555 -150.445 172.885 -150.115 ;
        RECT 172.555 -151.805 172.885 -151.475 ;
        RECT 172.555 -153.165 172.885 -152.835 ;
        RECT 172.555 -154.525 172.885 -154.195 ;
        RECT 172.555 -155.885 172.885 -155.555 ;
        RECT 172.555 -157.245 172.885 -156.915 ;
        RECT 172.555 -158.605 172.885 -158.275 ;
        RECT 172.555 -159.965 172.885 -159.635 ;
        RECT 172.555 -161.325 172.885 -160.995 ;
        RECT 172.555 -162.685 172.885 -162.355 ;
        RECT 172.555 -164.045 172.885 -163.715 ;
        RECT 172.555 -165.405 172.885 -165.075 ;
        RECT 172.555 -166.765 172.885 -166.435 ;
        RECT 172.555 -168.125 172.885 -167.795 ;
        RECT 172.555 -169.485 172.885 -169.155 ;
        RECT 172.555 -170.845 172.885 -170.515 ;
        RECT 172.555 -172.205 172.885 -171.875 ;
        RECT 172.555 -173.565 172.885 -173.235 ;
        RECT 172.555 -174.925 172.885 -174.595 ;
        RECT 172.555 -176.285 172.885 -175.955 ;
        RECT 172.555 -177.645 172.885 -177.315 ;
        RECT 172.555 -179.005 172.885 -178.675 ;
        RECT 172.555 -184.65 172.885 -183.52 ;
        RECT 172.56 -184.765 172.88 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 244.04 174.245 245.17 ;
        RECT 173.915 239.875 174.245 240.205 ;
        RECT 173.915 238.515 174.245 238.845 ;
        RECT 173.915 237.155 174.245 237.485 ;
        RECT 173.92 237.155 174.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 -0.845 174.245 -0.515 ;
        RECT 173.915 -2.205 174.245 -1.875 ;
        RECT 173.915 -3.565 174.245 -3.235 ;
        RECT 173.92 -3.565 174.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.915 -96.045 174.245 -95.715 ;
        RECT 173.915 -97.405 174.245 -97.075 ;
        RECT 173.915 -98.765 174.245 -98.435 ;
        RECT 173.915 -100.125 174.245 -99.795 ;
        RECT 173.915 -101.485 174.245 -101.155 ;
        RECT 173.915 -102.845 174.245 -102.515 ;
        RECT 173.915 -104.205 174.245 -103.875 ;
        RECT 173.915 -105.565 174.245 -105.235 ;
        RECT 173.915 -106.925 174.245 -106.595 ;
        RECT 173.915 -108.285 174.245 -107.955 ;
        RECT 173.915 -109.645 174.245 -109.315 ;
        RECT 173.915 -111.005 174.245 -110.675 ;
        RECT 173.915 -112.365 174.245 -112.035 ;
        RECT 173.915 -113.725 174.245 -113.395 ;
        RECT 173.915 -115.085 174.245 -114.755 ;
        RECT 173.915 -116.445 174.245 -116.115 ;
        RECT 173.915 -117.805 174.245 -117.475 ;
        RECT 173.915 -119.165 174.245 -118.835 ;
        RECT 173.915 -120.525 174.245 -120.195 ;
        RECT 173.915 -121.885 174.245 -121.555 ;
        RECT 173.915 -123.245 174.245 -122.915 ;
        RECT 173.915 -124.605 174.245 -124.275 ;
        RECT 173.915 -125.965 174.245 -125.635 ;
        RECT 173.915 -127.325 174.245 -126.995 ;
        RECT 173.915 -128.685 174.245 -128.355 ;
        RECT 173.915 -130.045 174.245 -129.715 ;
        RECT 173.915 -131.405 174.245 -131.075 ;
        RECT 173.915 -132.765 174.245 -132.435 ;
        RECT 173.915 -134.125 174.245 -133.795 ;
        RECT 173.915 -135.485 174.245 -135.155 ;
        RECT 173.915 -136.845 174.245 -136.515 ;
        RECT 173.915 -138.205 174.245 -137.875 ;
        RECT 173.915 -139.565 174.245 -139.235 ;
        RECT 173.915 -140.925 174.245 -140.595 ;
        RECT 173.915 -142.285 174.245 -141.955 ;
        RECT 173.915 -143.645 174.245 -143.315 ;
        RECT 173.915 -145.005 174.245 -144.675 ;
        RECT 173.915 -146.365 174.245 -146.035 ;
        RECT 173.915 -147.725 174.245 -147.395 ;
        RECT 173.915 -149.085 174.245 -148.755 ;
        RECT 173.915 -150.445 174.245 -150.115 ;
        RECT 173.915 -151.805 174.245 -151.475 ;
        RECT 173.915 -153.165 174.245 -152.835 ;
        RECT 173.915 -154.525 174.245 -154.195 ;
        RECT 173.915 -155.885 174.245 -155.555 ;
        RECT 173.915 -157.245 174.245 -156.915 ;
        RECT 173.915 -158.605 174.245 -158.275 ;
        RECT 173.915 -159.965 174.245 -159.635 ;
        RECT 173.915 -161.325 174.245 -160.995 ;
        RECT 173.915 -162.685 174.245 -162.355 ;
        RECT 173.915 -164.045 174.245 -163.715 ;
        RECT 173.915 -165.405 174.245 -165.075 ;
        RECT 173.915 -166.765 174.245 -166.435 ;
        RECT 173.915 -168.125 174.245 -167.795 ;
        RECT 173.915 -169.485 174.245 -169.155 ;
        RECT 173.915 -170.845 174.245 -170.515 ;
        RECT 173.915 -172.205 174.245 -171.875 ;
        RECT 173.915 -173.565 174.245 -173.235 ;
        RECT 173.915 -174.925 174.245 -174.595 ;
        RECT 173.915 -176.285 174.245 -175.955 ;
        RECT 173.915 -177.645 174.245 -177.315 ;
        RECT 173.915 -179.005 174.245 -178.675 ;
        RECT 173.915 -184.65 174.245 -183.52 ;
        RECT 173.92 -184.765 174.24 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 244.04 175.605 245.17 ;
        RECT 175.275 239.875 175.605 240.205 ;
        RECT 175.275 238.515 175.605 238.845 ;
        RECT 175.275 237.155 175.605 237.485 ;
        RECT 175.28 237.155 175.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 -0.845 175.605 -0.515 ;
        RECT 175.275 -2.205 175.605 -1.875 ;
        RECT 175.275 -3.565 175.605 -3.235 ;
        RECT 175.28 -3.565 175.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.275 -96.045 175.605 -95.715 ;
        RECT 175.275 -97.405 175.605 -97.075 ;
        RECT 175.275 -98.765 175.605 -98.435 ;
        RECT 175.275 -100.125 175.605 -99.795 ;
        RECT 175.275 -101.485 175.605 -101.155 ;
        RECT 175.275 -102.845 175.605 -102.515 ;
        RECT 175.275 -104.205 175.605 -103.875 ;
        RECT 175.275 -105.565 175.605 -105.235 ;
        RECT 175.275 -106.925 175.605 -106.595 ;
        RECT 175.275 -108.285 175.605 -107.955 ;
        RECT 175.275 -109.645 175.605 -109.315 ;
        RECT 175.275 -111.005 175.605 -110.675 ;
        RECT 175.275 -112.365 175.605 -112.035 ;
        RECT 175.275 -113.725 175.605 -113.395 ;
        RECT 175.275 -115.085 175.605 -114.755 ;
        RECT 175.275 -116.445 175.605 -116.115 ;
        RECT 175.275 -117.805 175.605 -117.475 ;
        RECT 175.275 -119.165 175.605 -118.835 ;
        RECT 175.275 -120.525 175.605 -120.195 ;
        RECT 175.275 -121.885 175.605 -121.555 ;
        RECT 175.275 -123.245 175.605 -122.915 ;
        RECT 175.275 -124.605 175.605 -124.275 ;
        RECT 175.275 -125.965 175.605 -125.635 ;
        RECT 175.275 -127.325 175.605 -126.995 ;
        RECT 175.275 -128.685 175.605 -128.355 ;
        RECT 175.275 -130.045 175.605 -129.715 ;
        RECT 175.275 -131.405 175.605 -131.075 ;
        RECT 175.275 -132.765 175.605 -132.435 ;
        RECT 175.275 -134.125 175.605 -133.795 ;
        RECT 175.275 -135.485 175.605 -135.155 ;
        RECT 175.275 -136.845 175.605 -136.515 ;
        RECT 175.275 -138.205 175.605 -137.875 ;
        RECT 175.275 -139.565 175.605 -139.235 ;
        RECT 175.275 -140.925 175.605 -140.595 ;
        RECT 175.275 -142.285 175.605 -141.955 ;
        RECT 175.275 -143.645 175.605 -143.315 ;
        RECT 175.275 -145.005 175.605 -144.675 ;
        RECT 175.275 -146.365 175.605 -146.035 ;
        RECT 175.275 -147.725 175.605 -147.395 ;
        RECT 175.275 -149.085 175.605 -148.755 ;
        RECT 175.275 -150.445 175.605 -150.115 ;
        RECT 175.275 -151.805 175.605 -151.475 ;
        RECT 175.275 -153.165 175.605 -152.835 ;
        RECT 175.275 -154.525 175.605 -154.195 ;
        RECT 175.275 -155.885 175.605 -155.555 ;
        RECT 175.275 -157.245 175.605 -156.915 ;
        RECT 175.275 -158.605 175.605 -158.275 ;
        RECT 175.275 -159.965 175.605 -159.635 ;
        RECT 175.275 -161.325 175.605 -160.995 ;
        RECT 175.275 -162.685 175.605 -162.355 ;
        RECT 175.275 -164.045 175.605 -163.715 ;
        RECT 175.275 -165.405 175.605 -165.075 ;
        RECT 175.275 -166.765 175.605 -166.435 ;
        RECT 175.275 -168.125 175.605 -167.795 ;
        RECT 175.275 -169.485 175.605 -169.155 ;
        RECT 175.275 -170.845 175.605 -170.515 ;
        RECT 175.275 -172.205 175.605 -171.875 ;
        RECT 175.275 -173.565 175.605 -173.235 ;
        RECT 175.275 -174.925 175.605 -174.595 ;
        RECT 175.275 -176.285 175.605 -175.955 ;
        RECT 175.275 -177.645 175.605 -177.315 ;
        RECT 175.275 -179.005 175.605 -178.675 ;
        RECT 175.275 -184.65 175.605 -183.52 ;
        RECT 175.28 -184.765 175.6 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 244.04 176.965 245.17 ;
        RECT 176.635 239.875 176.965 240.205 ;
        RECT 176.635 238.515 176.965 238.845 ;
        RECT 176.635 237.155 176.965 237.485 ;
        RECT 176.64 237.155 176.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 176.635 -98.765 176.965 -98.435 ;
        RECT 176.635 -100.125 176.965 -99.795 ;
        RECT 176.635 -101.485 176.965 -101.155 ;
        RECT 176.635 -102.845 176.965 -102.515 ;
        RECT 176.635 -104.205 176.965 -103.875 ;
        RECT 176.635 -105.565 176.965 -105.235 ;
        RECT 176.635 -106.925 176.965 -106.595 ;
        RECT 176.635 -108.285 176.965 -107.955 ;
        RECT 176.635 -109.645 176.965 -109.315 ;
        RECT 176.635 -111.005 176.965 -110.675 ;
        RECT 176.635 -112.365 176.965 -112.035 ;
        RECT 176.635 -113.725 176.965 -113.395 ;
        RECT 176.635 -115.085 176.965 -114.755 ;
        RECT 176.635 -116.445 176.965 -116.115 ;
        RECT 176.635 -117.805 176.965 -117.475 ;
        RECT 176.635 -119.165 176.965 -118.835 ;
        RECT 176.635 -120.525 176.965 -120.195 ;
        RECT 176.635 -121.885 176.965 -121.555 ;
        RECT 176.635 -123.245 176.965 -122.915 ;
        RECT 176.635 -124.605 176.965 -124.275 ;
        RECT 176.635 -125.965 176.965 -125.635 ;
        RECT 176.635 -127.325 176.965 -126.995 ;
        RECT 176.635 -128.685 176.965 -128.355 ;
        RECT 176.635 -130.045 176.965 -129.715 ;
        RECT 176.635 -131.405 176.965 -131.075 ;
        RECT 176.635 -132.765 176.965 -132.435 ;
        RECT 176.635 -134.125 176.965 -133.795 ;
        RECT 176.635 -135.485 176.965 -135.155 ;
        RECT 176.635 -136.845 176.965 -136.515 ;
        RECT 176.635 -138.205 176.965 -137.875 ;
        RECT 176.635 -139.565 176.965 -139.235 ;
        RECT 176.635 -140.925 176.965 -140.595 ;
        RECT 176.635 -142.285 176.965 -141.955 ;
        RECT 176.635 -143.645 176.965 -143.315 ;
        RECT 176.635 -145.005 176.965 -144.675 ;
        RECT 176.635 -146.365 176.965 -146.035 ;
        RECT 176.635 -147.725 176.965 -147.395 ;
        RECT 176.635 -149.085 176.965 -148.755 ;
        RECT 176.635 -150.445 176.965 -150.115 ;
        RECT 176.635 -151.805 176.965 -151.475 ;
        RECT 176.635 -153.165 176.965 -152.835 ;
        RECT 176.635 -154.525 176.965 -154.195 ;
        RECT 176.635 -155.885 176.965 -155.555 ;
        RECT 176.635 -157.245 176.965 -156.915 ;
        RECT 176.635 -158.605 176.965 -158.275 ;
        RECT 176.635 -159.965 176.965 -159.635 ;
        RECT 176.635 -161.325 176.965 -160.995 ;
        RECT 176.635 -162.685 176.965 -162.355 ;
        RECT 176.635 -164.045 176.965 -163.715 ;
        RECT 176.635 -165.405 176.965 -165.075 ;
        RECT 176.635 -166.765 176.965 -166.435 ;
        RECT 176.635 -168.125 176.965 -167.795 ;
        RECT 176.635 -169.485 176.965 -169.155 ;
        RECT 176.635 -170.845 176.965 -170.515 ;
        RECT 176.635 -172.205 176.965 -171.875 ;
        RECT 176.635 -173.565 176.965 -173.235 ;
        RECT 176.635 -174.925 176.965 -174.595 ;
        RECT 176.635 -176.285 176.965 -175.955 ;
        RECT 176.635 -177.645 176.965 -177.315 ;
        RECT 176.635 -179.005 176.965 -178.675 ;
        RECT 176.635 -184.65 176.965 -183.52 ;
        RECT 176.64 -184.765 176.96 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.06 -98.075 177.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.995 244.04 178.325 245.17 ;
        RECT 177.995 239.875 178.325 240.205 ;
        RECT 177.995 238.515 178.325 238.845 ;
        RECT 177.995 237.155 178.325 237.485 ;
        RECT 178 237.155 178.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 244.04 179.685 245.17 ;
        RECT 179.355 239.875 179.685 240.205 ;
        RECT 179.355 238.515 179.685 238.845 ;
        RECT 179.355 237.155 179.685 237.485 ;
        RECT 179.36 237.155 179.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 179.355 -0.845 179.685 -0.515 ;
        RECT 179.355 -2.205 179.685 -1.875 ;
        RECT 179.355 -3.565 179.685 -3.235 ;
        RECT 179.36 -3.565 179.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.715 244.04 181.045 245.17 ;
        RECT 180.715 239.875 181.045 240.205 ;
        RECT 180.715 238.515 181.045 238.845 ;
        RECT 180.715 237.155 181.045 237.485 ;
        RECT 180.72 237.155 181.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.715 -0.845 181.045 -0.515 ;
        RECT 180.715 -2.205 181.045 -1.875 ;
        RECT 180.715 -3.565 181.045 -3.235 ;
        RECT 180.72 -3.565 181.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 244.04 182.405 245.17 ;
        RECT 182.075 239.875 182.405 240.205 ;
        RECT 182.075 238.515 182.405 238.845 ;
        RECT 182.075 237.155 182.405 237.485 ;
        RECT 182.08 237.155 182.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 -0.845 182.405 -0.515 ;
        RECT 182.075 -2.205 182.405 -1.875 ;
        RECT 182.075 -3.565 182.405 -3.235 ;
        RECT 182.08 -3.565 182.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.075 -96.045 182.405 -95.715 ;
        RECT 182.075 -97.405 182.405 -97.075 ;
        RECT 182.075 -98.765 182.405 -98.435 ;
        RECT 182.075 -100.125 182.405 -99.795 ;
        RECT 182.075 -101.485 182.405 -101.155 ;
        RECT 182.075 -102.845 182.405 -102.515 ;
        RECT 182.075 -104.205 182.405 -103.875 ;
        RECT 182.075 -105.565 182.405 -105.235 ;
        RECT 182.075 -106.925 182.405 -106.595 ;
        RECT 182.075 -108.285 182.405 -107.955 ;
        RECT 182.075 -109.645 182.405 -109.315 ;
        RECT 182.075 -111.005 182.405 -110.675 ;
        RECT 182.075 -112.365 182.405 -112.035 ;
        RECT 182.075 -113.725 182.405 -113.395 ;
        RECT 182.075 -115.085 182.405 -114.755 ;
        RECT 182.075 -116.445 182.405 -116.115 ;
        RECT 182.075 -117.805 182.405 -117.475 ;
        RECT 182.075 -119.165 182.405 -118.835 ;
        RECT 182.075 -120.525 182.405 -120.195 ;
        RECT 182.075 -121.885 182.405 -121.555 ;
        RECT 182.075 -123.245 182.405 -122.915 ;
        RECT 182.075 -124.605 182.405 -124.275 ;
        RECT 182.075 -125.965 182.405 -125.635 ;
        RECT 182.075 -127.325 182.405 -126.995 ;
        RECT 182.075 -128.685 182.405 -128.355 ;
        RECT 182.075 -130.045 182.405 -129.715 ;
        RECT 182.075 -131.405 182.405 -131.075 ;
        RECT 182.075 -132.765 182.405 -132.435 ;
        RECT 182.075 -134.125 182.405 -133.795 ;
        RECT 182.075 -135.485 182.405 -135.155 ;
        RECT 182.075 -136.845 182.405 -136.515 ;
        RECT 182.075 -138.205 182.405 -137.875 ;
        RECT 182.075 -139.565 182.405 -139.235 ;
        RECT 182.075 -140.925 182.405 -140.595 ;
        RECT 182.075 -142.285 182.405 -141.955 ;
        RECT 182.075 -143.645 182.405 -143.315 ;
        RECT 182.075 -145.005 182.405 -144.675 ;
        RECT 182.075 -146.365 182.405 -146.035 ;
        RECT 182.075 -147.725 182.405 -147.395 ;
        RECT 182.075 -149.085 182.405 -148.755 ;
        RECT 182.075 -150.445 182.405 -150.115 ;
        RECT 182.075 -151.805 182.405 -151.475 ;
        RECT 182.075 -153.165 182.405 -152.835 ;
        RECT 182.075 -154.525 182.405 -154.195 ;
        RECT 182.075 -155.885 182.405 -155.555 ;
        RECT 182.075 -157.245 182.405 -156.915 ;
        RECT 182.075 -158.605 182.405 -158.275 ;
        RECT 182.075 -159.965 182.405 -159.635 ;
        RECT 182.075 -161.325 182.405 -160.995 ;
        RECT 182.075 -162.685 182.405 -162.355 ;
        RECT 182.075 -164.045 182.405 -163.715 ;
        RECT 182.075 -165.405 182.405 -165.075 ;
        RECT 182.075 -166.765 182.405 -166.435 ;
        RECT 182.075 -168.125 182.405 -167.795 ;
        RECT 182.075 -169.485 182.405 -169.155 ;
        RECT 182.075 -170.845 182.405 -170.515 ;
        RECT 182.075 -172.205 182.405 -171.875 ;
        RECT 182.075 -173.565 182.405 -173.235 ;
        RECT 182.075 -174.925 182.405 -174.595 ;
        RECT 182.075 -176.285 182.405 -175.955 ;
        RECT 182.075 -177.645 182.405 -177.315 ;
        RECT 182.075 -179.005 182.405 -178.675 ;
        RECT 182.075 -184.65 182.405 -183.52 ;
        RECT 182.08 -184.765 182.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 244.04 183.765 245.17 ;
        RECT 183.435 239.875 183.765 240.205 ;
        RECT 183.435 238.515 183.765 238.845 ;
        RECT 183.435 237.155 183.765 237.485 ;
        RECT 183.44 237.155 183.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 -0.845 183.765 -0.515 ;
        RECT 183.435 -2.205 183.765 -1.875 ;
        RECT 183.435 -3.565 183.765 -3.235 ;
        RECT 183.44 -3.565 183.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 183.435 -96.045 183.765 -95.715 ;
        RECT 183.435 -97.405 183.765 -97.075 ;
        RECT 183.435 -98.765 183.765 -98.435 ;
        RECT 183.435 -100.125 183.765 -99.795 ;
        RECT 183.435 -101.485 183.765 -101.155 ;
        RECT 183.435 -102.845 183.765 -102.515 ;
        RECT 183.435 -104.205 183.765 -103.875 ;
        RECT 183.435 -105.565 183.765 -105.235 ;
        RECT 183.435 -106.925 183.765 -106.595 ;
        RECT 183.435 -108.285 183.765 -107.955 ;
        RECT 183.435 -109.645 183.765 -109.315 ;
        RECT 183.435 -111.005 183.765 -110.675 ;
        RECT 183.435 -112.365 183.765 -112.035 ;
        RECT 183.435 -113.725 183.765 -113.395 ;
        RECT 183.435 -115.085 183.765 -114.755 ;
        RECT 183.435 -116.445 183.765 -116.115 ;
        RECT 183.435 -117.805 183.765 -117.475 ;
        RECT 183.435 -119.165 183.765 -118.835 ;
        RECT 183.435 -120.525 183.765 -120.195 ;
        RECT 183.435 -121.885 183.765 -121.555 ;
        RECT 183.435 -123.245 183.765 -122.915 ;
        RECT 183.435 -124.605 183.765 -124.275 ;
        RECT 183.435 -125.965 183.765 -125.635 ;
        RECT 183.435 -127.325 183.765 -126.995 ;
        RECT 183.435 -128.685 183.765 -128.355 ;
        RECT 183.435 -130.045 183.765 -129.715 ;
        RECT 183.435 -131.405 183.765 -131.075 ;
        RECT 183.435 -132.765 183.765 -132.435 ;
        RECT 183.435 -134.125 183.765 -133.795 ;
        RECT 183.435 -135.485 183.765 -135.155 ;
        RECT 183.435 -136.845 183.765 -136.515 ;
        RECT 183.435 -138.205 183.765 -137.875 ;
        RECT 183.435 -139.565 183.765 -139.235 ;
        RECT 183.435 -140.925 183.765 -140.595 ;
        RECT 183.435 -142.285 183.765 -141.955 ;
        RECT 183.435 -143.645 183.765 -143.315 ;
        RECT 183.435 -145.005 183.765 -144.675 ;
        RECT 183.435 -146.365 183.765 -146.035 ;
        RECT 183.435 -147.725 183.765 -147.395 ;
        RECT 183.435 -149.085 183.765 -148.755 ;
        RECT 183.435 -150.445 183.765 -150.115 ;
        RECT 183.435 -151.805 183.765 -151.475 ;
        RECT 183.435 -153.165 183.765 -152.835 ;
        RECT 183.435 -154.525 183.765 -154.195 ;
        RECT 183.435 -155.885 183.765 -155.555 ;
        RECT 183.435 -157.245 183.765 -156.915 ;
        RECT 183.435 -158.605 183.765 -158.275 ;
        RECT 183.435 -159.965 183.765 -159.635 ;
        RECT 183.435 -161.325 183.765 -160.995 ;
        RECT 183.435 -162.685 183.765 -162.355 ;
        RECT 183.435 -164.045 183.765 -163.715 ;
        RECT 183.435 -165.405 183.765 -165.075 ;
        RECT 183.435 -166.765 183.765 -166.435 ;
        RECT 183.435 -168.125 183.765 -167.795 ;
        RECT 183.435 -169.485 183.765 -169.155 ;
        RECT 183.435 -170.845 183.765 -170.515 ;
        RECT 183.435 -172.205 183.765 -171.875 ;
        RECT 183.435 -173.565 183.765 -173.235 ;
        RECT 183.435 -174.925 183.765 -174.595 ;
        RECT 183.435 -176.285 183.765 -175.955 ;
        RECT 183.435 -177.645 183.765 -177.315 ;
        RECT 183.435 -179.005 183.765 -178.675 ;
        RECT 183.435 -184.65 183.765 -183.52 ;
        RECT 183.44 -184.765 183.76 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 244.04 185.125 245.17 ;
        RECT 184.795 239.875 185.125 240.205 ;
        RECT 184.795 238.515 185.125 238.845 ;
        RECT 184.795 237.155 185.125 237.485 ;
        RECT 184.8 237.155 185.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 -0.845 185.125 -0.515 ;
        RECT 184.795 -2.205 185.125 -1.875 ;
        RECT 184.795 -3.565 185.125 -3.235 ;
        RECT 184.8 -3.565 185.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.795 -135.485 185.125 -135.155 ;
        RECT 184.795 -136.845 185.125 -136.515 ;
        RECT 184.795 -138.205 185.125 -137.875 ;
        RECT 184.795 -139.565 185.125 -139.235 ;
        RECT 184.795 -140.925 185.125 -140.595 ;
        RECT 184.795 -142.285 185.125 -141.955 ;
        RECT 184.795 -143.645 185.125 -143.315 ;
        RECT 184.795 -145.005 185.125 -144.675 ;
        RECT 184.795 -146.365 185.125 -146.035 ;
        RECT 184.795 -147.725 185.125 -147.395 ;
        RECT 184.795 -149.085 185.125 -148.755 ;
        RECT 184.795 -150.445 185.125 -150.115 ;
        RECT 184.795 -151.805 185.125 -151.475 ;
        RECT 184.795 -153.165 185.125 -152.835 ;
        RECT 184.795 -154.525 185.125 -154.195 ;
        RECT 184.795 -155.885 185.125 -155.555 ;
        RECT 184.795 -157.245 185.125 -156.915 ;
        RECT 184.795 -158.605 185.125 -158.275 ;
        RECT 184.795 -159.965 185.125 -159.635 ;
        RECT 184.795 -161.325 185.125 -160.995 ;
        RECT 184.795 -162.685 185.125 -162.355 ;
        RECT 184.795 -164.045 185.125 -163.715 ;
        RECT 184.795 -165.405 185.125 -165.075 ;
        RECT 184.795 -166.765 185.125 -166.435 ;
        RECT 184.795 -168.125 185.125 -167.795 ;
        RECT 184.795 -169.485 185.125 -169.155 ;
        RECT 184.795 -170.845 185.125 -170.515 ;
        RECT 184.795 -172.205 185.125 -171.875 ;
        RECT 184.795 -173.565 185.125 -173.235 ;
        RECT 184.795 -174.925 185.125 -174.595 ;
        RECT 184.795 -176.285 185.125 -175.955 ;
        RECT 184.795 -177.645 185.125 -177.315 ;
        RECT 184.795 -179.005 185.125 -178.675 ;
        RECT 184.795 -184.65 185.125 -183.52 ;
        RECT 184.8 -184.765 185.12 -95.04 ;
        RECT 184.795 -96.045 185.125 -95.715 ;
        RECT 184.795 -97.405 185.125 -97.075 ;
        RECT 184.795 -98.765 185.125 -98.435 ;
        RECT 184.795 -100.125 185.125 -99.795 ;
        RECT 184.795 -101.485 185.125 -101.155 ;
        RECT 184.795 -102.845 185.125 -102.515 ;
        RECT 184.795 -104.205 185.125 -103.875 ;
        RECT 184.795 -105.565 185.125 -105.235 ;
        RECT 184.795 -106.925 185.125 -106.595 ;
        RECT 184.795 -108.285 185.125 -107.955 ;
        RECT 184.795 -109.645 185.125 -109.315 ;
        RECT 184.795 -111.005 185.125 -110.675 ;
        RECT 184.795 -112.365 185.125 -112.035 ;
        RECT 184.795 -113.725 185.125 -113.395 ;
        RECT 184.795 -115.085 185.125 -114.755 ;
        RECT 184.795 -116.445 185.125 -116.115 ;
        RECT 184.795 -117.805 185.125 -117.475 ;
        RECT 184.795 -119.165 185.125 -118.835 ;
        RECT 184.795 -120.525 185.125 -120.195 ;
        RECT 184.795 -121.885 185.125 -121.555 ;
        RECT 184.795 -123.245 185.125 -122.915 ;
        RECT 184.795 -124.605 185.125 -124.275 ;
        RECT 184.795 -125.965 185.125 -125.635 ;
        RECT 184.795 -127.325 185.125 -126.995 ;
        RECT 184.795 -128.685 185.125 -128.355 ;
        RECT 184.795 -130.045 185.125 -129.715 ;
        RECT 184.795 -131.405 185.125 -131.075 ;
        RECT 184.795 -132.765 185.125 -132.435 ;
        RECT 184.795 -134.125 185.125 -133.795 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 -98.765 133.445 -98.435 ;
        RECT 133.115 -100.125 133.445 -99.795 ;
        RECT 133.115 -101.485 133.445 -101.155 ;
        RECT 133.115 -102.845 133.445 -102.515 ;
        RECT 133.115 -104.205 133.445 -103.875 ;
        RECT 133.115 -105.565 133.445 -105.235 ;
        RECT 133.115 -106.925 133.445 -106.595 ;
        RECT 133.115 -108.285 133.445 -107.955 ;
        RECT 133.115 -109.645 133.445 -109.315 ;
        RECT 133.115 -111.005 133.445 -110.675 ;
        RECT 133.115 -112.365 133.445 -112.035 ;
        RECT 133.115 -113.725 133.445 -113.395 ;
        RECT 133.115 -115.085 133.445 -114.755 ;
        RECT 133.115 -116.445 133.445 -116.115 ;
        RECT 133.115 -117.805 133.445 -117.475 ;
        RECT 133.115 -119.165 133.445 -118.835 ;
        RECT 133.115 -120.525 133.445 -120.195 ;
        RECT 133.115 -121.885 133.445 -121.555 ;
        RECT 133.115 -123.245 133.445 -122.915 ;
        RECT 133.115 -124.605 133.445 -124.275 ;
        RECT 133.115 -125.965 133.445 -125.635 ;
        RECT 133.115 -127.325 133.445 -126.995 ;
        RECT 133.115 -128.685 133.445 -128.355 ;
        RECT 133.115 -130.045 133.445 -129.715 ;
        RECT 133.115 -131.405 133.445 -131.075 ;
        RECT 133.115 -132.765 133.445 -132.435 ;
        RECT 133.115 -134.125 133.445 -133.795 ;
        RECT 133.115 -135.485 133.445 -135.155 ;
        RECT 133.115 -136.845 133.445 -136.515 ;
        RECT 133.115 -138.205 133.445 -137.875 ;
        RECT 133.115 -139.565 133.445 -139.235 ;
        RECT 133.115 -140.925 133.445 -140.595 ;
        RECT 133.115 -142.285 133.445 -141.955 ;
        RECT 133.115 -143.645 133.445 -143.315 ;
        RECT 133.115 -145.005 133.445 -144.675 ;
        RECT 133.115 -146.365 133.445 -146.035 ;
        RECT 133.115 -147.725 133.445 -147.395 ;
        RECT 133.115 -149.085 133.445 -148.755 ;
        RECT 133.115 -150.445 133.445 -150.115 ;
        RECT 133.115 -151.805 133.445 -151.475 ;
        RECT 133.115 -153.165 133.445 -152.835 ;
        RECT 133.115 -154.525 133.445 -154.195 ;
        RECT 133.115 -155.885 133.445 -155.555 ;
        RECT 133.115 -157.245 133.445 -156.915 ;
        RECT 133.115 -158.605 133.445 -158.275 ;
        RECT 133.115 -159.965 133.445 -159.635 ;
        RECT 133.115 -161.325 133.445 -160.995 ;
        RECT 133.115 -162.685 133.445 -162.355 ;
        RECT 133.115 -164.045 133.445 -163.715 ;
        RECT 133.115 -165.405 133.445 -165.075 ;
        RECT 133.115 -166.765 133.445 -166.435 ;
        RECT 133.115 -168.125 133.445 -167.795 ;
        RECT 133.115 -169.485 133.445 -169.155 ;
        RECT 133.115 -170.845 133.445 -170.515 ;
        RECT 133.115 -172.205 133.445 -171.875 ;
        RECT 133.115 -173.565 133.445 -173.235 ;
        RECT 133.115 -174.925 133.445 -174.595 ;
        RECT 133.115 -176.285 133.445 -175.955 ;
        RECT 133.115 -177.645 133.445 -177.315 ;
        RECT 133.115 -179.005 133.445 -178.675 ;
        RECT 133.115 -184.65 133.445 -183.52 ;
        RECT 133.12 -184.765 133.44 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.46 -98.075 133.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.475 244.04 134.805 245.17 ;
        RECT 134.475 239.875 134.805 240.205 ;
        RECT 134.475 238.515 134.805 238.845 ;
        RECT 134.475 237.155 134.805 237.485 ;
        RECT 134.48 237.155 134.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 244.04 136.165 245.17 ;
        RECT 135.835 239.875 136.165 240.205 ;
        RECT 135.835 238.515 136.165 238.845 ;
        RECT 135.835 237.155 136.165 237.485 ;
        RECT 135.84 237.155 136.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.835 -0.845 136.165 -0.515 ;
        RECT 135.835 -2.205 136.165 -1.875 ;
        RECT 135.835 -3.565 136.165 -3.235 ;
        RECT 135.84 -3.565 136.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 244.04 137.525 245.17 ;
        RECT 137.195 239.875 137.525 240.205 ;
        RECT 137.195 238.515 137.525 238.845 ;
        RECT 137.195 237.155 137.525 237.485 ;
        RECT 137.2 237.155 137.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 -0.845 137.525 -0.515 ;
        RECT 137.195 -2.205 137.525 -1.875 ;
        RECT 137.195 -3.565 137.525 -3.235 ;
        RECT 137.2 -3.565 137.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.195 -96.045 137.525 -95.715 ;
        RECT 137.195 -97.405 137.525 -97.075 ;
        RECT 137.195 -98.765 137.525 -98.435 ;
        RECT 137.195 -100.125 137.525 -99.795 ;
        RECT 137.195 -101.485 137.525 -101.155 ;
        RECT 137.195 -102.845 137.525 -102.515 ;
        RECT 137.195 -104.205 137.525 -103.875 ;
        RECT 137.195 -105.565 137.525 -105.235 ;
        RECT 137.195 -106.925 137.525 -106.595 ;
        RECT 137.195 -108.285 137.525 -107.955 ;
        RECT 137.195 -109.645 137.525 -109.315 ;
        RECT 137.195 -111.005 137.525 -110.675 ;
        RECT 137.195 -112.365 137.525 -112.035 ;
        RECT 137.195 -113.725 137.525 -113.395 ;
        RECT 137.195 -115.085 137.525 -114.755 ;
        RECT 137.195 -116.445 137.525 -116.115 ;
        RECT 137.195 -117.805 137.525 -117.475 ;
        RECT 137.195 -119.165 137.525 -118.835 ;
        RECT 137.195 -120.525 137.525 -120.195 ;
        RECT 137.195 -121.885 137.525 -121.555 ;
        RECT 137.195 -123.245 137.525 -122.915 ;
        RECT 137.195 -124.605 137.525 -124.275 ;
        RECT 137.195 -125.965 137.525 -125.635 ;
        RECT 137.195 -127.325 137.525 -126.995 ;
        RECT 137.195 -128.685 137.525 -128.355 ;
        RECT 137.195 -130.045 137.525 -129.715 ;
        RECT 137.195 -131.405 137.525 -131.075 ;
        RECT 137.195 -132.765 137.525 -132.435 ;
        RECT 137.195 -134.125 137.525 -133.795 ;
        RECT 137.195 -135.485 137.525 -135.155 ;
        RECT 137.195 -136.845 137.525 -136.515 ;
        RECT 137.195 -138.205 137.525 -137.875 ;
        RECT 137.195 -139.565 137.525 -139.235 ;
        RECT 137.195 -140.925 137.525 -140.595 ;
        RECT 137.195 -142.285 137.525 -141.955 ;
        RECT 137.195 -143.645 137.525 -143.315 ;
        RECT 137.195 -145.005 137.525 -144.675 ;
        RECT 137.195 -146.365 137.525 -146.035 ;
        RECT 137.195 -147.725 137.525 -147.395 ;
        RECT 137.195 -149.085 137.525 -148.755 ;
        RECT 137.195 -150.445 137.525 -150.115 ;
        RECT 137.195 -151.805 137.525 -151.475 ;
        RECT 137.195 -153.165 137.525 -152.835 ;
        RECT 137.195 -154.525 137.525 -154.195 ;
        RECT 137.195 -155.885 137.525 -155.555 ;
        RECT 137.195 -157.245 137.525 -156.915 ;
        RECT 137.195 -158.605 137.525 -158.275 ;
        RECT 137.195 -159.965 137.525 -159.635 ;
        RECT 137.195 -161.325 137.525 -160.995 ;
        RECT 137.195 -162.685 137.525 -162.355 ;
        RECT 137.195 -164.045 137.525 -163.715 ;
        RECT 137.195 -165.405 137.525 -165.075 ;
        RECT 137.195 -166.765 137.525 -166.435 ;
        RECT 137.195 -168.125 137.525 -167.795 ;
        RECT 137.195 -169.485 137.525 -169.155 ;
        RECT 137.195 -170.845 137.525 -170.515 ;
        RECT 137.195 -172.205 137.525 -171.875 ;
        RECT 137.195 -173.565 137.525 -173.235 ;
        RECT 137.195 -174.925 137.525 -174.595 ;
        RECT 137.195 -176.285 137.525 -175.955 ;
        RECT 137.195 -177.645 137.525 -177.315 ;
        RECT 137.195 -179.005 137.525 -178.675 ;
        RECT 137.195 -184.65 137.525 -183.52 ;
        RECT 137.2 -184.765 137.52 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 244.04 138.885 245.17 ;
        RECT 138.555 239.875 138.885 240.205 ;
        RECT 138.555 238.515 138.885 238.845 ;
        RECT 138.555 237.155 138.885 237.485 ;
        RECT 138.56 237.155 138.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 -0.845 138.885 -0.515 ;
        RECT 138.555 -2.205 138.885 -1.875 ;
        RECT 138.555 -3.565 138.885 -3.235 ;
        RECT 138.56 -3.565 138.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 138.555 -96.045 138.885 -95.715 ;
        RECT 138.555 -97.405 138.885 -97.075 ;
        RECT 138.555 -98.765 138.885 -98.435 ;
        RECT 138.555 -100.125 138.885 -99.795 ;
        RECT 138.555 -101.485 138.885 -101.155 ;
        RECT 138.555 -102.845 138.885 -102.515 ;
        RECT 138.555 -104.205 138.885 -103.875 ;
        RECT 138.555 -105.565 138.885 -105.235 ;
        RECT 138.555 -106.925 138.885 -106.595 ;
        RECT 138.555 -108.285 138.885 -107.955 ;
        RECT 138.555 -109.645 138.885 -109.315 ;
        RECT 138.555 -111.005 138.885 -110.675 ;
        RECT 138.555 -112.365 138.885 -112.035 ;
        RECT 138.555 -113.725 138.885 -113.395 ;
        RECT 138.555 -115.085 138.885 -114.755 ;
        RECT 138.555 -116.445 138.885 -116.115 ;
        RECT 138.555 -117.805 138.885 -117.475 ;
        RECT 138.555 -119.165 138.885 -118.835 ;
        RECT 138.555 -120.525 138.885 -120.195 ;
        RECT 138.555 -121.885 138.885 -121.555 ;
        RECT 138.555 -123.245 138.885 -122.915 ;
        RECT 138.555 -124.605 138.885 -124.275 ;
        RECT 138.555 -125.965 138.885 -125.635 ;
        RECT 138.555 -127.325 138.885 -126.995 ;
        RECT 138.555 -128.685 138.885 -128.355 ;
        RECT 138.555 -130.045 138.885 -129.715 ;
        RECT 138.555 -131.405 138.885 -131.075 ;
        RECT 138.555 -132.765 138.885 -132.435 ;
        RECT 138.555 -134.125 138.885 -133.795 ;
        RECT 138.555 -135.485 138.885 -135.155 ;
        RECT 138.555 -136.845 138.885 -136.515 ;
        RECT 138.555 -138.205 138.885 -137.875 ;
        RECT 138.555 -139.565 138.885 -139.235 ;
        RECT 138.555 -140.925 138.885 -140.595 ;
        RECT 138.555 -142.285 138.885 -141.955 ;
        RECT 138.555 -143.645 138.885 -143.315 ;
        RECT 138.555 -145.005 138.885 -144.675 ;
        RECT 138.555 -146.365 138.885 -146.035 ;
        RECT 138.555 -147.725 138.885 -147.395 ;
        RECT 138.555 -149.085 138.885 -148.755 ;
        RECT 138.555 -150.445 138.885 -150.115 ;
        RECT 138.555 -151.805 138.885 -151.475 ;
        RECT 138.555 -153.165 138.885 -152.835 ;
        RECT 138.555 -154.525 138.885 -154.195 ;
        RECT 138.555 -155.885 138.885 -155.555 ;
        RECT 138.555 -157.245 138.885 -156.915 ;
        RECT 138.555 -158.605 138.885 -158.275 ;
        RECT 138.555 -159.965 138.885 -159.635 ;
        RECT 138.555 -161.325 138.885 -160.995 ;
        RECT 138.555 -162.685 138.885 -162.355 ;
        RECT 138.555 -164.045 138.885 -163.715 ;
        RECT 138.555 -165.405 138.885 -165.075 ;
        RECT 138.555 -166.765 138.885 -166.435 ;
        RECT 138.555 -168.125 138.885 -167.795 ;
        RECT 138.555 -169.485 138.885 -169.155 ;
        RECT 138.555 -170.845 138.885 -170.515 ;
        RECT 138.555 -172.205 138.885 -171.875 ;
        RECT 138.555 -173.565 138.885 -173.235 ;
        RECT 138.555 -174.925 138.885 -174.595 ;
        RECT 138.555 -176.285 138.885 -175.955 ;
        RECT 138.555 -177.645 138.885 -177.315 ;
        RECT 138.555 -179.005 138.885 -178.675 ;
        RECT 138.555 -184.65 138.885 -183.52 ;
        RECT 138.56 -184.765 138.88 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 244.04 140.245 245.17 ;
        RECT 139.915 239.875 140.245 240.205 ;
        RECT 139.915 238.515 140.245 238.845 ;
        RECT 139.915 237.155 140.245 237.485 ;
        RECT 139.92 237.155 140.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 -0.845 140.245 -0.515 ;
        RECT 139.915 -2.205 140.245 -1.875 ;
        RECT 139.915 -3.565 140.245 -3.235 ;
        RECT 139.92 -3.565 140.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.915 -96.045 140.245 -95.715 ;
        RECT 139.915 -97.405 140.245 -97.075 ;
        RECT 139.915 -98.765 140.245 -98.435 ;
        RECT 139.915 -100.125 140.245 -99.795 ;
        RECT 139.915 -101.485 140.245 -101.155 ;
        RECT 139.915 -102.845 140.245 -102.515 ;
        RECT 139.915 -104.205 140.245 -103.875 ;
        RECT 139.915 -105.565 140.245 -105.235 ;
        RECT 139.915 -106.925 140.245 -106.595 ;
        RECT 139.915 -108.285 140.245 -107.955 ;
        RECT 139.915 -109.645 140.245 -109.315 ;
        RECT 139.915 -111.005 140.245 -110.675 ;
        RECT 139.915 -112.365 140.245 -112.035 ;
        RECT 139.915 -113.725 140.245 -113.395 ;
        RECT 139.915 -115.085 140.245 -114.755 ;
        RECT 139.915 -116.445 140.245 -116.115 ;
        RECT 139.915 -117.805 140.245 -117.475 ;
        RECT 139.915 -119.165 140.245 -118.835 ;
        RECT 139.915 -120.525 140.245 -120.195 ;
        RECT 139.915 -121.885 140.245 -121.555 ;
        RECT 139.915 -123.245 140.245 -122.915 ;
        RECT 139.915 -124.605 140.245 -124.275 ;
        RECT 139.915 -125.965 140.245 -125.635 ;
        RECT 139.915 -127.325 140.245 -126.995 ;
        RECT 139.915 -128.685 140.245 -128.355 ;
        RECT 139.915 -130.045 140.245 -129.715 ;
        RECT 139.915 -131.405 140.245 -131.075 ;
        RECT 139.915 -132.765 140.245 -132.435 ;
        RECT 139.915 -134.125 140.245 -133.795 ;
        RECT 139.915 -135.485 140.245 -135.155 ;
        RECT 139.915 -136.845 140.245 -136.515 ;
        RECT 139.915 -138.205 140.245 -137.875 ;
        RECT 139.915 -139.565 140.245 -139.235 ;
        RECT 139.915 -140.925 140.245 -140.595 ;
        RECT 139.915 -142.285 140.245 -141.955 ;
        RECT 139.915 -143.645 140.245 -143.315 ;
        RECT 139.915 -145.005 140.245 -144.675 ;
        RECT 139.915 -146.365 140.245 -146.035 ;
        RECT 139.915 -147.725 140.245 -147.395 ;
        RECT 139.915 -149.085 140.245 -148.755 ;
        RECT 139.915 -150.445 140.245 -150.115 ;
        RECT 139.915 -151.805 140.245 -151.475 ;
        RECT 139.915 -153.165 140.245 -152.835 ;
        RECT 139.915 -154.525 140.245 -154.195 ;
        RECT 139.915 -155.885 140.245 -155.555 ;
        RECT 139.915 -157.245 140.245 -156.915 ;
        RECT 139.915 -158.605 140.245 -158.275 ;
        RECT 139.915 -159.965 140.245 -159.635 ;
        RECT 139.915 -161.325 140.245 -160.995 ;
        RECT 139.915 -162.685 140.245 -162.355 ;
        RECT 139.915 -164.045 140.245 -163.715 ;
        RECT 139.915 -165.405 140.245 -165.075 ;
        RECT 139.915 -166.765 140.245 -166.435 ;
        RECT 139.915 -168.125 140.245 -167.795 ;
        RECT 139.915 -169.485 140.245 -169.155 ;
        RECT 139.915 -170.845 140.245 -170.515 ;
        RECT 139.915 -172.205 140.245 -171.875 ;
        RECT 139.915 -173.565 140.245 -173.235 ;
        RECT 139.915 -174.925 140.245 -174.595 ;
        RECT 139.915 -176.285 140.245 -175.955 ;
        RECT 139.915 -177.645 140.245 -177.315 ;
        RECT 139.915 -179.005 140.245 -178.675 ;
        RECT 139.915 -184.65 140.245 -183.52 ;
        RECT 139.92 -184.765 140.24 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 244.04 141.605 245.17 ;
        RECT 141.275 239.875 141.605 240.205 ;
        RECT 141.275 238.515 141.605 238.845 ;
        RECT 141.275 237.155 141.605 237.485 ;
        RECT 141.28 237.155 141.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 -0.845 141.605 -0.515 ;
        RECT 141.275 -2.205 141.605 -1.875 ;
        RECT 141.275 -3.565 141.605 -3.235 ;
        RECT 141.28 -3.565 141.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.275 -96.045 141.605 -95.715 ;
        RECT 141.275 -97.405 141.605 -97.075 ;
        RECT 141.275 -98.765 141.605 -98.435 ;
        RECT 141.275 -100.125 141.605 -99.795 ;
        RECT 141.275 -101.485 141.605 -101.155 ;
        RECT 141.275 -102.845 141.605 -102.515 ;
        RECT 141.275 -104.205 141.605 -103.875 ;
        RECT 141.275 -105.565 141.605 -105.235 ;
        RECT 141.275 -106.925 141.605 -106.595 ;
        RECT 141.275 -108.285 141.605 -107.955 ;
        RECT 141.275 -109.645 141.605 -109.315 ;
        RECT 141.275 -111.005 141.605 -110.675 ;
        RECT 141.275 -112.365 141.605 -112.035 ;
        RECT 141.275 -113.725 141.605 -113.395 ;
        RECT 141.275 -115.085 141.605 -114.755 ;
        RECT 141.275 -116.445 141.605 -116.115 ;
        RECT 141.275 -117.805 141.605 -117.475 ;
        RECT 141.275 -119.165 141.605 -118.835 ;
        RECT 141.275 -120.525 141.605 -120.195 ;
        RECT 141.275 -121.885 141.605 -121.555 ;
        RECT 141.275 -123.245 141.605 -122.915 ;
        RECT 141.275 -124.605 141.605 -124.275 ;
        RECT 141.275 -125.965 141.605 -125.635 ;
        RECT 141.275 -127.325 141.605 -126.995 ;
        RECT 141.275 -128.685 141.605 -128.355 ;
        RECT 141.275 -130.045 141.605 -129.715 ;
        RECT 141.275 -131.405 141.605 -131.075 ;
        RECT 141.275 -132.765 141.605 -132.435 ;
        RECT 141.275 -134.125 141.605 -133.795 ;
        RECT 141.275 -135.485 141.605 -135.155 ;
        RECT 141.275 -136.845 141.605 -136.515 ;
        RECT 141.275 -138.205 141.605 -137.875 ;
        RECT 141.275 -139.565 141.605 -139.235 ;
        RECT 141.275 -140.925 141.605 -140.595 ;
        RECT 141.275 -142.285 141.605 -141.955 ;
        RECT 141.275 -143.645 141.605 -143.315 ;
        RECT 141.275 -145.005 141.605 -144.675 ;
        RECT 141.275 -146.365 141.605 -146.035 ;
        RECT 141.275 -147.725 141.605 -147.395 ;
        RECT 141.275 -149.085 141.605 -148.755 ;
        RECT 141.275 -150.445 141.605 -150.115 ;
        RECT 141.275 -151.805 141.605 -151.475 ;
        RECT 141.275 -153.165 141.605 -152.835 ;
        RECT 141.275 -154.525 141.605 -154.195 ;
        RECT 141.275 -155.885 141.605 -155.555 ;
        RECT 141.275 -157.245 141.605 -156.915 ;
        RECT 141.275 -158.605 141.605 -158.275 ;
        RECT 141.275 -159.965 141.605 -159.635 ;
        RECT 141.275 -161.325 141.605 -160.995 ;
        RECT 141.275 -162.685 141.605 -162.355 ;
        RECT 141.275 -164.045 141.605 -163.715 ;
        RECT 141.275 -165.405 141.605 -165.075 ;
        RECT 141.275 -166.765 141.605 -166.435 ;
        RECT 141.275 -168.125 141.605 -167.795 ;
        RECT 141.275 -169.485 141.605 -169.155 ;
        RECT 141.275 -170.845 141.605 -170.515 ;
        RECT 141.275 -172.205 141.605 -171.875 ;
        RECT 141.275 -173.565 141.605 -173.235 ;
        RECT 141.275 -174.925 141.605 -174.595 ;
        RECT 141.275 -176.285 141.605 -175.955 ;
        RECT 141.275 -177.645 141.605 -177.315 ;
        RECT 141.275 -179.005 141.605 -178.675 ;
        RECT 141.275 -184.65 141.605 -183.52 ;
        RECT 141.28 -184.765 141.6 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 244.04 142.965 245.17 ;
        RECT 142.635 239.875 142.965 240.205 ;
        RECT 142.635 238.515 142.965 238.845 ;
        RECT 142.635 237.155 142.965 237.485 ;
        RECT 142.64 237.155 142.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 -0.845 142.965 -0.515 ;
        RECT 142.635 -2.205 142.965 -1.875 ;
        RECT 142.635 -3.565 142.965 -3.235 ;
        RECT 142.64 -3.565 142.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 142.635 -96.045 142.965 -95.715 ;
        RECT 142.635 -97.405 142.965 -97.075 ;
        RECT 142.635 -98.765 142.965 -98.435 ;
        RECT 142.635 -100.125 142.965 -99.795 ;
        RECT 142.635 -101.485 142.965 -101.155 ;
        RECT 142.635 -102.845 142.965 -102.515 ;
        RECT 142.635 -104.205 142.965 -103.875 ;
        RECT 142.635 -105.565 142.965 -105.235 ;
        RECT 142.635 -106.925 142.965 -106.595 ;
        RECT 142.635 -108.285 142.965 -107.955 ;
        RECT 142.635 -109.645 142.965 -109.315 ;
        RECT 142.635 -111.005 142.965 -110.675 ;
        RECT 142.635 -112.365 142.965 -112.035 ;
        RECT 142.635 -113.725 142.965 -113.395 ;
        RECT 142.635 -115.085 142.965 -114.755 ;
        RECT 142.635 -116.445 142.965 -116.115 ;
        RECT 142.635 -117.805 142.965 -117.475 ;
        RECT 142.635 -119.165 142.965 -118.835 ;
        RECT 142.635 -120.525 142.965 -120.195 ;
        RECT 142.635 -121.885 142.965 -121.555 ;
        RECT 142.635 -123.245 142.965 -122.915 ;
        RECT 142.635 -124.605 142.965 -124.275 ;
        RECT 142.635 -125.965 142.965 -125.635 ;
        RECT 142.635 -127.325 142.965 -126.995 ;
        RECT 142.635 -128.685 142.965 -128.355 ;
        RECT 142.635 -130.045 142.965 -129.715 ;
        RECT 142.635 -131.405 142.965 -131.075 ;
        RECT 142.635 -132.765 142.965 -132.435 ;
        RECT 142.635 -134.125 142.965 -133.795 ;
        RECT 142.635 -135.485 142.965 -135.155 ;
        RECT 142.635 -136.845 142.965 -136.515 ;
        RECT 142.635 -138.205 142.965 -137.875 ;
        RECT 142.635 -139.565 142.965 -139.235 ;
        RECT 142.635 -140.925 142.965 -140.595 ;
        RECT 142.635 -142.285 142.965 -141.955 ;
        RECT 142.635 -143.645 142.965 -143.315 ;
        RECT 142.635 -145.005 142.965 -144.675 ;
        RECT 142.635 -146.365 142.965 -146.035 ;
        RECT 142.635 -147.725 142.965 -147.395 ;
        RECT 142.635 -149.085 142.965 -148.755 ;
        RECT 142.635 -150.445 142.965 -150.115 ;
        RECT 142.635 -151.805 142.965 -151.475 ;
        RECT 142.635 -153.165 142.965 -152.835 ;
        RECT 142.635 -154.525 142.965 -154.195 ;
        RECT 142.635 -155.885 142.965 -155.555 ;
        RECT 142.635 -157.245 142.965 -156.915 ;
        RECT 142.635 -158.605 142.965 -158.275 ;
        RECT 142.635 -159.965 142.965 -159.635 ;
        RECT 142.635 -161.325 142.965 -160.995 ;
        RECT 142.635 -162.685 142.965 -162.355 ;
        RECT 142.635 -164.045 142.965 -163.715 ;
        RECT 142.635 -165.405 142.965 -165.075 ;
        RECT 142.635 -166.765 142.965 -166.435 ;
        RECT 142.635 -168.125 142.965 -167.795 ;
        RECT 142.635 -169.485 142.965 -169.155 ;
        RECT 142.635 -170.845 142.965 -170.515 ;
        RECT 142.635 -172.205 142.965 -171.875 ;
        RECT 142.635 -173.565 142.965 -173.235 ;
        RECT 142.635 -174.925 142.965 -174.595 ;
        RECT 142.635 -176.285 142.965 -175.955 ;
        RECT 142.635 -177.645 142.965 -177.315 ;
        RECT 142.635 -179.005 142.965 -178.675 ;
        RECT 142.635 -184.65 142.965 -183.52 ;
        RECT 142.64 -184.765 142.96 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.995 244.04 144.325 245.17 ;
        RECT 143.995 239.875 144.325 240.205 ;
        RECT 143.995 238.515 144.325 238.845 ;
        RECT 143.995 237.155 144.325 237.485 ;
        RECT 144 237.155 144.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.995 -98.765 144.325 -98.435 ;
        RECT 143.995 -100.125 144.325 -99.795 ;
        RECT 143.995 -101.485 144.325 -101.155 ;
        RECT 143.995 -102.845 144.325 -102.515 ;
        RECT 143.995 -104.205 144.325 -103.875 ;
        RECT 143.995 -105.565 144.325 -105.235 ;
        RECT 143.995 -106.925 144.325 -106.595 ;
        RECT 143.995 -108.285 144.325 -107.955 ;
        RECT 143.995 -109.645 144.325 -109.315 ;
        RECT 143.995 -111.005 144.325 -110.675 ;
        RECT 143.995 -112.365 144.325 -112.035 ;
        RECT 143.995 -113.725 144.325 -113.395 ;
        RECT 143.995 -115.085 144.325 -114.755 ;
        RECT 143.995 -116.445 144.325 -116.115 ;
        RECT 143.995 -117.805 144.325 -117.475 ;
        RECT 143.995 -119.165 144.325 -118.835 ;
        RECT 143.995 -120.525 144.325 -120.195 ;
        RECT 143.995 -121.885 144.325 -121.555 ;
        RECT 143.995 -123.245 144.325 -122.915 ;
        RECT 143.995 -124.605 144.325 -124.275 ;
        RECT 143.995 -125.965 144.325 -125.635 ;
        RECT 143.995 -127.325 144.325 -126.995 ;
        RECT 143.995 -128.685 144.325 -128.355 ;
        RECT 143.995 -130.045 144.325 -129.715 ;
        RECT 143.995 -131.405 144.325 -131.075 ;
        RECT 143.995 -132.765 144.325 -132.435 ;
        RECT 143.995 -134.125 144.325 -133.795 ;
        RECT 143.995 -135.485 144.325 -135.155 ;
        RECT 143.995 -136.845 144.325 -136.515 ;
        RECT 143.995 -138.205 144.325 -137.875 ;
        RECT 143.995 -139.565 144.325 -139.235 ;
        RECT 143.995 -140.925 144.325 -140.595 ;
        RECT 143.995 -142.285 144.325 -141.955 ;
        RECT 143.995 -143.645 144.325 -143.315 ;
        RECT 143.995 -145.005 144.325 -144.675 ;
        RECT 143.995 -146.365 144.325 -146.035 ;
        RECT 143.995 -147.725 144.325 -147.395 ;
        RECT 143.995 -149.085 144.325 -148.755 ;
        RECT 143.995 -150.445 144.325 -150.115 ;
        RECT 143.995 -151.805 144.325 -151.475 ;
        RECT 143.995 -153.165 144.325 -152.835 ;
        RECT 143.995 -154.525 144.325 -154.195 ;
        RECT 143.995 -155.885 144.325 -155.555 ;
        RECT 143.995 -157.245 144.325 -156.915 ;
        RECT 143.995 -158.605 144.325 -158.275 ;
        RECT 143.995 -159.965 144.325 -159.635 ;
        RECT 143.995 -161.325 144.325 -160.995 ;
        RECT 143.995 -162.685 144.325 -162.355 ;
        RECT 143.995 -164.045 144.325 -163.715 ;
        RECT 143.995 -165.405 144.325 -165.075 ;
        RECT 143.995 -166.765 144.325 -166.435 ;
        RECT 143.995 -168.125 144.325 -167.795 ;
        RECT 143.995 -169.485 144.325 -169.155 ;
        RECT 143.995 -170.845 144.325 -170.515 ;
        RECT 143.995 -172.205 144.325 -171.875 ;
        RECT 143.995 -173.565 144.325 -173.235 ;
        RECT 143.995 -174.925 144.325 -174.595 ;
        RECT 143.995 -176.285 144.325 -175.955 ;
        RECT 143.995 -177.645 144.325 -177.315 ;
        RECT 143.995 -179.005 144.325 -178.675 ;
        RECT 143.995 -184.65 144.325 -183.52 ;
        RECT 144 -184.765 144.32 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.36 -98.075 144.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.355 244.04 145.685 245.17 ;
        RECT 145.355 239.875 145.685 240.205 ;
        RECT 145.355 238.515 145.685 238.845 ;
        RECT 145.355 237.155 145.685 237.485 ;
        RECT 145.36 237.155 145.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 244.04 147.045 245.17 ;
        RECT 146.715 239.875 147.045 240.205 ;
        RECT 146.715 238.515 147.045 238.845 ;
        RECT 146.715 237.155 147.045 237.485 ;
        RECT 146.72 237.155 147.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.715 -0.845 147.045 -0.515 ;
        RECT 146.715 -2.205 147.045 -1.875 ;
        RECT 146.715 -3.565 147.045 -3.235 ;
        RECT 146.72 -3.565 147.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 244.04 148.405 245.17 ;
        RECT 148.075 239.875 148.405 240.205 ;
        RECT 148.075 238.515 148.405 238.845 ;
        RECT 148.075 237.155 148.405 237.485 ;
        RECT 148.08 237.155 148.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 -0.845 148.405 -0.515 ;
        RECT 148.075 -2.205 148.405 -1.875 ;
        RECT 148.075 -3.565 148.405 -3.235 ;
        RECT 148.08 -3.565 148.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.075 -96.045 148.405 -95.715 ;
        RECT 148.075 -97.405 148.405 -97.075 ;
        RECT 148.075 -98.765 148.405 -98.435 ;
        RECT 148.075 -100.125 148.405 -99.795 ;
        RECT 148.075 -101.485 148.405 -101.155 ;
        RECT 148.075 -102.845 148.405 -102.515 ;
        RECT 148.075 -104.205 148.405 -103.875 ;
        RECT 148.075 -105.565 148.405 -105.235 ;
        RECT 148.075 -106.925 148.405 -106.595 ;
        RECT 148.075 -108.285 148.405 -107.955 ;
        RECT 148.075 -109.645 148.405 -109.315 ;
        RECT 148.075 -111.005 148.405 -110.675 ;
        RECT 148.075 -112.365 148.405 -112.035 ;
        RECT 148.075 -113.725 148.405 -113.395 ;
        RECT 148.075 -115.085 148.405 -114.755 ;
        RECT 148.075 -116.445 148.405 -116.115 ;
        RECT 148.075 -117.805 148.405 -117.475 ;
        RECT 148.075 -119.165 148.405 -118.835 ;
        RECT 148.075 -120.525 148.405 -120.195 ;
        RECT 148.075 -121.885 148.405 -121.555 ;
        RECT 148.075 -123.245 148.405 -122.915 ;
        RECT 148.075 -124.605 148.405 -124.275 ;
        RECT 148.075 -125.965 148.405 -125.635 ;
        RECT 148.075 -127.325 148.405 -126.995 ;
        RECT 148.075 -128.685 148.405 -128.355 ;
        RECT 148.075 -130.045 148.405 -129.715 ;
        RECT 148.075 -131.405 148.405 -131.075 ;
        RECT 148.075 -132.765 148.405 -132.435 ;
        RECT 148.075 -134.125 148.405 -133.795 ;
        RECT 148.075 -135.485 148.405 -135.155 ;
        RECT 148.075 -136.845 148.405 -136.515 ;
        RECT 148.075 -138.205 148.405 -137.875 ;
        RECT 148.075 -139.565 148.405 -139.235 ;
        RECT 148.075 -140.925 148.405 -140.595 ;
        RECT 148.075 -142.285 148.405 -141.955 ;
        RECT 148.075 -143.645 148.405 -143.315 ;
        RECT 148.075 -145.005 148.405 -144.675 ;
        RECT 148.075 -146.365 148.405 -146.035 ;
        RECT 148.075 -147.725 148.405 -147.395 ;
        RECT 148.075 -149.085 148.405 -148.755 ;
        RECT 148.075 -150.445 148.405 -150.115 ;
        RECT 148.075 -151.805 148.405 -151.475 ;
        RECT 148.075 -153.165 148.405 -152.835 ;
        RECT 148.075 -154.525 148.405 -154.195 ;
        RECT 148.075 -155.885 148.405 -155.555 ;
        RECT 148.075 -157.245 148.405 -156.915 ;
        RECT 148.075 -158.605 148.405 -158.275 ;
        RECT 148.075 -159.965 148.405 -159.635 ;
        RECT 148.075 -161.325 148.405 -160.995 ;
        RECT 148.075 -162.685 148.405 -162.355 ;
        RECT 148.075 -164.045 148.405 -163.715 ;
        RECT 148.075 -165.405 148.405 -165.075 ;
        RECT 148.075 -166.765 148.405 -166.435 ;
        RECT 148.075 -168.125 148.405 -167.795 ;
        RECT 148.075 -169.485 148.405 -169.155 ;
        RECT 148.075 -170.845 148.405 -170.515 ;
        RECT 148.075 -172.205 148.405 -171.875 ;
        RECT 148.075 -173.565 148.405 -173.235 ;
        RECT 148.075 -174.925 148.405 -174.595 ;
        RECT 148.075 -176.285 148.405 -175.955 ;
        RECT 148.075 -177.645 148.405 -177.315 ;
        RECT 148.075 -179.005 148.405 -178.675 ;
        RECT 148.075 -184.65 148.405 -183.52 ;
        RECT 148.08 -184.765 148.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 244.04 149.765 245.17 ;
        RECT 149.435 239.875 149.765 240.205 ;
        RECT 149.435 238.515 149.765 238.845 ;
        RECT 149.435 237.155 149.765 237.485 ;
        RECT 149.44 237.155 149.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 -0.845 149.765 -0.515 ;
        RECT 149.435 -2.205 149.765 -1.875 ;
        RECT 149.435 -3.565 149.765 -3.235 ;
        RECT 149.44 -3.565 149.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 149.435 -96.045 149.765 -95.715 ;
        RECT 149.435 -97.405 149.765 -97.075 ;
        RECT 149.435 -98.765 149.765 -98.435 ;
        RECT 149.435 -100.125 149.765 -99.795 ;
        RECT 149.435 -101.485 149.765 -101.155 ;
        RECT 149.435 -102.845 149.765 -102.515 ;
        RECT 149.435 -104.205 149.765 -103.875 ;
        RECT 149.435 -105.565 149.765 -105.235 ;
        RECT 149.435 -106.925 149.765 -106.595 ;
        RECT 149.435 -108.285 149.765 -107.955 ;
        RECT 149.435 -109.645 149.765 -109.315 ;
        RECT 149.435 -111.005 149.765 -110.675 ;
        RECT 149.435 -112.365 149.765 -112.035 ;
        RECT 149.435 -113.725 149.765 -113.395 ;
        RECT 149.435 -115.085 149.765 -114.755 ;
        RECT 149.435 -116.445 149.765 -116.115 ;
        RECT 149.435 -117.805 149.765 -117.475 ;
        RECT 149.435 -119.165 149.765 -118.835 ;
        RECT 149.435 -120.525 149.765 -120.195 ;
        RECT 149.435 -121.885 149.765 -121.555 ;
        RECT 149.435 -123.245 149.765 -122.915 ;
        RECT 149.435 -124.605 149.765 -124.275 ;
        RECT 149.435 -125.965 149.765 -125.635 ;
        RECT 149.435 -127.325 149.765 -126.995 ;
        RECT 149.435 -128.685 149.765 -128.355 ;
        RECT 149.435 -130.045 149.765 -129.715 ;
        RECT 149.435 -131.405 149.765 -131.075 ;
        RECT 149.435 -132.765 149.765 -132.435 ;
        RECT 149.435 -134.125 149.765 -133.795 ;
        RECT 149.435 -135.485 149.765 -135.155 ;
        RECT 149.435 -136.845 149.765 -136.515 ;
        RECT 149.435 -138.205 149.765 -137.875 ;
        RECT 149.435 -139.565 149.765 -139.235 ;
        RECT 149.435 -140.925 149.765 -140.595 ;
        RECT 149.435 -142.285 149.765 -141.955 ;
        RECT 149.435 -143.645 149.765 -143.315 ;
        RECT 149.435 -145.005 149.765 -144.675 ;
        RECT 149.435 -146.365 149.765 -146.035 ;
        RECT 149.435 -147.725 149.765 -147.395 ;
        RECT 149.435 -149.085 149.765 -148.755 ;
        RECT 149.435 -150.445 149.765 -150.115 ;
        RECT 149.435 -151.805 149.765 -151.475 ;
        RECT 149.435 -153.165 149.765 -152.835 ;
        RECT 149.435 -154.525 149.765 -154.195 ;
        RECT 149.435 -155.885 149.765 -155.555 ;
        RECT 149.435 -157.245 149.765 -156.915 ;
        RECT 149.435 -158.605 149.765 -158.275 ;
        RECT 149.435 -159.965 149.765 -159.635 ;
        RECT 149.435 -161.325 149.765 -160.995 ;
        RECT 149.435 -162.685 149.765 -162.355 ;
        RECT 149.435 -164.045 149.765 -163.715 ;
        RECT 149.435 -165.405 149.765 -165.075 ;
        RECT 149.435 -166.765 149.765 -166.435 ;
        RECT 149.435 -168.125 149.765 -167.795 ;
        RECT 149.435 -169.485 149.765 -169.155 ;
        RECT 149.435 -170.845 149.765 -170.515 ;
        RECT 149.435 -172.205 149.765 -171.875 ;
        RECT 149.435 -173.565 149.765 -173.235 ;
        RECT 149.435 -174.925 149.765 -174.595 ;
        RECT 149.435 -176.285 149.765 -175.955 ;
        RECT 149.435 -177.645 149.765 -177.315 ;
        RECT 149.435 -179.005 149.765 -178.675 ;
        RECT 149.435 -184.65 149.765 -183.52 ;
        RECT 149.44 -184.765 149.76 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 244.04 151.125 245.17 ;
        RECT 150.795 239.875 151.125 240.205 ;
        RECT 150.795 238.515 151.125 238.845 ;
        RECT 150.795 237.155 151.125 237.485 ;
        RECT 150.8 237.155 151.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 -0.845 151.125 -0.515 ;
        RECT 150.795 -2.205 151.125 -1.875 ;
        RECT 150.795 -3.565 151.125 -3.235 ;
        RECT 150.8 -3.565 151.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.795 -96.045 151.125 -95.715 ;
        RECT 150.795 -97.405 151.125 -97.075 ;
        RECT 150.795 -98.765 151.125 -98.435 ;
        RECT 150.795 -100.125 151.125 -99.795 ;
        RECT 150.795 -101.485 151.125 -101.155 ;
        RECT 150.795 -102.845 151.125 -102.515 ;
        RECT 150.795 -104.205 151.125 -103.875 ;
        RECT 150.795 -105.565 151.125 -105.235 ;
        RECT 150.795 -106.925 151.125 -106.595 ;
        RECT 150.795 -108.285 151.125 -107.955 ;
        RECT 150.795 -109.645 151.125 -109.315 ;
        RECT 150.795 -111.005 151.125 -110.675 ;
        RECT 150.795 -112.365 151.125 -112.035 ;
        RECT 150.795 -113.725 151.125 -113.395 ;
        RECT 150.795 -115.085 151.125 -114.755 ;
        RECT 150.795 -116.445 151.125 -116.115 ;
        RECT 150.795 -117.805 151.125 -117.475 ;
        RECT 150.795 -119.165 151.125 -118.835 ;
        RECT 150.795 -120.525 151.125 -120.195 ;
        RECT 150.795 -121.885 151.125 -121.555 ;
        RECT 150.795 -123.245 151.125 -122.915 ;
        RECT 150.795 -124.605 151.125 -124.275 ;
        RECT 150.795 -125.965 151.125 -125.635 ;
        RECT 150.795 -127.325 151.125 -126.995 ;
        RECT 150.795 -128.685 151.125 -128.355 ;
        RECT 150.795 -130.045 151.125 -129.715 ;
        RECT 150.795 -131.405 151.125 -131.075 ;
        RECT 150.795 -132.765 151.125 -132.435 ;
        RECT 150.795 -134.125 151.125 -133.795 ;
        RECT 150.795 -135.485 151.125 -135.155 ;
        RECT 150.795 -136.845 151.125 -136.515 ;
        RECT 150.795 -138.205 151.125 -137.875 ;
        RECT 150.795 -139.565 151.125 -139.235 ;
        RECT 150.795 -140.925 151.125 -140.595 ;
        RECT 150.795 -142.285 151.125 -141.955 ;
        RECT 150.795 -143.645 151.125 -143.315 ;
        RECT 150.795 -145.005 151.125 -144.675 ;
        RECT 150.795 -146.365 151.125 -146.035 ;
        RECT 150.795 -147.725 151.125 -147.395 ;
        RECT 150.795 -149.085 151.125 -148.755 ;
        RECT 150.795 -150.445 151.125 -150.115 ;
        RECT 150.795 -151.805 151.125 -151.475 ;
        RECT 150.795 -153.165 151.125 -152.835 ;
        RECT 150.795 -154.525 151.125 -154.195 ;
        RECT 150.795 -155.885 151.125 -155.555 ;
        RECT 150.795 -157.245 151.125 -156.915 ;
        RECT 150.795 -158.605 151.125 -158.275 ;
        RECT 150.795 -159.965 151.125 -159.635 ;
        RECT 150.795 -161.325 151.125 -160.995 ;
        RECT 150.795 -162.685 151.125 -162.355 ;
        RECT 150.795 -164.045 151.125 -163.715 ;
        RECT 150.795 -165.405 151.125 -165.075 ;
        RECT 150.795 -166.765 151.125 -166.435 ;
        RECT 150.795 -168.125 151.125 -167.795 ;
        RECT 150.795 -169.485 151.125 -169.155 ;
        RECT 150.795 -170.845 151.125 -170.515 ;
        RECT 150.795 -172.205 151.125 -171.875 ;
        RECT 150.795 -173.565 151.125 -173.235 ;
        RECT 150.795 -174.925 151.125 -174.595 ;
        RECT 150.795 -176.285 151.125 -175.955 ;
        RECT 150.795 -177.645 151.125 -177.315 ;
        RECT 150.795 -179.005 151.125 -178.675 ;
        RECT 150.795 -184.65 151.125 -183.52 ;
        RECT 150.8 -184.765 151.12 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 244.04 152.485 245.17 ;
        RECT 152.155 239.875 152.485 240.205 ;
        RECT 152.155 238.515 152.485 238.845 ;
        RECT 152.155 237.155 152.485 237.485 ;
        RECT 152.16 237.155 152.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 -0.845 152.485 -0.515 ;
        RECT 152.155 -2.205 152.485 -1.875 ;
        RECT 152.155 -3.565 152.485 -3.235 ;
        RECT 152.16 -3.565 152.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.155 -96.045 152.485 -95.715 ;
        RECT 152.155 -97.405 152.485 -97.075 ;
        RECT 152.155 -98.765 152.485 -98.435 ;
        RECT 152.155 -100.125 152.485 -99.795 ;
        RECT 152.155 -101.485 152.485 -101.155 ;
        RECT 152.155 -102.845 152.485 -102.515 ;
        RECT 152.155 -104.205 152.485 -103.875 ;
        RECT 152.155 -105.565 152.485 -105.235 ;
        RECT 152.155 -106.925 152.485 -106.595 ;
        RECT 152.155 -108.285 152.485 -107.955 ;
        RECT 152.155 -109.645 152.485 -109.315 ;
        RECT 152.155 -111.005 152.485 -110.675 ;
        RECT 152.155 -112.365 152.485 -112.035 ;
        RECT 152.155 -113.725 152.485 -113.395 ;
        RECT 152.155 -115.085 152.485 -114.755 ;
        RECT 152.155 -116.445 152.485 -116.115 ;
        RECT 152.155 -117.805 152.485 -117.475 ;
        RECT 152.155 -119.165 152.485 -118.835 ;
        RECT 152.155 -120.525 152.485 -120.195 ;
        RECT 152.155 -121.885 152.485 -121.555 ;
        RECT 152.155 -123.245 152.485 -122.915 ;
        RECT 152.155 -124.605 152.485 -124.275 ;
        RECT 152.155 -125.965 152.485 -125.635 ;
        RECT 152.155 -127.325 152.485 -126.995 ;
        RECT 152.155 -128.685 152.485 -128.355 ;
        RECT 152.155 -130.045 152.485 -129.715 ;
        RECT 152.155 -131.405 152.485 -131.075 ;
        RECT 152.155 -132.765 152.485 -132.435 ;
        RECT 152.155 -134.125 152.485 -133.795 ;
        RECT 152.155 -135.485 152.485 -135.155 ;
        RECT 152.155 -136.845 152.485 -136.515 ;
        RECT 152.155 -138.205 152.485 -137.875 ;
        RECT 152.155 -139.565 152.485 -139.235 ;
        RECT 152.155 -140.925 152.485 -140.595 ;
        RECT 152.155 -142.285 152.485 -141.955 ;
        RECT 152.155 -143.645 152.485 -143.315 ;
        RECT 152.155 -145.005 152.485 -144.675 ;
        RECT 152.155 -146.365 152.485 -146.035 ;
        RECT 152.155 -147.725 152.485 -147.395 ;
        RECT 152.155 -149.085 152.485 -148.755 ;
        RECT 152.155 -150.445 152.485 -150.115 ;
        RECT 152.155 -151.805 152.485 -151.475 ;
        RECT 152.155 -153.165 152.485 -152.835 ;
        RECT 152.155 -154.525 152.485 -154.195 ;
        RECT 152.155 -155.885 152.485 -155.555 ;
        RECT 152.155 -157.245 152.485 -156.915 ;
        RECT 152.155 -158.605 152.485 -158.275 ;
        RECT 152.155 -159.965 152.485 -159.635 ;
        RECT 152.155 -161.325 152.485 -160.995 ;
        RECT 152.155 -162.685 152.485 -162.355 ;
        RECT 152.155 -164.045 152.485 -163.715 ;
        RECT 152.155 -165.405 152.485 -165.075 ;
        RECT 152.155 -166.765 152.485 -166.435 ;
        RECT 152.155 -168.125 152.485 -167.795 ;
        RECT 152.155 -169.485 152.485 -169.155 ;
        RECT 152.155 -170.845 152.485 -170.515 ;
        RECT 152.155 -172.205 152.485 -171.875 ;
        RECT 152.155 -173.565 152.485 -173.235 ;
        RECT 152.155 -174.925 152.485 -174.595 ;
        RECT 152.155 -176.285 152.485 -175.955 ;
        RECT 152.155 -177.645 152.485 -177.315 ;
        RECT 152.155 -179.005 152.485 -178.675 ;
        RECT 152.155 -184.65 152.485 -183.52 ;
        RECT 152.16 -184.765 152.48 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 244.04 153.845 245.17 ;
        RECT 153.515 239.875 153.845 240.205 ;
        RECT 153.515 238.515 153.845 238.845 ;
        RECT 153.515 237.155 153.845 237.485 ;
        RECT 153.52 237.155 153.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 -0.845 153.845 -0.515 ;
        RECT 153.515 -2.205 153.845 -1.875 ;
        RECT 153.515 -3.565 153.845 -3.235 ;
        RECT 153.52 -3.565 153.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 153.515 -96.045 153.845 -95.715 ;
        RECT 153.515 -97.405 153.845 -97.075 ;
        RECT 153.515 -98.765 153.845 -98.435 ;
        RECT 153.515 -100.125 153.845 -99.795 ;
        RECT 153.515 -101.485 153.845 -101.155 ;
        RECT 153.515 -102.845 153.845 -102.515 ;
        RECT 153.515 -104.205 153.845 -103.875 ;
        RECT 153.515 -105.565 153.845 -105.235 ;
        RECT 153.515 -106.925 153.845 -106.595 ;
        RECT 153.515 -108.285 153.845 -107.955 ;
        RECT 153.515 -109.645 153.845 -109.315 ;
        RECT 153.515 -111.005 153.845 -110.675 ;
        RECT 153.515 -112.365 153.845 -112.035 ;
        RECT 153.515 -113.725 153.845 -113.395 ;
        RECT 153.515 -115.085 153.845 -114.755 ;
        RECT 153.515 -116.445 153.845 -116.115 ;
        RECT 153.515 -117.805 153.845 -117.475 ;
        RECT 153.515 -119.165 153.845 -118.835 ;
        RECT 153.515 -120.525 153.845 -120.195 ;
        RECT 153.515 -121.885 153.845 -121.555 ;
        RECT 153.515 -123.245 153.845 -122.915 ;
        RECT 153.515 -124.605 153.845 -124.275 ;
        RECT 153.515 -125.965 153.845 -125.635 ;
        RECT 153.515 -127.325 153.845 -126.995 ;
        RECT 153.515 -128.685 153.845 -128.355 ;
        RECT 153.515 -130.045 153.845 -129.715 ;
        RECT 153.515 -131.405 153.845 -131.075 ;
        RECT 153.515 -132.765 153.845 -132.435 ;
        RECT 153.515 -134.125 153.845 -133.795 ;
        RECT 153.515 -135.485 153.845 -135.155 ;
        RECT 153.515 -136.845 153.845 -136.515 ;
        RECT 153.515 -138.205 153.845 -137.875 ;
        RECT 153.515 -139.565 153.845 -139.235 ;
        RECT 153.515 -140.925 153.845 -140.595 ;
        RECT 153.515 -142.285 153.845 -141.955 ;
        RECT 153.515 -143.645 153.845 -143.315 ;
        RECT 153.515 -145.005 153.845 -144.675 ;
        RECT 153.515 -146.365 153.845 -146.035 ;
        RECT 153.515 -147.725 153.845 -147.395 ;
        RECT 153.515 -149.085 153.845 -148.755 ;
        RECT 153.515 -150.445 153.845 -150.115 ;
        RECT 153.515 -151.805 153.845 -151.475 ;
        RECT 153.515 -153.165 153.845 -152.835 ;
        RECT 153.515 -154.525 153.845 -154.195 ;
        RECT 153.515 -155.885 153.845 -155.555 ;
        RECT 153.515 -157.245 153.845 -156.915 ;
        RECT 153.515 -158.605 153.845 -158.275 ;
        RECT 153.515 -159.965 153.845 -159.635 ;
        RECT 153.515 -161.325 153.845 -160.995 ;
        RECT 153.515 -162.685 153.845 -162.355 ;
        RECT 153.515 -164.045 153.845 -163.715 ;
        RECT 153.515 -165.405 153.845 -165.075 ;
        RECT 153.515 -166.765 153.845 -166.435 ;
        RECT 153.515 -168.125 153.845 -167.795 ;
        RECT 153.515 -169.485 153.845 -169.155 ;
        RECT 153.515 -170.845 153.845 -170.515 ;
        RECT 153.515 -172.205 153.845 -171.875 ;
        RECT 153.515 -173.565 153.845 -173.235 ;
        RECT 153.515 -174.925 153.845 -174.595 ;
        RECT 153.515 -176.285 153.845 -175.955 ;
        RECT 153.515 -177.645 153.845 -177.315 ;
        RECT 153.515 -179.005 153.845 -178.675 ;
        RECT 153.515 -184.65 153.845 -183.52 ;
        RECT 153.52 -184.765 153.84 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 244.04 155.205 245.17 ;
        RECT 154.875 239.875 155.205 240.205 ;
        RECT 154.875 238.515 155.205 238.845 ;
        RECT 154.875 237.155 155.205 237.485 ;
        RECT 154.88 237.155 155.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.875 -98.765 155.205 -98.435 ;
        RECT 154.875 -100.125 155.205 -99.795 ;
        RECT 154.875 -101.485 155.205 -101.155 ;
        RECT 154.875 -102.845 155.205 -102.515 ;
        RECT 154.875 -104.205 155.205 -103.875 ;
        RECT 154.875 -105.565 155.205 -105.235 ;
        RECT 154.875 -106.925 155.205 -106.595 ;
        RECT 154.875 -108.285 155.205 -107.955 ;
        RECT 154.875 -109.645 155.205 -109.315 ;
        RECT 154.875 -111.005 155.205 -110.675 ;
        RECT 154.875 -112.365 155.205 -112.035 ;
        RECT 154.875 -113.725 155.205 -113.395 ;
        RECT 154.875 -115.085 155.205 -114.755 ;
        RECT 154.875 -116.445 155.205 -116.115 ;
        RECT 154.875 -117.805 155.205 -117.475 ;
        RECT 154.875 -119.165 155.205 -118.835 ;
        RECT 154.875 -120.525 155.205 -120.195 ;
        RECT 154.875 -121.885 155.205 -121.555 ;
        RECT 154.875 -123.245 155.205 -122.915 ;
        RECT 154.875 -124.605 155.205 -124.275 ;
        RECT 154.875 -125.965 155.205 -125.635 ;
        RECT 154.875 -127.325 155.205 -126.995 ;
        RECT 154.875 -128.685 155.205 -128.355 ;
        RECT 154.875 -130.045 155.205 -129.715 ;
        RECT 154.875 -131.405 155.205 -131.075 ;
        RECT 154.875 -132.765 155.205 -132.435 ;
        RECT 154.875 -134.125 155.205 -133.795 ;
        RECT 154.875 -135.485 155.205 -135.155 ;
        RECT 154.875 -136.845 155.205 -136.515 ;
        RECT 154.875 -138.205 155.205 -137.875 ;
        RECT 154.875 -139.565 155.205 -139.235 ;
        RECT 154.875 -140.925 155.205 -140.595 ;
        RECT 154.875 -142.285 155.205 -141.955 ;
        RECT 154.875 -143.645 155.205 -143.315 ;
        RECT 154.875 -145.005 155.205 -144.675 ;
        RECT 154.875 -146.365 155.205 -146.035 ;
        RECT 154.875 -147.725 155.205 -147.395 ;
        RECT 154.875 -149.085 155.205 -148.755 ;
        RECT 154.875 -150.445 155.205 -150.115 ;
        RECT 154.875 -151.805 155.205 -151.475 ;
        RECT 154.875 -153.165 155.205 -152.835 ;
        RECT 154.875 -154.525 155.205 -154.195 ;
        RECT 154.875 -155.885 155.205 -155.555 ;
        RECT 154.875 -157.245 155.205 -156.915 ;
        RECT 154.875 -158.605 155.205 -158.275 ;
        RECT 154.875 -159.965 155.205 -159.635 ;
        RECT 154.875 -161.325 155.205 -160.995 ;
        RECT 154.875 -162.685 155.205 -162.355 ;
        RECT 154.875 -164.045 155.205 -163.715 ;
        RECT 154.875 -165.405 155.205 -165.075 ;
        RECT 154.875 -166.765 155.205 -166.435 ;
        RECT 154.875 -168.125 155.205 -167.795 ;
        RECT 154.875 -169.485 155.205 -169.155 ;
        RECT 154.875 -170.845 155.205 -170.515 ;
        RECT 154.875 -172.205 155.205 -171.875 ;
        RECT 154.875 -173.565 155.205 -173.235 ;
        RECT 154.875 -174.925 155.205 -174.595 ;
        RECT 154.875 -176.285 155.205 -175.955 ;
        RECT 154.875 -177.645 155.205 -177.315 ;
        RECT 154.875 -179.005 155.205 -178.675 ;
        RECT 154.875 -184.65 155.205 -183.52 ;
        RECT 154.88 -184.765 155.2 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.26 -98.075 155.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.235 244.04 156.565 245.17 ;
        RECT 156.235 239.875 156.565 240.205 ;
        RECT 156.235 238.515 156.565 238.845 ;
        RECT 156.235 237.155 156.565 237.485 ;
        RECT 156.24 237.155 156.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 244.04 157.925 245.17 ;
        RECT 157.595 239.875 157.925 240.205 ;
        RECT 157.595 238.515 157.925 238.845 ;
        RECT 157.595 237.155 157.925 237.485 ;
        RECT 157.6 237.155 157.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 157.595 -0.845 157.925 -0.515 ;
        RECT 157.595 -2.205 157.925 -1.875 ;
        RECT 157.595 -3.565 157.925 -3.235 ;
        RECT 157.6 -3.565 157.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 244.04 159.285 245.17 ;
        RECT 158.955 239.875 159.285 240.205 ;
        RECT 158.955 238.515 159.285 238.845 ;
        RECT 158.955 237.155 159.285 237.485 ;
        RECT 158.96 237.155 159.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 -0.845 159.285 -0.515 ;
        RECT 158.955 -2.205 159.285 -1.875 ;
        RECT 158.955 -3.565 159.285 -3.235 ;
        RECT 158.96 -3.565 159.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.955 -155.885 159.285 -155.555 ;
        RECT 158.955 -157.245 159.285 -156.915 ;
        RECT 158.955 -158.605 159.285 -158.275 ;
        RECT 158.955 -159.965 159.285 -159.635 ;
        RECT 158.955 -161.325 159.285 -160.995 ;
        RECT 158.955 -162.685 159.285 -162.355 ;
        RECT 158.955 -164.045 159.285 -163.715 ;
        RECT 158.955 -165.405 159.285 -165.075 ;
        RECT 158.955 -166.765 159.285 -166.435 ;
        RECT 158.955 -168.125 159.285 -167.795 ;
        RECT 158.955 -169.485 159.285 -169.155 ;
        RECT 158.955 -170.845 159.285 -170.515 ;
        RECT 158.955 -172.205 159.285 -171.875 ;
        RECT 158.955 -173.565 159.285 -173.235 ;
        RECT 158.955 -174.925 159.285 -174.595 ;
        RECT 158.955 -176.285 159.285 -175.955 ;
        RECT 158.955 -177.645 159.285 -177.315 ;
        RECT 158.955 -179.005 159.285 -178.675 ;
        RECT 158.955 -184.65 159.285 -183.52 ;
        RECT 158.96 -184.765 159.28 -95.04 ;
        RECT 158.955 -96.045 159.285 -95.715 ;
        RECT 158.955 -97.405 159.285 -97.075 ;
        RECT 158.955 -98.765 159.285 -98.435 ;
        RECT 158.955 -100.125 159.285 -99.795 ;
        RECT 158.955 -101.485 159.285 -101.155 ;
        RECT 158.955 -102.845 159.285 -102.515 ;
        RECT 158.955 -104.205 159.285 -103.875 ;
        RECT 158.955 -105.565 159.285 -105.235 ;
        RECT 158.955 -106.925 159.285 -106.595 ;
        RECT 158.955 -108.285 159.285 -107.955 ;
        RECT 158.955 -109.645 159.285 -109.315 ;
        RECT 158.955 -111.005 159.285 -110.675 ;
        RECT 158.955 -112.365 159.285 -112.035 ;
        RECT 158.955 -113.725 159.285 -113.395 ;
        RECT 158.955 -115.085 159.285 -114.755 ;
        RECT 158.955 -116.445 159.285 -116.115 ;
        RECT 158.955 -117.805 159.285 -117.475 ;
        RECT 158.955 -119.165 159.285 -118.835 ;
        RECT 158.955 -120.525 159.285 -120.195 ;
        RECT 158.955 -121.885 159.285 -121.555 ;
        RECT 158.955 -123.245 159.285 -122.915 ;
        RECT 158.955 -124.605 159.285 -124.275 ;
        RECT 158.955 -125.965 159.285 -125.635 ;
        RECT 158.955 -127.325 159.285 -126.995 ;
        RECT 158.955 -128.685 159.285 -128.355 ;
        RECT 158.955 -130.045 159.285 -129.715 ;
        RECT 158.955 -131.405 159.285 -131.075 ;
        RECT 158.955 -132.765 159.285 -132.435 ;
        RECT 158.955 -134.125 159.285 -133.795 ;
        RECT 158.955 -135.485 159.285 -135.155 ;
        RECT 158.955 -136.845 159.285 -136.515 ;
        RECT 158.955 -138.205 159.285 -137.875 ;
        RECT 158.955 -139.565 159.285 -139.235 ;
        RECT 158.955 -140.925 159.285 -140.595 ;
        RECT 158.955 -142.285 159.285 -141.955 ;
        RECT 158.955 -143.645 159.285 -143.315 ;
        RECT 158.955 -145.005 159.285 -144.675 ;
        RECT 158.955 -146.365 159.285 -146.035 ;
        RECT 158.955 -147.725 159.285 -147.395 ;
        RECT 158.955 -149.085 159.285 -148.755 ;
        RECT 158.955 -150.445 159.285 -150.115 ;
        RECT 158.955 -151.805 159.285 -151.475 ;
        RECT 158.955 -153.165 159.285 -152.835 ;
        RECT 158.955 -154.525 159.285 -154.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 244.04 110.325 245.17 ;
        RECT 109.995 239.875 110.325 240.205 ;
        RECT 109.995 238.515 110.325 238.845 ;
        RECT 109.995 237.155 110.325 237.485 ;
        RECT 110 237.155 110.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 -0.845 110.325 -0.515 ;
        RECT 109.995 -2.205 110.325 -1.875 ;
        RECT 109.995 -3.565 110.325 -3.235 ;
        RECT 110 -3.565 110.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.995 -96.045 110.325 -95.715 ;
        RECT 109.995 -97.405 110.325 -97.075 ;
        RECT 109.995 -98.765 110.325 -98.435 ;
        RECT 109.995 -100.125 110.325 -99.795 ;
        RECT 109.995 -101.485 110.325 -101.155 ;
        RECT 109.995 -102.845 110.325 -102.515 ;
        RECT 109.995 -104.205 110.325 -103.875 ;
        RECT 109.995 -105.565 110.325 -105.235 ;
        RECT 109.995 -106.925 110.325 -106.595 ;
        RECT 109.995 -108.285 110.325 -107.955 ;
        RECT 109.995 -109.645 110.325 -109.315 ;
        RECT 109.995 -111.005 110.325 -110.675 ;
        RECT 109.995 -112.365 110.325 -112.035 ;
        RECT 109.995 -113.725 110.325 -113.395 ;
        RECT 109.995 -115.085 110.325 -114.755 ;
        RECT 109.995 -116.445 110.325 -116.115 ;
        RECT 109.995 -117.805 110.325 -117.475 ;
        RECT 109.995 -119.165 110.325 -118.835 ;
        RECT 109.995 -120.525 110.325 -120.195 ;
        RECT 109.995 -121.885 110.325 -121.555 ;
        RECT 109.995 -123.245 110.325 -122.915 ;
        RECT 109.995 -124.605 110.325 -124.275 ;
        RECT 109.995 -125.965 110.325 -125.635 ;
        RECT 109.995 -127.325 110.325 -126.995 ;
        RECT 109.995 -128.685 110.325 -128.355 ;
        RECT 109.995 -130.045 110.325 -129.715 ;
        RECT 109.995 -131.405 110.325 -131.075 ;
        RECT 109.995 -132.765 110.325 -132.435 ;
        RECT 109.995 -134.125 110.325 -133.795 ;
        RECT 109.995 -135.485 110.325 -135.155 ;
        RECT 109.995 -136.845 110.325 -136.515 ;
        RECT 109.995 -138.205 110.325 -137.875 ;
        RECT 109.995 -139.565 110.325 -139.235 ;
        RECT 109.995 -140.925 110.325 -140.595 ;
        RECT 109.995 -142.285 110.325 -141.955 ;
        RECT 109.995 -143.645 110.325 -143.315 ;
        RECT 109.995 -145.005 110.325 -144.675 ;
        RECT 109.995 -146.365 110.325 -146.035 ;
        RECT 109.995 -147.725 110.325 -147.395 ;
        RECT 109.995 -149.085 110.325 -148.755 ;
        RECT 109.995 -150.445 110.325 -150.115 ;
        RECT 109.995 -151.805 110.325 -151.475 ;
        RECT 109.995 -153.165 110.325 -152.835 ;
        RECT 109.995 -154.525 110.325 -154.195 ;
        RECT 109.995 -155.885 110.325 -155.555 ;
        RECT 109.995 -157.245 110.325 -156.915 ;
        RECT 109.995 -158.605 110.325 -158.275 ;
        RECT 109.995 -159.965 110.325 -159.635 ;
        RECT 109.995 -161.325 110.325 -160.995 ;
        RECT 109.995 -162.685 110.325 -162.355 ;
        RECT 109.995 -164.045 110.325 -163.715 ;
        RECT 109.995 -165.405 110.325 -165.075 ;
        RECT 109.995 -166.765 110.325 -166.435 ;
        RECT 109.995 -168.125 110.325 -167.795 ;
        RECT 109.995 -169.485 110.325 -169.155 ;
        RECT 109.995 -170.845 110.325 -170.515 ;
        RECT 109.995 -172.205 110.325 -171.875 ;
        RECT 109.995 -173.565 110.325 -173.235 ;
        RECT 109.995 -174.925 110.325 -174.595 ;
        RECT 109.995 -176.285 110.325 -175.955 ;
        RECT 109.995 -177.645 110.325 -177.315 ;
        RECT 109.995 -179.005 110.325 -178.675 ;
        RECT 109.995 -184.65 110.325 -183.52 ;
        RECT 110 -184.765 110.32 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 244.04 111.685 245.17 ;
        RECT 111.355 239.875 111.685 240.205 ;
        RECT 111.355 238.515 111.685 238.845 ;
        RECT 111.355 237.155 111.685 237.485 ;
        RECT 111.36 237.155 111.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.355 -98.765 111.685 -98.435 ;
        RECT 111.355 -100.125 111.685 -99.795 ;
        RECT 111.355 -101.485 111.685 -101.155 ;
        RECT 111.355 -102.845 111.685 -102.515 ;
        RECT 111.355 -104.205 111.685 -103.875 ;
        RECT 111.355 -105.565 111.685 -105.235 ;
        RECT 111.355 -106.925 111.685 -106.595 ;
        RECT 111.355 -108.285 111.685 -107.955 ;
        RECT 111.355 -109.645 111.685 -109.315 ;
        RECT 111.355 -111.005 111.685 -110.675 ;
        RECT 111.355 -112.365 111.685 -112.035 ;
        RECT 111.355 -113.725 111.685 -113.395 ;
        RECT 111.355 -115.085 111.685 -114.755 ;
        RECT 111.355 -116.445 111.685 -116.115 ;
        RECT 111.355 -117.805 111.685 -117.475 ;
        RECT 111.355 -119.165 111.685 -118.835 ;
        RECT 111.355 -120.525 111.685 -120.195 ;
        RECT 111.355 -121.885 111.685 -121.555 ;
        RECT 111.355 -123.245 111.685 -122.915 ;
        RECT 111.355 -124.605 111.685 -124.275 ;
        RECT 111.355 -125.965 111.685 -125.635 ;
        RECT 111.355 -127.325 111.685 -126.995 ;
        RECT 111.355 -128.685 111.685 -128.355 ;
        RECT 111.355 -130.045 111.685 -129.715 ;
        RECT 111.355 -131.405 111.685 -131.075 ;
        RECT 111.355 -132.765 111.685 -132.435 ;
        RECT 111.355 -134.125 111.685 -133.795 ;
        RECT 111.355 -135.485 111.685 -135.155 ;
        RECT 111.355 -136.845 111.685 -136.515 ;
        RECT 111.355 -138.205 111.685 -137.875 ;
        RECT 111.355 -139.565 111.685 -139.235 ;
        RECT 111.355 -140.925 111.685 -140.595 ;
        RECT 111.355 -142.285 111.685 -141.955 ;
        RECT 111.355 -143.645 111.685 -143.315 ;
        RECT 111.355 -145.005 111.685 -144.675 ;
        RECT 111.355 -146.365 111.685 -146.035 ;
        RECT 111.355 -147.725 111.685 -147.395 ;
        RECT 111.355 -149.085 111.685 -148.755 ;
        RECT 111.355 -150.445 111.685 -150.115 ;
        RECT 111.355 -151.805 111.685 -151.475 ;
        RECT 111.355 -153.165 111.685 -152.835 ;
        RECT 111.355 -154.525 111.685 -154.195 ;
        RECT 111.355 -155.885 111.685 -155.555 ;
        RECT 111.355 -157.245 111.685 -156.915 ;
        RECT 111.355 -158.605 111.685 -158.275 ;
        RECT 111.355 -159.965 111.685 -159.635 ;
        RECT 111.355 -161.325 111.685 -160.995 ;
        RECT 111.355 -162.685 111.685 -162.355 ;
        RECT 111.355 -164.045 111.685 -163.715 ;
        RECT 111.355 -165.405 111.685 -165.075 ;
        RECT 111.355 -166.765 111.685 -166.435 ;
        RECT 111.355 -168.125 111.685 -167.795 ;
        RECT 111.355 -169.485 111.685 -169.155 ;
        RECT 111.355 -170.845 111.685 -170.515 ;
        RECT 111.355 -172.205 111.685 -171.875 ;
        RECT 111.355 -173.565 111.685 -173.235 ;
        RECT 111.355 -174.925 111.685 -174.595 ;
        RECT 111.355 -176.285 111.685 -175.955 ;
        RECT 111.355 -177.645 111.685 -177.315 ;
        RECT 111.355 -179.005 111.685 -178.675 ;
        RECT 111.355 -184.65 111.685 -183.52 ;
        RECT 111.36 -184.765 111.68 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 111.66 -98.075 111.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.715 244.04 113.045 245.17 ;
        RECT 112.715 239.875 113.045 240.205 ;
        RECT 112.715 238.515 113.045 238.845 ;
        RECT 112.715 237.155 113.045 237.485 ;
        RECT 112.72 237.155 113.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 244.04 114.405 245.17 ;
        RECT 114.075 239.875 114.405 240.205 ;
        RECT 114.075 238.515 114.405 238.845 ;
        RECT 114.075 237.155 114.405 237.485 ;
        RECT 114.08 237.155 114.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.075 -0.845 114.405 -0.515 ;
        RECT 114.075 -2.205 114.405 -1.875 ;
        RECT 114.075 -3.565 114.405 -3.235 ;
        RECT 114.08 -3.565 114.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 244.04 115.765 245.17 ;
        RECT 115.435 239.875 115.765 240.205 ;
        RECT 115.435 238.515 115.765 238.845 ;
        RECT 115.435 237.155 115.765 237.485 ;
        RECT 115.44 237.155 115.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 -0.845 115.765 -0.515 ;
        RECT 115.435 -2.205 115.765 -1.875 ;
        RECT 115.435 -3.565 115.765 -3.235 ;
        RECT 115.44 -3.565 115.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 115.435 -96.045 115.765 -95.715 ;
        RECT 115.435 -97.405 115.765 -97.075 ;
        RECT 115.435 -98.765 115.765 -98.435 ;
        RECT 115.435 -100.125 115.765 -99.795 ;
        RECT 115.435 -101.485 115.765 -101.155 ;
        RECT 115.435 -102.845 115.765 -102.515 ;
        RECT 115.435 -104.205 115.765 -103.875 ;
        RECT 115.435 -105.565 115.765 -105.235 ;
        RECT 115.435 -106.925 115.765 -106.595 ;
        RECT 115.435 -108.285 115.765 -107.955 ;
        RECT 115.435 -109.645 115.765 -109.315 ;
        RECT 115.435 -111.005 115.765 -110.675 ;
        RECT 115.435 -112.365 115.765 -112.035 ;
        RECT 115.435 -113.725 115.765 -113.395 ;
        RECT 115.435 -115.085 115.765 -114.755 ;
        RECT 115.435 -116.445 115.765 -116.115 ;
        RECT 115.435 -117.805 115.765 -117.475 ;
        RECT 115.435 -119.165 115.765 -118.835 ;
        RECT 115.435 -120.525 115.765 -120.195 ;
        RECT 115.435 -121.885 115.765 -121.555 ;
        RECT 115.435 -123.245 115.765 -122.915 ;
        RECT 115.435 -124.605 115.765 -124.275 ;
        RECT 115.435 -125.965 115.765 -125.635 ;
        RECT 115.435 -127.325 115.765 -126.995 ;
        RECT 115.435 -128.685 115.765 -128.355 ;
        RECT 115.435 -130.045 115.765 -129.715 ;
        RECT 115.435 -131.405 115.765 -131.075 ;
        RECT 115.435 -132.765 115.765 -132.435 ;
        RECT 115.435 -134.125 115.765 -133.795 ;
        RECT 115.435 -135.485 115.765 -135.155 ;
        RECT 115.435 -136.845 115.765 -136.515 ;
        RECT 115.435 -138.205 115.765 -137.875 ;
        RECT 115.435 -139.565 115.765 -139.235 ;
        RECT 115.435 -140.925 115.765 -140.595 ;
        RECT 115.435 -142.285 115.765 -141.955 ;
        RECT 115.435 -143.645 115.765 -143.315 ;
        RECT 115.435 -145.005 115.765 -144.675 ;
        RECT 115.435 -146.365 115.765 -146.035 ;
        RECT 115.435 -147.725 115.765 -147.395 ;
        RECT 115.435 -149.085 115.765 -148.755 ;
        RECT 115.435 -150.445 115.765 -150.115 ;
        RECT 115.435 -151.805 115.765 -151.475 ;
        RECT 115.435 -153.165 115.765 -152.835 ;
        RECT 115.435 -154.525 115.765 -154.195 ;
        RECT 115.435 -155.885 115.765 -155.555 ;
        RECT 115.435 -157.245 115.765 -156.915 ;
        RECT 115.435 -158.605 115.765 -158.275 ;
        RECT 115.435 -159.965 115.765 -159.635 ;
        RECT 115.435 -161.325 115.765 -160.995 ;
        RECT 115.435 -162.685 115.765 -162.355 ;
        RECT 115.435 -164.045 115.765 -163.715 ;
        RECT 115.435 -165.405 115.765 -165.075 ;
        RECT 115.435 -166.765 115.765 -166.435 ;
        RECT 115.435 -168.125 115.765 -167.795 ;
        RECT 115.435 -169.485 115.765 -169.155 ;
        RECT 115.435 -170.845 115.765 -170.515 ;
        RECT 115.435 -172.205 115.765 -171.875 ;
        RECT 115.435 -173.565 115.765 -173.235 ;
        RECT 115.435 -174.925 115.765 -174.595 ;
        RECT 115.435 -176.285 115.765 -175.955 ;
        RECT 115.435 -177.645 115.765 -177.315 ;
        RECT 115.435 -179.005 115.765 -178.675 ;
        RECT 115.435 -184.65 115.765 -183.52 ;
        RECT 115.44 -184.765 115.76 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 244.04 117.125 245.17 ;
        RECT 116.795 239.875 117.125 240.205 ;
        RECT 116.795 238.515 117.125 238.845 ;
        RECT 116.795 237.155 117.125 237.485 ;
        RECT 116.8 237.155 117.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 -0.845 117.125 -0.515 ;
        RECT 116.795 -2.205 117.125 -1.875 ;
        RECT 116.795 -3.565 117.125 -3.235 ;
        RECT 116.8 -3.565 117.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.795 -96.045 117.125 -95.715 ;
        RECT 116.795 -97.405 117.125 -97.075 ;
        RECT 116.795 -98.765 117.125 -98.435 ;
        RECT 116.795 -100.125 117.125 -99.795 ;
        RECT 116.795 -101.485 117.125 -101.155 ;
        RECT 116.795 -102.845 117.125 -102.515 ;
        RECT 116.795 -104.205 117.125 -103.875 ;
        RECT 116.795 -105.565 117.125 -105.235 ;
        RECT 116.795 -106.925 117.125 -106.595 ;
        RECT 116.795 -108.285 117.125 -107.955 ;
        RECT 116.795 -109.645 117.125 -109.315 ;
        RECT 116.795 -111.005 117.125 -110.675 ;
        RECT 116.795 -112.365 117.125 -112.035 ;
        RECT 116.795 -113.725 117.125 -113.395 ;
        RECT 116.795 -115.085 117.125 -114.755 ;
        RECT 116.795 -116.445 117.125 -116.115 ;
        RECT 116.795 -117.805 117.125 -117.475 ;
        RECT 116.795 -119.165 117.125 -118.835 ;
        RECT 116.795 -120.525 117.125 -120.195 ;
        RECT 116.795 -121.885 117.125 -121.555 ;
        RECT 116.795 -123.245 117.125 -122.915 ;
        RECT 116.795 -124.605 117.125 -124.275 ;
        RECT 116.795 -125.965 117.125 -125.635 ;
        RECT 116.795 -127.325 117.125 -126.995 ;
        RECT 116.795 -128.685 117.125 -128.355 ;
        RECT 116.795 -130.045 117.125 -129.715 ;
        RECT 116.795 -131.405 117.125 -131.075 ;
        RECT 116.795 -132.765 117.125 -132.435 ;
        RECT 116.795 -134.125 117.125 -133.795 ;
        RECT 116.795 -135.485 117.125 -135.155 ;
        RECT 116.795 -136.845 117.125 -136.515 ;
        RECT 116.795 -138.205 117.125 -137.875 ;
        RECT 116.795 -139.565 117.125 -139.235 ;
        RECT 116.795 -140.925 117.125 -140.595 ;
        RECT 116.795 -142.285 117.125 -141.955 ;
        RECT 116.795 -143.645 117.125 -143.315 ;
        RECT 116.795 -145.005 117.125 -144.675 ;
        RECT 116.795 -146.365 117.125 -146.035 ;
        RECT 116.795 -147.725 117.125 -147.395 ;
        RECT 116.795 -149.085 117.125 -148.755 ;
        RECT 116.795 -150.445 117.125 -150.115 ;
        RECT 116.795 -151.805 117.125 -151.475 ;
        RECT 116.795 -153.165 117.125 -152.835 ;
        RECT 116.795 -154.525 117.125 -154.195 ;
        RECT 116.795 -155.885 117.125 -155.555 ;
        RECT 116.795 -157.245 117.125 -156.915 ;
        RECT 116.795 -158.605 117.125 -158.275 ;
        RECT 116.795 -159.965 117.125 -159.635 ;
        RECT 116.795 -161.325 117.125 -160.995 ;
        RECT 116.795 -162.685 117.125 -162.355 ;
        RECT 116.795 -164.045 117.125 -163.715 ;
        RECT 116.795 -165.405 117.125 -165.075 ;
        RECT 116.795 -166.765 117.125 -166.435 ;
        RECT 116.795 -168.125 117.125 -167.795 ;
        RECT 116.795 -169.485 117.125 -169.155 ;
        RECT 116.795 -170.845 117.125 -170.515 ;
        RECT 116.795 -172.205 117.125 -171.875 ;
        RECT 116.795 -173.565 117.125 -173.235 ;
        RECT 116.795 -174.925 117.125 -174.595 ;
        RECT 116.795 -176.285 117.125 -175.955 ;
        RECT 116.795 -177.645 117.125 -177.315 ;
        RECT 116.795 -179.005 117.125 -178.675 ;
        RECT 116.795 -184.65 117.125 -183.52 ;
        RECT 116.8 -184.765 117.12 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 244.04 118.485 245.17 ;
        RECT 118.155 239.875 118.485 240.205 ;
        RECT 118.155 238.515 118.485 238.845 ;
        RECT 118.155 237.155 118.485 237.485 ;
        RECT 118.16 237.155 118.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 -0.845 118.485 -0.515 ;
        RECT 118.155 -2.205 118.485 -1.875 ;
        RECT 118.155 -3.565 118.485 -3.235 ;
        RECT 118.16 -3.565 118.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.155 -96.045 118.485 -95.715 ;
        RECT 118.155 -97.405 118.485 -97.075 ;
        RECT 118.155 -98.765 118.485 -98.435 ;
        RECT 118.155 -100.125 118.485 -99.795 ;
        RECT 118.155 -101.485 118.485 -101.155 ;
        RECT 118.155 -102.845 118.485 -102.515 ;
        RECT 118.155 -104.205 118.485 -103.875 ;
        RECT 118.155 -105.565 118.485 -105.235 ;
        RECT 118.155 -106.925 118.485 -106.595 ;
        RECT 118.155 -108.285 118.485 -107.955 ;
        RECT 118.155 -109.645 118.485 -109.315 ;
        RECT 118.155 -111.005 118.485 -110.675 ;
        RECT 118.155 -112.365 118.485 -112.035 ;
        RECT 118.155 -113.725 118.485 -113.395 ;
        RECT 118.155 -115.085 118.485 -114.755 ;
        RECT 118.155 -116.445 118.485 -116.115 ;
        RECT 118.155 -117.805 118.485 -117.475 ;
        RECT 118.155 -119.165 118.485 -118.835 ;
        RECT 118.155 -120.525 118.485 -120.195 ;
        RECT 118.155 -121.885 118.485 -121.555 ;
        RECT 118.155 -123.245 118.485 -122.915 ;
        RECT 118.155 -124.605 118.485 -124.275 ;
        RECT 118.155 -125.965 118.485 -125.635 ;
        RECT 118.155 -127.325 118.485 -126.995 ;
        RECT 118.155 -128.685 118.485 -128.355 ;
        RECT 118.155 -130.045 118.485 -129.715 ;
        RECT 118.155 -131.405 118.485 -131.075 ;
        RECT 118.155 -132.765 118.485 -132.435 ;
        RECT 118.155 -134.125 118.485 -133.795 ;
        RECT 118.155 -135.485 118.485 -135.155 ;
        RECT 118.155 -136.845 118.485 -136.515 ;
        RECT 118.155 -138.205 118.485 -137.875 ;
        RECT 118.155 -139.565 118.485 -139.235 ;
        RECT 118.155 -140.925 118.485 -140.595 ;
        RECT 118.155 -142.285 118.485 -141.955 ;
        RECT 118.155 -143.645 118.485 -143.315 ;
        RECT 118.155 -145.005 118.485 -144.675 ;
        RECT 118.155 -146.365 118.485 -146.035 ;
        RECT 118.155 -147.725 118.485 -147.395 ;
        RECT 118.155 -149.085 118.485 -148.755 ;
        RECT 118.155 -150.445 118.485 -150.115 ;
        RECT 118.155 -151.805 118.485 -151.475 ;
        RECT 118.155 -153.165 118.485 -152.835 ;
        RECT 118.155 -154.525 118.485 -154.195 ;
        RECT 118.155 -155.885 118.485 -155.555 ;
        RECT 118.155 -157.245 118.485 -156.915 ;
        RECT 118.155 -158.605 118.485 -158.275 ;
        RECT 118.155 -159.965 118.485 -159.635 ;
        RECT 118.155 -161.325 118.485 -160.995 ;
        RECT 118.155 -162.685 118.485 -162.355 ;
        RECT 118.155 -164.045 118.485 -163.715 ;
        RECT 118.155 -165.405 118.485 -165.075 ;
        RECT 118.155 -166.765 118.485 -166.435 ;
        RECT 118.155 -168.125 118.485 -167.795 ;
        RECT 118.155 -169.485 118.485 -169.155 ;
        RECT 118.155 -170.845 118.485 -170.515 ;
        RECT 118.155 -172.205 118.485 -171.875 ;
        RECT 118.155 -173.565 118.485 -173.235 ;
        RECT 118.155 -174.925 118.485 -174.595 ;
        RECT 118.155 -176.285 118.485 -175.955 ;
        RECT 118.155 -177.645 118.485 -177.315 ;
        RECT 118.155 -179.005 118.485 -178.675 ;
        RECT 118.155 -184.65 118.485 -183.52 ;
        RECT 118.16 -184.765 118.48 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.515 244.04 119.845 245.17 ;
        RECT 119.515 239.875 119.845 240.205 ;
        RECT 119.515 238.515 119.845 238.845 ;
        RECT 119.515 237.155 119.845 237.485 ;
        RECT 119.52 237.155 119.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.515 -0.845 119.845 -0.515 ;
        RECT 119.515 -2.205 119.845 -1.875 ;
        RECT 119.515 -3.565 119.845 -3.235 ;
        RECT 119.52 -3.565 119.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 119.515 -96.045 119.845 -95.715 ;
        RECT 119.515 -97.405 119.845 -97.075 ;
        RECT 119.515 -98.765 119.845 -98.435 ;
        RECT 119.515 -100.125 119.845 -99.795 ;
        RECT 119.515 -101.485 119.845 -101.155 ;
        RECT 119.515 -102.845 119.845 -102.515 ;
        RECT 119.515 -104.205 119.845 -103.875 ;
        RECT 119.515 -105.565 119.845 -105.235 ;
        RECT 119.515 -106.925 119.845 -106.595 ;
        RECT 119.515 -108.285 119.845 -107.955 ;
        RECT 119.515 -109.645 119.845 -109.315 ;
        RECT 119.515 -111.005 119.845 -110.675 ;
        RECT 119.515 -112.365 119.845 -112.035 ;
        RECT 119.515 -113.725 119.845 -113.395 ;
        RECT 119.515 -115.085 119.845 -114.755 ;
        RECT 119.515 -116.445 119.845 -116.115 ;
        RECT 119.515 -117.805 119.845 -117.475 ;
        RECT 119.515 -119.165 119.845 -118.835 ;
        RECT 119.515 -120.525 119.845 -120.195 ;
        RECT 119.515 -121.885 119.845 -121.555 ;
        RECT 119.515 -123.245 119.845 -122.915 ;
        RECT 119.515 -124.605 119.845 -124.275 ;
        RECT 119.515 -125.965 119.845 -125.635 ;
        RECT 119.515 -127.325 119.845 -126.995 ;
        RECT 119.515 -128.685 119.845 -128.355 ;
        RECT 119.515 -130.045 119.845 -129.715 ;
        RECT 119.515 -131.405 119.845 -131.075 ;
        RECT 119.515 -132.765 119.845 -132.435 ;
        RECT 119.515 -134.125 119.845 -133.795 ;
        RECT 119.515 -135.485 119.845 -135.155 ;
        RECT 119.515 -136.845 119.845 -136.515 ;
        RECT 119.515 -138.205 119.845 -137.875 ;
        RECT 119.515 -139.565 119.845 -139.235 ;
        RECT 119.515 -140.925 119.845 -140.595 ;
        RECT 119.515 -142.285 119.845 -141.955 ;
        RECT 119.515 -143.645 119.845 -143.315 ;
        RECT 119.515 -145.005 119.845 -144.675 ;
        RECT 119.515 -146.365 119.845 -146.035 ;
        RECT 119.515 -147.725 119.845 -147.395 ;
        RECT 119.515 -149.085 119.845 -148.755 ;
        RECT 119.515 -150.445 119.845 -150.115 ;
        RECT 119.515 -151.805 119.845 -151.475 ;
        RECT 119.515 -153.165 119.845 -152.835 ;
        RECT 119.515 -154.525 119.845 -154.195 ;
        RECT 119.515 -155.885 119.845 -155.555 ;
        RECT 119.515 -157.245 119.845 -156.915 ;
        RECT 119.515 -158.605 119.845 -158.275 ;
        RECT 119.515 -159.965 119.845 -159.635 ;
        RECT 119.515 -161.325 119.845 -160.995 ;
        RECT 119.515 -162.685 119.845 -162.355 ;
        RECT 119.515 -164.045 119.845 -163.715 ;
        RECT 119.515 -165.405 119.845 -165.075 ;
        RECT 119.515 -166.765 119.845 -166.435 ;
        RECT 119.515 -168.125 119.845 -167.795 ;
        RECT 119.515 -169.485 119.845 -169.155 ;
        RECT 119.515 -170.845 119.845 -170.515 ;
        RECT 119.515 -172.205 119.845 -171.875 ;
        RECT 119.515 -173.565 119.845 -173.235 ;
        RECT 119.515 -174.925 119.845 -174.595 ;
        RECT 119.515 -176.285 119.845 -175.955 ;
        RECT 119.515 -177.645 119.845 -177.315 ;
        RECT 119.515 -179.005 119.845 -178.675 ;
        RECT 119.515 -184.65 119.845 -183.52 ;
        RECT 119.52 -184.765 119.84 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 244.04 121.205 245.17 ;
        RECT 120.875 239.875 121.205 240.205 ;
        RECT 120.875 238.515 121.205 238.845 ;
        RECT 120.875 237.155 121.205 237.485 ;
        RECT 120.88 237.155 121.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 -0.845 121.205 -0.515 ;
        RECT 120.875 -2.205 121.205 -1.875 ;
        RECT 120.875 -3.565 121.205 -3.235 ;
        RECT 120.88 -3.565 121.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.875 -96.045 121.205 -95.715 ;
        RECT 120.875 -97.405 121.205 -97.075 ;
        RECT 120.875 -98.765 121.205 -98.435 ;
        RECT 120.875 -100.125 121.205 -99.795 ;
        RECT 120.875 -101.485 121.205 -101.155 ;
        RECT 120.875 -102.845 121.205 -102.515 ;
        RECT 120.875 -104.205 121.205 -103.875 ;
        RECT 120.875 -105.565 121.205 -105.235 ;
        RECT 120.875 -106.925 121.205 -106.595 ;
        RECT 120.875 -108.285 121.205 -107.955 ;
        RECT 120.875 -109.645 121.205 -109.315 ;
        RECT 120.875 -111.005 121.205 -110.675 ;
        RECT 120.875 -112.365 121.205 -112.035 ;
        RECT 120.875 -113.725 121.205 -113.395 ;
        RECT 120.875 -115.085 121.205 -114.755 ;
        RECT 120.875 -116.445 121.205 -116.115 ;
        RECT 120.875 -117.805 121.205 -117.475 ;
        RECT 120.875 -119.165 121.205 -118.835 ;
        RECT 120.875 -120.525 121.205 -120.195 ;
        RECT 120.875 -121.885 121.205 -121.555 ;
        RECT 120.875 -123.245 121.205 -122.915 ;
        RECT 120.875 -124.605 121.205 -124.275 ;
        RECT 120.875 -125.965 121.205 -125.635 ;
        RECT 120.875 -127.325 121.205 -126.995 ;
        RECT 120.875 -128.685 121.205 -128.355 ;
        RECT 120.875 -130.045 121.205 -129.715 ;
        RECT 120.875 -131.405 121.205 -131.075 ;
        RECT 120.875 -132.765 121.205 -132.435 ;
        RECT 120.875 -134.125 121.205 -133.795 ;
        RECT 120.875 -135.485 121.205 -135.155 ;
        RECT 120.875 -136.845 121.205 -136.515 ;
        RECT 120.875 -138.205 121.205 -137.875 ;
        RECT 120.875 -139.565 121.205 -139.235 ;
        RECT 120.875 -140.925 121.205 -140.595 ;
        RECT 120.875 -142.285 121.205 -141.955 ;
        RECT 120.875 -143.645 121.205 -143.315 ;
        RECT 120.875 -145.005 121.205 -144.675 ;
        RECT 120.875 -146.365 121.205 -146.035 ;
        RECT 120.875 -147.725 121.205 -147.395 ;
        RECT 120.875 -149.085 121.205 -148.755 ;
        RECT 120.875 -150.445 121.205 -150.115 ;
        RECT 120.875 -151.805 121.205 -151.475 ;
        RECT 120.875 -153.165 121.205 -152.835 ;
        RECT 120.875 -154.525 121.205 -154.195 ;
        RECT 120.875 -155.885 121.205 -155.555 ;
        RECT 120.875 -157.245 121.205 -156.915 ;
        RECT 120.875 -158.605 121.205 -158.275 ;
        RECT 120.875 -159.965 121.205 -159.635 ;
        RECT 120.875 -161.325 121.205 -160.995 ;
        RECT 120.875 -162.685 121.205 -162.355 ;
        RECT 120.875 -164.045 121.205 -163.715 ;
        RECT 120.875 -165.405 121.205 -165.075 ;
        RECT 120.875 -166.765 121.205 -166.435 ;
        RECT 120.875 -168.125 121.205 -167.795 ;
        RECT 120.875 -169.485 121.205 -169.155 ;
        RECT 120.875 -170.845 121.205 -170.515 ;
        RECT 120.875 -172.205 121.205 -171.875 ;
        RECT 120.875 -173.565 121.205 -173.235 ;
        RECT 120.875 -174.925 121.205 -174.595 ;
        RECT 120.875 -176.285 121.205 -175.955 ;
        RECT 120.875 -177.645 121.205 -177.315 ;
        RECT 120.875 -179.005 121.205 -178.675 ;
        RECT 120.875 -184.65 121.205 -183.52 ;
        RECT 120.88 -184.765 121.2 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 244.04 122.565 245.17 ;
        RECT 122.235 239.875 122.565 240.205 ;
        RECT 122.235 238.515 122.565 238.845 ;
        RECT 122.235 237.155 122.565 237.485 ;
        RECT 122.24 237.155 122.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.235 -98.765 122.565 -98.435 ;
        RECT 122.235 -100.125 122.565 -99.795 ;
        RECT 122.235 -101.485 122.565 -101.155 ;
        RECT 122.235 -102.845 122.565 -102.515 ;
        RECT 122.235 -104.205 122.565 -103.875 ;
        RECT 122.235 -105.565 122.565 -105.235 ;
        RECT 122.235 -106.925 122.565 -106.595 ;
        RECT 122.235 -108.285 122.565 -107.955 ;
        RECT 122.235 -109.645 122.565 -109.315 ;
        RECT 122.235 -111.005 122.565 -110.675 ;
        RECT 122.235 -112.365 122.565 -112.035 ;
        RECT 122.235 -113.725 122.565 -113.395 ;
        RECT 122.235 -115.085 122.565 -114.755 ;
        RECT 122.235 -116.445 122.565 -116.115 ;
        RECT 122.235 -117.805 122.565 -117.475 ;
        RECT 122.235 -119.165 122.565 -118.835 ;
        RECT 122.235 -120.525 122.565 -120.195 ;
        RECT 122.235 -121.885 122.565 -121.555 ;
        RECT 122.235 -123.245 122.565 -122.915 ;
        RECT 122.235 -124.605 122.565 -124.275 ;
        RECT 122.235 -125.965 122.565 -125.635 ;
        RECT 122.235 -127.325 122.565 -126.995 ;
        RECT 122.235 -128.685 122.565 -128.355 ;
        RECT 122.235 -130.045 122.565 -129.715 ;
        RECT 122.235 -131.405 122.565 -131.075 ;
        RECT 122.235 -132.765 122.565 -132.435 ;
        RECT 122.235 -134.125 122.565 -133.795 ;
        RECT 122.235 -135.485 122.565 -135.155 ;
        RECT 122.235 -136.845 122.565 -136.515 ;
        RECT 122.235 -138.205 122.565 -137.875 ;
        RECT 122.235 -139.565 122.565 -139.235 ;
        RECT 122.235 -140.925 122.565 -140.595 ;
        RECT 122.235 -142.285 122.565 -141.955 ;
        RECT 122.235 -143.645 122.565 -143.315 ;
        RECT 122.235 -145.005 122.565 -144.675 ;
        RECT 122.235 -146.365 122.565 -146.035 ;
        RECT 122.235 -147.725 122.565 -147.395 ;
        RECT 122.235 -149.085 122.565 -148.755 ;
        RECT 122.235 -150.445 122.565 -150.115 ;
        RECT 122.235 -151.805 122.565 -151.475 ;
        RECT 122.235 -153.165 122.565 -152.835 ;
        RECT 122.235 -154.525 122.565 -154.195 ;
        RECT 122.235 -155.885 122.565 -155.555 ;
        RECT 122.235 -157.245 122.565 -156.915 ;
        RECT 122.235 -158.605 122.565 -158.275 ;
        RECT 122.235 -159.965 122.565 -159.635 ;
        RECT 122.235 -161.325 122.565 -160.995 ;
        RECT 122.235 -162.685 122.565 -162.355 ;
        RECT 122.235 -164.045 122.565 -163.715 ;
        RECT 122.235 -165.405 122.565 -165.075 ;
        RECT 122.235 -166.765 122.565 -166.435 ;
        RECT 122.235 -168.125 122.565 -167.795 ;
        RECT 122.235 -169.485 122.565 -169.155 ;
        RECT 122.235 -170.845 122.565 -170.515 ;
        RECT 122.235 -172.205 122.565 -171.875 ;
        RECT 122.235 -173.565 122.565 -173.235 ;
        RECT 122.235 -174.925 122.565 -174.595 ;
        RECT 122.235 -176.285 122.565 -175.955 ;
        RECT 122.235 -177.645 122.565 -177.315 ;
        RECT 122.235 -179.005 122.565 -178.675 ;
        RECT 122.235 -184.65 122.565 -183.52 ;
        RECT 122.24 -184.765 122.56 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.56 -98.075 122.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.595 244.04 123.925 245.17 ;
        RECT 123.595 239.875 123.925 240.205 ;
        RECT 123.595 238.515 123.925 238.845 ;
        RECT 123.595 237.155 123.925 237.485 ;
        RECT 123.6 237.155 123.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 244.04 125.285 245.17 ;
        RECT 124.955 239.875 125.285 240.205 ;
        RECT 124.955 238.515 125.285 238.845 ;
        RECT 124.955 237.155 125.285 237.485 ;
        RECT 124.96 237.155 125.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.955 -0.845 125.285 -0.515 ;
        RECT 124.955 -2.205 125.285 -1.875 ;
        RECT 124.955 -3.565 125.285 -3.235 ;
        RECT 124.96 -3.565 125.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 244.04 126.645 245.17 ;
        RECT 126.315 239.875 126.645 240.205 ;
        RECT 126.315 238.515 126.645 238.845 ;
        RECT 126.315 237.155 126.645 237.485 ;
        RECT 126.32 237.155 126.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 -0.845 126.645 -0.515 ;
        RECT 126.315 -2.205 126.645 -1.875 ;
        RECT 126.315 -3.565 126.645 -3.235 ;
        RECT 126.32 -3.565 126.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.315 -96.045 126.645 -95.715 ;
        RECT 126.315 -97.405 126.645 -97.075 ;
        RECT 126.315 -98.765 126.645 -98.435 ;
        RECT 126.315 -100.125 126.645 -99.795 ;
        RECT 126.315 -101.485 126.645 -101.155 ;
        RECT 126.315 -102.845 126.645 -102.515 ;
        RECT 126.315 -104.205 126.645 -103.875 ;
        RECT 126.315 -105.565 126.645 -105.235 ;
        RECT 126.315 -106.925 126.645 -106.595 ;
        RECT 126.315 -108.285 126.645 -107.955 ;
        RECT 126.315 -109.645 126.645 -109.315 ;
        RECT 126.315 -111.005 126.645 -110.675 ;
        RECT 126.315 -112.365 126.645 -112.035 ;
        RECT 126.315 -113.725 126.645 -113.395 ;
        RECT 126.315 -115.085 126.645 -114.755 ;
        RECT 126.315 -116.445 126.645 -116.115 ;
        RECT 126.315 -117.805 126.645 -117.475 ;
        RECT 126.315 -119.165 126.645 -118.835 ;
        RECT 126.315 -120.525 126.645 -120.195 ;
        RECT 126.315 -121.885 126.645 -121.555 ;
        RECT 126.315 -123.245 126.645 -122.915 ;
        RECT 126.315 -124.605 126.645 -124.275 ;
        RECT 126.315 -125.965 126.645 -125.635 ;
        RECT 126.315 -127.325 126.645 -126.995 ;
        RECT 126.315 -128.685 126.645 -128.355 ;
        RECT 126.315 -130.045 126.645 -129.715 ;
        RECT 126.315 -131.405 126.645 -131.075 ;
        RECT 126.315 -132.765 126.645 -132.435 ;
        RECT 126.315 -134.125 126.645 -133.795 ;
        RECT 126.315 -135.485 126.645 -135.155 ;
        RECT 126.315 -136.845 126.645 -136.515 ;
        RECT 126.315 -138.205 126.645 -137.875 ;
        RECT 126.315 -139.565 126.645 -139.235 ;
        RECT 126.315 -140.925 126.645 -140.595 ;
        RECT 126.315 -142.285 126.645 -141.955 ;
        RECT 126.315 -143.645 126.645 -143.315 ;
        RECT 126.315 -145.005 126.645 -144.675 ;
        RECT 126.315 -146.365 126.645 -146.035 ;
        RECT 126.315 -147.725 126.645 -147.395 ;
        RECT 126.315 -149.085 126.645 -148.755 ;
        RECT 126.315 -150.445 126.645 -150.115 ;
        RECT 126.315 -151.805 126.645 -151.475 ;
        RECT 126.315 -153.165 126.645 -152.835 ;
        RECT 126.315 -154.525 126.645 -154.195 ;
        RECT 126.315 -155.885 126.645 -155.555 ;
        RECT 126.315 -157.245 126.645 -156.915 ;
        RECT 126.315 -158.605 126.645 -158.275 ;
        RECT 126.315 -159.965 126.645 -159.635 ;
        RECT 126.315 -161.325 126.645 -160.995 ;
        RECT 126.315 -162.685 126.645 -162.355 ;
        RECT 126.315 -164.045 126.645 -163.715 ;
        RECT 126.315 -165.405 126.645 -165.075 ;
        RECT 126.315 -166.765 126.645 -166.435 ;
        RECT 126.315 -168.125 126.645 -167.795 ;
        RECT 126.315 -169.485 126.645 -169.155 ;
        RECT 126.315 -170.845 126.645 -170.515 ;
        RECT 126.315 -172.205 126.645 -171.875 ;
        RECT 126.315 -173.565 126.645 -173.235 ;
        RECT 126.315 -174.925 126.645 -174.595 ;
        RECT 126.315 -176.285 126.645 -175.955 ;
        RECT 126.315 -177.645 126.645 -177.315 ;
        RECT 126.315 -179.005 126.645 -178.675 ;
        RECT 126.315 -184.65 126.645 -183.52 ;
        RECT 126.32 -184.765 126.64 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 244.04 128.005 245.17 ;
        RECT 127.675 239.875 128.005 240.205 ;
        RECT 127.675 238.515 128.005 238.845 ;
        RECT 127.675 237.155 128.005 237.485 ;
        RECT 127.68 237.155 128 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 -0.845 128.005 -0.515 ;
        RECT 127.675 -2.205 128.005 -1.875 ;
        RECT 127.675 -3.565 128.005 -3.235 ;
        RECT 127.68 -3.565 128 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.675 -96.045 128.005 -95.715 ;
        RECT 127.675 -97.405 128.005 -97.075 ;
        RECT 127.675 -98.765 128.005 -98.435 ;
        RECT 127.675 -100.125 128.005 -99.795 ;
        RECT 127.675 -101.485 128.005 -101.155 ;
        RECT 127.675 -102.845 128.005 -102.515 ;
        RECT 127.675 -104.205 128.005 -103.875 ;
        RECT 127.675 -105.565 128.005 -105.235 ;
        RECT 127.675 -106.925 128.005 -106.595 ;
        RECT 127.675 -108.285 128.005 -107.955 ;
        RECT 127.675 -109.645 128.005 -109.315 ;
        RECT 127.675 -111.005 128.005 -110.675 ;
        RECT 127.675 -112.365 128.005 -112.035 ;
        RECT 127.675 -113.725 128.005 -113.395 ;
        RECT 127.675 -115.085 128.005 -114.755 ;
        RECT 127.675 -116.445 128.005 -116.115 ;
        RECT 127.675 -117.805 128.005 -117.475 ;
        RECT 127.675 -119.165 128.005 -118.835 ;
        RECT 127.675 -120.525 128.005 -120.195 ;
        RECT 127.675 -121.885 128.005 -121.555 ;
        RECT 127.675 -123.245 128.005 -122.915 ;
        RECT 127.675 -124.605 128.005 -124.275 ;
        RECT 127.675 -125.965 128.005 -125.635 ;
        RECT 127.675 -127.325 128.005 -126.995 ;
        RECT 127.675 -128.685 128.005 -128.355 ;
        RECT 127.675 -130.045 128.005 -129.715 ;
        RECT 127.675 -131.405 128.005 -131.075 ;
        RECT 127.675 -132.765 128.005 -132.435 ;
        RECT 127.675 -134.125 128.005 -133.795 ;
        RECT 127.675 -135.485 128.005 -135.155 ;
        RECT 127.675 -136.845 128.005 -136.515 ;
        RECT 127.675 -138.205 128.005 -137.875 ;
        RECT 127.675 -139.565 128.005 -139.235 ;
        RECT 127.675 -140.925 128.005 -140.595 ;
        RECT 127.675 -142.285 128.005 -141.955 ;
        RECT 127.675 -143.645 128.005 -143.315 ;
        RECT 127.675 -145.005 128.005 -144.675 ;
        RECT 127.675 -146.365 128.005 -146.035 ;
        RECT 127.675 -147.725 128.005 -147.395 ;
        RECT 127.675 -149.085 128.005 -148.755 ;
        RECT 127.675 -150.445 128.005 -150.115 ;
        RECT 127.675 -151.805 128.005 -151.475 ;
        RECT 127.675 -153.165 128.005 -152.835 ;
        RECT 127.675 -154.525 128.005 -154.195 ;
        RECT 127.675 -155.885 128.005 -155.555 ;
        RECT 127.675 -157.245 128.005 -156.915 ;
        RECT 127.675 -158.605 128.005 -158.275 ;
        RECT 127.675 -159.965 128.005 -159.635 ;
        RECT 127.675 -161.325 128.005 -160.995 ;
        RECT 127.675 -162.685 128.005 -162.355 ;
        RECT 127.675 -164.045 128.005 -163.715 ;
        RECT 127.675 -165.405 128.005 -165.075 ;
        RECT 127.675 -166.765 128.005 -166.435 ;
        RECT 127.675 -168.125 128.005 -167.795 ;
        RECT 127.675 -169.485 128.005 -169.155 ;
        RECT 127.675 -170.845 128.005 -170.515 ;
        RECT 127.675 -172.205 128.005 -171.875 ;
        RECT 127.675 -173.565 128.005 -173.235 ;
        RECT 127.675 -174.925 128.005 -174.595 ;
        RECT 127.675 -176.285 128.005 -175.955 ;
        RECT 127.675 -177.645 128.005 -177.315 ;
        RECT 127.675 -179.005 128.005 -178.675 ;
        RECT 127.675 -184.65 128.005 -183.52 ;
        RECT 127.68 -184.765 128 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 244.04 129.365 245.17 ;
        RECT 129.035 239.875 129.365 240.205 ;
        RECT 129.035 238.515 129.365 238.845 ;
        RECT 129.035 237.155 129.365 237.485 ;
        RECT 129.04 237.155 129.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 -0.845 129.365 -0.515 ;
        RECT 129.035 -2.205 129.365 -1.875 ;
        RECT 129.035 -3.565 129.365 -3.235 ;
        RECT 129.04 -3.565 129.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.035 -96.045 129.365 -95.715 ;
        RECT 129.035 -97.405 129.365 -97.075 ;
        RECT 129.035 -98.765 129.365 -98.435 ;
        RECT 129.035 -100.125 129.365 -99.795 ;
        RECT 129.035 -101.485 129.365 -101.155 ;
        RECT 129.035 -102.845 129.365 -102.515 ;
        RECT 129.035 -104.205 129.365 -103.875 ;
        RECT 129.035 -105.565 129.365 -105.235 ;
        RECT 129.035 -106.925 129.365 -106.595 ;
        RECT 129.035 -108.285 129.365 -107.955 ;
        RECT 129.035 -109.645 129.365 -109.315 ;
        RECT 129.035 -111.005 129.365 -110.675 ;
        RECT 129.035 -112.365 129.365 -112.035 ;
        RECT 129.035 -113.725 129.365 -113.395 ;
        RECT 129.035 -115.085 129.365 -114.755 ;
        RECT 129.035 -116.445 129.365 -116.115 ;
        RECT 129.035 -117.805 129.365 -117.475 ;
        RECT 129.035 -119.165 129.365 -118.835 ;
        RECT 129.035 -120.525 129.365 -120.195 ;
        RECT 129.035 -121.885 129.365 -121.555 ;
        RECT 129.035 -123.245 129.365 -122.915 ;
        RECT 129.035 -124.605 129.365 -124.275 ;
        RECT 129.035 -125.965 129.365 -125.635 ;
        RECT 129.035 -127.325 129.365 -126.995 ;
        RECT 129.035 -128.685 129.365 -128.355 ;
        RECT 129.035 -130.045 129.365 -129.715 ;
        RECT 129.035 -131.405 129.365 -131.075 ;
        RECT 129.035 -132.765 129.365 -132.435 ;
        RECT 129.035 -134.125 129.365 -133.795 ;
        RECT 129.035 -135.485 129.365 -135.155 ;
        RECT 129.035 -136.845 129.365 -136.515 ;
        RECT 129.035 -138.205 129.365 -137.875 ;
        RECT 129.035 -139.565 129.365 -139.235 ;
        RECT 129.035 -140.925 129.365 -140.595 ;
        RECT 129.035 -142.285 129.365 -141.955 ;
        RECT 129.035 -143.645 129.365 -143.315 ;
        RECT 129.035 -145.005 129.365 -144.675 ;
        RECT 129.035 -146.365 129.365 -146.035 ;
        RECT 129.035 -147.725 129.365 -147.395 ;
        RECT 129.035 -149.085 129.365 -148.755 ;
        RECT 129.035 -150.445 129.365 -150.115 ;
        RECT 129.035 -151.805 129.365 -151.475 ;
        RECT 129.035 -153.165 129.365 -152.835 ;
        RECT 129.035 -154.525 129.365 -154.195 ;
        RECT 129.035 -155.885 129.365 -155.555 ;
        RECT 129.035 -157.245 129.365 -156.915 ;
        RECT 129.035 -158.605 129.365 -158.275 ;
        RECT 129.035 -159.965 129.365 -159.635 ;
        RECT 129.035 -161.325 129.365 -160.995 ;
        RECT 129.035 -162.685 129.365 -162.355 ;
        RECT 129.035 -164.045 129.365 -163.715 ;
        RECT 129.035 -165.405 129.365 -165.075 ;
        RECT 129.035 -166.765 129.365 -166.435 ;
        RECT 129.035 -168.125 129.365 -167.795 ;
        RECT 129.035 -169.485 129.365 -169.155 ;
        RECT 129.035 -170.845 129.365 -170.515 ;
        RECT 129.035 -172.205 129.365 -171.875 ;
        RECT 129.035 -173.565 129.365 -173.235 ;
        RECT 129.035 -174.925 129.365 -174.595 ;
        RECT 129.035 -176.285 129.365 -175.955 ;
        RECT 129.035 -177.645 129.365 -177.315 ;
        RECT 129.035 -179.005 129.365 -178.675 ;
        RECT 129.035 -184.65 129.365 -183.52 ;
        RECT 129.04 -184.765 129.36 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 244.04 130.725 245.17 ;
        RECT 130.395 239.875 130.725 240.205 ;
        RECT 130.395 238.515 130.725 238.845 ;
        RECT 130.395 237.155 130.725 237.485 ;
        RECT 130.4 237.155 130.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 -0.845 130.725 -0.515 ;
        RECT 130.395 -2.205 130.725 -1.875 ;
        RECT 130.395 -3.565 130.725 -3.235 ;
        RECT 130.4 -3.565 130.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 130.395 -96.045 130.725 -95.715 ;
        RECT 130.395 -97.405 130.725 -97.075 ;
        RECT 130.395 -98.765 130.725 -98.435 ;
        RECT 130.395 -100.125 130.725 -99.795 ;
        RECT 130.395 -101.485 130.725 -101.155 ;
        RECT 130.395 -102.845 130.725 -102.515 ;
        RECT 130.395 -104.205 130.725 -103.875 ;
        RECT 130.395 -105.565 130.725 -105.235 ;
        RECT 130.395 -106.925 130.725 -106.595 ;
        RECT 130.395 -108.285 130.725 -107.955 ;
        RECT 130.395 -109.645 130.725 -109.315 ;
        RECT 130.395 -111.005 130.725 -110.675 ;
        RECT 130.395 -112.365 130.725 -112.035 ;
        RECT 130.395 -113.725 130.725 -113.395 ;
        RECT 130.395 -115.085 130.725 -114.755 ;
        RECT 130.395 -116.445 130.725 -116.115 ;
        RECT 130.395 -117.805 130.725 -117.475 ;
        RECT 130.395 -119.165 130.725 -118.835 ;
        RECT 130.395 -120.525 130.725 -120.195 ;
        RECT 130.395 -121.885 130.725 -121.555 ;
        RECT 130.395 -123.245 130.725 -122.915 ;
        RECT 130.395 -124.605 130.725 -124.275 ;
        RECT 130.395 -125.965 130.725 -125.635 ;
        RECT 130.395 -127.325 130.725 -126.995 ;
        RECT 130.395 -128.685 130.725 -128.355 ;
        RECT 130.395 -130.045 130.725 -129.715 ;
        RECT 130.395 -131.405 130.725 -131.075 ;
        RECT 130.395 -132.765 130.725 -132.435 ;
        RECT 130.395 -134.125 130.725 -133.795 ;
        RECT 130.395 -135.485 130.725 -135.155 ;
        RECT 130.395 -136.845 130.725 -136.515 ;
        RECT 130.395 -138.205 130.725 -137.875 ;
        RECT 130.395 -139.565 130.725 -139.235 ;
        RECT 130.395 -140.925 130.725 -140.595 ;
        RECT 130.395 -142.285 130.725 -141.955 ;
        RECT 130.395 -143.645 130.725 -143.315 ;
        RECT 130.395 -145.005 130.725 -144.675 ;
        RECT 130.395 -146.365 130.725 -146.035 ;
        RECT 130.395 -147.725 130.725 -147.395 ;
        RECT 130.395 -149.085 130.725 -148.755 ;
        RECT 130.395 -150.445 130.725 -150.115 ;
        RECT 130.395 -151.805 130.725 -151.475 ;
        RECT 130.395 -153.165 130.725 -152.835 ;
        RECT 130.395 -154.525 130.725 -154.195 ;
        RECT 130.395 -155.885 130.725 -155.555 ;
        RECT 130.395 -157.245 130.725 -156.915 ;
        RECT 130.395 -158.605 130.725 -158.275 ;
        RECT 130.395 -159.965 130.725 -159.635 ;
        RECT 130.395 -161.325 130.725 -160.995 ;
        RECT 130.395 -162.685 130.725 -162.355 ;
        RECT 130.395 -164.045 130.725 -163.715 ;
        RECT 130.395 -165.405 130.725 -165.075 ;
        RECT 130.395 -166.765 130.725 -166.435 ;
        RECT 130.395 -168.125 130.725 -167.795 ;
        RECT 130.395 -169.485 130.725 -169.155 ;
        RECT 130.395 -170.845 130.725 -170.515 ;
        RECT 130.395 -172.205 130.725 -171.875 ;
        RECT 130.395 -173.565 130.725 -173.235 ;
        RECT 130.395 -174.925 130.725 -174.595 ;
        RECT 130.395 -176.285 130.725 -175.955 ;
        RECT 130.395 -177.645 130.725 -177.315 ;
        RECT 130.395 -179.005 130.725 -178.675 ;
        RECT 130.395 -184.65 130.725 -183.52 ;
        RECT 130.4 -184.765 130.72 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.755 244.04 132.085 245.17 ;
        RECT 131.755 239.875 132.085 240.205 ;
        RECT 131.755 238.515 132.085 238.845 ;
        RECT 131.755 237.155 132.085 237.485 ;
        RECT 131.76 237.155 132.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.755 -0.845 132.085 -0.515 ;
        RECT 131.755 -2.205 132.085 -1.875 ;
        RECT 131.755 -3.565 132.085 -3.235 ;
        RECT 131.76 -3.565 132.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.755 -96.045 132.085 -95.715 ;
        RECT 131.755 -97.405 132.085 -97.075 ;
        RECT 131.755 -98.765 132.085 -98.435 ;
        RECT 131.755 -100.125 132.085 -99.795 ;
        RECT 131.755 -101.485 132.085 -101.155 ;
        RECT 131.755 -102.845 132.085 -102.515 ;
        RECT 131.755 -104.205 132.085 -103.875 ;
        RECT 131.755 -105.565 132.085 -105.235 ;
        RECT 131.755 -106.925 132.085 -106.595 ;
        RECT 131.755 -108.285 132.085 -107.955 ;
        RECT 131.755 -109.645 132.085 -109.315 ;
        RECT 131.755 -111.005 132.085 -110.675 ;
        RECT 131.755 -112.365 132.085 -112.035 ;
        RECT 131.755 -113.725 132.085 -113.395 ;
        RECT 131.755 -115.085 132.085 -114.755 ;
        RECT 131.755 -116.445 132.085 -116.115 ;
        RECT 131.755 -117.805 132.085 -117.475 ;
        RECT 131.755 -119.165 132.085 -118.835 ;
        RECT 131.755 -120.525 132.085 -120.195 ;
        RECT 131.755 -121.885 132.085 -121.555 ;
        RECT 131.755 -123.245 132.085 -122.915 ;
        RECT 131.755 -124.605 132.085 -124.275 ;
        RECT 131.755 -125.965 132.085 -125.635 ;
        RECT 131.755 -127.325 132.085 -126.995 ;
        RECT 131.755 -128.685 132.085 -128.355 ;
        RECT 131.755 -130.045 132.085 -129.715 ;
        RECT 131.755 -131.405 132.085 -131.075 ;
        RECT 131.755 -132.765 132.085 -132.435 ;
        RECT 131.755 -134.125 132.085 -133.795 ;
        RECT 131.755 -135.485 132.085 -135.155 ;
        RECT 131.755 -136.845 132.085 -136.515 ;
        RECT 131.755 -138.205 132.085 -137.875 ;
        RECT 131.755 -139.565 132.085 -139.235 ;
        RECT 131.755 -140.925 132.085 -140.595 ;
        RECT 131.755 -142.285 132.085 -141.955 ;
        RECT 131.755 -143.645 132.085 -143.315 ;
        RECT 131.755 -145.005 132.085 -144.675 ;
        RECT 131.755 -146.365 132.085 -146.035 ;
        RECT 131.755 -147.725 132.085 -147.395 ;
        RECT 131.755 -149.085 132.085 -148.755 ;
        RECT 131.755 -150.445 132.085 -150.115 ;
        RECT 131.755 -151.805 132.085 -151.475 ;
        RECT 131.755 -153.165 132.085 -152.835 ;
        RECT 131.755 -154.525 132.085 -154.195 ;
        RECT 131.755 -155.885 132.085 -155.555 ;
        RECT 131.755 -157.245 132.085 -156.915 ;
        RECT 131.755 -158.605 132.085 -158.275 ;
        RECT 131.755 -159.965 132.085 -159.635 ;
        RECT 131.755 -161.325 132.085 -160.995 ;
        RECT 131.755 -162.685 132.085 -162.355 ;
        RECT 131.755 -164.045 132.085 -163.715 ;
        RECT 131.755 -165.405 132.085 -165.075 ;
        RECT 131.755 -166.765 132.085 -166.435 ;
        RECT 131.755 -168.125 132.085 -167.795 ;
        RECT 131.755 -169.485 132.085 -169.155 ;
        RECT 131.755 -170.845 132.085 -170.515 ;
        RECT 131.755 -172.205 132.085 -171.875 ;
        RECT 131.755 -173.565 132.085 -173.235 ;
        RECT 131.755 -174.925 132.085 -174.595 ;
        RECT 131.755 -176.285 132.085 -175.955 ;
        RECT 131.755 -177.645 132.085 -177.315 ;
        RECT 131.755 -179.005 132.085 -178.675 ;
        RECT 131.755 -184.65 132.085 -183.52 ;
        RECT 131.76 -184.765 132.08 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.115 244.04 133.445 245.17 ;
        RECT 133.115 239.875 133.445 240.205 ;
        RECT 133.115 238.515 133.445 238.845 ;
        RECT 133.115 237.155 133.445 237.485 ;
        RECT 133.12 237.155 133.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 244.04 87.205 245.17 ;
        RECT 86.875 239.875 87.205 240.205 ;
        RECT 86.875 238.515 87.205 238.845 ;
        RECT 86.875 237.155 87.205 237.485 ;
        RECT 86.88 237.155 87.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 -0.845 87.205 -0.515 ;
        RECT 86.875 -2.205 87.205 -1.875 ;
        RECT 86.875 -3.565 87.205 -3.235 ;
        RECT 86.88 -3.565 87.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.875 -96.045 87.205 -95.715 ;
        RECT 86.875 -97.405 87.205 -97.075 ;
        RECT 86.875 -98.765 87.205 -98.435 ;
        RECT 86.875 -100.125 87.205 -99.795 ;
        RECT 86.875 -101.485 87.205 -101.155 ;
        RECT 86.875 -102.845 87.205 -102.515 ;
        RECT 86.875 -104.205 87.205 -103.875 ;
        RECT 86.875 -105.565 87.205 -105.235 ;
        RECT 86.875 -106.925 87.205 -106.595 ;
        RECT 86.875 -108.285 87.205 -107.955 ;
        RECT 86.875 -109.645 87.205 -109.315 ;
        RECT 86.875 -111.005 87.205 -110.675 ;
        RECT 86.875 -112.365 87.205 -112.035 ;
        RECT 86.875 -113.725 87.205 -113.395 ;
        RECT 86.875 -115.085 87.205 -114.755 ;
        RECT 86.875 -116.445 87.205 -116.115 ;
        RECT 86.875 -117.805 87.205 -117.475 ;
        RECT 86.875 -119.165 87.205 -118.835 ;
        RECT 86.875 -120.525 87.205 -120.195 ;
        RECT 86.875 -121.885 87.205 -121.555 ;
        RECT 86.875 -123.245 87.205 -122.915 ;
        RECT 86.875 -124.605 87.205 -124.275 ;
        RECT 86.875 -125.965 87.205 -125.635 ;
        RECT 86.875 -127.325 87.205 -126.995 ;
        RECT 86.875 -128.685 87.205 -128.355 ;
        RECT 86.875 -130.045 87.205 -129.715 ;
        RECT 86.875 -131.405 87.205 -131.075 ;
        RECT 86.875 -132.765 87.205 -132.435 ;
        RECT 86.875 -134.125 87.205 -133.795 ;
        RECT 86.875 -135.485 87.205 -135.155 ;
        RECT 86.875 -136.845 87.205 -136.515 ;
        RECT 86.875 -138.205 87.205 -137.875 ;
        RECT 86.875 -139.565 87.205 -139.235 ;
        RECT 86.875 -140.925 87.205 -140.595 ;
        RECT 86.875 -142.285 87.205 -141.955 ;
        RECT 86.875 -143.645 87.205 -143.315 ;
        RECT 86.875 -145.005 87.205 -144.675 ;
        RECT 86.875 -146.365 87.205 -146.035 ;
        RECT 86.875 -147.725 87.205 -147.395 ;
        RECT 86.875 -149.085 87.205 -148.755 ;
        RECT 86.875 -150.445 87.205 -150.115 ;
        RECT 86.875 -151.805 87.205 -151.475 ;
        RECT 86.875 -153.165 87.205 -152.835 ;
        RECT 86.875 -154.525 87.205 -154.195 ;
        RECT 86.875 -155.885 87.205 -155.555 ;
        RECT 86.875 -157.245 87.205 -156.915 ;
        RECT 86.875 -158.605 87.205 -158.275 ;
        RECT 86.875 -159.965 87.205 -159.635 ;
        RECT 86.875 -161.325 87.205 -160.995 ;
        RECT 86.875 -162.685 87.205 -162.355 ;
        RECT 86.875 -164.045 87.205 -163.715 ;
        RECT 86.875 -165.405 87.205 -165.075 ;
        RECT 86.875 -166.765 87.205 -166.435 ;
        RECT 86.875 -168.125 87.205 -167.795 ;
        RECT 86.875 -169.485 87.205 -169.155 ;
        RECT 86.875 -170.845 87.205 -170.515 ;
        RECT 86.875 -172.205 87.205 -171.875 ;
        RECT 86.875 -173.565 87.205 -173.235 ;
        RECT 86.875 -174.925 87.205 -174.595 ;
        RECT 86.875 -176.285 87.205 -175.955 ;
        RECT 86.875 -177.645 87.205 -177.315 ;
        RECT 86.875 -179.005 87.205 -178.675 ;
        RECT 86.875 -184.65 87.205 -183.52 ;
        RECT 86.88 -184.765 87.2 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 244.04 88.565 245.17 ;
        RECT 88.235 239.875 88.565 240.205 ;
        RECT 88.235 238.515 88.565 238.845 ;
        RECT 88.235 237.155 88.565 237.485 ;
        RECT 88.24 237.155 88.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 -0.845 88.565 -0.515 ;
        RECT 88.235 -2.205 88.565 -1.875 ;
        RECT 88.235 -3.565 88.565 -3.235 ;
        RECT 88.24 -3.565 88.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.235 -96.045 88.565 -95.715 ;
        RECT 88.235 -97.405 88.565 -97.075 ;
        RECT 88.235 -98.765 88.565 -98.435 ;
        RECT 88.235 -100.125 88.565 -99.795 ;
        RECT 88.235 -101.485 88.565 -101.155 ;
        RECT 88.235 -102.845 88.565 -102.515 ;
        RECT 88.235 -104.205 88.565 -103.875 ;
        RECT 88.235 -105.565 88.565 -105.235 ;
        RECT 88.235 -106.925 88.565 -106.595 ;
        RECT 88.235 -108.285 88.565 -107.955 ;
        RECT 88.235 -109.645 88.565 -109.315 ;
        RECT 88.235 -111.005 88.565 -110.675 ;
        RECT 88.235 -112.365 88.565 -112.035 ;
        RECT 88.235 -113.725 88.565 -113.395 ;
        RECT 88.235 -115.085 88.565 -114.755 ;
        RECT 88.235 -116.445 88.565 -116.115 ;
        RECT 88.235 -117.805 88.565 -117.475 ;
        RECT 88.235 -119.165 88.565 -118.835 ;
        RECT 88.235 -120.525 88.565 -120.195 ;
        RECT 88.235 -121.885 88.565 -121.555 ;
        RECT 88.235 -123.245 88.565 -122.915 ;
        RECT 88.235 -124.605 88.565 -124.275 ;
        RECT 88.235 -125.965 88.565 -125.635 ;
        RECT 88.235 -127.325 88.565 -126.995 ;
        RECT 88.235 -128.685 88.565 -128.355 ;
        RECT 88.235 -130.045 88.565 -129.715 ;
        RECT 88.235 -131.405 88.565 -131.075 ;
        RECT 88.235 -132.765 88.565 -132.435 ;
        RECT 88.235 -134.125 88.565 -133.795 ;
        RECT 88.235 -135.485 88.565 -135.155 ;
        RECT 88.235 -136.845 88.565 -136.515 ;
        RECT 88.235 -138.205 88.565 -137.875 ;
        RECT 88.235 -139.565 88.565 -139.235 ;
        RECT 88.235 -140.925 88.565 -140.595 ;
        RECT 88.235 -142.285 88.565 -141.955 ;
        RECT 88.235 -143.645 88.565 -143.315 ;
        RECT 88.235 -145.005 88.565 -144.675 ;
        RECT 88.235 -146.365 88.565 -146.035 ;
        RECT 88.235 -147.725 88.565 -147.395 ;
        RECT 88.235 -149.085 88.565 -148.755 ;
        RECT 88.235 -150.445 88.565 -150.115 ;
        RECT 88.235 -151.805 88.565 -151.475 ;
        RECT 88.235 -153.165 88.565 -152.835 ;
        RECT 88.235 -154.525 88.565 -154.195 ;
        RECT 88.235 -155.885 88.565 -155.555 ;
        RECT 88.235 -157.245 88.565 -156.915 ;
        RECT 88.235 -158.605 88.565 -158.275 ;
        RECT 88.235 -159.965 88.565 -159.635 ;
        RECT 88.235 -161.325 88.565 -160.995 ;
        RECT 88.235 -162.685 88.565 -162.355 ;
        RECT 88.235 -164.045 88.565 -163.715 ;
        RECT 88.235 -165.405 88.565 -165.075 ;
        RECT 88.235 -166.765 88.565 -166.435 ;
        RECT 88.235 -168.125 88.565 -167.795 ;
        RECT 88.235 -169.485 88.565 -169.155 ;
        RECT 88.235 -170.845 88.565 -170.515 ;
        RECT 88.235 -172.205 88.565 -171.875 ;
        RECT 88.235 -173.565 88.565 -173.235 ;
        RECT 88.235 -174.925 88.565 -174.595 ;
        RECT 88.235 -176.285 88.565 -175.955 ;
        RECT 88.235 -177.645 88.565 -177.315 ;
        RECT 88.235 -179.005 88.565 -178.675 ;
        RECT 88.235 -184.65 88.565 -183.52 ;
        RECT 88.24 -184.765 88.56 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 244.04 89.925 245.17 ;
        RECT 89.595 239.875 89.925 240.205 ;
        RECT 89.595 238.515 89.925 238.845 ;
        RECT 89.595 237.155 89.925 237.485 ;
        RECT 89.6 237.155 89.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.595 -98.765 89.925 -98.435 ;
        RECT 89.595 -100.125 89.925 -99.795 ;
        RECT 89.595 -101.485 89.925 -101.155 ;
        RECT 89.595 -102.845 89.925 -102.515 ;
        RECT 89.595 -104.205 89.925 -103.875 ;
        RECT 89.595 -105.565 89.925 -105.235 ;
        RECT 89.595 -106.925 89.925 -106.595 ;
        RECT 89.595 -108.285 89.925 -107.955 ;
        RECT 89.595 -109.645 89.925 -109.315 ;
        RECT 89.595 -111.005 89.925 -110.675 ;
        RECT 89.595 -112.365 89.925 -112.035 ;
        RECT 89.595 -113.725 89.925 -113.395 ;
        RECT 89.595 -115.085 89.925 -114.755 ;
        RECT 89.595 -116.445 89.925 -116.115 ;
        RECT 89.595 -117.805 89.925 -117.475 ;
        RECT 89.595 -119.165 89.925 -118.835 ;
        RECT 89.595 -120.525 89.925 -120.195 ;
        RECT 89.595 -121.885 89.925 -121.555 ;
        RECT 89.595 -123.245 89.925 -122.915 ;
        RECT 89.595 -124.605 89.925 -124.275 ;
        RECT 89.595 -125.965 89.925 -125.635 ;
        RECT 89.595 -127.325 89.925 -126.995 ;
        RECT 89.595 -128.685 89.925 -128.355 ;
        RECT 89.595 -130.045 89.925 -129.715 ;
        RECT 89.595 -131.405 89.925 -131.075 ;
        RECT 89.595 -132.765 89.925 -132.435 ;
        RECT 89.595 -134.125 89.925 -133.795 ;
        RECT 89.595 -135.485 89.925 -135.155 ;
        RECT 89.595 -136.845 89.925 -136.515 ;
        RECT 89.595 -138.205 89.925 -137.875 ;
        RECT 89.595 -139.565 89.925 -139.235 ;
        RECT 89.595 -140.925 89.925 -140.595 ;
        RECT 89.595 -142.285 89.925 -141.955 ;
        RECT 89.595 -143.645 89.925 -143.315 ;
        RECT 89.595 -145.005 89.925 -144.675 ;
        RECT 89.595 -146.365 89.925 -146.035 ;
        RECT 89.595 -147.725 89.925 -147.395 ;
        RECT 89.595 -149.085 89.925 -148.755 ;
        RECT 89.595 -150.445 89.925 -150.115 ;
        RECT 89.595 -151.805 89.925 -151.475 ;
        RECT 89.595 -153.165 89.925 -152.835 ;
        RECT 89.595 -154.525 89.925 -154.195 ;
        RECT 89.595 -155.885 89.925 -155.555 ;
        RECT 89.595 -157.245 89.925 -156.915 ;
        RECT 89.595 -158.605 89.925 -158.275 ;
        RECT 89.595 -159.965 89.925 -159.635 ;
        RECT 89.595 -161.325 89.925 -160.995 ;
        RECT 89.595 -162.685 89.925 -162.355 ;
        RECT 89.595 -164.045 89.925 -163.715 ;
        RECT 89.595 -165.405 89.925 -165.075 ;
        RECT 89.595 -166.765 89.925 -166.435 ;
        RECT 89.595 -168.125 89.925 -167.795 ;
        RECT 89.595 -169.485 89.925 -169.155 ;
        RECT 89.595 -170.845 89.925 -170.515 ;
        RECT 89.595 -172.205 89.925 -171.875 ;
        RECT 89.595 -173.565 89.925 -173.235 ;
        RECT 89.595 -174.925 89.925 -174.595 ;
        RECT 89.595 -176.285 89.925 -175.955 ;
        RECT 89.595 -177.645 89.925 -177.315 ;
        RECT 89.595 -179.005 89.925 -178.675 ;
        RECT 89.595 -184.65 89.925 -183.52 ;
        RECT 89.6 -184.765 89.92 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 89.86 -98.075 90.19 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.955 244.04 91.285 245.17 ;
        RECT 90.955 239.875 91.285 240.205 ;
        RECT 90.955 238.515 91.285 238.845 ;
        RECT 90.955 237.155 91.285 237.485 ;
        RECT 90.96 237.155 91.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 244.04 92.645 245.17 ;
        RECT 92.315 239.875 92.645 240.205 ;
        RECT 92.315 238.515 92.645 238.845 ;
        RECT 92.315 237.155 92.645 237.485 ;
        RECT 92.32 237.155 92.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.315 -0.845 92.645 -0.515 ;
        RECT 92.315 -2.205 92.645 -1.875 ;
        RECT 92.315 -3.565 92.645 -3.235 ;
        RECT 92.32 -3.565 92.64 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 244.04 94.005 245.17 ;
        RECT 93.675 239.875 94.005 240.205 ;
        RECT 93.675 238.515 94.005 238.845 ;
        RECT 93.675 237.155 94.005 237.485 ;
        RECT 93.68 237.155 94 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 -0.845 94.005 -0.515 ;
        RECT 93.675 -2.205 94.005 -1.875 ;
        RECT 93.675 -3.565 94.005 -3.235 ;
        RECT 93.68 -3.565 94 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 93.675 -96.045 94.005 -95.715 ;
        RECT 93.675 -97.405 94.005 -97.075 ;
        RECT 93.675 -98.765 94.005 -98.435 ;
        RECT 93.675 -100.125 94.005 -99.795 ;
        RECT 93.675 -101.485 94.005 -101.155 ;
        RECT 93.675 -102.845 94.005 -102.515 ;
        RECT 93.675 -104.205 94.005 -103.875 ;
        RECT 93.675 -105.565 94.005 -105.235 ;
        RECT 93.675 -106.925 94.005 -106.595 ;
        RECT 93.675 -108.285 94.005 -107.955 ;
        RECT 93.675 -109.645 94.005 -109.315 ;
        RECT 93.675 -111.005 94.005 -110.675 ;
        RECT 93.675 -112.365 94.005 -112.035 ;
        RECT 93.675 -113.725 94.005 -113.395 ;
        RECT 93.675 -115.085 94.005 -114.755 ;
        RECT 93.675 -116.445 94.005 -116.115 ;
        RECT 93.675 -117.805 94.005 -117.475 ;
        RECT 93.675 -119.165 94.005 -118.835 ;
        RECT 93.675 -120.525 94.005 -120.195 ;
        RECT 93.675 -121.885 94.005 -121.555 ;
        RECT 93.675 -123.245 94.005 -122.915 ;
        RECT 93.675 -124.605 94.005 -124.275 ;
        RECT 93.675 -125.965 94.005 -125.635 ;
        RECT 93.675 -127.325 94.005 -126.995 ;
        RECT 93.675 -128.685 94.005 -128.355 ;
        RECT 93.675 -130.045 94.005 -129.715 ;
        RECT 93.675 -131.405 94.005 -131.075 ;
        RECT 93.675 -132.765 94.005 -132.435 ;
        RECT 93.675 -134.125 94.005 -133.795 ;
        RECT 93.675 -135.485 94.005 -135.155 ;
        RECT 93.675 -136.845 94.005 -136.515 ;
        RECT 93.675 -138.205 94.005 -137.875 ;
        RECT 93.675 -139.565 94.005 -139.235 ;
        RECT 93.675 -140.925 94.005 -140.595 ;
        RECT 93.675 -142.285 94.005 -141.955 ;
        RECT 93.675 -143.645 94.005 -143.315 ;
        RECT 93.675 -145.005 94.005 -144.675 ;
        RECT 93.675 -146.365 94.005 -146.035 ;
        RECT 93.675 -147.725 94.005 -147.395 ;
        RECT 93.675 -149.085 94.005 -148.755 ;
        RECT 93.675 -150.445 94.005 -150.115 ;
        RECT 93.675 -151.805 94.005 -151.475 ;
        RECT 93.675 -153.165 94.005 -152.835 ;
        RECT 93.675 -154.525 94.005 -154.195 ;
        RECT 93.675 -155.885 94.005 -155.555 ;
        RECT 93.675 -157.245 94.005 -156.915 ;
        RECT 93.675 -158.605 94.005 -158.275 ;
        RECT 93.675 -159.965 94.005 -159.635 ;
        RECT 93.675 -161.325 94.005 -160.995 ;
        RECT 93.675 -162.685 94.005 -162.355 ;
        RECT 93.675 -164.045 94.005 -163.715 ;
        RECT 93.675 -165.405 94.005 -165.075 ;
        RECT 93.675 -166.765 94.005 -166.435 ;
        RECT 93.675 -168.125 94.005 -167.795 ;
        RECT 93.675 -169.485 94.005 -169.155 ;
        RECT 93.675 -170.845 94.005 -170.515 ;
        RECT 93.675 -172.205 94.005 -171.875 ;
        RECT 93.675 -173.565 94.005 -173.235 ;
        RECT 93.675 -174.925 94.005 -174.595 ;
        RECT 93.675 -176.285 94.005 -175.955 ;
        RECT 93.675 -177.645 94.005 -177.315 ;
        RECT 93.675 -179.005 94.005 -178.675 ;
        RECT 93.675 -184.65 94.005 -183.52 ;
        RECT 93.68 -184.765 94 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.035 244.04 95.365 245.17 ;
        RECT 95.035 239.875 95.365 240.205 ;
        RECT 95.035 238.515 95.365 238.845 ;
        RECT 95.035 237.155 95.365 237.485 ;
        RECT 95.04 237.155 95.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.035 -0.845 95.365 -0.515 ;
        RECT 95.035 -2.205 95.365 -1.875 ;
        RECT 95.035 -3.565 95.365 -3.235 ;
        RECT 95.04 -3.565 95.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.035 -96.045 95.365 -95.715 ;
        RECT 95.035 -97.405 95.365 -97.075 ;
        RECT 95.035 -98.765 95.365 -98.435 ;
        RECT 95.035 -100.125 95.365 -99.795 ;
        RECT 95.035 -101.485 95.365 -101.155 ;
        RECT 95.035 -102.845 95.365 -102.515 ;
        RECT 95.035 -104.205 95.365 -103.875 ;
        RECT 95.035 -105.565 95.365 -105.235 ;
        RECT 95.035 -106.925 95.365 -106.595 ;
        RECT 95.035 -108.285 95.365 -107.955 ;
        RECT 95.035 -109.645 95.365 -109.315 ;
        RECT 95.035 -111.005 95.365 -110.675 ;
        RECT 95.035 -112.365 95.365 -112.035 ;
        RECT 95.035 -113.725 95.365 -113.395 ;
        RECT 95.035 -115.085 95.365 -114.755 ;
        RECT 95.035 -116.445 95.365 -116.115 ;
        RECT 95.035 -117.805 95.365 -117.475 ;
        RECT 95.035 -119.165 95.365 -118.835 ;
        RECT 95.035 -120.525 95.365 -120.195 ;
        RECT 95.035 -121.885 95.365 -121.555 ;
        RECT 95.035 -123.245 95.365 -122.915 ;
        RECT 95.035 -124.605 95.365 -124.275 ;
        RECT 95.035 -125.965 95.365 -125.635 ;
        RECT 95.035 -127.325 95.365 -126.995 ;
        RECT 95.035 -128.685 95.365 -128.355 ;
        RECT 95.035 -130.045 95.365 -129.715 ;
        RECT 95.035 -131.405 95.365 -131.075 ;
        RECT 95.035 -132.765 95.365 -132.435 ;
        RECT 95.035 -134.125 95.365 -133.795 ;
        RECT 95.035 -135.485 95.365 -135.155 ;
        RECT 95.035 -136.845 95.365 -136.515 ;
        RECT 95.035 -138.205 95.365 -137.875 ;
        RECT 95.035 -139.565 95.365 -139.235 ;
        RECT 95.035 -140.925 95.365 -140.595 ;
        RECT 95.035 -142.285 95.365 -141.955 ;
        RECT 95.035 -143.645 95.365 -143.315 ;
        RECT 95.035 -145.005 95.365 -144.675 ;
        RECT 95.035 -146.365 95.365 -146.035 ;
        RECT 95.035 -147.725 95.365 -147.395 ;
        RECT 95.035 -149.085 95.365 -148.755 ;
        RECT 95.035 -150.445 95.365 -150.115 ;
        RECT 95.035 -151.805 95.365 -151.475 ;
        RECT 95.035 -153.165 95.365 -152.835 ;
        RECT 95.035 -154.525 95.365 -154.195 ;
        RECT 95.035 -155.885 95.365 -155.555 ;
        RECT 95.035 -157.245 95.365 -156.915 ;
        RECT 95.035 -158.605 95.365 -158.275 ;
        RECT 95.035 -159.965 95.365 -159.635 ;
        RECT 95.035 -161.325 95.365 -160.995 ;
        RECT 95.035 -162.685 95.365 -162.355 ;
        RECT 95.035 -164.045 95.365 -163.715 ;
        RECT 95.035 -165.405 95.365 -165.075 ;
        RECT 95.035 -166.765 95.365 -166.435 ;
        RECT 95.035 -168.125 95.365 -167.795 ;
        RECT 95.035 -169.485 95.365 -169.155 ;
        RECT 95.035 -170.845 95.365 -170.515 ;
        RECT 95.035 -172.205 95.365 -171.875 ;
        RECT 95.035 -173.565 95.365 -173.235 ;
        RECT 95.035 -174.925 95.365 -174.595 ;
        RECT 95.035 -176.285 95.365 -175.955 ;
        RECT 95.035 -177.645 95.365 -177.315 ;
        RECT 95.035 -179.005 95.365 -178.675 ;
        RECT 95.035 -184.65 95.365 -183.52 ;
        RECT 95.04 -184.765 95.36 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 244.04 96.725 245.17 ;
        RECT 96.395 239.875 96.725 240.205 ;
        RECT 96.395 238.515 96.725 238.845 ;
        RECT 96.395 237.155 96.725 237.485 ;
        RECT 96.4 237.155 96.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 -0.845 96.725 -0.515 ;
        RECT 96.395 -2.205 96.725 -1.875 ;
        RECT 96.395 -3.565 96.725 -3.235 ;
        RECT 96.4 -3.565 96.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 96.395 -96.045 96.725 -95.715 ;
        RECT 96.395 -97.405 96.725 -97.075 ;
        RECT 96.395 -98.765 96.725 -98.435 ;
        RECT 96.395 -100.125 96.725 -99.795 ;
        RECT 96.395 -101.485 96.725 -101.155 ;
        RECT 96.395 -102.845 96.725 -102.515 ;
        RECT 96.395 -104.205 96.725 -103.875 ;
        RECT 96.395 -105.565 96.725 -105.235 ;
        RECT 96.395 -106.925 96.725 -106.595 ;
        RECT 96.395 -108.285 96.725 -107.955 ;
        RECT 96.395 -109.645 96.725 -109.315 ;
        RECT 96.395 -111.005 96.725 -110.675 ;
        RECT 96.395 -112.365 96.725 -112.035 ;
        RECT 96.395 -113.725 96.725 -113.395 ;
        RECT 96.395 -115.085 96.725 -114.755 ;
        RECT 96.395 -116.445 96.725 -116.115 ;
        RECT 96.395 -117.805 96.725 -117.475 ;
        RECT 96.395 -119.165 96.725 -118.835 ;
        RECT 96.395 -120.525 96.725 -120.195 ;
        RECT 96.395 -121.885 96.725 -121.555 ;
        RECT 96.395 -123.245 96.725 -122.915 ;
        RECT 96.395 -124.605 96.725 -124.275 ;
        RECT 96.395 -125.965 96.725 -125.635 ;
        RECT 96.395 -127.325 96.725 -126.995 ;
        RECT 96.395 -128.685 96.725 -128.355 ;
        RECT 96.395 -130.045 96.725 -129.715 ;
        RECT 96.395 -131.405 96.725 -131.075 ;
        RECT 96.395 -132.765 96.725 -132.435 ;
        RECT 96.395 -134.125 96.725 -133.795 ;
        RECT 96.395 -135.485 96.725 -135.155 ;
        RECT 96.395 -136.845 96.725 -136.515 ;
        RECT 96.395 -138.205 96.725 -137.875 ;
        RECT 96.395 -139.565 96.725 -139.235 ;
        RECT 96.395 -140.925 96.725 -140.595 ;
        RECT 96.395 -142.285 96.725 -141.955 ;
        RECT 96.395 -143.645 96.725 -143.315 ;
        RECT 96.395 -145.005 96.725 -144.675 ;
        RECT 96.395 -146.365 96.725 -146.035 ;
        RECT 96.395 -147.725 96.725 -147.395 ;
        RECT 96.395 -149.085 96.725 -148.755 ;
        RECT 96.395 -150.445 96.725 -150.115 ;
        RECT 96.395 -151.805 96.725 -151.475 ;
        RECT 96.395 -153.165 96.725 -152.835 ;
        RECT 96.395 -154.525 96.725 -154.195 ;
        RECT 96.395 -155.885 96.725 -155.555 ;
        RECT 96.395 -157.245 96.725 -156.915 ;
        RECT 96.395 -158.605 96.725 -158.275 ;
        RECT 96.395 -159.965 96.725 -159.635 ;
        RECT 96.395 -161.325 96.725 -160.995 ;
        RECT 96.395 -162.685 96.725 -162.355 ;
        RECT 96.395 -164.045 96.725 -163.715 ;
        RECT 96.395 -165.405 96.725 -165.075 ;
        RECT 96.395 -166.765 96.725 -166.435 ;
        RECT 96.395 -168.125 96.725 -167.795 ;
        RECT 96.395 -169.485 96.725 -169.155 ;
        RECT 96.395 -170.845 96.725 -170.515 ;
        RECT 96.395 -172.205 96.725 -171.875 ;
        RECT 96.395 -173.565 96.725 -173.235 ;
        RECT 96.395 -174.925 96.725 -174.595 ;
        RECT 96.395 -176.285 96.725 -175.955 ;
        RECT 96.395 -177.645 96.725 -177.315 ;
        RECT 96.395 -179.005 96.725 -178.675 ;
        RECT 96.395 -184.65 96.725 -183.52 ;
        RECT 96.4 -184.765 96.72 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 244.04 98.085 245.17 ;
        RECT 97.755 239.875 98.085 240.205 ;
        RECT 97.755 238.515 98.085 238.845 ;
        RECT 97.755 237.155 98.085 237.485 ;
        RECT 97.76 237.155 98.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 -0.845 98.085 -0.515 ;
        RECT 97.755 -2.205 98.085 -1.875 ;
        RECT 97.755 -3.565 98.085 -3.235 ;
        RECT 97.76 -3.565 98.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.755 -96.045 98.085 -95.715 ;
        RECT 97.755 -97.405 98.085 -97.075 ;
        RECT 97.755 -98.765 98.085 -98.435 ;
        RECT 97.755 -100.125 98.085 -99.795 ;
        RECT 97.755 -101.485 98.085 -101.155 ;
        RECT 97.755 -102.845 98.085 -102.515 ;
        RECT 97.755 -104.205 98.085 -103.875 ;
        RECT 97.755 -105.565 98.085 -105.235 ;
        RECT 97.755 -106.925 98.085 -106.595 ;
        RECT 97.755 -108.285 98.085 -107.955 ;
        RECT 97.755 -109.645 98.085 -109.315 ;
        RECT 97.755 -111.005 98.085 -110.675 ;
        RECT 97.755 -112.365 98.085 -112.035 ;
        RECT 97.755 -113.725 98.085 -113.395 ;
        RECT 97.755 -115.085 98.085 -114.755 ;
        RECT 97.755 -116.445 98.085 -116.115 ;
        RECT 97.755 -117.805 98.085 -117.475 ;
        RECT 97.755 -119.165 98.085 -118.835 ;
        RECT 97.755 -120.525 98.085 -120.195 ;
        RECT 97.755 -121.885 98.085 -121.555 ;
        RECT 97.755 -123.245 98.085 -122.915 ;
        RECT 97.755 -124.605 98.085 -124.275 ;
        RECT 97.755 -125.965 98.085 -125.635 ;
        RECT 97.755 -127.325 98.085 -126.995 ;
        RECT 97.755 -128.685 98.085 -128.355 ;
        RECT 97.755 -130.045 98.085 -129.715 ;
        RECT 97.755 -131.405 98.085 -131.075 ;
        RECT 97.755 -132.765 98.085 -132.435 ;
        RECT 97.755 -134.125 98.085 -133.795 ;
        RECT 97.755 -135.485 98.085 -135.155 ;
        RECT 97.755 -136.845 98.085 -136.515 ;
        RECT 97.755 -138.205 98.085 -137.875 ;
        RECT 97.755 -139.565 98.085 -139.235 ;
        RECT 97.755 -140.925 98.085 -140.595 ;
        RECT 97.755 -142.285 98.085 -141.955 ;
        RECT 97.755 -143.645 98.085 -143.315 ;
        RECT 97.755 -145.005 98.085 -144.675 ;
        RECT 97.755 -146.365 98.085 -146.035 ;
        RECT 97.755 -147.725 98.085 -147.395 ;
        RECT 97.755 -149.085 98.085 -148.755 ;
        RECT 97.755 -150.445 98.085 -150.115 ;
        RECT 97.755 -151.805 98.085 -151.475 ;
        RECT 97.755 -153.165 98.085 -152.835 ;
        RECT 97.755 -154.525 98.085 -154.195 ;
        RECT 97.755 -155.885 98.085 -155.555 ;
        RECT 97.755 -157.245 98.085 -156.915 ;
        RECT 97.755 -158.605 98.085 -158.275 ;
        RECT 97.755 -159.965 98.085 -159.635 ;
        RECT 97.755 -161.325 98.085 -160.995 ;
        RECT 97.755 -162.685 98.085 -162.355 ;
        RECT 97.755 -164.045 98.085 -163.715 ;
        RECT 97.755 -165.405 98.085 -165.075 ;
        RECT 97.755 -166.765 98.085 -166.435 ;
        RECT 97.755 -168.125 98.085 -167.795 ;
        RECT 97.755 -169.485 98.085 -169.155 ;
        RECT 97.755 -170.845 98.085 -170.515 ;
        RECT 97.755 -172.205 98.085 -171.875 ;
        RECT 97.755 -173.565 98.085 -173.235 ;
        RECT 97.755 -174.925 98.085 -174.595 ;
        RECT 97.755 -176.285 98.085 -175.955 ;
        RECT 97.755 -177.645 98.085 -177.315 ;
        RECT 97.755 -179.005 98.085 -178.675 ;
        RECT 97.755 -184.65 98.085 -183.52 ;
        RECT 97.76 -184.765 98.08 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 244.04 99.445 245.17 ;
        RECT 99.115 239.875 99.445 240.205 ;
        RECT 99.115 238.515 99.445 238.845 ;
        RECT 99.115 237.155 99.445 237.485 ;
        RECT 99.12 237.155 99.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 -0.845 99.445 -0.515 ;
        RECT 99.115 -2.205 99.445 -1.875 ;
        RECT 99.115 -3.565 99.445 -3.235 ;
        RECT 99.12 -3.565 99.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.115 -96.045 99.445 -95.715 ;
        RECT 99.115 -97.405 99.445 -97.075 ;
        RECT 99.115 -98.765 99.445 -98.435 ;
        RECT 99.115 -100.125 99.445 -99.795 ;
        RECT 99.115 -101.485 99.445 -101.155 ;
        RECT 99.115 -102.845 99.445 -102.515 ;
        RECT 99.115 -104.205 99.445 -103.875 ;
        RECT 99.115 -105.565 99.445 -105.235 ;
        RECT 99.115 -106.925 99.445 -106.595 ;
        RECT 99.115 -108.285 99.445 -107.955 ;
        RECT 99.115 -109.645 99.445 -109.315 ;
        RECT 99.115 -111.005 99.445 -110.675 ;
        RECT 99.115 -112.365 99.445 -112.035 ;
        RECT 99.115 -113.725 99.445 -113.395 ;
        RECT 99.115 -115.085 99.445 -114.755 ;
        RECT 99.115 -116.445 99.445 -116.115 ;
        RECT 99.115 -117.805 99.445 -117.475 ;
        RECT 99.115 -119.165 99.445 -118.835 ;
        RECT 99.115 -120.525 99.445 -120.195 ;
        RECT 99.115 -121.885 99.445 -121.555 ;
        RECT 99.115 -123.245 99.445 -122.915 ;
        RECT 99.115 -124.605 99.445 -124.275 ;
        RECT 99.115 -125.965 99.445 -125.635 ;
        RECT 99.115 -127.325 99.445 -126.995 ;
        RECT 99.115 -128.685 99.445 -128.355 ;
        RECT 99.115 -130.045 99.445 -129.715 ;
        RECT 99.115 -131.405 99.445 -131.075 ;
        RECT 99.115 -132.765 99.445 -132.435 ;
        RECT 99.115 -134.125 99.445 -133.795 ;
        RECT 99.115 -135.485 99.445 -135.155 ;
        RECT 99.115 -136.845 99.445 -136.515 ;
        RECT 99.115 -138.205 99.445 -137.875 ;
        RECT 99.115 -139.565 99.445 -139.235 ;
        RECT 99.115 -140.925 99.445 -140.595 ;
        RECT 99.115 -142.285 99.445 -141.955 ;
        RECT 99.115 -143.645 99.445 -143.315 ;
        RECT 99.115 -145.005 99.445 -144.675 ;
        RECT 99.115 -146.365 99.445 -146.035 ;
        RECT 99.115 -147.725 99.445 -147.395 ;
        RECT 99.115 -149.085 99.445 -148.755 ;
        RECT 99.115 -150.445 99.445 -150.115 ;
        RECT 99.115 -151.805 99.445 -151.475 ;
        RECT 99.115 -153.165 99.445 -152.835 ;
        RECT 99.115 -154.525 99.445 -154.195 ;
        RECT 99.115 -155.885 99.445 -155.555 ;
        RECT 99.115 -157.245 99.445 -156.915 ;
        RECT 99.115 -158.605 99.445 -158.275 ;
        RECT 99.115 -159.965 99.445 -159.635 ;
        RECT 99.115 -161.325 99.445 -160.995 ;
        RECT 99.115 -162.685 99.445 -162.355 ;
        RECT 99.115 -164.045 99.445 -163.715 ;
        RECT 99.115 -165.405 99.445 -165.075 ;
        RECT 99.115 -166.765 99.445 -166.435 ;
        RECT 99.115 -168.125 99.445 -167.795 ;
        RECT 99.115 -169.485 99.445 -169.155 ;
        RECT 99.115 -170.845 99.445 -170.515 ;
        RECT 99.115 -172.205 99.445 -171.875 ;
        RECT 99.115 -173.565 99.445 -173.235 ;
        RECT 99.115 -174.925 99.445 -174.595 ;
        RECT 99.115 -176.285 99.445 -175.955 ;
        RECT 99.115 -177.645 99.445 -177.315 ;
        RECT 99.115 -179.005 99.445 -178.675 ;
        RECT 99.115 -184.65 99.445 -183.52 ;
        RECT 99.12 -184.765 99.44 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 244.04 100.805 245.17 ;
        RECT 100.475 239.875 100.805 240.205 ;
        RECT 100.475 238.515 100.805 238.845 ;
        RECT 100.475 237.155 100.805 237.485 ;
        RECT 100.48 237.155 100.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.475 -98.765 100.805 -98.435 ;
        RECT 100.475 -100.125 100.805 -99.795 ;
        RECT 100.475 -101.485 100.805 -101.155 ;
        RECT 100.475 -102.845 100.805 -102.515 ;
        RECT 100.475 -104.205 100.805 -103.875 ;
        RECT 100.475 -105.565 100.805 -105.235 ;
        RECT 100.475 -106.925 100.805 -106.595 ;
        RECT 100.475 -108.285 100.805 -107.955 ;
        RECT 100.475 -109.645 100.805 -109.315 ;
        RECT 100.475 -111.005 100.805 -110.675 ;
        RECT 100.475 -112.365 100.805 -112.035 ;
        RECT 100.475 -113.725 100.805 -113.395 ;
        RECT 100.475 -115.085 100.805 -114.755 ;
        RECT 100.475 -116.445 100.805 -116.115 ;
        RECT 100.475 -117.805 100.805 -117.475 ;
        RECT 100.475 -119.165 100.805 -118.835 ;
        RECT 100.475 -120.525 100.805 -120.195 ;
        RECT 100.475 -121.885 100.805 -121.555 ;
        RECT 100.475 -123.245 100.805 -122.915 ;
        RECT 100.475 -124.605 100.805 -124.275 ;
        RECT 100.475 -125.965 100.805 -125.635 ;
        RECT 100.475 -127.325 100.805 -126.995 ;
        RECT 100.475 -128.685 100.805 -128.355 ;
        RECT 100.475 -130.045 100.805 -129.715 ;
        RECT 100.475 -131.405 100.805 -131.075 ;
        RECT 100.475 -132.765 100.805 -132.435 ;
        RECT 100.475 -134.125 100.805 -133.795 ;
        RECT 100.475 -135.485 100.805 -135.155 ;
        RECT 100.475 -136.845 100.805 -136.515 ;
        RECT 100.475 -138.205 100.805 -137.875 ;
        RECT 100.475 -139.565 100.805 -139.235 ;
        RECT 100.475 -140.925 100.805 -140.595 ;
        RECT 100.475 -142.285 100.805 -141.955 ;
        RECT 100.475 -143.645 100.805 -143.315 ;
        RECT 100.475 -145.005 100.805 -144.675 ;
        RECT 100.475 -146.365 100.805 -146.035 ;
        RECT 100.475 -147.725 100.805 -147.395 ;
        RECT 100.475 -149.085 100.805 -148.755 ;
        RECT 100.475 -150.445 100.805 -150.115 ;
        RECT 100.475 -151.805 100.805 -151.475 ;
        RECT 100.475 -153.165 100.805 -152.835 ;
        RECT 100.475 -154.525 100.805 -154.195 ;
        RECT 100.475 -155.885 100.805 -155.555 ;
        RECT 100.475 -157.245 100.805 -156.915 ;
        RECT 100.475 -158.605 100.805 -158.275 ;
        RECT 100.475 -159.965 100.805 -159.635 ;
        RECT 100.475 -161.325 100.805 -160.995 ;
        RECT 100.475 -162.685 100.805 -162.355 ;
        RECT 100.475 -164.045 100.805 -163.715 ;
        RECT 100.475 -165.405 100.805 -165.075 ;
        RECT 100.475 -166.765 100.805 -166.435 ;
        RECT 100.475 -168.125 100.805 -167.795 ;
        RECT 100.475 -169.485 100.805 -169.155 ;
        RECT 100.475 -170.845 100.805 -170.515 ;
        RECT 100.475 -172.205 100.805 -171.875 ;
        RECT 100.475 -173.565 100.805 -173.235 ;
        RECT 100.475 -174.925 100.805 -174.595 ;
        RECT 100.475 -176.285 100.805 -175.955 ;
        RECT 100.475 -177.645 100.805 -177.315 ;
        RECT 100.475 -179.005 100.805 -178.675 ;
        RECT 100.475 -184.65 100.805 -183.52 ;
        RECT 100.48 -184.765 100.8 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 100.76 -98.075 101.09 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.835 244.04 102.165 245.17 ;
        RECT 101.835 239.875 102.165 240.205 ;
        RECT 101.835 238.515 102.165 238.845 ;
        RECT 101.835 237.155 102.165 237.485 ;
        RECT 101.84 237.155 102.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 244.04 103.525 245.17 ;
        RECT 103.195 239.875 103.525 240.205 ;
        RECT 103.195 238.515 103.525 238.845 ;
        RECT 103.195 237.155 103.525 237.485 ;
        RECT 103.2 237.155 103.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.195 -0.845 103.525 -0.515 ;
        RECT 103.195 -2.205 103.525 -1.875 ;
        RECT 103.195 -3.565 103.525 -3.235 ;
        RECT 103.2 -3.565 103.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 244.04 104.885 245.17 ;
        RECT 104.555 239.875 104.885 240.205 ;
        RECT 104.555 238.515 104.885 238.845 ;
        RECT 104.555 237.155 104.885 237.485 ;
        RECT 104.56 237.155 104.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 -0.845 104.885 -0.515 ;
        RECT 104.555 -2.205 104.885 -1.875 ;
        RECT 104.555 -3.565 104.885 -3.235 ;
        RECT 104.56 -3.565 104.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 104.555 -96.045 104.885 -95.715 ;
        RECT 104.555 -97.405 104.885 -97.075 ;
        RECT 104.555 -98.765 104.885 -98.435 ;
        RECT 104.555 -100.125 104.885 -99.795 ;
        RECT 104.555 -101.485 104.885 -101.155 ;
        RECT 104.555 -102.845 104.885 -102.515 ;
        RECT 104.555 -104.205 104.885 -103.875 ;
        RECT 104.555 -105.565 104.885 -105.235 ;
        RECT 104.555 -106.925 104.885 -106.595 ;
        RECT 104.555 -108.285 104.885 -107.955 ;
        RECT 104.555 -109.645 104.885 -109.315 ;
        RECT 104.555 -111.005 104.885 -110.675 ;
        RECT 104.555 -112.365 104.885 -112.035 ;
        RECT 104.555 -113.725 104.885 -113.395 ;
        RECT 104.555 -115.085 104.885 -114.755 ;
        RECT 104.555 -116.445 104.885 -116.115 ;
        RECT 104.555 -117.805 104.885 -117.475 ;
        RECT 104.555 -119.165 104.885 -118.835 ;
        RECT 104.555 -120.525 104.885 -120.195 ;
        RECT 104.555 -121.885 104.885 -121.555 ;
        RECT 104.555 -123.245 104.885 -122.915 ;
        RECT 104.555 -124.605 104.885 -124.275 ;
        RECT 104.555 -125.965 104.885 -125.635 ;
        RECT 104.555 -127.325 104.885 -126.995 ;
        RECT 104.555 -128.685 104.885 -128.355 ;
        RECT 104.555 -130.045 104.885 -129.715 ;
        RECT 104.555 -131.405 104.885 -131.075 ;
        RECT 104.555 -132.765 104.885 -132.435 ;
        RECT 104.555 -134.125 104.885 -133.795 ;
        RECT 104.555 -135.485 104.885 -135.155 ;
        RECT 104.555 -136.845 104.885 -136.515 ;
        RECT 104.555 -138.205 104.885 -137.875 ;
        RECT 104.555 -139.565 104.885 -139.235 ;
        RECT 104.555 -140.925 104.885 -140.595 ;
        RECT 104.555 -142.285 104.885 -141.955 ;
        RECT 104.555 -143.645 104.885 -143.315 ;
        RECT 104.555 -145.005 104.885 -144.675 ;
        RECT 104.555 -146.365 104.885 -146.035 ;
        RECT 104.555 -147.725 104.885 -147.395 ;
        RECT 104.555 -149.085 104.885 -148.755 ;
        RECT 104.555 -150.445 104.885 -150.115 ;
        RECT 104.555 -151.805 104.885 -151.475 ;
        RECT 104.555 -153.165 104.885 -152.835 ;
        RECT 104.555 -154.525 104.885 -154.195 ;
        RECT 104.555 -155.885 104.885 -155.555 ;
        RECT 104.555 -157.245 104.885 -156.915 ;
        RECT 104.555 -158.605 104.885 -158.275 ;
        RECT 104.555 -159.965 104.885 -159.635 ;
        RECT 104.555 -161.325 104.885 -160.995 ;
        RECT 104.555 -162.685 104.885 -162.355 ;
        RECT 104.555 -164.045 104.885 -163.715 ;
        RECT 104.555 -165.405 104.885 -165.075 ;
        RECT 104.555 -166.765 104.885 -166.435 ;
        RECT 104.555 -168.125 104.885 -167.795 ;
        RECT 104.555 -169.485 104.885 -169.155 ;
        RECT 104.555 -170.845 104.885 -170.515 ;
        RECT 104.555 -172.205 104.885 -171.875 ;
        RECT 104.555 -173.565 104.885 -173.235 ;
        RECT 104.555 -174.925 104.885 -174.595 ;
        RECT 104.555 -176.285 104.885 -175.955 ;
        RECT 104.555 -177.645 104.885 -177.315 ;
        RECT 104.555 -179.005 104.885 -178.675 ;
        RECT 104.555 -184.65 104.885 -183.52 ;
        RECT 104.56 -184.765 104.88 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 244.04 106.245 245.17 ;
        RECT 105.915 239.875 106.245 240.205 ;
        RECT 105.915 238.515 106.245 238.845 ;
        RECT 105.915 237.155 106.245 237.485 ;
        RECT 105.92 237.155 106.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 -0.845 106.245 -0.515 ;
        RECT 105.915 -2.205 106.245 -1.875 ;
        RECT 105.915 -3.565 106.245 -3.235 ;
        RECT 105.92 -3.565 106.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.915 -96.045 106.245 -95.715 ;
        RECT 105.915 -97.405 106.245 -97.075 ;
        RECT 105.915 -98.765 106.245 -98.435 ;
        RECT 105.915 -100.125 106.245 -99.795 ;
        RECT 105.915 -101.485 106.245 -101.155 ;
        RECT 105.915 -102.845 106.245 -102.515 ;
        RECT 105.915 -104.205 106.245 -103.875 ;
        RECT 105.915 -105.565 106.245 -105.235 ;
        RECT 105.915 -106.925 106.245 -106.595 ;
        RECT 105.915 -108.285 106.245 -107.955 ;
        RECT 105.915 -109.645 106.245 -109.315 ;
        RECT 105.915 -111.005 106.245 -110.675 ;
        RECT 105.915 -112.365 106.245 -112.035 ;
        RECT 105.915 -113.725 106.245 -113.395 ;
        RECT 105.915 -115.085 106.245 -114.755 ;
        RECT 105.915 -116.445 106.245 -116.115 ;
        RECT 105.915 -117.805 106.245 -117.475 ;
        RECT 105.915 -119.165 106.245 -118.835 ;
        RECT 105.915 -120.525 106.245 -120.195 ;
        RECT 105.915 -121.885 106.245 -121.555 ;
        RECT 105.915 -123.245 106.245 -122.915 ;
        RECT 105.915 -124.605 106.245 -124.275 ;
        RECT 105.915 -125.965 106.245 -125.635 ;
        RECT 105.915 -127.325 106.245 -126.995 ;
        RECT 105.915 -128.685 106.245 -128.355 ;
        RECT 105.915 -130.045 106.245 -129.715 ;
        RECT 105.915 -131.405 106.245 -131.075 ;
        RECT 105.915 -132.765 106.245 -132.435 ;
        RECT 105.915 -134.125 106.245 -133.795 ;
        RECT 105.915 -135.485 106.245 -135.155 ;
        RECT 105.915 -136.845 106.245 -136.515 ;
        RECT 105.915 -138.205 106.245 -137.875 ;
        RECT 105.915 -139.565 106.245 -139.235 ;
        RECT 105.915 -140.925 106.245 -140.595 ;
        RECT 105.915 -142.285 106.245 -141.955 ;
        RECT 105.915 -143.645 106.245 -143.315 ;
        RECT 105.915 -145.005 106.245 -144.675 ;
        RECT 105.915 -146.365 106.245 -146.035 ;
        RECT 105.915 -147.725 106.245 -147.395 ;
        RECT 105.915 -149.085 106.245 -148.755 ;
        RECT 105.915 -150.445 106.245 -150.115 ;
        RECT 105.915 -151.805 106.245 -151.475 ;
        RECT 105.915 -153.165 106.245 -152.835 ;
        RECT 105.915 -154.525 106.245 -154.195 ;
        RECT 105.915 -155.885 106.245 -155.555 ;
        RECT 105.915 -157.245 106.245 -156.915 ;
        RECT 105.915 -158.605 106.245 -158.275 ;
        RECT 105.915 -159.965 106.245 -159.635 ;
        RECT 105.915 -161.325 106.245 -160.995 ;
        RECT 105.915 -162.685 106.245 -162.355 ;
        RECT 105.915 -164.045 106.245 -163.715 ;
        RECT 105.915 -165.405 106.245 -165.075 ;
        RECT 105.915 -166.765 106.245 -166.435 ;
        RECT 105.915 -168.125 106.245 -167.795 ;
        RECT 105.915 -169.485 106.245 -169.155 ;
        RECT 105.915 -170.845 106.245 -170.515 ;
        RECT 105.915 -172.205 106.245 -171.875 ;
        RECT 105.915 -173.565 106.245 -173.235 ;
        RECT 105.915 -174.925 106.245 -174.595 ;
        RECT 105.915 -176.285 106.245 -175.955 ;
        RECT 105.915 -177.645 106.245 -177.315 ;
        RECT 105.915 -179.005 106.245 -178.675 ;
        RECT 105.915 -184.65 106.245 -183.52 ;
        RECT 105.92 -184.765 106.24 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 244.04 107.605 245.17 ;
        RECT 107.275 239.875 107.605 240.205 ;
        RECT 107.275 238.515 107.605 238.845 ;
        RECT 107.275 237.155 107.605 237.485 ;
        RECT 107.28 237.155 107.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 -0.845 107.605 -0.515 ;
        RECT 107.275 -2.205 107.605 -1.875 ;
        RECT 107.275 -3.565 107.605 -3.235 ;
        RECT 107.28 -3.565 107.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.275 -96.045 107.605 -95.715 ;
        RECT 107.275 -97.405 107.605 -97.075 ;
        RECT 107.275 -98.765 107.605 -98.435 ;
        RECT 107.275 -100.125 107.605 -99.795 ;
        RECT 107.275 -101.485 107.605 -101.155 ;
        RECT 107.275 -102.845 107.605 -102.515 ;
        RECT 107.275 -104.205 107.605 -103.875 ;
        RECT 107.275 -105.565 107.605 -105.235 ;
        RECT 107.275 -106.925 107.605 -106.595 ;
        RECT 107.275 -108.285 107.605 -107.955 ;
        RECT 107.275 -109.645 107.605 -109.315 ;
        RECT 107.275 -111.005 107.605 -110.675 ;
        RECT 107.275 -112.365 107.605 -112.035 ;
        RECT 107.275 -113.725 107.605 -113.395 ;
        RECT 107.275 -115.085 107.605 -114.755 ;
        RECT 107.275 -116.445 107.605 -116.115 ;
        RECT 107.275 -117.805 107.605 -117.475 ;
        RECT 107.275 -119.165 107.605 -118.835 ;
        RECT 107.275 -120.525 107.605 -120.195 ;
        RECT 107.275 -121.885 107.605 -121.555 ;
        RECT 107.275 -123.245 107.605 -122.915 ;
        RECT 107.275 -124.605 107.605 -124.275 ;
        RECT 107.275 -125.965 107.605 -125.635 ;
        RECT 107.275 -127.325 107.605 -126.995 ;
        RECT 107.275 -128.685 107.605 -128.355 ;
        RECT 107.275 -130.045 107.605 -129.715 ;
        RECT 107.275 -131.405 107.605 -131.075 ;
        RECT 107.275 -132.765 107.605 -132.435 ;
        RECT 107.275 -134.125 107.605 -133.795 ;
        RECT 107.275 -135.485 107.605 -135.155 ;
        RECT 107.275 -136.845 107.605 -136.515 ;
        RECT 107.275 -138.205 107.605 -137.875 ;
        RECT 107.275 -139.565 107.605 -139.235 ;
        RECT 107.275 -140.925 107.605 -140.595 ;
        RECT 107.275 -142.285 107.605 -141.955 ;
        RECT 107.275 -143.645 107.605 -143.315 ;
        RECT 107.275 -145.005 107.605 -144.675 ;
        RECT 107.275 -146.365 107.605 -146.035 ;
        RECT 107.275 -147.725 107.605 -147.395 ;
        RECT 107.275 -149.085 107.605 -148.755 ;
        RECT 107.275 -150.445 107.605 -150.115 ;
        RECT 107.275 -151.805 107.605 -151.475 ;
        RECT 107.275 -153.165 107.605 -152.835 ;
        RECT 107.275 -154.525 107.605 -154.195 ;
        RECT 107.275 -155.885 107.605 -155.555 ;
        RECT 107.275 -157.245 107.605 -156.915 ;
        RECT 107.275 -158.605 107.605 -158.275 ;
        RECT 107.275 -159.965 107.605 -159.635 ;
        RECT 107.275 -161.325 107.605 -160.995 ;
        RECT 107.275 -162.685 107.605 -162.355 ;
        RECT 107.275 -164.045 107.605 -163.715 ;
        RECT 107.275 -165.405 107.605 -165.075 ;
        RECT 107.275 -166.765 107.605 -166.435 ;
        RECT 107.275 -168.125 107.605 -167.795 ;
        RECT 107.275 -169.485 107.605 -169.155 ;
        RECT 107.275 -170.845 107.605 -170.515 ;
        RECT 107.275 -172.205 107.605 -171.875 ;
        RECT 107.275 -173.565 107.605 -173.235 ;
        RECT 107.275 -174.925 107.605 -174.595 ;
        RECT 107.275 -176.285 107.605 -175.955 ;
        RECT 107.275 -177.645 107.605 -177.315 ;
        RECT 107.275 -179.005 107.605 -178.675 ;
        RECT 107.275 -184.65 107.605 -183.52 ;
        RECT 107.28 -184.765 107.6 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 244.04 108.965 245.17 ;
        RECT 108.635 239.875 108.965 240.205 ;
        RECT 108.635 238.515 108.965 238.845 ;
        RECT 108.635 237.155 108.965 237.485 ;
        RECT 108.64 237.155 108.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 -0.845 108.965 -0.515 ;
        RECT 108.635 -2.205 108.965 -1.875 ;
        RECT 108.635 -3.565 108.965 -3.235 ;
        RECT 108.64 -3.565 108.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 108.635 -134.125 108.965 -133.795 ;
        RECT 108.635 -135.485 108.965 -135.155 ;
        RECT 108.635 -136.845 108.965 -136.515 ;
        RECT 108.635 -138.205 108.965 -137.875 ;
        RECT 108.635 -139.565 108.965 -139.235 ;
        RECT 108.635 -140.925 108.965 -140.595 ;
        RECT 108.635 -142.285 108.965 -141.955 ;
        RECT 108.635 -143.645 108.965 -143.315 ;
        RECT 108.635 -145.005 108.965 -144.675 ;
        RECT 108.635 -146.365 108.965 -146.035 ;
        RECT 108.635 -147.725 108.965 -147.395 ;
        RECT 108.635 -149.085 108.965 -148.755 ;
        RECT 108.635 -150.445 108.965 -150.115 ;
        RECT 108.635 -151.805 108.965 -151.475 ;
        RECT 108.635 -153.165 108.965 -152.835 ;
        RECT 108.635 -154.525 108.965 -154.195 ;
        RECT 108.635 -155.885 108.965 -155.555 ;
        RECT 108.635 -157.245 108.965 -156.915 ;
        RECT 108.635 -158.605 108.965 -158.275 ;
        RECT 108.635 -159.965 108.965 -159.635 ;
        RECT 108.635 -161.325 108.965 -160.995 ;
        RECT 108.635 -162.685 108.965 -162.355 ;
        RECT 108.635 -164.045 108.965 -163.715 ;
        RECT 108.635 -165.405 108.965 -165.075 ;
        RECT 108.635 -166.765 108.965 -166.435 ;
        RECT 108.635 -168.125 108.965 -167.795 ;
        RECT 108.635 -169.485 108.965 -169.155 ;
        RECT 108.635 -170.845 108.965 -170.515 ;
        RECT 108.635 -172.205 108.965 -171.875 ;
        RECT 108.635 -173.565 108.965 -173.235 ;
        RECT 108.635 -174.925 108.965 -174.595 ;
        RECT 108.635 -176.285 108.965 -175.955 ;
        RECT 108.635 -177.645 108.965 -177.315 ;
        RECT 108.635 -179.005 108.965 -178.675 ;
        RECT 108.635 -184.65 108.965 -183.52 ;
        RECT 108.64 -184.765 108.96 -95.04 ;
        RECT 108.635 -96.045 108.965 -95.715 ;
        RECT 108.635 -97.405 108.965 -97.075 ;
        RECT 108.635 -98.765 108.965 -98.435 ;
        RECT 108.635 -100.125 108.965 -99.795 ;
        RECT 108.635 -101.485 108.965 -101.155 ;
        RECT 108.635 -102.845 108.965 -102.515 ;
        RECT 108.635 -104.205 108.965 -103.875 ;
        RECT 108.635 -105.565 108.965 -105.235 ;
        RECT 108.635 -106.925 108.965 -106.595 ;
        RECT 108.635 -108.285 108.965 -107.955 ;
        RECT 108.635 -109.645 108.965 -109.315 ;
        RECT 108.635 -111.005 108.965 -110.675 ;
        RECT 108.635 -112.365 108.965 -112.035 ;
        RECT 108.635 -113.725 108.965 -113.395 ;
        RECT 108.635 -115.085 108.965 -114.755 ;
        RECT 108.635 -116.445 108.965 -116.115 ;
        RECT 108.635 -117.805 108.965 -117.475 ;
        RECT 108.635 -119.165 108.965 -118.835 ;
        RECT 108.635 -120.525 108.965 -120.195 ;
        RECT 108.635 -121.885 108.965 -121.555 ;
        RECT 108.635 -123.245 108.965 -122.915 ;
        RECT 108.635 -124.605 108.965 -124.275 ;
        RECT 108.635 -125.965 108.965 -125.635 ;
        RECT 108.635 -127.325 108.965 -126.995 ;
        RECT 108.635 -128.685 108.965 -128.355 ;
        RECT 108.635 -130.045 108.965 -129.715 ;
        RECT 108.635 -131.405 108.965 -131.075 ;
        RECT 108.635 -132.765 108.965 -132.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 244.04 62.725 245.17 ;
        RECT 62.395 239.875 62.725 240.205 ;
        RECT 62.395 238.515 62.725 238.845 ;
        RECT 62.395 237.155 62.725 237.485 ;
        RECT 62.4 237.155 62.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 -0.845 62.725 -0.515 ;
        RECT 62.395 -2.205 62.725 -1.875 ;
        RECT 62.395 -3.565 62.725 -3.235 ;
        RECT 62.4 -3.565 62.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 62.395 -96.045 62.725 -95.715 ;
        RECT 62.395 -97.405 62.725 -97.075 ;
        RECT 62.395 -98.765 62.725 -98.435 ;
        RECT 62.395 -100.125 62.725 -99.795 ;
        RECT 62.395 -101.485 62.725 -101.155 ;
        RECT 62.395 -102.845 62.725 -102.515 ;
        RECT 62.395 -104.205 62.725 -103.875 ;
        RECT 62.395 -105.565 62.725 -105.235 ;
        RECT 62.395 -106.925 62.725 -106.595 ;
        RECT 62.395 -108.285 62.725 -107.955 ;
        RECT 62.395 -109.645 62.725 -109.315 ;
        RECT 62.395 -111.005 62.725 -110.675 ;
        RECT 62.395 -112.365 62.725 -112.035 ;
        RECT 62.395 -113.725 62.725 -113.395 ;
        RECT 62.395 -115.085 62.725 -114.755 ;
        RECT 62.395 -116.445 62.725 -116.115 ;
        RECT 62.395 -117.805 62.725 -117.475 ;
        RECT 62.395 -119.165 62.725 -118.835 ;
        RECT 62.395 -120.525 62.725 -120.195 ;
        RECT 62.395 -121.885 62.725 -121.555 ;
        RECT 62.395 -123.245 62.725 -122.915 ;
        RECT 62.395 -124.605 62.725 -124.275 ;
        RECT 62.395 -125.965 62.725 -125.635 ;
        RECT 62.395 -127.325 62.725 -126.995 ;
        RECT 62.395 -128.685 62.725 -128.355 ;
        RECT 62.395 -130.045 62.725 -129.715 ;
        RECT 62.395 -131.405 62.725 -131.075 ;
        RECT 62.395 -132.765 62.725 -132.435 ;
        RECT 62.395 -134.125 62.725 -133.795 ;
        RECT 62.395 -135.485 62.725 -135.155 ;
        RECT 62.395 -136.845 62.725 -136.515 ;
        RECT 62.395 -138.205 62.725 -137.875 ;
        RECT 62.395 -139.565 62.725 -139.235 ;
        RECT 62.395 -140.925 62.725 -140.595 ;
        RECT 62.395 -142.285 62.725 -141.955 ;
        RECT 62.395 -143.645 62.725 -143.315 ;
        RECT 62.395 -145.005 62.725 -144.675 ;
        RECT 62.395 -146.365 62.725 -146.035 ;
        RECT 62.395 -147.725 62.725 -147.395 ;
        RECT 62.395 -149.085 62.725 -148.755 ;
        RECT 62.395 -150.445 62.725 -150.115 ;
        RECT 62.395 -151.805 62.725 -151.475 ;
        RECT 62.395 -153.165 62.725 -152.835 ;
        RECT 62.395 -154.525 62.725 -154.195 ;
        RECT 62.395 -155.885 62.725 -155.555 ;
        RECT 62.395 -157.245 62.725 -156.915 ;
        RECT 62.395 -158.605 62.725 -158.275 ;
        RECT 62.395 -159.965 62.725 -159.635 ;
        RECT 62.395 -161.325 62.725 -160.995 ;
        RECT 62.395 -162.685 62.725 -162.355 ;
        RECT 62.395 -164.045 62.725 -163.715 ;
        RECT 62.395 -165.405 62.725 -165.075 ;
        RECT 62.395 -166.765 62.725 -166.435 ;
        RECT 62.395 -168.125 62.725 -167.795 ;
        RECT 62.395 -169.485 62.725 -169.155 ;
        RECT 62.395 -170.845 62.725 -170.515 ;
        RECT 62.395 -172.205 62.725 -171.875 ;
        RECT 62.395 -173.565 62.725 -173.235 ;
        RECT 62.395 -174.925 62.725 -174.595 ;
        RECT 62.395 -176.285 62.725 -175.955 ;
        RECT 62.395 -177.645 62.725 -177.315 ;
        RECT 62.395 -179.005 62.725 -178.675 ;
        RECT 62.395 -184.65 62.725 -183.52 ;
        RECT 62.4 -184.765 62.72 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 244.04 64.085 245.17 ;
        RECT 63.755 239.875 64.085 240.205 ;
        RECT 63.755 238.515 64.085 238.845 ;
        RECT 63.755 237.155 64.085 237.485 ;
        RECT 63.76 237.155 64.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 -0.845 64.085 -0.515 ;
        RECT 63.755 -2.205 64.085 -1.875 ;
        RECT 63.755 -3.565 64.085 -3.235 ;
        RECT 63.76 -3.565 64.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.755 -96.045 64.085 -95.715 ;
        RECT 63.755 -97.405 64.085 -97.075 ;
        RECT 63.755 -98.765 64.085 -98.435 ;
        RECT 63.755 -100.125 64.085 -99.795 ;
        RECT 63.755 -101.485 64.085 -101.155 ;
        RECT 63.755 -102.845 64.085 -102.515 ;
        RECT 63.755 -104.205 64.085 -103.875 ;
        RECT 63.755 -105.565 64.085 -105.235 ;
        RECT 63.755 -106.925 64.085 -106.595 ;
        RECT 63.755 -108.285 64.085 -107.955 ;
        RECT 63.755 -109.645 64.085 -109.315 ;
        RECT 63.755 -111.005 64.085 -110.675 ;
        RECT 63.755 -112.365 64.085 -112.035 ;
        RECT 63.755 -113.725 64.085 -113.395 ;
        RECT 63.755 -115.085 64.085 -114.755 ;
        RECT 63.755 -116.445 64.085 -116.115 ;
        RECT 63.755 -117.805 64.085 -117.475 ;
        RECT 63.755 -119.165 64.085 -118.835 ;
        RECT 63.755 -120.525 64.085 -120.195 ;
        RECT 63.755 -121.885 64.085 -121.555 ;
        RECT 63.755 -123.245 64.085 -122.915 ;
        RECT 63.755 -124.605 64.085 -124.275 ;
        RECT 63.755 -125.965 64.085 -125.635 ;
        RECT 63.755 -127.325 64.085 -126.995 ;
        RECT 63.755 -128.685 64.085 -128.355 ;
        RECT 63.755 -130.045 64.085 -129.715 ;
        RECT 63.755 -131.405 64.085 -131.075 ;
        RECT 63.755 -132.765 64.085 -132.435 ;
        RECT 63.755 -134.125 64.085 -133.795 ;
        RECT 63.755 -135.485 64.085 -135.155 ;
        RECT 63.755 -136.845 64.085 -136.515 ;
        RECT 63.755 -138.205 64.085 -137.875 ;
        RECT 63.755 -139.565 64.085 -139.235 ;
        RECT 63.755 -140.925 64.085 -140.595 ;
        RECT 63.755 -142.285 64.085 -141.955 ;
        RECT 63.755 -143.645 64.085 -143.315 ;
        RECT 63.755 -145.005 64.085 -144.675 ;
        RECT 63.755 -146.365 64.085 -146.035 ;
        RECT 63.755 -147.725 64.085 -147.395 ;
        RECT 63.755 -149.085 64.085 -148.755 ;
        RECT 63.755 -150.445 64.085 -150.115 ;
        RECT 63.755 -151.805 64.085 -151.475 ;
        RECT 63.755 -153.165 64.085 -152.835 ;
        RECT 63.755 -154.525 64.085 -154.195 ;
        RECT 63.755 -155.885 64.085 -155.555 ;
        RECT 63.755 -157.245 64.085 -156.915 ;
        RECT 63.755 -158.605 64.085 -158.275 ;
        RECT 63.755 -159.965 64.085 -159.635 ;
        RECT 63.755 -161.325 64.085 -160.995 ;
        RECT 63.755 -162.685 64.085 -162.355 ;
        RECT 63.755 -164.045 64.085 -163.715 ;
        RECT 63.755 -165.405 64.085 -165.075 ;
        RECT 63.755 -166.765 64.085 -166.435 ;
        RECT 63.755 -168.125 64.085 -167.795 ;
        RECT 63.755 -169.485 64.085 -169.155 ;
        RECT 63.755 -170.845 64.085 -170.515 ;
        RECT 63.755 -172.205 64.085 -171.875 ;
        RECT 63.755 -173.565 64.085 -173.235 ;
        RECT 63.755 -174.925 64.085 -174.595 ;
        RECT 63.755 -176.285 64.085 -175.955 ;
        RECT 63.755 -177.645 64.085 -177.315 ;
        RECT 63.755 -179.005 64.085 -178.675 ;
        RECT 63.755 -184.65 64.085 -183.52 ;
        RECT 63.76 -184.765 64.08 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 244.04 65.445 245.17 ;
        RECT 65.115 239.875 65.445 240.205 ;
        RECT 65.115 238.515 65.445 238.845 ;
        RECT 65.115 237.155 65.445 237.485 ;
        RECT 65.12 237.155 65.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 -0.845 65.445 -0.515 ;
        RECT 65.115 -2.205 65.445 -1.875 ;
        RECT 65.115 -3.565 65.445 -3.235 ;
        RECT 65.12 -3.565 65.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.115 -96.045 65.445 -95.715 ;
        RECT 65.115 -97.405 65.445 -97.075 ;
        RECT 65.115 -98.765 65.445 -98.435 ;
        RECT 65.115 -100.125 65.445 -99.795 ;
        RECT 65.115 -101.485 65.445 -101.155 ;
        RECT 65.115 -102.845 65.445 -102.515 ;
        RECT 65.115 -104.205 65.445 -103.875 ;
        RECT 65.115 -105.565 65.445 -105.235 ;
        RECT 65.115 -106.925 65.445 -106.595 ;
        RECT 65.115 -108.285 65.445 -107.955 ;
        RECT 65.115 -109.645 65.445 -109.315 ;
        RECT 65.115 -111.005 65.445 -110.675 ;
        RECT 65.115 -112.365 65.445 -112.035 ;
        RECT 65.115 -113.725 65.445 -113.395 ;
        RECT 65.115 -115.085 65.445 -114.755 ;
        RECT 65.115 -116.445 65.445 -116.115 ;
        RECT 65.115 -117.805 65.445 -117.475 ;
        RECT 65.115 -119.165 65.445 -118.835 ;
        RECT 65.115 -120.525 65.445 -120.195 ;
        RECT 65.115 -121.885 65.445 -121.555 ;
        RECT 65.115 -123.245 65.445 -122.915 ;
        RECT 65.115 -124.605 65.445 -124.275 ;
        RECT 65.115 -125.965 65.445 -125.635 ;
        RECT 65.115 -127.325 65.445 -126.995 ;
        RECT 65.115 -128.685 65.445 -128.355 ;
        RECT 65.115 -130.045 65.445 -129.715 ;
        RECT 65.115 -131.405 65.445 -131.075 ;
        RECT 65.115 -132.765 65.445 -132.435 ;
        RECT 65.115 -134.125 65.445 -133.795 ;
        RECT 65.115 -135.485 65.445 -135.155 ;
        RECT 65.115 -136.845 65.445 -136.515 ;
        RECT 65.115 -138.205 65.445 -137.875 ;
        RECT 65.115 -139.565 65.445 -139.235 ;
        RECT 65.115 -140.925 65.445 -140.595 ;
        RECT 65.115 -142.285 65.445 -141.955 ;
        RECT 65.115 -143.645 65.445 -143.315 ;
        RECT 65.115 -145.005 65.445 -144.675 ;
        RECT 65.115 -146.365 65.445 -146.035 ;
        RECT 65.115 -147.725 65.445 -147.395 ;
        RECT 65.115 -149.085 65.445 -148.755 ;
        RECT 65.115 -150.445 65.445 -150.115 ;
        RECT 65.115 -151.805 65.445 -151.475 ;
        RECT 65.115 -153.165 65.445 -152.835 ;
        RECT 65.115 -154.525 65.445 -154.195 ;
        RECT 65.115 -155.885 65.445 -155.555 ;
        RECT 65.115 -157.245 65.445 -156.915 ;
        RECT 65.115 -158.605 65.445 -158.275 ;
        RECT 65.115 -159.965 65.445 -159.635 ;
        RECT 65.115 -161.325 65.445 -160.995 ;
        RECT 65.115 -162.685 65.445 -162.355 ;
        RECT 65.115 -164.045 65.445 -163.715 ;
        RECT 65.115 -165.405 65.445 -165.075 ;
        RECT 65.115 -166.765 65.445 -166.435 ;
        RECT 65.115 -168.125 65.445 -167.795 ;
        RECT 65.115 -169.485 65.445 -169.155 ;
        RECT 65.115 -170.845 65.445 -170.515 ;
        RECT 65.115 -172.205 65.445 -171.875 ;
        RECT 65.115 -173.565 65.445 -173.235 ;
        RECT 65.115 -174.925 65.445 -174.595 ;
        RECT 65.115 -176.285 65.445 -175.955 ;
        RECT 65.115 -177.645 65.445 -177.315 ;
        RECT 65.115 -179.005 65.445 -178.675 ;
        RECT 65.115 -184.65 65.445 -183.52 ;
        RECT 65.12 -184.765 65.44 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 244.04 66.805 245.17 ;
        RECT 66.475 239.875 66.805 240.205 ;
        RECT 66.475 238.515 66.805 238.845 ;
        RECT 66.475 237.155 66.805 237.485 ;
        RECT 66.48 237.155 66.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 -0.845 66.805 -0.515 ;
        RECT 66.475 -2.205 66.805 -1.875 ;
        RECT 66.475 -3.565 66.805 -3.235 ;
        RECT 66.48 -3.565 66.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 66.475 -96.045 66.805 -95.715 ;
        RECT 66.475 -97.405 66.805 -97.075 ;
        RECT 66.475 -98.765 66.805 -98.435 ;
        RECT 66.475 -100.125 66.805 -99.795 ;
        RECT 66.475 -101.485 66.805 -101.155 ;
        RECT 66.475 -102.845 66.805 -102.515 ;
        RECT 66.475 -104.205 66.805 -103.875 ;
        RECT 66.475 -105.565 66.805 -105.235 ;
        RECT 66.475 -106.925 66.805 -106.595 ;
        RECT 66.475 -108.285 66.805 -107.955 ;
        RECT 66.475 -109.645 66.805 -109.315 ;
        RECT 66.475 -111.005 66.805 -110.675 ;
        RECT 66.475 -112.365 66.805 -112.035 ;
        RECT 66.475 -113.725 66.805 -113.395 ;
        RECT 66.475 -115.085 66.805 -114.755 ;
        RECT 66.475 -116.445 66.805 -116.115 ;
        RECT 66.475 -117.805 66.805 -117.475 ;
        RECT 66.475 -119.165 66.805 -118.835 ;
        RECT 66.475 -120.525 66.805 -120.195 ;
        RECT 66.475 -121.885 66.805 -121.555 ;
        RECT 66.475 -123.245 66.805 -122.915 ;
        RECT 66.475 -124.605 66.805 -124.275 ;
        RECT 66.475 -125.965 66.805 -125.635 ;
        RECT 66.475 -127.325 66.805 -126.995 ;
        RECT 66.475 -128.685 66.805 -128.355 ;
        RECT 66.475 -130.045 66.805 -129.715 ;
        RECT 66.475 -131.405 66.805 -131.075 ;
        RECT 66.475 -132.765 66.805 -132.435 ;
        RECT 66.475 -134.125 66.805 -133.795 ;
        RECT 66.475 -135.485 66.805 -135.155 ;
        RECT 66.475 -136.845 66.805 -136.515 ;
        RECT 66.475 -138.205 66.805 -137.875 ;
        RECT 66.475 -139.565 66.805 -139.235 ;
        RECT 66.475 -140.925 66.805 -140.595 ;
        RECT 66.475 -142.285 66.805 -141.955 ;
        RECT 66.475 -143.645 66.805 -143.315 ;
        RECT 66.475 -145.005 66.805 -144.675 ;
        RECT 66.475 -146.365 66.805 -146.035 ;
        RECT 66.475 -147.725 66.805 -147.395 ;
        RECT 66.475 -149.085 66.805 -148.755 ;
        RECT 66.475 -150.445 66.805 -150.115 ;
        RECT 66.475 -151.805 66.805 -151.475 ;
        RECT 66.475 -153.165 66.805 -152.835 ;
        RECT 66.475 -154.525 66.805 -154.195 ;
        RECT 66.475 -155.885 66.805 -155.555 ;
        RECT 66.475 -157.245 66.805 -156.915 ;
        RECT 66.475 -158.605 66.805 -158.275 ;
        RECT 66.475 -159.965 66.805 -159.635 ;
        RECT 66.475 -161.325 66.805 -160.995 ;
        RECT 66.475 -162.685 66.805 -162.355 ;
        RECT 66.475 -164.045 66.805 -163.715 ;
        RECT 66.475 -165.405 66.805 -165.075 ;
        RECT 66.475 -166.765 66.805 -166.435 ;
        RECT 66.475 -168.125 66.805 -167.795 ;
        RECT 66.475 -169.485 66.805 -169.155 ;
        RECT 66.475 -170.845 66.805 -170.515 ;
        RECT 66.475 -172.205 66.805 -171.875 ;
        RECT 66.475 -173.565 66.805 -173.235 ;
        RECT 66.475 -174.925 66.805 -174.595 ;
        RECT 66.475 -176.285 66.805 -175.955 ;
        RECT 66.475 -177.645 66.805 -177.315 ;
        RECT 66.475 -179.005 66.805 -178.675 ;
        RECT 66.475 -184.65 66.805 -183.52 ;
        RECT 66.48 -184.765 66.8 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 244.04 68.165 245.17 ;
        RECT 67.835 239.875 68.165 240.205 ;
        RECT 67.835 238.515 68.165 238.845 ;
        RECT 67.835 237.155 68.165 237.485 ;
        RECT 67.84 237.155 68.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.835 -98.765 68.165 -98.435 ;
        RECT 67.835 -100.125 68.165 -99.795 ;
        RECT 67.835 -101.485 68.165 -101.155 ;
        RECT 67.835 -102.845 68.165 -102.515 ;
        RECT 67.835 -104.205 68.165 -103.875 ;
        RECT 67.835 -105.565 68.165 -105.235 ;
        RECT 67.835 -106.925 68.165 -106.595 ;
        RECT 67.835 -108.285 68.165 -107.955 ;
        RECT 67.835 -109.645 68.165 -109.315 ;
        RECT 67.835 -111.005 68.165 -110.675 ;
        RECT 67.835 -112.365 68.165 -112.035 ;
        RECT 67.835 -113.725 68.165 -113.395 ;
        RECT 67.835 -115.085 68.165 -114.755 ;
        RECT 67.835 -116.445 68.165 -116.115 ;
        RECT 67.835 -117.805 68.165 -117.475 ;
        RECT 67.835 -119.165 68.165 -118.835 ;
        RECT 67.835 -120.525 68.165 -120.195 ;
        RECT 67.835 -121.885 68.165 -121.555 ;
        RECT 67.835 -123.245 68.165 -122.915 ;
        RECT 67.835 -124.605 68.165 -124.275 ;
        RECT 67.835 -125.965 68.165 -125.635 ;
        RECT 67.835 -127.325 68.165 -126.995 ;
        RECT 67.835 -128.685 68.165 -128.355 ;
        RECT 67.835 -130.045 68.165 -129.715 ;
        RECT 67.835 -131.405 68.165 -131.075 ;
        RECT 67.835 -132.765 68.165 -132.435 ;
        RECT 67.835 -134.125 68.165 -133.795 ;
        RECT 67.835 -135.485 68.165 -135.155 ;
        RECT 67.835 -136.845 68.165 -136.515 ;
        RECT 67.835 -138.205 68.165 -137.875 ;
        RECT 67.835 -139.565 68.165 -139.235 ;
        RECT 67.835 -140.925 68.165 -140.595 ;
        RECT 67.835 -142.285 68.165 -141.955 ;
        RECT 67.835 -143.645 68.165 -143.315 ;
        RECT 67.835 -145.005 68.165 -144.675 ;
        RECT 67.835 -146.365 68.165 -146.035 ;
        RECT 67.835 -147.725 68.165 -147.395 ;
        RECT 67.835 -149.085 68.165 -148.755 ;
        RECT 67.835 -150.445 68.165 -150.115 ;
        RECT 67.835 -151.805 68.165 -151.475 ;
        RECT 67.835 -153.165 68.165 -152.835 ;
        RECT 67.835 -154.525 68.165 -154.195 ;
        RECT 67.835 -155.885 68.165 -155.555 ;
        RECT 67.835 -157.245 68.165 -156.915 ;
        RECT 67.835 -158.605 68.165 -158.275 ;
        RECT 67.835 -159.965 68.165 -159.635 ;
        RECT 67.835 -161.325 68.165 -160.995 ;
        RECT 67.835 -162.685 68.165 -162.355 ;
        RECT 67.835 -164.045 68.165 -163.715 ;
        RECT 67.835 -165.405 68.165 -165.075 ;
        RECT 67.835 -166.765 68.165 -166.435 ;
        RECT 67.835 -168.125 68.165 -167.795 ;
        RECT 67.835 -169.485 68.165 -169.155 ;
        RECT 67.835 -170.845 68.165 -170.515 ;
        RECT 67.835 -172.205 68.165 -171.875 ;
        RECT 67.835 -173.565 68.165 -173.235 ;
        RECT 67.835 -174.925 68.165 -174.595 ;
        RECT 67.835 -176.285 68.165 -175.955 ;
        RECT 67.835 -177.645 68.165 -177.315 ;
        RECT 67.835 -179.005 68.165 -178.675 ;
        RECT 67.835 -184.65 68.165 -183.52 ;
        RECT 67.84 -184.765 68.16 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.06 -98.075 68.39 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.195 244.04 69.525 245.17 ;
        RECT 69.195 239.875 69.525 240.205 ;
        RECT 69.195 238.515 69.525 238.845 ;
        RECT 69.195 237.155 69.525 237.485 ;
        RECT 69.2 237.155 69.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.555 244.04 70.885 245.17 ;
        RECT 70.555 239.875 70.885 240.205 ;
        RECT 70.555 238.515 70.885 238.845 ;
        RECT 70.555 237.155 70.885 237.485 ;
        RECT 70.56 237.155 70.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 70.555 -0.845 70.885 -0.515 ;
        RECT 70.555 -2.205 70.885 -1.875 ;
        RECT 70.555 -3.565 70.885 -3.235 ;
        RECT 70.56 -3.565 70.88 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 244.04 72.245 245.17 ;
        RECT 71.915 239.875 72.245 240.205 ;
        RECT 71.915 238.515 72.245 238.845 ;
        RECT 71.915 237.155 72.245 237.485 ;
        RECT 71.92 237.155 72.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 -0.845 72.245 -0.515 ;
        RECT 71.915 -2.205 72.245 -1.875 ;
        RECT 71.915 -3.565 72.245 -3.235 ;
        RECT 71.92 -3.565 72.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.915 -96.045 72.245 -95.715 ;
        RECT 71.915 -97.405 72.245 -97.075 ;
        RECT 71.915 -98.765 72.245 -98.435 ;
        RECT 71.915 -100.125 72.245 -99.795 ;
        RECT 71.915 -101.485 72.245 -101.155 ;
        RECT 71.915 -102.845 72.245 -102.515 ;
        RECT 71.915 -104.205 72.245 -103.875 ;
        RECT 71.915 -105.565 72.245 -105.235 ;
        RECT 71.915 -106.925 72.245 -106.595 ;
        RECT 71.915 -108.285 72.245 -107.955 ;
        RECT 71.915 -109.645 72.245 -109.315 ;
        RECT 71.915 -111.005 72.245 -110.675 ;
        RECT 71.915 -112.365 72.245 -112.035 ;
        RECT 71.915 -113.725 72.245 -113.395 ;
        RECT 71.915 -115.085 72.245 -114.755 ;
        RECT 71.915 -116.445 72.245 -116.115 ;
        RECT 71.915 -117.805 72.245 -117.475 ;
        RECT 71.915 -119.165 72.245 -118.835 ;
        RECT 71.915 -120.525 72.245 -120.195 ;
        RECT 71.915 -121.885 72.245 -121.555 ;
        RECT 71.915 -123.245 72.245 -122.915 ;
        RECT 71.915 -124.605 72.245 -124.275 ;
        RECT 71.915 -125.965 72.245 -125.635 ;
        RECT 71.915 -127.325 72.245 -126.995 ;
        RECT 71.915 -128.685 72.245 -128.355 ;
        RECT 71.915 -130.045 72.245 -129.715 ;
        RECT 71.915 -131.405 72.245 -131.075 ;
        RECT 71.915 -132.765 72.245 -132.435 ;
        RECT 71.915 -134.125 72.245 -133.795 ;
        RECT 71.915 -135.485 72.245 -135.155 ;
        RECT 71.915 -136.845 72.245 -136.515 ;
        RECT 71.915 -138.205 72.245 -137.875 ;
        RECT 71.915 -139.565 72.245 -139.235 ;
        RECT 71.915 -140.925 72.245 -140.595 ;
        RECT 71.915 -142.285 72.245 -141.955 ;
        RECT 71.915 -143.645 72.245 -143.315 ;
        RECT 71.915 -145.005 72.245 -144.675 ;
        RECT 71.915 -146.365 72.245 -146.035 ;
        RECT 71.915 -147.725 72.245 -147.395 ;
        RECT 71.915 -149.085 72.245 -148.755 ;
        RECT 71.915 -150.445 72.245 -150.115 ;
        RECT 71.915 -151.805 72.245 -151.475 ;
        RECT 71.915 -153.165 72.245 -152.835 ;
        RECT 71.915 -154.525 72.245 -154.195 ;
        RECT 71.915 -155.885 72.245 -155.555 ;
        RECT 71.915 -157.245 72.245 -156.915 ;
        RECT 71.915 -158.605 72.245 -158.275 ;
        RECT 71.915 -159.965 72.245 -159.635 ;
        RECT 71.915 -161.325 72.245 -160.995 ;
        RECT 71.915 -162.685 72.245 -162.355 ;
        RECT 71.915 -164.045 72.245 -163.715 ;
        RECT 71.915 -165.405 72.245 -165.075 ;
        RECT 71.915 -166.765 72.245 -166.435 ;
        RECT 71.915 -168.125 72.245 -167.795 ;
        RECT 71.915 -169.485 72.245 -169.155 ;
        RECT 71.915 -170.845 72.245 -170.515 ;
        RECT 71.915 -172.205 72.245 -171.875 ;
        RECT 71.915 -173.565 72.245 -173.235 ;
        RECT 71.915 -174.925 72.245 -174.595 ;
        RECT 71.915 -176.285 72.245 -175.955 ;
        RECT 71.915 -177.645 72.245 -177.315 ;
        RECT 71.915 -179.005 72.245 -178.675 ;
        RECT 71.915 -184.65 72.245 -183.52 ;
        RECT 71.92 -184.765 72.24 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 244.04 73.605 245.17 ;
        RECT 73.275 239.875 73.605 240.205 ;
        RECT 73.275 238.515 73.605 238.845 ;
        RECT 73.275 237.155 73.605 237.485 ;
        RECT 73.28 237.155 73.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 -0.845 73.605 -0.515 ;
        RECT 73.275 -2.205 73.605 -1.875 ;
        RECT 73.275 -3.565 73.605 -3.235 ;
        RECT 73.28 -3.565 73.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.275 -96.045 73.605 -95.715 ;
        RECT 73.275 -97.405 73.605 -97.075 ;
        RECT 73.275 -98.765 73.605 -98.435 ;
        RECT 73.275 -100.125 73.605 -99.795 ;
        RECT 73.275 -101.485 73.605 -101.155 ;
        RECT 73.275 -102.845 73.605 -102.515 ;
        RECT 73.275 -104.205 73.605 -103.875 ;
        RECT 73.275 -105.565 73.605 -105.235 ;
        RECT 73.275 -106.925 73.605 -106.595 ;
        RECT 73.275 -108.285 73.605 -107.955 ;
        RECT 73.275 -109.645 73.605 -109.315 ;
        RECT 73.275 -111.005 73.605 -110.675 ;
        RECT 73.275 -112.365 73.605 -112.035 ;
        RECT 73.275 -113.725 73.605 -113.395 ;
        RECT 73.275 -115.085 73.605 -114.755 ;
        RECT 73.275 -116.445 73.605 -116.115 ;
        RECT 73.275 -117.805 73.605 -117.475 ;
        RECT 73.275 -119.165 73.605 -118.835 ;
        RECT 73.275 -120.525 73.605 -120.195 ;
        RECT 73.275 -121.885 73.605 -121.555 ;
        RECT 73.275 -123.245 73.605 -122.915 ;
        RECT 73.275 -124.605 73.605 -124.275 ;
        RECT 73.275 -125.965 73.605 -125.635 ;
        RECT 73.275 -127.325 73.605 -126.995 ;
        RECT 73.275 -128.685 73.605 -128.355 ;
        RECT 73.275 -130.045 73.605 -129.715 ;
        RECT 73.275 -131.405 73.605 -131.075 ;
        RECT 73.275 -132.765 73.605 -132.435 ;
        RECT 73.275 -134.125 73.605 -133.795 ;
        RECT 73.275 -135.485 73.605 -135.155 ;
        RECT 73.275 -136.845 73.605 -136.515 ;
        RECT 73.275 -138.205 73.605 -137.875 ;
        RECT 73.275 -139.565 73.605 -139.235 ;
        RECT 73.275 -140.925 73.605 -140.595 ;
        RECT 73.275 -142.285 73.605 -141.955 ;
        RECT 73.275 -143.645 73.605 -143.315 ;
        RECT 73.275 -145.005 73.605 -144.675 ;
        RECT 73.275 -146.365 73.605 -146.035 ;
        RECT 73.275 -147.725 73.605 -147.395 ;
        RECT 73.275 -149.085 73.605 -148.755 ;
        RECT 73.275 -150.445 73.605 -150.115 ;
        RECT 73.275 -151.805 73.605 -151.475 ;
        RECT 73.275 -153.165 73.605 -152.835 ;
        RECT 73.275 -154.525 73.605 -154.195 ;
        RECT 73.275 -155.885 73.605 -155.555 ;
        RECT 73.275 -157.245 73.605 -156.915 ;
        RECT 73.275 -158.605 73.605 -158.275 ;
        RECT 73.275 -159.965 73.605 -159.635 ;
        RECT 73.275 -161.325 73.605 -160.995 ;
        RECT 73.275 -162.685 73.605 -162.355 ;
        RECT 73.275 -164.045 73.605 -163.715 ;
        RECT 73.275 -165.405 73.605 -165.075 ;
        RECT 73.275 -166.765 73.605 -166.435 ;
        RECT 73.275 -168.125 73.605 -167.795 ;
        RECT 73.275 -169.485 73.605 -169.155 ;
        RECT 73.275 -170.845 73.605 -170.515 ;
        RECT 73.275 -172.205 73.605 -171.875 ;
        RECT 73.275 -173.565 73.605 -173.235 ;
        RECT 73.275 -174.925 73.605 -174.595 ;
        RECT 73.275 -176.285 73.605 -175.955 ;
        RECT 73.275 -177.645 73.605 -177.315 ;
        RECT 73.275 -179.005 73.605 -178.675 ;
        RECT 73.275 -184.65 73.605 -183.52 ;
        RECT 73.28 -184.765 73.6 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 244.04 74.965 245.17 ;
        RECT 74.635 239.875 74.965 240.205 ;
        RECT 74.635 238.515 74.965 238.845 ;
        RECT 74.635 237.155 74.965 237.485 ;
        RECT 74.64 237.155 74.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 -0.845 74.965 -0.515 ;
        RECT 74.635 -2.205 74.965 -1.875 ;
        RECT 74.635 -3.565 74.965 -3.235 ;
        RECT 74.64 -3.565 74.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 74.635 -96.045 74.965 -95.715 ;
        RECT 74.635 -97.405 74.965 -97.075 ;
        RECT 74.635 -98.765 74.965 -98.435 ;
        RECT 74.635 -100.125 74.965 -99.795 ;
        RECT 74.635 -101.485 74.965 -101.155 ;
        RECT 74.635 -102.845 74.965 -102.515 ;
        RECT 74.635 -104.205 74.965 -103.875 ;
        RECT 74.635 -105.565 74.965 -105.235 ;
        RECT 74.635 -106.925 74.965 -106.595 ;
        RECT 74.635 -108.285 74.965 -107.955 ;
        RECT 74.635 -109.645 74.965 -109.315 ;
        RECT 74.635 -111.005 74.965 -110.675 ;
        RECT 74.635 -112.365 74.965 -112.035 ;
        RECT 74.635 -113.725 74.965 -113.395 ;
        RECT 74.635 -115.085 74.965 -114.755 ;
        RECT 74.635 -116.445 74.965 -116.115 ;
        RECT 74.635 -117.805 74.965 -117.475 ;
        RECT 74.635 -119.165 74.965 -118.835 ;
        RECT 74.635 -120.525 74.965 -120.195 ;
        RECT 74.635 -121.885 74.965 -121.555 ;
        RECT 74.635 -123.245 74.965 -122.915 ;
        RECT 74.635 -124.605 74.965 -124.275 ;
        RECT 74.635 -125.965 74.965 -125.635 ;
        RECT 74.635 -127.325 74.965 -126.995 ;
        RECT 74.635 -128.685 74.965 -128.355 ;
        RECT 74.635 -130.045 74.965 -129.715 ;
        RECT 74.635 -131.405 74.965 -131.075 ;
        RECT 74.635 -132.765 74.965 -132.435 ;
        RECT 74.635 -134.125 74.965 -133.795 ;
        RECT 74.635 -135.485 74.965 -135.155 ;
        RECT 74.635 -136.845 74.965 -136.515 ;
        RECT 74.635 -138.205 74.965 -137.875 ;
        RECT 74.635 -139.565 74.965 -139.235 ;
        RECT 74.635 -140.925 74.965 -140.595 ;
        RECT 74.635 -142.285 74.965 -141.955 ;
        RECT 74.635 -143.645 74.965 -143.315 ;
        RECT 74.635 -145.005 74.965 -144.675 ;
        RECT 74.635 -146.365 74.965 -146.035 ;
        RECT 74.635 -147.725 74.965 -147.395 ;
        RECT 74.635 -149.085 74.965 -148.755 ;
        RECT 74.635 -150.445 74.965 -150.115 ;
        RECT 74.635 -151.805 74.965 -151.475 ;
        RECT 74.635 -153.165 74.965 -152.835 ;
        RECT 74.635 -154.525 74.965 -154.195 ;
        RECT 74.635 -155.885 74.965 -155.555 ;
        RECT 74.635 -157.245 74.965 -156.915 ;
        RECT 74.635 -158.605 74.965 -158.275 ;
        RECT 74.635 -159.965 74.965 -159.635 ;
        RECT 74.635 -161.325 74.965 -160.995 ;
        RECT 74.635 -162.685 74.965 -162.355 ;
        RECT 74.635 -164.045 74.965 -163.715 ;
        RECT 74.635 -165.405 74.965 -165.075 ;
        RECT 74.635 -166.765 74.965 -166.435 ;
        RECT 74.635 -168.125 74.965 -167.795 ;
        RECT 74.635 -169.485 74.965 -169.155 ;
        RECT 74.635 -170.845 74.965 -170.515 ;
        RECT 74.635 -172.205 74.965 -171.875 ;
        RECT 74.635 -173.565 74.965 -173.235 ;
        RECT 74.635 -174.925 74.965 -174.595 ;
        RECT 74.635 -176.285 74.965 -175.955 ;
        RECT 74.635 -177.645 74.965 -177.315 ;
        RECT 74.635 -179.005 74.965 -178.675 ;
        RECT 74.635 -184.65 74.965 -183.52 ;
        RECT 74.64 -184.765 74.96 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 244.04 76.325 245.17 ;
        RECT 75.995 239.875 76.325 240.205 ;
        RECT 75.995 238.515 76.325 238.845 ;
        RECT 75.995 237.155 76.325 237.485 ;
        RECT 76 237.155 76.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 -0.845 76.325 -0.515 ;
        RECT 75.995 -2.205 76.325 -1.875 ;
        RECT 75.995 -3.565 76.325 -3.235 ;
        RECT 76 -3.565 76.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.995 -96.045 76.325 -95.715 ;
        RECT 75.995 -97.405 76.325 -97.075 ;
        RECT 75.995 -98.765 76.325 -98.435 ;
        RECT 75.995 -100.125 76.325 -99.795 ;
        RECT 75.995 -101.485 76.325 -101.155 ;
        RECT 75.995 -102.845 76.325 -102.515 ;
        RECT 75.995 -104.205 76.325 -103.875 ;
        RECT 75.995 -105.565 76.325 -105.235 ;
        RECT 75.995 -106.925 76.325 -106.595 ;
        RECT 75.995 -108.285 76.325 -107.955 ;
        RECT 75.995 -109.645 76.325 -109.315 ;
        RECT 75.995 -111.005 76.325 -110.675 ;
        RECT 75.995 -112.365 76.325 -112.035 ;
        RECT 75.995 -113.725 76.325 -113.395 ;
        RECT 75.995 -115.085 76.325 -114.755 ;
        RECT 75.995 -116.445 76.325 -116.115 ;
        RECT 75.995 -117.805 76.325 -117.475 ;
        RECT 75.995 -119.165 76.325 -118.835 ;
        RECT 75.995 -120.525 76.325 -120.195 ;
        RECT 75.995 -121.885 76.325 -121.555 ;
        RECT 75.995 -123.245 76.325 -122.915 ;
        RECT 75.995 -124.605 76.325 -124.275 ;
        RECT 75.995 -125.965 76.325 -125.635 ;
        RECT 75.995 -127.325 76.325 -126.995 ;
        RECT 75.995 -128.685 76.325 -128.355 ;
        RECT 75.995 -130.045 76.325 -129.715 ;
        RECT 75.995 -131.405 76.325 -131.075 ;
        RECT 75.995 -132.765 76.325 -132.435 ;
        RECT 75.995 -134.125 76.325 -133.795 ;
        RECT 75.995 -135.485 76.325 -135.155 ;
        RECT 75.995 -136.845 76.325 -136.515 ;
        RECT 75.995 -138.205 76.325 -137.875 ;
        RECT 75.995 -139.565 76.325 -139.235 ;
        RECT 75.995 -140.925 76.325 -140.595 ;
        RECT 75.995 -142.285 76.325 -141.955 ;
        RECT 75.995 -143.645 76.325 -143.315 ;
        RECT 75.995 -145.005 76.325 -144.675 ;
        RECT 75.995 -146.365 76.325 -146.035 ;
        RECT 75.995 -147.725 76.325 -147.395 ;
        RECT 75.995 -149.085 76.325 -148.755 ;
        RECT 75.995 -150.445 76.325 -150.115 ;
        RECT 75.995 -151.805 76.325 -151.475 ;
        RECT 75.995 -153.165 76.325 -152.835 ;
        RECT 75.995 -154.525 76.325 -154.195 ;
        RECT 75.995 -155.885 76.325 -155.555 ;
        RECT 75.995 -157.245 76.325 -156.915 ;
        RECT 75.995 -158.605 76.325 -158.275 ;
        RECT 75.995 -159.965 76.325 -159.635 ;
        RECT 75.995 -161.325 76.325 -160.995 ;
        RECT 75.995 -162.685 76.325 -162.355 ;
        RECT 75.995 -164.045 76.325 -163.715 ;
        RECT 75.995 -165.405 76.325 -165.075 ;
        RECT 75.995 -166.765 76.325 -166.435 ;
        RECT 75.995 -168.125 76.325 -167.795 ;
        RECT 75.995 -169.485 76.325 -169.155 ;
        RECT 75.995 -170.845 76.325 -170.515 ;
        RECT 75.995 -172.205 76.325 -171.875 ;
        RECT 75.995 -173.565 76.325 -173.235 ;
        RECT 75.995 -174.925 76.325 -174.595 ;
        RECT 75.995 -176.285 76.325 -175.955 ;
        RECT 75.995 -177.645 76.325 -177.315 ;
        RECT 75.995 -179.005 76.325 -178.675 ;
        RECT 75.995 -184.65 76.325 -183.52 ;
        RECT 76 -184.765 76.32 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 244.04 77.685 245.17 ;
        RECT 77.355 239.875 77.685 240.205 ;
        RECT 77.355 238.515 77.685 238.845 ;
        RECT 77.355 237.155 77.685 237.485 ;
        RECT 77.36 237.155 77.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 -0.845 77.685 -0.515 ;
        RECT 77.355 -2.205 77.685 -1.875 ;
        RECT 77.355 -3.565 77.685 -3.235 ;
        RECT 77.36 -3.565 77.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 77.355 -96.045 77.685 -95.715 ;
        RECT 77.355 -97.405 77.685 -97.075 ;
        RECT 77.355 -98.765 77.685 -98.435 ;
        RECT 77.355 -100.125 77.685 -99.795 ;
        RECT 77.355 -101.485 77.685 -101.155 ;
        RECT 77.355 -102.845 77.685 -102.515 ;
        RECT 77.355 -104.205 77.685 -103.875 ;
        RECT 77.355 -105.565 77.685 -105.235 ;
        RECT 77.355 -106.925 77.685 -106.595 ;
        RECT 77.355 -108.285 77.685 -107.955 ;
        RECT 77.355 -109.645 77.685 -109.315 ;
        RECT 77.355 -111.005 77.685 -110.675 ;
        RECT 77.355 -112.365 77.685 -112.035 ;
        RECT 77.355 -113.725 77.685 -113.395 ;
        RECT 77.355 -115.085 77.685 -114.755 ;
        RECT 77.355 -116.445 77.685 -116.115 ;
        RECT 77.355 -117.805 77.685 -117.475 ;
        RECT 77.355 -119.165 77.685 -118.835 ;
        RECT 77.355 -120.525 77.685 -120.195 ;
        RECT 77.355 -121.885 77.685 -121.555 ;
        RECT 77.355 -123.245 77.685 -122.915 ;
        RECT 77.355 -124.605 77.685 -124.275 ;
        RECT 77.355 -125.965 77.685 -125.635 ;
        RECT 77.355 -127.325 77.685 -126.995 ;
        RECT 77.355 -128.685 77.685 -128.355 ;
        RECT 77.355 -130.045 77.685 -129.715 ;
        RECT 77.355 -131.405 77.685 -131.075 ;
        RECT 77.355 -132.765 77.685 -132.435 ;
        RECT 77.355 -134.125 77.685 -133.795 ;
        RECT 77.355 -135.485 77.685 -135.155 ;
        RECT 77.355 -136.845 77.685 -136.515 ;
        RECT 77.355 -138.205 77.685 -137.875 ;
        RECT 77.355 -139.565 77.685 -139.235 ;
        RECT 77.355 -140.925 77.685 -140.595 ;
        RECT 77.355 -142.285 77.685 -141.955 ;
        RECT 77.355 -143.645 77.685 -143.315 ;
        RECT 77.355 -145.005 77.685 -144.675 ;
        RECT 77.355 -146.365 77.685 -146.035 ;
        RECT 77.355 -147.725 77.685 -147.395 ;
        RECT 77.355 -149.085 77.685 -148.755 ;
        RECT 77.355 -150.445 77.685 -150.115 ;
        RECT 77.355 -151.805 77.685 -151.475 ;
        RECT 77.355 -153.165 77.685 -152.835 ;
        RECT 77.355 -154.525 77.685 -154.195 ;
        RECT 77.355 -155.885 77.685 -155.555 ;
        RECT 77.355 -157.245 77.685 -156.915 ;
        RECT 77.355 -158.605 77.685 -158.275 ;
        RECT 77.355 -159.965 77.685 -159.635 ;
        RECT 77.355 -161.325 77.685 -160.995 ;
        RECT 77.355 -162.685 77.685 -162.355 ;
        RECT 77.355 -164.045 77.685 -163.715 ;
        RECT 77.355 -165.405 77.685 -165.075 ;
        RECT 77.355 -166.765 77.685 -166.435 ;
        RECT 77.355 -168.125 77.685 -167.795 ;
        RECT 77.355 -169.485 77.685 -169.155 ;
        RECT 77.355 -170.845 77.685 -170.515 ;
        RECT 77.355 -172.205 77.685 -171.875 ;
        RECT 77.355 -173.565 77.685 -173.235 ;
        RECT 77.355 -174.925 77.685 -174.595 ;
        RECT 77.355 -176.285 77.685 -175.955 ;
        RECT 77.355 -177.645 77.685 -177.315 ;
        RECT 77.355 -179.005 77.685 -178.675 ;
        RECT 77.355 -184.65 77.685 -183.52 ;
        RECT 77.36 -184.765 77.68 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 244.04 79.045 245.17 ;
        RECT 78.715 239.875 79.045 240.205 ;
        RECT 78.715 238.515 79.045 238.845 ;
        RECT 78.715 237.155 79.045 237.485 ;
        RECT 78.72 237.155 79.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.715 -98.765 79.045 -98.435 ;
        RECT 78.715 -100.125 79.045 -99.795 ;
        RECT 78.715 -101.485 79.045 -101.155 ;
        RECT 78.715 -102.845 79.045 -102.515 ;
        RECT 78.715 -104.205 79.045 -103.875 ;
        RECT 78.715 -105.565 79.045 -105.235 ;
        RECT 78.715 -106.925 79.045 -106.595 ;
        RECT 78.715 -108.285 79.045 -107.955 ;
        RECT 78.715 -109.645 79.045 -109.315 ;
        RECT 78.715 -111.005 79.045 -110.675 ;
        RECT 78.715 -112.365 79.045 -112.035 ;
        RECT 78.715 -113.725 79.045 -113.395 ;
        RECT 78.715 -115.085 79.045 -114.755 ;
        RECT 78.715 -116.445 79.045 -116.115 ;
        RECT 78.715 -117.805 79.045 -117.475 ;
        RECT 78.715 -119.165 79.045 -118.835 ;
        RECT 78.715 -120.525 79.045 -120.195 ;
        RECT 78.715 -121.885 79.045 -121.555 ;
        RECT 78.715 -123.245 79.045 -122.915 ;
        RECT 78.715 -124.605 79.045 -124.275 ;
        RECT 78.715 -125.965 79.045 -125.635 ;
        RECT 78.715 -127.325 79.045 -126.995 ;
        RECT 78.715 -128.685 79.045 -128.355 ;
        RECT 78.715 -130.045 79.045 -129.715 ;
        RECT 78.715 -131.405 79.045 -131.075 ;
        RECT 78.715 -132.765 79.045 -132.435 ;
        RECT 78.715 -134.125 79.045 -133.795 ;
        RECT 78.715 -135.485 79.045 -135.155 ;
        RECT 78.715 -136.845 79.045 -136.515 ;
        RECT 78.715 -138.205 79.045 -137.875 ;
        RECT 78.715 -139.565 79.045 -139.235 ;
        RECT 78.715 -140.925 79.045 -140.595 ;
        RECT 78.715 -142.285 79.045 -141.955 ;
        RECT 78.715 -143.645 79.045 -143.315 ;
        RECT 78.715 -145.005 79.045 -144.675 ;
        RECT 78.715 -146.365 79.045 -146.035 ;
        RECT 78.715 -147.725 79.045 -147.395 ;
        RECT 78.715 -149.085 79.045 -148.755 ;
        RECT 78.715 -150.445 79.045 -150.115 ;
        RECT 78.715 -151.805 79.045 -151.475 ;
        RECT 78.715 -153.165 79.045 -152.835 ;
        RECT 78.715 -154.525 79.045 -154.195 ;
        RECT 78.715 -155.885 79.045 -155.555 ;
        RECT 78.715 -157.245 79.045 -156.915 ;
        RECT 78.715 -158.605 79.045 -158.275 ;
        RECT 78.715 -159.965 79.045 -159.635 ;
        RECT 78.715 -161.325 79.045 -160.995 ;
        RECT 78.715 -162.685 79.045 -162.355 ;
        RECT 78.715 -164.045 79.045 -163.715 ;
        RECT 78.715 -165.405 79.045 -165.075 ;
        RECT 78.715 -166.765 79.045 -166.435 ;
        RECT 78.715 -168.125 79.045 -167.795 ;
        RECT 78.715 -169.485 79.045 -169.155 ;
        RECT 78.715 -170.845 79.045 -170.515 ;
        RECT 78.715 -172.205 79.045 -171.875 ;
        RECT 78.715 -173.565 79.045 -173.235 ;
        RECT 78.715 -174.925 79.045 -174.595 ;
        RECT 78.715 -176.285 79.045 -175.955 ;
        RECT 78.715 -177.645 79.045 -177.315 ;
        RECT 78.715 -179.005 79.045 -178.675 ;
        RECT 78.715 -184.65 79.045 -183.52 ;
        RECT 78.72 -184.765 79.04 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.96 -98.075 79.29 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.075 244.04 80.405 245.17 ;
        RECT 80.075 239.875 80.405 240.205 ;
        RECT 80.075 238.515 80.405 238.845 ;
        RECT 80.075 237.155 80.405 237.485 ;
        RECT 80.08 237.155 80.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 244.04 81.765 245.17 ;
        RECT 81.435 239.875 81.765 240.205 ;
        RECT 81.435 238.515 81.765 238.845 ;
        RECT 81.435 237.155 81.765 237.485 ;
        RECT 81.44 237.155 81.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 81.435 -0.845 81.765 -0.515 ;
        RECT 81.435 -2.205 81.765 -1.875 ;
        RECT 81.435 -3.565 81.765 -3.235 ;
        RECT 81.44 -3.565 81.76 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.795 244.04 83.125 245.17 ;
        RECT 82.795 239.875 83.125 240.205 ;
        RECT 82.795 238.515 83.125 238.845 ;
        RECT 82.795 237.155 83.125 237.485 ;
        RECT 82.8 237.155 83.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.795 -0.845 83.125 -0.515 ;
        RECT 82.795 -2.205 83.125 -1.875 ;
        RECT 82.795 -3.565 83.125 -3.235 ;
        RECT 82.8 -3.565 83.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.795 -96.045 83.125 -95.715 ;
        RECT 82.795 -97.405 83.125 -97.075 ;
        RECT 82.795 -98.765 83.125 -98.435 ;
        RECT 82.795 -100.125 83.125 -99.795 ;
        RECT 82.795 -101.485 83.125 -101.155 ;
        RECT 82.795 -102.845 83.125 -102.515 ;
        RECT 82.795 -104.205 83.125 -103.875 ;
        RECT 82.795 -105.565 83.125 -105.235 ;
        RECT 82.795 -106.925 83.125 -106.595 ;
        RECT 82.795 -108.285 83.125 -107.955 ;
        RECT 82.795 -109.645 83.125 -109.315 ;
        RECT 82.795 -111.005 83.125 -110.675 ;
        RECT 82.795 -112.365 83.125 -112.035 ;
        RECT 82.795 -113.725 83.125 -113.395 ;
        RECT 82.795 -115.085 83.125 -114.755 ;
        RECT 82.795 -116.445 83.125 -116.115 ;
        RECT 82.795 -117.805 83.125 -117.475 ;
        RECT 82.795 -119.165 83.125 -118.835 ;
        RECT 82.795 -120.525 83.125 -120.195 ;
        RECT 82.795 -121.885 83.125 -121.555 ;
        RECT 82.795 -123.245 83.125 -122.915 ;
        RECT 82.795 -124.605 83.125 -124.275 ;
        RECT 82.795 -125.965 83.125 -125.635 ;
        RECT 82.795 -127.325 83.125 -126.995 ;
        RECT 82.795 -128.685 83.125 -128.355 ;
        RECT 82.795 -130.045 83.125 -129.715 ;
        RECT 82.795 -131.405 83.125 -131.075 ;
        RECT 82.795 -132.765 83.125 -132.435 ;
        RECT 82.795 -134.125 83.125 -133.795 ;
        RECT 82.795 -135.485 83.125 -135.155 ;
        RECT 82.795 -136.845 83.125 -136.515 ;
        RECT 82.795 -138.205 83.125 -137.875 ;
        RECT 82.795 -139.565 83.125 -139.235 ;
        RECT 82.795 -140.925 83.125 -140.595 ;
        RECT 82.795 -142.285 83.125 -141.955 ;
        RECT 82.795 -143.645 83.125 -143.315 ;
        RECT 82.795 -145.005 83.125 -144.675 ;
        RECT 82.795 -146.365 83.125 -146.035 ;
        RECT 82.795 -147.725 83.125 -147.395 ;
        RECT 82.795 -149.085 83.125 -148.755 ;
        RECT 82.795 -150.445 83.125 -150.115 ;
        RECT 82.795 -151.805 83.125 -151.475 ;
        RECT 82.795 -153.165 83.125 -152.835 ;
        RECT 82.795 -154.525 83.125 -154.195 ;
        RECT 82.795 -155.885 83.125 -155.555 ;
        RECT 82.795 -157.245 83.125 -156.915 ;
        RECT 82.795 -158.605 83.125 -158.275 ;
        RECT 82.795 -159.965 83.125 -159.635 ;
        RECT 82.795 -161.325 83.125 -160.995 ;
        RECT 82.795 -162.685 83.125 -162.355 ;
        RECT 82.795 -164.045 83.125 -163.715 ;
        RECT 82.795 -165.405 83.125 -165.075 ;
        RECT 82.795 -166.765 83.125 -166.435 ;
        RECT 82.795 -168.125 83.125 -167.795 ;
        RECT 82.795 -169.485 83.125 -169.155 ;
        RECT 82.795 -170.845 83.125 -170.515 ;
        RECT 82.795 -172.205 83.125 -171.875 ;
        RECT 82.795 -173.565 83.125 -173.235 ;
        RECT 82.795 -174.925 83.125 -174.595 ;
        RECT 82.795 -176.285 83.125 -175.955 ;
        RECT 82.795 -177.645 83.125 -177.315 ;
        RECT 82.795 -179.005 83.125 -178.675 ;
        RECT 82.795 -184.65 83.125 -183.52 ;
        RECT 82.8 -184.765 83.12 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 244.04 84.485 245.17 ;
        RECT 84.155 239.875 84.485 240.205 ;
        RECT 84.155 238.515 84.485 238.845 ;
        RECT 84.155 237.155 84.485 237.485 ;
        RECT 84.16 237.155 84.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 -0.845 84.485 -0.515 ;
        RECT 84.155 -2.205 84.485 -1.875 ;
        RECT 84.155 -3.565 84.485 -3.235 ;
        RECT 84.16 -3.565 84.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.155 -96.045 84.485 -95.715 ;
        RECT 84.155 -97.405 84.485 -97.075 ;
        RECT 84.155 -98.765 84.485 -98.435 ;
        RECT 84.155 -100.125 84.485 -99.795 ;
        RECT 84.155 -101.485 84.485 -101.155 ;
        RECT 84.155 -102.845 84.485 -102.515 ;
        RECT 84.155 -104.205 84.485 -103.875 ;
        RECT 84.155 -105.565 84.485 -105.235 ;
        RECT 84.155 -106.925 84.485 -106.595 ;
        RECT 84.155 -108.285 84.485 -107.955 ;
        RECT 84.155 -109.645 84.485 -109.315 ;
        RECT 84.155 -111.005 84.485 -110.675 ;
        RECT 84.155 -112.365 84.485 -112.035 ;
        RECT 84.155 -113.725 84.485 -113.395 ;
        RECT 84.155 -115.085 84.485 -114.755 ;
        RECT 84.155 -116.445 84.485 -116.115 ;
        RECT 84.155 -117.805 84.485 -117.475 ;
        RECT 84.155 -119.165 84.485 -118.835 ;
        RECT 84.155 -120.525 84.485 -120.195 ;
        RECT 84.155 -121.885 84.485 -121.555 ;
        RECT 84.155 -123.245 84.485 -122.915 ;
        RECT 84.155 -124.605 84.485 -124.275 ;
        RECT 84.155 -125.965 84.485 -125.635 ;
        RECT 84.155 -127.325 84.485 -126.995 ;
        RECT 84.155 -128.685 84.485 -128.355 ;
        RECT 84.155 -130.045 84.485 -129.715 ;
        RECT 84.155 -131.405 84.485 -131.075 ;
        RECT 84.155 -132.765 84.485 -132.435 ;
        RECT 84.155 -134.125 84.485 -133.795 ;
        RECT 84.155 -135.485 84.485 -135.155 ;
        RECT 84.155 -136.845 84.485 -136.515 ;
        RECT 84.155 -138.205 84.485 -137.875 ;
        RECT 84.155 -139.565 84.485 -139.235 ;
        RECT 84.155 -140.925 84.485 -140.595 ;
        RECT 84.155 -142.285 84.485 -141.955 ;
        RECT 84.155 -143.645 84.485 -143.315 ;
        RECT 84.155 -145.005 84.485 -144.675 ;
        RECT 84.155 -146.365 84.485 -146.035 ;
        RECT 84.155 -147.725 84.485 -147.395 ;
        RECT 84.155 -149.085 84.485 -148.755 ;
        RECT 84.155 -150.445 84.485 -150.115 ;
        RECT 84.155 -151.805 84.485 -151.475 ;
        RECT 84.155 -153.165 84.485 -152.835 ;
        RECT 84.155 -154.525 84.485 -154.195 ;
        RECT 84.155 -155.885 84.485 -155.555 ;
        RECT 84.155 -157.245 84.485 -156.915 ;
        RECT 84.155 -158.605 84.485 -158.275 ;
        RECT 84.155 -159.965 84.485 -159.635 ;
        RECT 84.155 -161.325 84.485 -160.995 ;
        RECT 84.155 -162.685 84.485 -162.355 ;
        RECT 84.155 -164.045 84.485 -163.715 ;
        RECT 84.155 -165.405 84.485 -165.075 ;
        RECT 84.155 -166.765 84.485 -166.435 ;
        RECT 84.155 -168.125 84.485 -167.795 ;
        RECT 84.155 -169.485 84.485 -169.155 ;
        RECT 84.155 -170.845 84.485 -170.515 ;
        RECT 84.155 -172.205 84.485 -171.875 ;
        RECT 84.155 -173.565 84.485 -173.235 ;
        RECT 84.155 -174.925 84.485 -174.595 ;
        RECT 84.155 -176.285 84.485 -175.955 ;
        RECT 84.155 -177.645 84.485 -177.315 ;
        RECT 84.155 -179.005 84.485 -178.675 ;
        RECT 84.155 -184.65 84.485 -183.52 ;
        RECT 84.16 -184.765 84.48 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 244.04 85.845 245.17 ;
        RECT 85.515 239.875 85.845 240.205 ;
        RECT 85.515 238.515 85.845 238.845 ;
        RECT 85.515 237.155 85.845 237.485 ;
        RECT 85.52 237.155 85.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 -0.845 85.845 -0.515 ;
        RECT 85.515 -2.205 85.845 -1.875 ;
        RECT 85.515 -3.565 85.845 -3.235 ;
        RECT 85.52 -3.565 85.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 85.515 -179.005 85.845 -178.675 ;
        RECT 85.515 -184.65 85.845 -183.52 ;
        RECT 85.52 -184.765 85.84 -95.04 ;
        RECT 85.515 -96.045 85.845 -95.715 ;
        RECT 85.515 -97.405 85.845 -97.075 ;
        RECT 85.515 -98.765 85.845 -98.435 ;
        RECT 85.515 -100.125 85.845 -99.795 ;
        RECT 85.515 -101.485 85.845 -101.155 ;
        RECT 85.515 -102.845 85.845 -102.515 ;
        RECT 85.515 -104.205 85.845 -103.875 ;
        RECT 85.515 -105.565 85.845 -105.235 ;
        RECT 85.515 -106.925 85.845 -106.595 ;
        RECT 85.515 -108.285 85.845 -107.955 ;
        RECT 85.515 -109.645 85.845 -109.315 ;
        RECT 85.515 -111.005 85.845 -110.675 ;
        RECT 85.515 -112.365 85.845 -112.035 ;
        RECT 85.515 -113.725 85.845 -113.395 ;
        RECT 85.515 -115.085 85.845 -114.755 ;
        RECT 85.515 -116.445 85.845 -116.115 ;
        RECT 85.515 -117.805 85.845 -117.475 ;
        RECT 85.515 -119.165 85.845 -118.835 ;
        RECT 85.515 -120.525 85.845 -120.195 ;
        RECT 85.515 -121.885 85.845 -121.555 ;
        RECT 85.515 -123.245 85.845 -122.915 ;
        RECT 85.515 -124.605 85.845 -124.275 ;
        RECT 85.515 -125.965 85.845 -125.635 ;
        RECT 85.515 -127.325 85.845 -126.995 ;
        RECT 85.515 -128.685 85.845 -128.355 ;
        RECT 85.515 -130.045 85.845 -129.715 ;
        RECT 85.515 -131.405 85.845 -131.075 ;
        RECT 85.515 -132.765 85.845 -132.435 ;
        RECT 85.515 -134.125 85.845 -133.795 ;
        RECT 85.515 -135.485 85.845 -135.155 ;
        RECT 85.515 -136.845 85.845 -136.515 ;
        RECT 85.515 -138.205 85.845 -137.875 ;
        RECT 85.515 -139.565 85.845 -139.235 ;
        RECT 85.515 -140.925 85.845 -140.595 ;
        RECT 85.515 -142.285 85.845 -141.955 ;
        RECT 85.515 -143.645 85.845 -143.315 ;
        RECT 85.515 -145.005 85.845 -144.675 ;
        RECT 85.515 -146.365 85.845 -146.035 ;
        RECT 85.515 -147.725 85.845 -147.395 ;
        RECT 85.515 -149.085 85.845 -148.755 ;
        RECT 85.515 -150.445 85.845 -150.115 ;
        RECT 85.515 -151.805 85.845 -151.475 ;
        RECT 85.515 -153.165 85.845 -152.835 ;
        RECT 85.515 -154.525 85.845 -154.195 ;
        RECT 85.515 -155.885 85.845 -155.555 ;
        RECT 85.515 -157.245 85.845 -156.915 ;
        RECT 85.515 -158.605 85.845 -158.275 ;
        RECT 85.515 -159.965 85.845 -159.635 ;
        RECT 85.515 -161.325 85.845 -160.995 ;
        RECT 85.515 -162.685 85.845 -162.355 ;
        RECT 85.515 -164.045 85.845 -163.715 ;
        RECT 85.515 -165.405 85.845 -165.075 ;
        RECT 85.515 -166.765 85.845 -166.435 ;
        RECT 85.515 -168.125 85.845 -167.795 ;
        RECT 85.515 -169.485 85.845 -169.155 ;
        RECT 85.515 -170.845 85.845 -170.515 ;
        RECT 85.515 -172.205 85.845 -171.875 ;
        RECT 85.515 -173.565 85.845 -173.235 ;
        RECT 85.515 -174.925 85.845 -174.595 ;
        RECT 85.515 -176.285 85.845 -175.955 ;
        RECT 85.515 -177.645 85.845 -177.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.36 -98.075 35.69 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.555 244.04 36.885 245.17 ;
        RECT 36.555 239.875 36.885 240.205 ;
        RECT 36.555 238.515 36.885 238.845 ;
        RECT 36.555 237.155 36.885 237.485 ;
        RECT 36.56 237.155 36.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 244.04 38.245 245.17 ;
        RECT 37.915 239.875 38.245 240.205 ;
        RECT 37.915 238.515 38.245 238.845 ;
        RECT 37.915 237.155 38.245 237.485 ;
        RECT 37.92 237.155 38.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.915 -0.845 38.245 -0.515 ;
        RECT 37.915 -2.205 38.245 -1.875 ;
        RECT 37.915 -3.565 38.245 -3.235 ;
        RECT 37.92 -3.565 38.24 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 244.04 39.605 245.17 ;
        RECT 39.275 239.875 39.605 240.205 ;
        RECT 39.275 238.515 39.605 238.845 ;
        RECT 39.275 237.155 39.605 237.485 ;
        RECT 39.28 237.155 39.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 -0.845 39.605 -0.515 ;
        RECT 39.275 -2.205 39.605 -1.875 ;
        RECT 39.275 -3.565 39.605 -3.235 ;
        RECT 39.28 -3.565 39.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.275 -96.045 39.605 -95.715 ;
        RECT 39.275 -97.405 39.605 -97.075 ;
        RECT 39.275 -98.765 39.605 -98.435 ;
        RECT 39.275 -100.125 39.605 -99.795 ;
        RECT 39.275 -101.485 39.605 -101.155 ;
        RECT 39.275 -102.845 39.605 -102.515 ;
        RECT 39.275 -104.205 39.605 -103.875 ;
        RECT 39.275 -105.565 39.605 -105.235 ;
        RECT 39.275 -106.925 39.605 -106.595 ;
        RECT 39.275 -108.285 39.605 -107.955 ;
        RECT 39.275 -109.645 39.605 -109.315 ;
        RECT 39.275 -111.005 39.605 -110.675 ;
        RECT 39.275 -112.365 39.605 -112.035 ;
        RECT 39.275 -113.725 39.605 -113.395 ;
        RECT 39.275 -115.085 39.605 -114.755 ;
        RECT 39.275 -116.445 39.605 -116.115 ;
        RECT 39.275 -117.805 39.605 -117.475 ;
        RECT 39.275 -119.165 39.605 -118.835 ;
        RECT 39.275 -120.525 39.605 -120.195 ;
        RECT 39.275 -121.885 39.605 -121.555 ;
        RECT 39.275 -123.245 39.605 -122.915 ;
        RECT 39.275 -124.605 39.605 -124.275 ;
        RECT 39.275 -125.965 39.605 -125.635 ;
        RECT 39.275 -127.325 39.605 -126.995 ;
        RECT 39.275 -128.685 39.605 -128.355 ;
        RECT 39.275 -130.045 39.605 -129.715 ;
        RECT 39.275 -131.405 39.605 -131.075 ;
        RECT 39.275 -132.765 39.605 -132.435 ;
        RECT 39.275 -134.125 39.605 -133.795 ;
        RECT 39.275 -135.485 39.605 -135.155 ;
        RECT 39.275 -136.845 39.605 -136.515 ;
        RECT 39.275 -138.205 39.605 -137.875 ;
        RECT 39.275 -139.565 39.605 -139.235 ;
        RECT 39.275 -140.925 39.605 -140.595 ;
        RECT 39.275 -142.285 39.605 -141.955 ;
        RECT 39.275 -143.645 39.605 -143.315 ;
        RECT 39.275 -145.005 39.605 -144.675 ;
        RECT 39.275 -146.365 39.605 -146.035 ;
        RECT 39.275 -147.725 39.605 -147.395 ;
        RECT 39.275 -149.085 39.605 -148.755 ;
        RECT 39.275 -150.445 39.605 -150.115 ;
        RECT 39.275 -151.805 39.605 -151.475 ;
        RECT 39.275 -153.165 39.605 -152.835 ;
        RECT 39.275 -154.525 39.605 -154.195 ;
        RECT 39.275 -155.885 39.605 -155.555 ;
        RECT 39.275 -157.245 39.605 -156.915 ;
        RECT 39.275 -158.605 39.605 -158.275 ;
        RECT 39.275 -159.965 39.605 -159.635 ;
        RECT 39.275 -161.325 39.605 -160.995 ;
        RECT 39.275 -162.685 39.605 -162.355 ;
        RECT 39.275 -164.045 39.605 -163.715 ;
        RECT 39.275 -165.405 39.605 -165.075 ;
        RECT 39.275 -166.765 39.605 -166.435 ;
        RECT 39.275 -168.125 39.605 -167.795 ;
        RECT 39.275 -169.485 39.605 -169.155 ;
        RECT 39.275 -170.845 39.605 -170.515 ;
        RECT 39.275 -172.205 39.605 -171.875 ;
        RECT 39.275 -173.565 39.605 -173.235 ;
        RECT 39.275 -174.925 39.605 -174.595 ;
        RECT 39.275 -176.285 39.605 -175.955 ;
        RECT 39.275 -177.645 39.605 -177.315 ;
        RECT 39.275 -179.005 39.605 -178.675 ;
        RECT 39.275 -184.65 39.605 -183.52 ;
        RECT 39.28 -184.765 39.6 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 244.04 40.965 245.17 ;
        RECT 40.635 239.875 40.965 240.205 ;
        RECT 40.635 238.515 40.965 238.845 ;
        RECT 40.635 237.155 40.965 237.485 ;
        RECT 40.64 237.155 40.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 -0.845 40.965 -0.515 ;
        RECT 40.635 -2.205 40.965 -1.875 ;
        RECT 40.635 -3.565 40.965 -3.235 ;
        RECT 40.64 -3.565 40.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 40.635 -96.045 40.965 -95.715 ;
        RECT 40.635 -97.405 40.965 -97.075 ;
        RECT 40.635 -98.765 40.965 -98.435 ;
        RECT 40.635 -100.125 40.965 -99.795 ;
        RECT 40.635 -101.485 40.965 -101.155 ;
        RECT 40.635 -102.845 40.965 -102.515 ;
        RECT 40.635 -104.205 40.965 -103.875 ;
        RECT 40.635 -105.565 40.965 -105.235 ;
        RECT 40.635 -106.925 40.965 -106.595 ;
        RECT 40.635 -108.285 40.965 -107.955 ;
        RECT 40.635 -109.645 40.965 -109.315 ;
        RECT 40.635 -111.005 40.965 -110.675 ;
        RECT 40.635 -112.365 40.965 -112.035 ;
        RECT 40.635 -113.725 40.965 -113.395 ;
        RECT 40.635 -115.085 40.965 -114.755 ;
        RECT 40.635 -116.445 40.965 -116.115 ;
        RECT 40.635 -117.805 40.965 -117.475 ;
        RECT 40.635 -119.165 40.965 -118.835 ;
        RECT 40.635 -120.525 40.965 -120.195 ;
        RECT 40.635 -121.885 40.965 -121.555 ;
        RECT 40.635 -123.245 40.965 -122.915 ;
        RECT 40.635 -124.605 40.965 -124.275 ;
        RECT 40.635 -125.965 40.965 -125.635 ;
        RECT 40.635 -127.325 40.965 -126.995 ;
        RECT 40.635 -128.685 40.965 -128.355 ;
        RECT 40.635 -130.045 40.965 -129.715 ;
        RECT 40.635 -131.405 40.965 -131.075 ;
        RECT 40.635 -132.765 40.965 -132.435 ;
        RECT 40.635 -134.125 40.965 -133.795 ;
        RECT 40.635 -135.485 40.965 -135.155 ;
        RECT 40.635 -136.845 40.965 -136.515 ;
        RECT 40.635 -138.205 40.965 -137.875 ;
        RECT 40.635 -139.565 40.965 -139.235 ;
        RECT 40.635 -140.925 40.965 -140.595 ;
        RECT 40.635 -142.285 40.965 -141.955 ;
        RECT 40.635 -143.645 40.965 -143.315 ;
        RECT 40.635 -145.005 40.965 -144.675 ;
        RECT 40.635 -146.365 40.965 -146.035 ;
        RECT 40.635 -147.725 40.965 -147.395 ;
        RECT 40.635 -149.085 40.965 -148.755 ;
        RECT 40.635 -150.445 40.965 -150.115 ;
        RECT 40.635 -151.805 40.965 -151.475 ;
        RECT 40.635 -153.165 40.965 -152.835 ;
        RECT 40.635 -154.525 40.965 -154.195 ;
        RECT 40.635 -155.885 40.965 -155.555 ;
        RECT 40.635 -157.245 40.965 -156.915 ;
        RECT 40.635 -158.605 40.965 -158.275 ;
        RECT 40.635 -159.965 40.965 -159.635 ;
        RECT 40.635 -161.325 40.965 -160.995 ;
        RECT 40.635 -162.685 40.965 -162.355 ;
        RECT 40.635 -164.045 40.965 -163.715 ;
        RECT 40.635 -165.405 40.965 -165.075 ;
        RECT 40.635 -166.765 40.965 -166.435 ;
        RECT 40.635 -168.125 40.965 -167.795 ;
        RECT 40.635 -169.485 40.965 -169.155 ;
        RECT 40.635 -170.845 40.965 -170.515 ;
        RECT 40.635 -172.205 40.965 -171.875 ;
        RECT 40.635 -173.565 40.965 -173.235 ;
        RECT 40.635 -174.925 40.965 -174.595 ;
        RECT 40.635 -176.285 40.965 -175.955 ;
        RECT 40.635 -177.645 40.965 -177.315 ;
        RECT 40.635 -179.005 40.965 -178.675 ;
        RECT 40.635 -184.65 40.965 -183.52 ;
        RECT 40.64 -184.765 40.96 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 244.04 42.325 245.17 ;
        RECT 41.995 239.875 42.325 240.205 ;
        RECT 41.995 238.515 42.325 238.845 ;
        RECT 41.995 237.155 42.325 237.485 ;
        RECT 42 237.155 42.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 -0.845 42.325 -0.515 ;
        RECT 41.995 -2.205 42.325 -1.875 ;
        RECT 41.995 -3.565 42.325 -3.235 ;
        RECT 42 -3.565 42.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.995 -96.045 42.325 -95.715 ;
        RECT 41.995 -97.405 42.325 -97.075 ;
        RECT 41.995 -98.765 42.325 -98.435 ;
        RECT 41.995 -100.125 42.325 -99.795 ;
        RECT 41.995 -101.485 42.325 -101.155 ;
        RECT 41.995 -102.845 42.325 -102.515 ;
        RECT 41.995 -104.205 42.325 -103.875 ;
        RECT 41.995 -105.565 42.325 -105.235 ;
        RECT 41.995 -106.925 42.325 -106.595 ;
        RECT 41.995 -108.285 42.325 -107.955 ;
        RECT 41.995 -109.645 42.325 -109.315 ;
        RECT 41.995 -111.005 42.325 -110.675 ;
        RECT 41.995 -112.365 42.325 -112.035 ;
        RECT 41.995 -113.725 42.325 -113.395 ;
        RECT 41.995 -115.085 42.325 -114.755 ;
        RECT 41.995 -116.445 42.325 -116.115 ;
        RECT 41.995 -117.805 42.325 -117.475 ;
        RECT 41.995 -119.165 42.325 -118.835 ;
        RECT 41.995 -120.525 42.325 -120.195 ;
        RECT 41.995 -121.885 42.325 -121.555 ;
        RECT 41.995 -123.245 42.325 -122.915 ;
        RECT 41.995 -124.605 42.325 -124.275 ;
        RECT 41.995 -125.965 42.325 -125.635 ;
        RECT 41.995 -127.325 42.325 -126.995 ;
        RECT 41.995 -128.685 42.325 -128.355 ;
        RECT 41.995 -130.045 42.325 -129.715 ;
        RECT 41.995 -131.405 42.325 -131.075 ;
        RECT 41.995 -132.765 42.325 -132.435 ;
        RECT 41.995 -134.125 42.325 -133.795 ;
        RECT 41.995 -135.485 42.325 -135.155 ;
        RECT 41.995 -136.845 42.325 -136.515 ;
        RECT 41.995 -138.205 42.325 -137.875 ;
        RECT 41.995 -139.565 42.325 -139.235 ;
        RECT 41.995 -140.925 42.325 -140.595 ;
        RECT 41.995 -142.285 42.325 -141.955 ;
        RECT 41.995 -143.645 42.325 -143.315 ;
        RECT 41.995 -145.005 42.325 -144.675 ;
        RECT 41.995 -146.365 42.325 -146.035 ;
        RECT 41.995 -147.725 42.325 -147.395 ;
        RECT 41.995 -149.085 42.325 -148.755 ;
        RECT 41.995 -150.445 42.325 -150.115 ;
        RECT 41.995 -151.805 42.325 -151.475 ;
        RECT 41.995 -153.165 42.325 -152.835 ;
        RECT 41.995 -154.525 42.325 -154.195 ;
        RECT 41.995 -155.885 42.325 -155.555 ;
        RECT 41.995 -157.245 42.325 -156.915 ;
        RECT 41.995 -158.605 42.325 -158.275 ;
        RECT 41.995 -159.965 42.325 -159.635 ;
        RECT 41.995 -161.325 42.325 -160.995 ;
        RECT 41.995 -162.685 42.325 -162.355 ;
        RECT 41.995 -164.045 42.325 -163.715 ;
        RECT 41.995 -165.405 42.325 -165.075 ;
        RECT 41.995 -166.765 42.325 -166.435 ;
        RECT 41.995 -168.125 42.325 -167.795 ;
        RECT 41.995 -169.485 42.325 -169.155 ;
        RECT 41.995 -170.845 42.325 -170.515 ;
        RECT 41.995 -172.205 42.325 -171.875 ;
        RECT 41.995 -173.565 42.325 -173.235 ;
        RECT 41.995 -174.925 42.325 -174.595 ;
        RECT 41.995 -176.285 42.325 -175.955 ;
        RECT 41.995 -177.645 42.325 -177.315 ;
        RECT 41.995 -179.005 42.325 -178.675 ;
        RECT 41.995 -184.65 42.325 -183.52 ;
        RECT 42 -184.765 42.32 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 244.04 43.685 245.17 ;
        RECT 43.355 239.875 43.685 240.205 ;
        RECT 43.355 238.515 43.685 238.845 ;
        RECT 43.355 237.155 43.685 237.485 ;
        RECT 43.36 237.155 43.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 -0.845 43.685 -0.515 ;
        RECT 43.355 -2.205 43.685 -1.875 ;
        RECT 43.355 -3.565 43.685 -3.235 ;
        RECT 43.36 -3.565 43.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 43.355 -96.045 43.685 -95.715 ;
        RECT 43.355 -97.405 43.685 -97.075 ;
        RECT 43.355 -98.765 43.685 -98.435 ;
        RECT 43.355 -100.125 43.685 -99.795 ;
        RECT 43.355 -101.485 43.685 -101.155 ;
        RECT 43.355 -102.845 43.685 -102.515 ;
        RECT 43.355 -104.205 43.685 -103.875 ;
        RECT 43.355 -105.565 43.685 -105.235 ;
        RECT 43.355 -106.925 43.685 -106.595 ;
        RECT 43.355 -108.285 43.685 -107.955 ;
        RECT 43.355 -109.645 43.685 -109.315 ;
        RECT 43.355 -111.005 43.685 -110.675 ;
        RECT 43.355 -112.365 43.685 -112.035 ;
        RECT 43.355 -113.725 43.685 -113.395 ;
        RECT 43.355 -115.085 43.685 -114.755 ;
        RECT 43.355 -116.445 43.685 -116.115 ;
        RECT 43.355 -117.805 43.685 -117.475 ;
        RECT 43.355 -119.165 43.685 -118.835 ;
        RECT 43.355 -120.525 43.685 -120.195 ;
        RECT 43.355 -121.885 43.685 -121.555 ;
        RECT 43.355 -123.245 43.685 -122.915 ;
        RECT 43.355 -124.605 43.685 -124.275 ;
        RECT 43.355 -125.965 43.685 -125.635 ;
        RECT 43.355 -127.325 43.685 -126.995 ;
        RECT 43.355 -128.685 43.685 -128.355 ;
        RECT 43.355 -130.045 43.685 -129.715 ;
        RECT 43.355 -131.405 43.685 -131.075 ;
        RECT 43.355 -132.765 43.685 -132.435 ;
        RECT 43.355 -134.125 43.685 -133.795 ;
        RECT 43.355 -135.485 43.685 -135.155 ;
        RECT 43.355 -136.845 43.685 -136.515 ;
        RECT 43.355 -138.205 43.685 -137.875 ;
        RECT 43.355 -139.565 43.685 -139.235 ;
        RECT 43.355 -140.925 43.685 -140.595 ;
        RECT 43.355 -142.285 43.685 -141.955 ;
        RECT 43.355 -143.645 43.685 -143.315 ;
        RECT 43.355 -145.005 43.685 -144.675 ;
        RECT 43.355 -146.365 43.685 -146.035 ;
        RECT 43.355 -147.725 43.685 -147.395 ;
        RECT 43.355 -149.085 43.685 -148.755 ;
        RECT 43.355 -150.445 43.685 -150.115 ;
        RECT 43.355 -151.805 43.685 -151.475 ;
        RECT 43.355 -153.165 43.685 -152.835 ;
        RECT 43.355 -154.525 43.685 -154.195 ;
        RECT 43.355 -155.885 43.685 -155.555 ;
        RECT 43.355 -157.245 43.685 -156.915 ;
        RECT 43.355 -158.605 43.685 -158.275 ;
        RECT 43.355 -159.965 43.685 -159.635 ;
        RECT 43.355 -161.325 43.685 -160.995 ;
        RECT 43.355 -162.685 43.685 -162.355 ;
        RECT 43.355 -164.045 43.685 -163.715 ;
        RECT 43.355 -165.405 43.685 -165.075 ;
        RECT 43.355 -166.765 43.685 -166.435 ;
        RECT 43.355 -168.125 43.685 -167.795 ;
        RECT 43.355 -169.485 43.685 -169.155 ;
        RECT 43.355 -170.845 43.685 -170.515 ;
        RECT 43.355 -172.205 43.685 -171.875 ;
        RECT 43.355 -173.565 43.685 -173.235 ;
        RECT 43.355 -174.925 43.685 -174.595 ;
        RECT 43.355 -176.285 43.685 -175.955 ;
        RECT 43.355 -177.645 43.685 -177.315 ;
        RECT 43.355 -179.005 43.685 -178.675 ;
        RECT 43.355 -184.65 43.685 -183.52 ;
        RECT 43.36 -184.765 43.68 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 244.04 45.045 245.17 ;
        RECT 44.715 239.875 45.045 240.205 ;
        RECT 44.715 238.515 45.045 238.845 ;
        RECT 44.715 237.155 45.045 237.485 ;
        RECT 44.72 237.155 45.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 -0.845 45.045 -0.515 ;
        RECT 44.715 -2.205 45.045 -1.875 ;
        RECT 44.715 -3.565 45.045 -3.235 ;
        RECT 44.72 -3.565 45.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.715 -96.045 45.045 -95.715 ;
        RECT 44.715 -97.405 45.045 -97.075 ;
        RECT 44.715 -98.765 45.045 -98.435 ;
        RECT 44.715 -100.125 45.045 -99.795 ;
        RECT 44.715 -101.485 45.045 -101.155 ;
        RECT 44.715 -102.845 45.045 -102.515 ;
        RECT 44.715 -104.205 45.045 -103.875 ;
        RECT 44.715 -105.565 45.045 -105.235 ;
        RECT 44.715 -106.925 45.045 -106.595 ;
        RECT 44.715 -108.285 45.045 -107.955 ;
        RECT 44.715 -109.645 45.045 -109.315 ;
        RECT 44.715 -111.005 45.045 -110.675 ;
        RECT 44.715 -112.365 45.045 -112.035 ;
        RECT 44.715 -113.725 45.045 -113.395 ;
        RECT 44.715 -115.085 45.045 -114.755 ;
        RECT 44.715 -116.445 45.045 -116.115 ;
        RECT 44.715 -117.805 45.045 -117.475 ;
        RECT 44.715 -119.165 45.045 -118.835 ;
        RECT 44.715 -120.525 45.045 -120.195 ;
        RECT 44.715 -121.885 45.045 -121.555 ;
        RECT 44.715 -123.245 45.045 -122.915 ;
        RECT 44.715 -124.605 45.045 -124.275 ;
        RECT 44.715 -125.965 45.045 -125.635 ;
        RECT 44.715 -127.325 45.045 -126.995 ;
        RECT 44.715 -128.685 45.045 -128.355 ;
        RECT 44.715 -130.045 45.045 -129.715 ;
        RECT 44.715 -131.405 45.045 -131.075 ;
        RECT 44.715 -132.765 45.045 -132.435 ;
        RECT 44.715 -134.125 45.045 -133.795 ;
        RECT 44.715 -135.485 45.045 -135.155 ;
        RECT 44.715 -136.845 45.045 -136.515 ;
        RECT 44.715 -138.205 45.045 -137.875 ;
        RECT 44.715 -139.565 45.045 -139.235 ;
        RECT 44.715 -140.925 45.045 -140.595 ;
        RECT 44.715 -142.285 45.045 -141.955 ;
        RECT 44.715 -143.645 45.045 -143.315 ;
        RECT 44.715 -145.005 45.045 -144.675 ;
        RECT 44.715 -146.365 45.045 -146.035 ;
        RECT 44.715 -147.725 45.045 -147.395 ;
        RECT 44.715 -149.085 45.045 -148.755 ;
        RECT 44.715 -150.445 45.045 -150.115 ;
        RECT 44.715 -151.805 45.045 -151.475 ;
        RECT 44.715 -153.165 45.045 -152.835 ;
        RECT 44.715 -154.525 45.045 -154.195 ;
        RECT 44.715 -155.885 45.045 -155.555 ;
        RECT 44.715 -157.245 45.045 -156.915 ;
        RECT 44.715 -158.605 45.045 -158.275 ;
        RECT 44.715 -159.965 45.045 -159.635 ;
        RECT 44.715 -161.325 45.045 -160.995 ;
        RECT 44.715 -162.685 45.045 -162.355 ;
        RECT 44.715 -164.045 45.045 -163.715 ;
        RECT 44.715 -165.405 45.045 -165.075 ;
        RECT 44.715 -166.765 45.045 -166.435 ;
        RECT 44.715 -168.125 45.045 -167.795 ;
        RECT 44.715 -169.485 45.045 -169.155 ;
        RECT 44.715 -170.845 45.045 -170.515 ;
        RECT 44.715 -172.205 45.045 -171.875 ;
        RECT 44.715 -173.565 45.045 -173.235 ;
        RECT 44.715 -174.925 45.045 -174.595 ;
        RECT 44.715 -176.285 45.045 -175.955 ;
        RECT 44.715 -177.645 45.045 -177.315 ;
        RECT 44.715 -179.005 45.045 -178.675 ;
        RECT 44.715 -184.65 45.045 -183.52 ;
        RECT 44.72 -184.765 45.04 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.075 244.04 46.405 245.17 ;
        RECT 46.075 239.875 46.405 240.205 ;
        RECT 46.075 238.515 46.405 238.845 ;
        RECT 46.075 237.155 46.405 237.485 ;
        RECT 46.08 237.155 46.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.075 -98.765 46.405 -98.435 ;
        RECT 46.075 -100.125 46.405 -99.795 ;
        RECT 46.075 -101.485 46.405 -101.155 ;
        RECT 46.075 -102.845 46.405 -102.515 ;
        RECT 46.075 -104.205 46.405 -103.875 ;
        RECT 46.075 -105.565 46.405 -105.235 ;
        RECT 46.075 -106.925 46.405 -106.595 ;
        RECT 46.075 -108.285 46.405 -107.955 ;
        RECT 46.075 -109.645 46.405 -109.315 ;
        RECT 46.075 -111.005 46.405 -110.675 ;
        RECT 46.075 -112.365 46.405 -112.035 ;
        RECT 46.075 -113.725 46.405 -113.395 ;
        RECT 46.075 -115.085 46.405 -114.755 ;
        RECT 46.075 -116.445 46.405 -116.115 ;
        RECT 46.075 -117.805 46.405 -117.475 ;
        RECT 46.075 -119.165 46.405 -118.835 ;
        RECT 46.075 -120.525 46.405 -120.195 ;
        RECT 46.075 -121.885 46.405 -121.555 ;
        RECT 46.075 -123.245 46.405 -122.915 ;
        RECT 46.075 -124.605 46.405 -124.275 ;
        RECT 46.075 -125.965 46.405 -125.635 ;
        RECT 46.075 -127.325 46.405 -126.995 ;
        RECT 46.075 -128.685 46.405 -128.355 ;
        RECT 46.075 -130.045 46.405 -129.715 ;
        RECT 46.075 -131.405 46.405 -131.075 ;
        RECT 46.075 -132.765 46.405 -132.435 ;
        RECT 46.075 -134.125 46.405 -133.795 ;
        RECT 46.075 -135.485 46.405 -135.155 ;
        RECT 46.075 -136.845 46.405 -136.515 ;
        RECT 46.075 -138.205 46.405 -137.875 ;
        RECT 46.075 -139.565 46.405 -139.235 ;
        RECT 46.075 -140.925 46.405 -140.595 ;
        RECT 46.075 -142.285 46.405 -141.955 ;
        RECT 46.075 -143.645 46.405 -143.315 ;
        RECT 46.075 -145.005 46.405 -144.675 ;
        RECT 46.075 -146.365 46.405 -146.035 ;
        RECT 46.075 -147.725 46.405 -147.395 ;
        RECT 46.075 -149.085 46.405 -148.755 ;
        RECT 46.075 -150.445 46.405 -150.115 ;
        RECT 46.075 -151.805 46.405 -151.475 ;
        RECT 46.075 -153.165 46.405 -152.835 ;
        RECT 46.075 -154.525 46.405 -154.195 ;
        RECT 46.075 -155.885 46.405 -155.555 ;
        RECT 46.075 -157.245 46.405 -156.915 ;
        RECT 46.075 -158.605 46.405 -158.275 ;
        RECT 46.075 -159.965 46.405 -159.635 ;
        RECT 46.075 -161.325 46.405 -160.995 ;
        RECT 46.075 -162.685 46.405 -162.355 ;
        RECT 46.075 -164.045 46.405 -163.715 ;
        RECT 46.075 -165.405 46.405 -165.075 ;
        RECT 46.075 -166.765 46.405 -166.435 ;
        RECT 46.075 -168.125 46.405 -167.795 ;
        RECT 46.075 -169.485 46.405 -169.155 ;
        RECT 46.075 -170.845 46.405 -170.515 ;
        RECT 46.075 -172.205 46.405 -171.875 ;
        RECT 46.075 -173.565 46.405 -173.235 ;
        RECT 46.075 -174.925 46.405 -174.595 ;
        RECT 46.075 -176.285 46.405 -175.955 ;
        RECT 46.075 -177.645 46.405 -177.315 ;
        RECT 46.075 -179.005 46.405 -178.675 ;
        RECT 46.075 -184.65 46.405 -183.52 ;
        RECT 46.08 -184.765 46.4 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.26 -98.075 46.59 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 47.435 244.04 47.765 245.17 ;
        RECT 47.435 239.875 47.765 240.205 ;
        RECT 47.435 238.515 47.765 238.845 ;
        RECT 47.435 237.155 47.765 237.485 ;
        RECT 47.44 237.155 47.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 244.04 49.125 245.17 ;
        RECT 48.795 239.875 49.125 240.205 ;
        RECT 48.795 238.515 49.125 238.845 ;
        RECT 48.795 237.155 49.125 237.485 ;
        RECT 48.8 237.155 49.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.795 -0.845 49.125 -0.515 ;
        RECT 48.795 -2.205 49.125 -1.875 ;
        RECT 48.795 -3.565 49.125 -3.235 ;
        RECT 48.8 -3.565 49.12 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 244.04 50.485 245.17 ;
        RECT 50.155 239.875 50.485 240.205 ;
        RECT 50.155 238.515 50.485 238.845 ;
        RECT 50.155 237.155 50.485 237.485 ;
        RECT 50.16 237.155 50.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 -0.845 50.485 -0.515 ;
        RECT 50.155 -2.205 50.485 -1.875 ;
        RECT 50.155 -3.565 50.485 -3.235 ;
        RECT 50.16 -3.565 50.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.155 -96.045 50.485 -95.715 ;
        RECT 50.155 -97.405 50.485 -97.075 ;
        RECT 50.155 -98.765 50.485 -98.435 ;
        RECT 50.155 -100.125 50.485 -99.795 ;
        RECT 50.155 -101.485 50.485 -101.155 ;
        RECT 50.155 -102.845 50.485 -102.515 ;
        RECT 50.155 -104.205 50.485 -103.875 ;
        RECT 50.155 -105.565 50.485 -105.235 ;
        RECT 50.155 -106.925 50.485 -106.595 ;
        RECT 50.155 -108.285 50.485 -107.955 ;
        RECT 50.155 -109.645 50.485 -109.315 ;
        RECT 50.155 -111.005 50.485 -110.675 ;
        RECT 50.155 -112.365 50.485 -112.035 ;
        RECT 50.155 -113.725 50.485 -113.395 ;
        RECT 50.155 -115.085 50.485 -114.755 ;
        RECT 50.155 -116.445 50.485 -116.115 ;
        RECT 50.155 -117.805 50.485 -117.475 ;
        RECT 50.155 -119.165 50.485 -118.835 ;
        RECT 50.155 -120.525 50.485 -120.195 ;
        RECT 50.155 -121.885 50.485 -121.555 ;
        RECT 50.155 -123.245 50.485 -122.915 ;
        RECT 50.155 -124.605 50.485 -124.275 ;
        RECT 50.155 -125.965 50.485 -125.635 ;
        RECT 50.155 -127.325 50.485 -126.995 ;
        RECT 50.155 -128.685 50.485 -128.355 ;
        RECT 50.155 -130.045 50.485 -129.715 ;
        RECT 50.155 -131.405 50.485 -131.075 ;
        RECT 50.155 -132.765 50.485 -132.435 ;
        RECT 50.155 -134.125 50.485 -133.795 ;
        RECT 50.155 -135.485 50.485 -135.155 ;
        RECT 50.155 -136.845 50.485 -136.515 ;
        RECT 50.155 -138.205 50.485 -137.875 ;
        RECT 50.155 -139.565 50.485 -139.235 ;
        RECT 50.155 -140.925 50.485 -140.595 ;
        RECT 50.155 -142.285 50.485 -141.955 ;
        RECT 50.155 -143.645 50.485 -143.315 ;
        RECT 50.155 -145.005 50.485 -144.675 ;
        RECT 50.155 -146.365 50.485 -146.035 ;
        RECT 50.155 -147.725 50.485 -147.395 ;
        RECT 50.155 -149.085 50.485 -148.755 ;
        RECT 50.155 -150.445 50.485 -150.115 ;
        RECT 50.155 -151.805 50.485 -151.475 ;
        RECT 50.155 -153.165 50.485 -152.835 ;
        RECT 50.155 -154.525 50.485 -154.195 ;
        RECT 50.155 -155.885 50.485 -155.555 ;
        RECT 50.155 -157.245 50.485 -156.915 ;
        RECT 50.155 -158.605 50.485 -158.275 ;
        RECT 50.155 -159.965 50.485 -159.635 ;
        RECT 50.155 -161.325 50.485 -160.995 ;
        RECT 50.155 -162.685 50.485 -162.355 ;
        RECT 50.155 -164.045 50.485 -163.715 ;
        RECT 50.155 -165.405 50.485 -165.075 ;
        RECT 50.155 -166.765 50.485 -166.435 ;
        RECT 50.155 -168.125 50.485 -167.795 ;
        RECT 50.155 -169.485 50.485 -169.155 ;
        RECT 50.155 -170.845 50.485 -170.515 ;
        RECT 50.155 -172.205 50.485 -171.875 ;
        RECT 50.155 -173.565 50.485 -173.235 ;
        RECT 50.155 -174.925 50.485 -174.595 ;
        RECT 50.155 -176.285 50.485 -175.955 ;
        RECT 50.155 -177.645 50.485 -177.315 ;
        RECT 50.155 -179.005 50.485 -178.675 ;
        RECT 50.155 -184.65 50.485 -183.52 ;
        RECT 50.16 -184.765 50.48 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 244.04 51.845 245.17 ;
        RECT 51.515 239.875 51.845 240.205 ;
        RECT 51.515 238.515 51.845 238.845 ;
        RECT 51.515 237.155 51.845 237.485 ;
        RECT 51.52 237.155 51.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 -0.845 51.845 -0.515 ;
        RECT 51.515 -2.205 51.845 -1.875 ;
        RECT 51.515 -3.565 51.845 -3.235 ;
        RECT 51.52 -3.565 51.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 51.515 -96.045 51.845 -95.715 ;
        RECT 51.515 -97.405 51.845 -97.075 ;
        RECT 51.515 -98.765 51.845 -98.435 ;
        RECT 51.515 -100.125 51.845 -99.795 ;
        RECT 51.515 -101.485 51.845 -101.155 ;
        RECT 51.515 -102.845 51.845 -102.515 ;
        RECT 51.515 -104.205 51.845 -103.875 ;
        RECT 51.515 -105.565 51.845 -105.235 ;
        RECT 51.515 -106.925 51.845 -106.595 ;
        RECT 51.515 -108.285 51.845 -107.955 ;
        RECT 51.515 -109.645 51.845 -109.315 ;
        RECT 51.515 -111.005 51.845 -110.675 ;
        RECT 51.515 -112.365 51.845 -112.035 ;
        RECT 51.515 -113.725 51.845 -113.395 ;
        RECT 51.515 -115.085 51.845 -114.755 ;
        RECT 51.515 -116.445 51.845 -116.115 ;
        RECT 51.515 -117.805 51.845 -117.475 ;
        RECT 51.515 -119.165 51.845 -118.835 ;
        RECT 51.515 -120.525 51.845 -120.195 ;
        RECT 51.515 -121.885 51.845 -121.555 ;
        RECT 51.515 -123.245 51.845 -122.915 ;
        RECT 51.515 -124.605 51.845 -124.275 ;
        RECT 51.515 -125.965 51.845 -125.635 ;
        RECT 51.515 -127.325 51.845 -126.995 ;
        RECT 51.515 -128.685 51.845 -128.355 ;
        RECT 51.515 -130.045 51.845 -129.715 ;
        RECT 51.515 -131.405 51.845 -131.075 ;
        RECT 51.515 -132.765 51.845 -132.435 ;
        RECT 51.515 -134.125 51.845 -133.795 ;
        RECT 51.515 -135.485 51.845 -135.155 ;
        RECT 51.515 -136.845 51.845 -136.515 ;
        RECT 51.515 -138.205 51.845 -137.875 ;
        RECT 51.515 -139.565 51.845 -139.235 ;
        RECT 51.515 -140.925 51.845 -140.595 ;
        RECT 51.515 -142.285 51.845 -141.955 ;
        RECT 51.515 -143.645 51.845 -143.315 ;
        RECT 51.515 -145.005 51.845 -144.675 ;
        RECT 51.515 -146.365 51.845 -146.035 ;
        RECT 51.515 -147.725 51.845 -147.395 ;
        RECT 51.515 -149.085 51.845 -148.755 ;
        RECT 51.515 -150.445 51.845 -150.115 ;
        RECT 51.515 -151.805 51.845 -151.475 ;
        RECT 51.515 -153.165 51.845 -152.835 ;
        RECT 51.515 -154.525 51.845 -154.195 ;
        RECT 51.515 -155.885 51.845 -155.555 ;
        RECT 51.515 -157.245 51.845 -156.915 ;
        RECT 51.515 -158.605 51.845 -158.275 ;
        RECT 51.515 -159.965 51.845 -159.635 ;
        RECT 51.515 -161.325 51.845 -160.995 ;
        RECT 51.515 -162.685 51.845 -162.355 ;
        RECT 51.515 -164.045 51.845 -163.715 ;
        RECT 51.515 -165.405 51.845 -165.075 ;
        RECT 51.515 -166.765 51.845 -166.435 ;
        RECT 51.515 -168.125 51.845 -167.795 ;
        RECT 51.515 -169.485 51.845 -169.155 ;
        RECT 51.515 -170.845 51.845 -170.515 ;
        RECT 51.515 -172.205 51.845 -171.875 ;
        RECT 51.515 -173.565 51.845 -173.235 ;
        RECT 51.515 -174.925 51.845 -174.595 ;
        RECT 51.515 -176.285 51.845 -175.955 ;
        RECT 51.515 -177.645 51.845 -177.315 ;
        RECT 51.515 -179.005 51.845 -178.675 ;
        RECT 51.515 -184.65 51.845 -183.52 ;
        RECT 51.52 -184.765 51.84 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 244.04 53.205 245.17 ;
        RECT 52.875 239.875 53.205 240.205 ;
        RECT 52.875 238.515 53.205 238.845 ;
        RECT 52.875 237.155 53.205 237.485 ;
        RECT 52.88 237.155 53.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 -0.845 53.205 -0.515 ;
        RECT 52.875 -2.205 53.205 -1.875 ;
        RECT 52.875 -3.565 53.205 -3.235 ;
        RECT 52.88 -3.565 53.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.875 -96.045 53.205 -95.715 ;
        RECT 52.875 -97.405 53.205 -97.075 ;
        RECT 52.875 -98.765 53.205 -98.435 ;
        RECT 52.875 -100.125 53.205 -99.795 ;
        RECT 52.875 -101.485 53.205 -101.155 ;
        RECT 52.875 -102.845 53.205 -102.515 ;
        RECT 52.875 -104.205 53.205 -103.875 ;
        RECT 52.875 -105.565 53.205 -105.235 ;
        RECT 52.875 -106.925 53.205 -106.595 ;
        RECT 52.875 -108.285 53.205 -107.955 ;
        RECT 52.875 -109.645 53.205 -109.315 ;
        RECT 52.875 -111.005 53.205 -110.675 ;
        RECT 52.875 -112.365 53.205 -112.035 ;
        RECT 52.875 -113.725 53.205 -113.395 ;
        RECT 52.875 -115.085 53.205 -114.755 ;
        RECT 52.875 -116.445 53.205 -116.115 ;
        RECT 52.875 -117.805 53.205 -117.475 ;
        RECT 52.875 -119.165 53.205 -118.835 ;
        RECT 52.875 -120.525 53.205 -120.195 ;
        RECT 52.875 -121.885 53.205 -121.555 ;
        RECT 52.875 -123.245 53.205 -122.915 ;
        RECT 52.875 -124.605 53.205 -124.275 ;
        RECT 52.875 -125.965 53.205 -125.635 ;
        RECT 52.875 -127.325 53.205 -126.995 ;
        RECT 52.875 -128.685 53.205 -128.355 ;
        RECT 52.875 -130.045 53.205 -129.715 ;
        RECT 52.875 -131.405 53.205 -131.075 ;
        RECT 52.875 -132.765 53.205 -132.435 ;
        RECT 52.875 -134.125 53.205 -133.795 ;
        RECT 52.875 -135.485 53.205 -135.155 ;
        RECT 52.875 -136.845 53.205 -136.515 ;
        RECT 52.875 -138.205 53.205 -137.875 ;
        RECT 52.875 -139.565 53.205 -139.235 ;
        RECT 52.875 -140.925 53.205 -140.595 ;
        RECT 52.875 -142.285 53.205 -141.955 ;
        RECT 52.875 -143.645 53.205 -143.315 ;
        RECT 52.875 -145.005 53.205 -144.675 ;
        RECT 52.875 -146.365 53.205 -146.035 ;
        RECT 52.875 -147.725 53.205 -147.395 ;
        RECT 52.875 -149.085 53.205 -148.755 ;
        RECT 52.875 -150.445 53.205 -150.115 ;
        RECT 52.875 -151.805 53.205 -151.475 ;
        RECT 52.875 -153.165 53.205 -152.835 ;
        RECT 52.875 -154.525 53.205 -154.195 ;
        RECT 52.875 -155.885 53.205 -155.555 ;
        RECT 52.875 -157.245 53.205 -156.915 ;
        RECT 52.875 -158.605 53.205 -158.275 ;
        RECT 52.875 -159.965 53.205 -159.635 ;
        RECT 52.875 -161.325 53.205 -160.995 ;
        RECT 52.875 -162.685 53.205 -162.355 ;
        RECT 52.875 -164.045 53.205 -163.715 ;
        RECT 52.875 -165.405 53.205 -165.075 ;
        RECT 52.875 -166.765 53.205 -166.435 ;
        RECT 52.875 -168.125 53.205 -167.795 ;
        RECT 52.875 -169.485 53.205 -169.155 ;
        RECT 52.875 -170.845 53.205 -170.515 ;
        RECT 52.875 -172.205 53.205 -171.875 ;
        RECT 52.875 -173.565 53.205 -173.235 ;
        RECT 52.875 -174.925 53.205 -174.595 ;
        RECT 52.875 -176.285 53.205 -175.955 ;
        RECT 52.875 -177.645 53.205 -177.315 ;
        RECT 52.875 -179.005 53.205 -178.675 ;
        RECT 52.875 -184.65 53.205 -183.52 ;
        RECT 52.88 -184.765 53.2 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 244.04 54.565 245.17 ;
        RECT 54.235 239.875 54.565 240.205 ;
        RECT 54.235 238.515 54.565 238.845 ;
        RECT 54.235 237.155 54.565 237.485 ;
        RECT 54.24 237.155 54.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 -0.845 54.565 -0.515 ;
        RECT 54.235 -2.205 54.565 -1.875 ;
        RECT 54.235 -3.565 54.565 -3.235 ;
        RECT 54.24 -3.565 54.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.235 -96.045 54.565 -95.715 ;
        RECT 54.235 -97.405 54.565 -97.075 ;
        RECT 54.235 -98.765 54.565 -98.435 ;
        RECT 54.235 -100.125 54.565 -99.795 ;
        RECT 54.235 -101.485 54.565 -101.155 ;
        RECT 54.235 -102.845 54.565 -102.515 ;
        RECT 54.235 -104.205 54.565 -103.875 ;
        RECT 54.235 -105.565 54.565 -105.235 ;
        RECT 54.235 -106.925 54.565 -106.595 ;
        RECT 54.235 -108.285 54.565 -107.955 ;
        RECT 54.235 -109.645 54.565 -109.315 ;
        RECT 54.235 -111.005 54.565 -110.675 ;
        RECT 54.235 -112.365 54.565 -112.035 ;
        RECT 54.235 -113.725 54.565 -113.395 ;
        RECT 54.235 -115.085 54.565 -114.755 ;
        RECT 54.235 -116.445 54.565 -116.115 ;
        RECT 54.235 -117.805 54.565 -117.475 ;
        RECT 54.235 -119.165 54.565 -118.835 ;
        RECT 54.235 -120.525 54.565 -120.195 ;
        RECT 54.235 -121.885 54.565 -121.555 ;
        RECT 54.235 -123.245 54.565 -122.915 ;
        RECT 54.235 -124.605 54.565 -124.275 ;
        RECT 54.235 -125.965 54.565 -125.635 ;
        RECT 54.235 -127.325 54.565 -126.995 ;
        RECT 54.235 -128.685 54.565 -128.355 ;
        RECT 54.235 -130.045 54.565 -129.715 ;
        RECT 54.235 -131.405 54.565 -131.075 ;
        RECT 54.235 -132.765 54.565 -132.435 ;
        RECT 54.235 -134.125 54.565 -133.795 ;
        RECT 54.235 -135.485 54.565 -135.155 ;
        RECT 54.235 -136.845 54.565 -136.515 ;
        RECT 54.235 -138.205 54.565 -137.875 ;
        RECT 54.235 -139.565 54.565 -139.235 ;
        RECT 54.235 -140.925 54.565 -140.595 ;
        RECT 54.235 -142.285 54.565 -141.955 ;
        RECT 54.235 -143.645 54.565 -143.315 ;
        RECT 54.235 -145.005 54.565 -144.675 ;
        RECT 54.235 -146.365 54.565 -146.035 ;
        RECT 54.235 -147.725 54.565 -147.395 ;
        RECT 54.235 -149.085 54.565 -148.755 ;
        RECT 54.235 -150.445 54.565 -150.115 ;
        RECT 54.235 -151.805 54.565 -151.475 ;
        RECT 54.235 -153.165 54.565 -152.835 ;
        RECT 54.235 -154.525 54.565 -154.195 ;
        RECT 54.235 -155.885 54.565 -155.555 ;
        RECT 54.235 -157.245 54.565 -156.915 ;
        RECT 54.235 -158.605 54.565 -158.275 ;
        RECT 54.235 -159.965 54.565 -159.635 ;
        RECT 54.235 -161.325 54.565 -160.995 ;
        RECT 54.235 -162.685 54.565 -162.355 ;
        RECT 54.235 -164.045 54.565 -163.715 ;
        RECT 54.235 -165.405 54.565 -165.075 ;
        RECT 54.235 -166.765 54.565 -166.435 ;
        RECT 54.235 -168.125 54.565 -167.795 ;
        RECT 54.235 -169.485 54.565 -169.155 ;
        RECT 54.235 -170.845 54.565 -170.515 ;
        RECT 54.235 -172.205 54.565 -171.875 ;
        RECT 54.235 -173.565 54.565 -173.235 ;
        RECT 54.235 -174.925 54.565 -174.595 ;
        RECT 54.235 -176.285 54.565 -175.955 ;
        RECT 54.235 -177.645 54.565 -177.315 ;
        RECT 54.235 -179.005 54.565 -178.675 ;
        RECT 54.235 -184.65 54.565 -183.52 ;
        RECT 54.24 -184.765 54.56 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 244.04 55.925 245.17 ;
        RECT 55.595 239.875 55.925 240.205 ;
        RECT 55.595 238.515 55.925 238.845 ;
        RECT 55.595 237.155 55.925 237.485 ;
        RECT 55.6 237.155 55.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 -0.845 55.925 -0.515 ;
        RECT 55.595 -2.205 55.925 -1.875 ;
        RECT 55.595 -3.565 55.925 -3.235 ;
        RECT 55.6 -3.565 55.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 55.595 -96.045 55.925 -95.715 ;
        RECT 55.595 -97.405 55.925 -97.075 ;
        RECT 55.595 -98.765 55.925 -98.435 ;
        RECT 55.595 -100.125 55.925 -99.795 ;
        RECT 55.595 -101.485 55.925 -101.155 ;
        RECT 55.595 -102.845 55.925 -102.515 ;
        RECT 55.595 -104.205 55.925 -103.875 ;
        RECT 55.595 -105.565 55.925 -105.235 ;
        RECT 55.595 -106.925 55.925 -106.595 ;
        RECT 55.595 -108.285 55.925 -107.955 ;
        RECT 55.595 -109.645 55.925 -109.315 ;
        RECT 55.595 -111.005 55.925 -110.675 ;
        RECT 55.595 -112.365 55.925 -112.035 ;
        RECT 55.595 -113.725 55.925 -113.395 ;
        RECT 55.595 -115.085 55.925 -114.755 ;
        RECT 55.595 -116.445 55.925 -116.115 ;
        RECT 55.595 -117.805 55.925 -117.475 ;
        RECT 55.595 -119.165 55.925 -118.835 ;
        RECT 55.595 -120.525 55.925 -120.195 ;
        RECT 55.595 -121.885 55.925 -121.555 ;
        RECT 55.595 -123.245 55.925 -122.915 ;
        RECT 55.595 -124.605 55.925 -124.275 ;
        RECT 55.595 -125.965 55.925 -125.635 ;
        RECT 55.595 -127.325 55.925 -126.995 ;
        RECT 55.595 -128.685 55.925 -128.355 ;
        RECT 55.595 -130.045 55.925 -129.715 ;
        RECT 55.595 -131.405 55.925 -131.075 ;
        RECT 55.595 -132.765 55.925 -132.435 ;
        RECT 55.595 -134.125 55.925 -133.795 ;
        RECT 55.595 -135.485 55.925 -135.155 ;
        RECT 55.595 -136.845 55.925 -136.515 ;
        RECT 55.595 -138.205 55.925 -137.875 ;
        RECT 55.595 -139.565 55.925 -139.235 ;
        RECT 55.595 -140.925 55.925 -140.595 ;
        RECT 55.595 -142.285 55.925 -141.955 ;
        RECT 55.595 -143.645 55.925 -143.315 ;
        RECT 55.595 -145.005 55.925 -144.675 ;
        RECT 55.595 -146.365 55.925 -146.035 ;
        RECT 55.595 -147.725 55.925 -147.395 ;
        RECT 55.595 -149.085 55.925 -148.755 ;
        RECT 55.595 -150.445 55.925 -150.115 ;
        RECT 55.595 -151.805 55.925 -151.475 ;
        RECT 55.595 -153.165 55.925 -152.835 ;
        RECT 55.595 -154.525 55.925 -154.195 ;
        RECT 55.595 -155.885 55.925 -155.555 ;
        RECT 55.595 -157.245 55.925 -156.915 ;
        RECT 55.595 -158.605 55.925 -158.275 ;
        RECT 55.595 -159.965 55.925 -159.635 ;
        RECT 55.595 -161.325 55.925 -160.995 ;
        RECT 55.595 -162.685 55.925 -162.355 ;
        RECT 55.595 -164.045 55.925 -163.715 ;
        RECT 55.595 -165.405 55.925 -165.075 ;
        RECT 55.595 -166.765 55.925 -166.435 ;
        RECT 55.595 -168.125 55.925 -167.795 ;
        RECT 55.595 -169.485 55.925 -169.155 ;
        RECT 55.595 -170.845 55.925 -170.515 ;
        RECT 55.595 -172.205 55.925 -171.875 ;
        RECT 55.595 -173.565 55.925 -173.235 ;
        RECT 55.595 -174.925 55.925 -174.595 ;
        RECT 55.595 -176.285 55.925 -175.955 ;
        RECT 55.595 -177.645 55.925 -177.315 ;
        RECT 55.595 -179.005 55.925 -178.675 ;
        RECT 55.595 -184.65 55.925 -183.52 ;
        RECT 55.6 -184.765 55.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 244.04 57.285 245.17 ;
        RECT 56.955 239.875 57.285 240.205 ;
        RECT 56.955 238.515 57.285 238.845 ;
        RECT 56.955 237.155 57.285 237.485 ;
        RECT 56.96 237.155 57.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.955 -98.765 57.285 -98.435 ;
        RECT 56.955 -100.125 57.285 -99.795 ;
        RECT 56.955 -101.485 57.285 -101.155 ;
        RECT 56.955 -102.845 57.285 -102.515 ;
        RECT 56.955 -104.205 57.285 -103.875 ;
        RECT 56.955 -105.565 57.285 -105.235 ;
        RECT 56.955 -106.925 57.285 -106.595 ;
        RECT 56.955 -108.285 57.285 -107.955 ;
        RECT 56.955 -109.645 57.285 -109.315 ;
        RECT 56.955 -111.005 57.285 -110.675 ;
        RECT 56.955 -112.365 57.285 -112.035 ;
        RECT 56.955 -113.725 57.285 -113.395 ;
        RECT 56.955 -115.085 57.285 -114.755 ;
        RECT 56.955 -116.445 57.285 -116.115 ;
        RECT 56.955 -117.805 57.285 -117.475 ;
        RECT 56.955 -119.165 57.285 -118.835 ;
        RECT 56.955 -120.525 57.285 -120.195 ;
        RECT 56.955 -121.885 57.285 -121.555 ;
        RECT 56.955 -123.245 57.285 -122.915 ;
        RECT 56.955 -124.605 57.285 -124.275 ;
        RECT 56.955 -125.965 57.285 -125.635 ;
        RECT 56.955 -127.325 57.285 -126.995 ;
        RECT 56.955 -128.685 57.285 -128.355 ;
        RECT 56.955 -130.045 57.285 -129.715 ;
        RECT 56.955 -131.405 57.285 -131.075 ;
        RECT 56.955 -132.765 57.285 -132.435 ;
        RECT 56.955 -134.125 57.285 -133.795 ;
        RECT 56.955 -135.485 57.285 -135.155 ;
        RECT 56.955 -136.845 57.285 -136.515 ;
        RECT 56.955 -138.205 57.285 -137.875 ;
        RECT 56.955 -139.565 57.285 -139.235 ;
        RECT 56.955 -140.925 57.285 -140.595 ;
        RECT 56.955 -142.285 57.285 -141.955 ;
        RECT 56.955 -143.645 57.285 -143.315 ;
        RECT 56.955 -145.005 57.285 -144.675 ;
        RECT 56.955 -146.365 57.285 -146.035 ;
        RECT 56.955 -147.725 57.285 -147.395 ;
        RECT 56.955 -149.085 57.285 -148.755 ;
        RECT 56.955 -150.445 57.285 -150.115 ;
        RECT 56.955 -151.805 57.285 -151.475 ;
        RECT 56.955 -153.165 57.285 -152.835 ;
        RECT 56.955 -154.525 57.285 -154.195 ;
        RECT 56.955 -155.885 57.285 -155.555 ;
        RECT 56.955 -157.245 57.285 -156.915 ;
        RECT 56.955 -158.605 57.285 -158.275 ;
        RECT 56.955 -159.965 57.285 -159.635 ;
        RECT 56.955 -161.325 57.285 -160.995 ;
        RECT 56.955 -162.685 57.285 -162.355 ;
        RECT 56.955 -164.045 57.285 -163.715 ;
        RECT 56.955 -165.405 57.285 -165.075 ;
        RECT 56.955 -166.765 57.285 -166.435 ;
        RECT 56.955 -168.125 57.285 -167.795 ;
        RECT 56.955 -169.485 57.285 -169.155 ;
        RECT 56.955 -170.845 57.285 -170.515 ;
        RECT 56.955 -172.205 57.285 -171.875 ;
        RECT 56.955 -173.565 57.285 -173.235 ;
        RECT 56.955 -174.925 57.285 -174.595 ;
        RECT 56.955 -176.285 57.285 -175.955 ;
        RECT 56.955 -177.645 57.285 -177.315 ;
        RECT 56.955 -179.005 57.285 -178.675 ;
        RECT 56.955 -184.65 57.285 -183.52 ;
        RECT 56.96 -184.765 57.28 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.16 -98.075 57.49 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.315 244.04 58.645 245.17 ;
        RECT 58.315 239.875 58.645 240.205 ;
        RECT 58.315 238.515 58.645 238.845 ;
        RECT 58.315 237.155 58.645 237.485 ;
        RECT 58.32 237.155 58.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 244.04 60.005 245.17 ;
        RECT 59.675 239.875 60.005 240.205 ;
        RECT 59.675 238.515 60.005 238.845 ;
        RECT 59.675 237.155 60.005 237.485 ;
        RECT 59.68 237.155 60 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 59.675 -0.845 60.005 -0.515 ;
        RECT 59.675 -2.205 60.005 -1.875 ;
        RECT 59.675 -3.565 60.005 -3.235 ;
        RECT 59.68 -3.565 60 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 244.04 61.365 245.17 ;
        RECT 61.035 239.875 61.365 240.205 ;
        RECT 61.035 238.515 61.365 238.845 ;
        RECT 61.035 237.155 61.365 237.485 ;
        RECT 61.04 237.155 61.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 -0.845 61.365 -0.515 ;
        RECT 61.035 -2.205 61.365 -1.875 ;
        RECT 61.035 -3.565 61.365 -3.235 ;
        RECT 61.04 -3.565 61.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.035 -124.605 61.365 -124.275 ;
        RECT 61.035 -125.965 61.365 -125.635 ;
        RECT 61.035 -127.325 61.365 -126.995 ;
        RECT 61.035 -128.685 61.365 -128.355 ;
        RECT 61.035 -130.045 61.365 -129.715 ;
        RECT 61.035 -131.405 61.365 -131.075 ;
        RECT 61.035 -132.765 61.365 -132.435 ;
        RECT 61.035 -134.125 61.365 -133.795 ;
        RECT 61.035 -135.485 61.365 -135.155 ;
        RECT 61.035 -136.845 61.365 -136.515 ;
        RECT 61.035 -138.205 61.365 -137.875 ;
        RECT 61.035 -139.565 61.365 -139.235 ;
        RECT 61.035 -140.925 61.365 -140.595 ;
        RECT 61.035 -142.285 61.365 -141.955 ;
        RECT 61.035 -143.645 61.365 -143.315 ;
        RECT 61.035 -145.005 61.365 -144.675 ;
        RECT 61.035 -146.365 61.365 -146.035 ;
        RECT 61.035 -147.725 61.365 -147.395 ;
        RECT 61.035 -149.085 61.365 -148.755 ;
        RECT 61.035 -150.445 61.365 -150.115 ;
        RECT 61.035 -151.805 61.365 -151.475 ;
        RECT 61.035 -153.165 61.365 -152.835 ;
        RECT 61.035 -154.525 61.365 -154.195 ;
        RECT 61.035 -155.885 61.365 -155.555 ;
        RECT 61.035 -157.245 61.365 -156.915 ;
        RECT 61.035 -158.605 61.365 -158.275 ;
        RECT 61.035 -159.965 61.365 -159.635 ;
        RECT 61.035 -161.325 61.365 -160.995 ;
        RECT 61.035 -162.685 61.365 -162.355 ;
        RECT 61.035 -164.045 61.365 -163.715 ;
        RECT 61.035 -165.405 61.365 -165.075 ;
        RECT 61.035 -166.765 61.365 -166.435 ;
        RECT 61.035 -168.125 61.365 -167.795 ;
        RECT 61.035 -169.485 61.365 -169.155 ;
        RECT 61.035 -170.845 61.365 -170.515 ;
        RECT 61.035 -172.205 61.365 -171.875 ;
        RECT 61.035 -173.565 61.365 -173.235 ;
        RECT 61.035 -174.925 61.365 -174.595 ;
        RECT 61.035 -176.285 61.365 -175.955 ;
        RECT 61.035 -177.645 61.365 -177.315 ;
        RECT 61.035 -179.005 61.365 -178.675 ;
        RECT 61.035 -184.65 61.365 -183.52 ;
        RECT 61.04 -184.765 61.36 -95.04 ;
        RECT 61.035 -96.045 61.365 -95.715 ;
        RECT 61.035 -97.405 61.365 -97.075 ;
        RECT 61.035 -98.765 61.365 -98.435 ;
        RECT 61.035 -100.125 61.365 -99.795 ;
        RECT 61.035 -101.485 61.365 -101.155 ;
        RECT 61.035 -102.845 61.365 -102.515 ;
        RECT 61.035 -104.205 61.365 -103.875 ;
        RECT 61.035 -105.565 61.365 -105.235 ;
        RECT 61.035 -106.925 61.365 -106.595 ;
        RECT 61.035 -108.285 61.365 -107.955 ;
        RECT 61.035 -109.645 61.365 -109.315 ;
        RECT 61.035 -111.005 61.365 -110.675 ;
        RECT 61.035 -112.365 61.365 -112.035 ;
        RECT 61.035 -113.725 61.365 -113.395 ;
        RECT 61.035 -115.085 61.365 -114.755 ;
        RECT 61.035 -116.445 61.365 -116.115 ;
        RECT 61.035 -117.805 61.365 -117.475 ;
        RECT 61.035 -119.165 61.365 -118.835 ;
        RECT 61.035 -120.525 61.365 -120.195 ;
        RECT 61.035 -121.885 61.365 -121.555 ;
        RECT 61.035 -123.245 61.365 -122.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 244.04 12.405 245.17 ;
        RECT 12.075 239.875 12.405 240.205 ;
        RECT 12.075 238.515 12.405 238.845 ;
        RECT 12.075 237.155 12.405 237.485 ;
        RECT 12.08 237.155 12.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 -0.845 12.405 -0.515 ;
        RECT 12.075 -2.205 12.405 -1.875 ;
        RECT 12.075 -3.565 12.405 -3.235 ;
        RECT 12.08 -3.565 12.4 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.075 -96.045 12.405 -95.715 ;
        RECT 12.075 -97.405 12.405 -97.075 ;
        RECT 12.075 -98.765 12.405 -98.435 ;
        RECT 12.075 -100.125 12.405 -99.795 ;
        RECT 12.075 -101.485 12.405 -101.155 ;
        RECT 12.075 -102.845 12.405 -102.515 ;
        RECT 12.075 -104.205 12.405 -103.875 ;
        RECT 12.075 -105.565 12.405 -105.235 ;
        RECT 12.075 -106.925 12.405 -106.595 ;
        RECT 12.075 -108.285 12.405 -107.955 ;
        RECT 12.075 -109.645 12.405 -109.315 ;
        RECT 12.075 -111.005 12.405 -110.675 ;
        RECT 12.075 -112.365 12.405 -112.035 ;
        RECT 12.075 -113.725 12.405 -113.395 ;
        RECT 12.075 -115.085 12.405 -114.755 ;
        RECT 12.075 -116.445 12.405 -116.115 ;
        RECT 12.075 -117.805 12.405 -117.475 ;
        RECT 12.075 -119.165 12.405 -118.835 ;
        RECT 12.075 -120.525 12.405 -120.195 ;
        RECT 12.075 -121.885 12.405 -121.555 ;
        RECT 12.075 -123.245 12.405 -122.915 ;
        RECT 12.075 -124.605 12.405 -124.275 ;
        RECT 12.075 -125.965 12.405 -125.635 ;
        RECT 12.075 -127.325 12.405 -126.995 ;
        RECT 12.075 -128.685 12.405 -128.355 ;
        RECT 12.075 -130.045 12.405 -129.715 ;
        RECT 12.075 -131.405 12.405 -131.075 ;
        RECT 12.075 -132.765 12.405 -132.435 ;
        RECT 12.075 -134.125 12.405 -133.795 ;
        RECT 12.075 -135.485 12.405 -135.155 ;
        RECT 12.075 -136.845 12.405 -136.515 ;
        RECT 12.075 -138.205 12.405 -137.875 ;
        RECT 12.075 -139.565 12.405 -139.235 ;
        RECT 12.075 -140.925 12.405 -140.595 ;
        RECT 12.075 -142.285 12.405 -141.955 ;
        RECT 12.075 -143.645 12.405 -143.315 ;
        RECT 12.075 -145.005 12.405 -144.675 ;
        RECT 12.075 -146.365 12.405 -146.035 ;
        RECT 12.075 -147.725 12.405 -147.395 ;
        RECT 12.075 -149.085 12.405 -148.755 ;
        RECT 12.075 -150.445 12.405 -150.115 ;
        RECT 12.075 -151.805 12.405 -151.475 ;
        RECT 12.075 -153.165 12.405 -152.835 ;
        RECT 12.075 -154.525 12.405 -154.195 ;
        RECT 12.075 -155.885 12.405 -155.555 ;
        RECT 12.075 -157.245 12.405 -156.915 ;
        RECT 12.075 -158.605 12.405 -158.275 ;
        RECT 12.075 -159.965 12.405 -159.635 ;
        RECT 12.075 -161.325 12.405 -160.995 ;
        RECT 12.075 -162.685 12.405 -162.355 ;
        RECT 12.075 -164.045 12.405 -163.715 ;
        RECT 12.075 -165.405 12.405 -165.075 ;
        RECT 12.075 -166.765 12.405 -166.435 ;
        RECT 12.075 -168.125 12.405 -167.795 ;
        RECT 12.075 -169.485 12.405 -169.155 ;
        RECT 12.075 -170.845 12.405 -170.515 ;
        RECT 12.075 -172.205 12.405 -171.875 ;
        RECT 12.075 -173.565 12.405 -173.235 ;
        RECT 12.075 -174.925 12.405 -174.595 ;
        RECT 12.075 -176.285 12.405 -175.955 ;
        RECT 12.075 -177.645 12.405 -177.315 ;
        RECT 12.075 -179.005 12.405 -178.675 ;
        RECT 12.075 -184.65 12.405 -183.52 ;
        RECT 12.08 -184.765 12.4 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 244.04 13.765 245.17 ;
        RECT 13.435 239.875 13.765 240.205 ;
        RECT 13.435 238.515 13.765 238.845 ;
        RECT 13.435 237.155 13.765 237.485 ;
        RECT 13.44 237.155 13.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.435 -98.765 13.765 -98.435 ;
        RECT 13.435 -100.125 13.765 -99.795 ;
        RECT 13.435 -101.485 13.765 -101.155 ;
        RECT 13.435 -102.845 13.765 -102.515 ;
        RECT 13.435 -104.205 13.765 -103.875 ;
        RECT 13.435 -105.565 13.765 -105.235 ;
        RECT 13.435 -106.925 13.765 -106.595 ;
        RECT 13.435 -108.285 13.765 -107.955 ;
        RECT 13.435 -109.645 13.765 -109.315 ;
        RECT 13.435 -111.005 13.765 -110.675 ;
        RECT 13.435 -112.365 13.765 -112.035 ;
        RECT 13.435 -113.725 13.765 -113.395 ;
        RECT 13.435 -115.085 13.765 -114.755 ;
        RECT 13.435 -116.445 13.765 -116.115 ;
        RECT 13.435 -117.805 13.765 -117.475 ;
        RECT 13.435 -119.165 13.765 -118.835 ;
        RECT 13.435 -120.525 13.765 -120.195 ;
        RECT 13.435 -121.885 13.765 -121.555 ;
        RECT 13.435 -123.245 13.765 -122.915 ;
        RECT 13.435 -124.605 13.765 -124.275 ;
        RECT 13.435 -125.965 13.765 -125.635 ;
        RECT 13.435 -127.325 13.765 -126.995 ;
        RECT 13.435 -128.685 13.765 -128.355 ;
        RECT 13.435 -130.045 13.765 -129.715 ;
        RECT 13.435 -131.405 13.765 -131.075 ;
        RECT 13.435 -132.765 13.765 -132.435 ;
        RECT 13.435 -134.125 13.765 -133.795 ;
        RECT 13.435 -135.485 13.765 -135.155 ;
        RECT 13.435 -136.845 13.765 -136.515 ;
        RECT 13.435 -138.205 13.765 -137.875 ;
        RECT 13.435 -139.565 13.765 -139.235 ;
        RECT 13.435 -140.925 13.765 -140.595 ;
        RECT 13.435 -142.285 13.765 -141.955 ;
        RECT 13.435 -143.645 13.765 -143.315 ;
        RECT 13.435 -145.005 13.765 -144.675 ;
        RECT 13.435 -146.365 13.765 -146.035 ;
        RECT 13.435 -147.725 13.765 -147.395 ;
        RECT 13.435 -149.085 13.765 -148.755 ;
        RECT 13.435 -150.445 13.765 -150.115 ;
        RECT 13.435 -151.805 13.765 -151.475 ;
        RECT 13.435 -153.165 13.765 -152.835 ;
        RECT 13.435 -154.525 13.765 -154.195 ;
        RECT 13.435 -155.885 13.765 -155.555 ;
        RECT 13.435 -157.245 13.765 -156.915 ;
        RECT 13.435 -158.605 13.765 -158.275 ;
        RECT 13.435 -159.965 13.765 -159.635 ;
        RECT 13.435 -161.325 13.765 -160.995 ;
        RECT 13.435 -162.685 13.765 -162.355 ;
        RECT 13.435 -164.045 13.765 -163.715 ;
        RECT 13.435 -165.405 13.765 -165.075 ;
        RECT 13.435 -166.765 13.765 -166.435 ;
        RECT 13.435 -168.125 13.765 -167.795 ;
        RECT 13.435 -169.485 13.765 -169.155 ;
        RECT 13.435 -170.845 13.765 -170.515 ;
        RECT 13.435 -172.205 13.765 -171.875 ;
        RECT 13.435 -173.565 13.765 -173.235 ;
        RECT 13.435 -174.925 13.765 -174.595 ;
        RECT 13.435 -176.285 13.765 -175.955 ;
        RECT 13.435 -177.645 13.765 -177.315 ;
        RECT 13.435 -179.005 13.765 -178.675 ;
        RECT 13.435 -184.65 13.765 -183.52 ;
        RECT 13.44 -184.765 13.76 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 13.56 -98.075 13.89 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.795 244.04 15.125 245.17 ;
        RECT 14.795 239.875 15.125 240.205 ;
        RECT 14.795 238.515 15.125 238.845 ;
        RECT 14.795 237.155 15.125 237.485 ;
        RECT 14.8 237.155 15.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.155 244.04 16.485 245.17 ;
        RECT 16.155 239.875 16.485 240.205 ;
        RECT 16.155 238.515 16.485 238.845 ;
        RECT 16.155 237.155 16.485 237.485 ;
        RECT 16.16 237.155 16.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.155 -0.845 16.485 -0.515 ;
        RECT 16.155 -2.205 16.485 -1.875 ;
        RECT 16.155 -3.565 16.485 -3.235 ;
        RECT 16.16 -3.565 16.48 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 244.04 17.845 245.17 ;
        RECT 17.515 239.875 17.845 240.205 ;
        RECT 17.515 238.515 17.845 238.845 ;
        RECT 17.515 237.155 17.845 237.485 ;
        RECT 17.52 237.155 17.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 -0.845 17.845 -0.515 ;
        RECT 17.515 -2.205 17.845 -1.875 ;
        RECT 17.515 -3.565 17.845 -3.235 ;
        RECT 17.52 -3.565 17.84 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 17.515 -96.045 17.845 -95.715 ;
        RECT 17.515 -97.405 17.845 -97.075 ;
        RECT 17.515 -98.765 17.845 -98.435 ;
        RECT 17.515 -100.125 17.845 -99.795 ;
        RECT 17.515 -101.485 17.845 -101.155 ;
        RECT 17.515 -102.845 17.845 -102.515 ;
        RECT 17.515 -104.205 17.845 -103.875 ;
        RECT 17.515 -105.565 17.845 -105.235 ;
        RECT 17.515 -106.925 17.845 -106.595 ;
        RECT 17.515 -108.285 17.845 -107.955 ;
        RECT 17.515 -109.645 17.845 -109.315 ;
        RECT 17.515 -111.005 17.845 -110.675 ;
        RECT 17.515 -112.365 17.845 -112.035 ;
        RECT 17.515 -113.725 17.845 -113.395 ;
        RECT 17.515 -115.085 17.845 -114.755 ;
        RECT 17.515 -116.445 17.845 -116.115 ;
        RECT 17.515 -117.805 17.845 -117.475 ;
        RECT 17.515 -119.165 17.845 -118.835 ;
        RECT 17.515 -120.525 17.845 -120.195 ;
        RECT 17.515 -121.885 17.845 -121.555 ;
        RECT 17.515 -123.245 17.845 -122.915 ;
        RECT 17.515 -124.605 17.845 -124.275 ;
        RECT 17.515 -125.965 17.845 -125.635 ;
        RECT 17.515 -127.325 17.845 -126.995 ;
        RECT 17.515 -128.685 17.845 -128.355 ;
        RECT 17.515 -130.045 17.845 -129.715 ;
        RECT 17.515 -131.405 17.845 -131.075 ;
        RECT 17.515 -132.765 17.845 -132.435 ;
        RECT 17.515 -134.125 17.845 -133.795 ;
        RECT 17.515 -135.485 17.845 -135.155 ;
        RECT 17.515 -136.845 17.845 -136.515 ;
        RECT 17.515 -138.205 17.845 -137.875 ;
        RECT 17.515 -139.565 17.845 -139.235 ;
        RECT 17.515 -140.925 17.845 -140.595 ;
        RECT 17.515 -142.285 17.845 -141.955 ;
        RECT 17.515 -143.645 17.845 -143.315 ;
        RECT 17.515 -145.005 17.845 -144.675 ;
        RECT 17.515 -146.365 17.845 -146.035 ;
        RECT 17.515 -147.725 17.845 -147.395 ;
        RECT 17.515 -149.085 17.845 -148.755 ;
        RECT 17.515 -150.445 17.845 -150.115 ;
        RECT 17.515 -151.805 17.845 -151.475 ;
        RECT 17.515 -153.165 17.845 -152.835 ;
        RECT 17.515 -154.525 17.845 -154.195 ;
        RECT 17.515 -155.885 17.845 -155.555 ;
        RECT 17.515 -157.245 17.845 -156.915 ;
        RECT 17.515 -158.605 17.845 -158.275 ;
        RECT 17.515 -159.965 17.845 -159.635 ;
        RECT 17.515 -161.325 17.845 -160.995 ;
        RECT 17.515 -162.685 17.845 -162.355 ;
        RECT 17.515 -164.045 17.845 -163.715 ;
        RECT 17.515 -165.405 17.845 -165.075 ;
        RECT 17.515 -166.765 17.845 -166.435 ;
        RECT 17.515 -168.125 17.845 -167.795 ;
        RECT 17.515 -169.485 17.845 -169.155 ;
        RECT 17.515 -170.845 17.845 -170.515 ;
        RECT 17.515 -172.205 17.845 -171.875 ;
        RECT 17.515 -173.565 17.845 -173.235 ;
        RECT 17.515 -174.925 17.845 -174.595 ;
        RECT 17.515 -176.285 17.845 -175.955 ;
        RECT 17.515 -177.645 17.845 -177.315 ;
        RECT 17.515 -179.005 17.845 -178.675 ;
        RECT 17.515 -184.65 17.845 -183.52 ;
        RECT 17.52 -184.765 17.84 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 244.04 19.205 245.17 ;
        RECT 18.875 239.875 19.205 240.205 ;
        RECT 18.875 238.515 19.205 238.845 ;
        RECT 18.875 237.155 19.205 237.485 ;
        RECT 18.88 237.155 19.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 -0.845 19.205 -0.515 ;
        RECT 18.875 -2.205 19.205 -1.875 ;
        RECT 18.875 -3.565 19.205 -3.235 ;
        RECT 18.88 -3.565 19.2 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.875 -96.045 19.205 -95.715 ;
        RECT 18.875 -97.405 19.205 -97.075 ;
        RECT 18.875 -98.765 19.205 -98.435 ;
        RECT 18.875 -100.125 19.205 -99.795 ;
        RECT 18.875 -101.485 19.205 -101.155 ;
        RECT 18.875 -102.845 19.205 -102.515 ;
        RECT 18.875 -104.205 19.205 -103.875 ;
        RECT 18.875 -105.565 19.205 -105.235 ;
        RECT 18.875 -106.925 19.205 -106.595 ;
        RECT 18.875 -108.285 19.205 -107.955 ;
        RECT 18.875 -109.645 19.205 -109.315 ;
        RECT 18.875 -111.005 19.205 -110.675 ;
        RECT 18.875 -112.365 19.205 -112.035 ;
        RECT 18.875 -113.725 19.205 -113.395 ;
        RECT 18.875 -115.085 19.205 -114.755 ;
        RECT 18.875 -116.445 19.205 -116.115 ;
        RECT 18.875 -117.805 19.205 -117.475 ;
        RECT 18.875 -119.165 19.205 -118.835 ;
        RECT 18.875 -120.525 19.205 -120.195 ;
        RECT 18.875 -121.885 19.205 -121.555 ;
        RECT 18.875 -123.245 19.205 -122.915 ;
        RECT 18.875 -124.605 19.205 -124.275 ;
        RECT 18.875 -125.965 19.205 -125.635 ;
        RECT 18.875 -127.325 19.205 -126.995 ;
        RECT 18.875 -128.685 19.205 -128.355 ;
        RECT 18.875 -130.045 19.205 -129.715 ;
        RECT 18.875 -131.405 19.205 -131.075 ;
        RECT 18.875 -132.765 19.205 -132.435 ;
        RECT 18.875 -134.125 19.205 -133.795 ;
        RECT 18.875 -135.485 19.205 -135.155 ;
        RECT 18.875 -136.845 19.205 -136.515 ;
        RECT 18.875 -138.205 19.205 -137.875 ;
        RECT 18.875 -139.565 19.205 -139.235 ;
        RECT 18.875 -140.925 19.205 -140.595 ;
        RECT 18.875 -142.285 19.205 -141.955 ;
        RECT 18.875 -143.645 19.205 -143.315 ;
        RECT 18.875 -145.005 19.205 -144.675 ;
        RECT 18.875 -146.365 19.205 -146.035 ;
        RECT 18.875 -147.725 19.205 -147.395 ;
        RECT 18.875 -149.085 19.205 -148.755 ;
        RECT 18.875 -150.445 19.205 -150.115 ;
        RECT 18.875 -151.805 19.205 -151.475 ;
        RECT 18.875 -153.165 19.205 -152.835 ;
        RECT 18.875 -154.525 19.205 -154.195 ;
        RECT 18.875 -155.885 19.205 -155.555 ;
        RECT 18.875 -157.245 19.205 -156.915 ;
        RECT 18.875 -158.605 19.205 -158.275 ;
        RECT 18.875 -159.965 19.205 -159.635 ;
        RECT 18.875 -161.325 19.205 -160.995 ;
        RECT 18.875 -162.685 19.205 -162.355 ;
        RECT 18.875 -164.045 19.205 -163.715 ;
        RECT 18.875 -165.405 19.205 -165.075 ;
        RECT 18.875 -166.765 19.205 -166.435 ;
        RECT 18.875 -168.125 19.205 -167.795 ;
        RECT 18.875 -169.485 19.205 -169.155 ;
        RECT 18.875 -170.845 19.205 -170.515 ;
        RECT 18.875 -172.205 19.205 -171.875 ;
        RECT 18.875 -173.565 19.205 -173.235 ;
        RECT 18.875 -174.925 19.205 -174.595 ;
        RECT 18.875 -176.285 19.205 -175.955 ;
        RECT 18.875 -177.645 19.205 -177.315 ;
        RECT 18.875 -179.005 19.205 -178.675 ;
        RECT 18.875 -184.65 19.205 -183.52 ;
        RECT 18.88 -184.765 19.2 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 244.04 20.565 245.17 ;
        RECT 20.235 239.875 20.565 240.205 ;
        RECT 20.235 238.515 20.565 238.845 ;
        RECT 20.235 237.155 20.565 237.485 ;
        RECT 20.24 237.155 20.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 -0.845 20.565 -0.515 ;
        RECT 20.235 -2.205 20.565 -1.875 ;
        RECT 20.235 -3.565 20.565 -3.235 ;
        RECT 20.24 -3.565 20.56 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.235 -96.045 20.565 -95.715 ;
        RECT 20.235 -97.405 20.565 -97.075 ;
        RECT 20.235 -98.765 20.565 -98.435 ;
        RECT 20.235 -100.125 20.565 -99.795 ;
        RECT 20.235 -101.485 20.565 -101.155 ;
        RECT 20.235 -102.845 20.565 -102.515 ;
        RECT 20.235 -104.205 20.565 -103.875 ;
        RECT 20.235 -105.565 20.565 -105.235 ;
        RECT 20.235 -106.925 20.565 -106.595 ;
        RECT 20.235 -108.285 20.565 -107.955 ;
        RECT 20.235 -109.645 20.565 -109.315 ;
        RECT 20.235 -111.005 20.565 -110.675 ;
        RECT 20.235 -112.365 20.565 -112.035 ;
        RECT 20.235 -113.725 20.565 -113.395 ;
        RECT 20.235 -115.085 20.565 -114.755 ;
        RECT 20.235 -116.445 20.565 -116.115 ;
        RECT 20.235 -117.805 20.565 -117.475 ;
        RECT 20.235 -119.165 20.565 -118.835 ;
        RECT 20.235 -120.525 20.565 -120.195 ;
        RECT 20.235 -121.885 20.565 -121.555 ;
        RECT 20.235 -123.245 20.565 -122.915 ;
        RECT 20.235 -124.605 20.565 -124.275 ;
        RECT 20.235 -125.965 20.565 -125.635 ;
        RECT 20.235 -127.325 20.565 -126.995 ;
        RECT 20.235 -128.685 20.565 -128.355 ;
        RECT 20.235 -130.045 20.565 -129.715 ;
        RECT 20.235 -131.405 20.565 -131.075 ;
        RECT 20.235 -132.765 20.565 -132.435 ;
        RECT 20.235 -134.125 20.565 -133.795 ;
        RECT 20.235 -135.485 20.565 -135.155 ;
        RECT 20.235 -136.845 20.565 -136.515 ;
        RECT 20.235 -138.205 20.565 -137.875 ;
        RECT 20.235 -139.565 20.565 -139.235 ;
        RECT 20.235 -140.925 20.565 -140.595 ;
        RECT 20.235 -142.285 20.565 -141.955 ;
        RECT 20.235 -143.645 20.565 -143.315 ;
        RECT 20.235 -145.005 20.565 -144.675 ;
        RECT 20.235 -146.365 20.565 -146.035 ;
        RECT 20.235 -147.725 20.565 -147.395 ;
        RECT 20.235 -149.085 20.565 -148.755 ;
        RECT 20.235 -150.445 20.565 -150.115 ;
        RECT 20.235 -151.805 20.565 -151.475 ;
        RECT 20.235 -153.165 20.565 -152.835 ;
        RECT 20.235 -154.525 20.565 -154.195 ;
        RECT 20.235 -155.885 20.565 -155.555 ;
        RECT 20.235 -157.245 20.565 -156.915 ;
        RECT 20.235 -158.605 20.565 -158.275 ;
        RECT 20.235 -159.965 20.565 -159.635 ;
        RECT 20.235 -161.325 20.565 -160.995 ;
        RECT 20.235 -162.685 20.565 -162.355 ;
        RECT 20.235 -164.045 20.565 -163.715 ;
        RECT 20.235 -165.405 20.565 -165.075 ;
        RECT 20.235 -166.765 20.565 -166.435 ;
        RECT 20.235 -168.125 20.565 -167.795 ;
        RECT 20.235 -169.485 20.565 -169.155 ;
        RECT 20.235 -170.845 20.565 -170.515 ;
        RECT 20.235 -172.205 20.565 -171.875 ;
        RECT 20.235 -173.565 20.565 -173.235 ;
        RECT 20.235 -174.925 20.565 -174.595 ;
        RECT 20.235 -176.285 20.565 -175.955 ;
        RECT 20.235 -177.645 20.565 -177.315 ;
        RECT 20.235 -179.005 20.565 -178.675 ;
        RECT 20.235 -184.65 20.565 -183.52 ;
        RECT 20.24 -184.765 20.56 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 244.04 21.925 245.17 ;
        RECT 21.595 239.875 21.925 240.205 ;
        RECT 21.595 238.515 21.925 238.845 ;
        RECT 21.595 237.155 21.925 237.485 ;
        RECT 21.6 237.155 21.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 -0.845 21.925 -0.515 ;
        RECT 21.595 -2.205 21.925 -1.875 ;
        RECT 21.595 -3.565 21.925 -3.235 ;
        RECT 21.6 -3.565 21.92 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 21.595 -96.045 21.925 -95.715 ;
        RECT 21.595 -97.405 21.925 -97.075 ;
        RECT 21.595 -98.765 21.925 -98.435 ;
        RECT 21.595 -100.125 21.925 -99.795 ;
        RECT 21.595 -101.485 21.925 -101.155 ;
        RECT 21.595 -102.845 21.925 -102.515 ;
        RECT 21.595 -104.205 21.925 -103.875 ;
        RECT 21.595 -105.565 21.925 -105.235 ;
        RECT 21.595 -106.925 21.925 -106.595 ;
        RECT 21.595 -108.285 21.925 -107.955 ;
        RECT 21.595 -109.645 21.925 -109.315 ;
        RECT 21.595 -111.005 21.925 -110.675 ;
        RECT 21.595 -112.365 21.925 -112.035 ;
        RECT 21.595 -113.725 21.925 -113.395 ;
        RECT 21.595 -115.085 21.925 -114.755 ;
        RECT 21.595 -116.445 21.925 -116.115 ;
        RECT 21.595 -117.805 21.925 -117.475 ;
        RECT 21.595 -119.165 21.925 -118.835 ;
        RECT 21.595 -120.525 21.925 -120.195 ;
        RECT 21.595 -121.885 21.925 -121.555 ;
        RECT 21.595 -123.245 21.925 -122.915 ;
        RECT 21.595 -124.605 21.925 -124.275 ;
        RECT 21.595 -125.965 21.925 -125.635 ;
        RECT 21.595 -127.325 21.925 -126.995 ;
        RECT 21.595 -128.685 21.925 -128.355 ;
        RECT 21.595 -130.045 21.925 -129.715 ;
        RECT 21.595 -131.405 21.925 -131.075 ;
        RECT 21.595 -132.765 21.925 -132.435 ;
        RECT 21.595 -134.125 21.925 -133.795 ;
        RECT 21.595 -135.485 21.925 -135.155 ;
        RECT 21.595 -136.845 21.925 -136.515 ;
        RECT 21.595 -138.205 21.925 -137.875 ;
        RECT 21.595 -139.565 21.925 -139.235 ;
        RECT 21.595 -140.925 21.925 -140.595 ;
        RECT 21.595 -142.285 21.925 -141.955 ;
        RECT 21.595 -143.645 21.925 -143.315 ;
        RECT 21.595 -145.005 21.925 -144.675 ;
        RECT 21.595 -146.365 21.925 -146.035 ;
        RECT 21.595 -147.725 21.925 -147.395 ;
        RECT 21.595 -149.085 21.925 -148.755 ;
        RECT 21.595 -150.445 21.925 -150.115 ;
        RECT 21.595 -151.805 21.925 -151.475 ;
        RECT 21.595 -153.165 21.925 -152.835 ;
        RECT 21.595 -154.525 21.925 -154.195 ;
        RECT 21.595 -155.885 21.925 -155.555 ;
        RECT 21.595 -157.245 21.925 -156.915 ;
        RECT 21.595 -158.605 21.925 -158.275 ;
        RECT 21.595 -159.965 21.925 -159.635 ;
        RECT 21.595 -161.325 21.925 -160.995 ;
        RECT 21.595 -162.685 21.925 -162.355 ;
        RECT 21.595 -164.045 21.925 -163.715 ;
        RECT 21.595 -165.405 21.925 -165.075 ;
        RECT 21.595 -166.765 21.925 -166.435 ;
        RECT 21.595 -168.125 21.925 -167.795 ;
        RECT 21.595 -169.485 21.925 -169.155 ;
        RECT 21.595 -170.845 21.925 -170.515 ;
        RECT 21.595 -172.205 21.925 -171.875 ;
        RECT 21.595 -173.565 21.925 -173.235 ;
        RECT 21.595 -174.925 21.925 -174.595 ;
        RECT 21.595 -176.285 21.925 -175.955 ;
        RECT 21.595 -177.645 21.925 -177.315 ;
        RECT 21.595 -179.005 21.925 -178.675 ;
        RECT 21.595 -184.65 21.925 -183.52 ;
        RECT 21.6 -184.765 21.92 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 244.04 23.285 245.17 ;
        RECT 22.955 239.875 23.285 240.205 ;
        RECT 22.955 238.515 23.285 238.845 ;
        RECT 22.955 237.155 23.285 237.485 ;
        RECT 22.96 237.155 23.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 -0.845 23.285 -0.515 ;
        RECT 22.955 -2.205 23.285 -1.875 ;
        RECT 22.955 -3.565 23.285 -3.235 ;
        RECT 22.96 -3.565 23.28 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.955 -96.045 23.285 -95.715 ;
        RECT 22.955 -97.405 23.285 -97.075 ;
        RECT 22.955 -98.765 23.285 -98.435 ;
        RECT 22.955 -100.125 23.285 -99.795 ;
        RECT 22.955 -101.485 23.285 -101.155 ;
        RECT 22.955 -102.845 23.285 -102.515 ;
        RECT 22.955 -104.205 23.285 -103.875 ;
        RECT 22.955 -105.565 23.285 -105.235 ;
        RECT 22.955 -106.925 23.285 -106.595 ;
        RECT 22.955 -108.285 23.285 -107.955 ;
        RECT 22.955 -109.645 23.285 -109.315 ;
        RECT 22.955 -111.005 23.285 -110.675 ;
        RECT 22.955 -112.365 23.285 -112.035 ;
        RECT 22.955 -113.725 23.285 -113.395 ;
        RECT 22.955 -115.085 23.285 -114.755 ;
        RECT 22.955 -116.445 23.285 -116.115 ;
        RECT 22.955 -117.805 23.285 -117.475 ;
        RECT 22.955 -119.165 23.285 -118.835 ;
        RECT 22.955 -120.525 23.285 -120.195 ;
        RECT 22.955 -121.885 23.285 -121.555 ;
        RECT 22.955 -123.245 23.285 -122.915 ;
        RECT 22.955 -124.605 23.285 -124.275 ;
        RECT 22.955 -125.965 23.285 -125.635 ;
        RECT 22.955 -127.325 23.285 -126.995 ;
        RECT 22.955 -128.685 23.285 -128.355 ;
        RECT 22.955 -130.045 23.285 -129.715 ;
        RECT 22.955 -131.405 23.285 -131.075 ;
        RECT 22.955 -132.765 23.285 -132.435 ;
        RECT 22.955 -134.125 23.285 -133.795 ;
        RECT 22.955 -135.485 23.285 -135.155 ;
        RECT 22.955 -136.845 23.285 -136.515 ;
        RECT 22.955 -138.205 23.285 -137.875 ;
        RECT 22.955 -139.565 23.285 -139.235 ;
        RECT 22.955 -140.925 23.285 -140.595 ;
        RECT 22.955 -142.285 23.285 -141.955 ;
        RECT 22.955 -143.645 23.285 -143.315 ;
        RECT 22.955 -145.005 23.285 -144.675 ;
        RECT 22.955 -146.365 23.285 -146.035 ;
        RECT 22.955 -147.725 23.285 -147.395 ;
        RECT 22.955 -149.085 23.285 -148.755 ;
        RECT 22.955 -150.445 23.285 -150.115 ;
        RECT 22.955 -151.805 23.285 -151.475 ;
        RECT 22.955 -153.165 23.285 -152.835 ;
        RECT 22.955 -154.525 23.285 -154.195 ;
        RECT 22.955 -155.885 23.285 -155.555 ;
        RECT 22.955 -157.245 23.285 -156.915 ;
        RECT 22.955 -158.605 23.285 -158.275 ;
        RECT 22.955 -159.965 23.285 -159.635 ;
        RECT 22.955 -161.325 23.285 -160.995 ;
        RECT 22.955 -162.685 23.285 -162.355 ;
        RECT 22.955 -164.045 23.285 -163.715 ;
        RECT 22.955 -165.405 23.285 -165.075 ;
        RECT 22.955 -166.765 23.285 -166.435 ;
        RECT 22.955 -168.125 23.285 -167.795 ;
        RECT 22.955 -169.485 23.285 -169.155 ;
        RECT 22.955 -170.845 23.285 -170.515 ;
        RECT 22.955 -172.205 23.285 -171.875 ;
        RECT 22.955 -173.565 23.285 -173.235 ;
        RECT 22.955 -174.925 23.285 -174.595 ;
        RECT 22.955 -176.285 23.285 -175.955 ;
        RECT 22.955 -177.645 23.285 -177.315 ;
        RECT 22.955 -179.005 23.285 -178.675 ;
        RECT 22.955 -184.65 23.285 -183.52 ;
        RECT 22.96 -184.765 23.28 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 244.04 24.645 245.17 ;
        RECT 24.315 239.875 24.645 240.205 ;
        RECT 24.315 238.515 24.645 238.845 ;
        RECT 24.315 237.155 24.645 237.485 ;
        RECT 24.32 237.155 24.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.315 -98.765 24.645 -98.435 ;
        RECT 24.315 -100.125 24.645 -99.795 ;
        RECT 24.315 -101.485 24.645 -101.155 ;
        RECT 24.315 -102.845 24.645 -102.515 ;
        RECT 24.315 -104.205 24.645 -103.875 ;
        RECT 24.315 -105.565 24.645 -105.235 ;
        RECT 24.315 -106.925 24.645 -106.595 ;
        RECT 24.315 -108.285 24.645 -107.955 ;
        RECT 24.315 -109.645 24.645 -109.315 ;
        RECT 24.315 -111.005 24.645 -110.675 ;
        RECT 24.315 -112.365 24.645 -112.035 ;
        RECT 24.315 -113.725 24.645 -113.395 ;
        RECT 24.315 -115.085 24.645 -114.755 ;
        RECT 24.315 -116.445 24.645 -116.115 ;
        RECT 24.315 -117.805 24.645 -117.475 ;
        RECT 24.315 -119.165 24.645 -118.835 ;
        RECT 24.315 -120.525 24.645 -120.195 ;
        RECT 24.315 -121.885 24.645 -121.555 ;
        RECT 24.315 -123.245 24.645 -122.915 ;
        RECT 24.315 -124.605 24.645 -124.275 ;
        RECT 24.315 -125.965 24.645 -125.635 ;
        RECT 24.315 -127.325 24.645 -126.995 ;
        RECT 24.315 -128.685 24.645 -128.355 ;
        RECT 24.315 -130.045 24.645 -129.715 ;
        RECT 24.315 -131.405 24.645 -131.075 ;
        RECT 24.315 -132.765 24.645 -132.435 ;
        RECT 24.315 -134.125 24.645 -133.795 ;
        RECT 24.315 -135.485 24.645 -135.155 ;
        RECT 24.315 -136.845 24.645 -136.515 ;
        RECT 24.315 -138.205 24.645 -137.875 ;
        RECT 24.315 -139.565 24.645 -139.235 ;
        RECT 24.315 -140.925 24.645 -140.595 ;
        RECT 24.315 -142.285 24.645 -141.955 ;
        RECT 24.315 -143.645 24.645 -143.315 ;
        RECT 24.315 -145.005 24.645 -144.675 ;
        RECT 24.315 -146.365 24.645 -146.035 ;
        RECT 24.315 -147.725 24.645 -147.395 ;
        RECT 24.315 -149.085 24.645 -148.755 ;
        RECT 24.315 -150.445 24.645 -150.115 ;
        RECT 24.315 -151.805 24.645 -151.475 ;
        RECT 24.315 -153.165 24.645 -152.835 ;
        RECT 24.315 -154.525 24.645 -154.195 ;
        RECT 24.315 -155.885 24.645 -155.555 ;
        RECT 24.315 -157.245 24.645 -156.915 ;
        RECT 24.315 -158.605 24.645 -158.275 ;
        RECT 24.315 -159.965 24.645 -159.635 ;
        RECT 24.315 -161.325 24.645 -160.995 ;
        RECT 24.315 -162.685 24.645 -162.355 ;
        RECT 24.315 -164.045 24.645 -163.715 ;
        RECT 24.315 -165.405 24.645 -165.075 ;
        RECT 24.315 -166.765 24.645 -166.435 ;
        RECT 24.315 -168.125 24.645 -167.795 ;
        RECT 24.315 -169.485 24.645 -169.155 ;
        RECT 24.315 -170.845 24.645 -170.515 ;
        RECT 24.315 -172.205 24.645 -171.875 ;
        RECT 24.315 -173.565 24.645 -173.235 ;
        RECT 24.315 -174.925 24.645 -174.595 ;
        RECT 24.315 -176.285 24.645 -175.955 ;
        RECT 24.315 -177.645 24.645 -177.315 ;
        RECT 24.315 -179.005 24.645 -178.675 ;
        RECT 24.315 -184.65 24.645 -183.52 ;
        RECT 24.32 -184.765 24.64 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.46 -98.075 24.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.675 244.04 26.005 245.17 ;
        RECT 25.675 239.875 26.005 240.205 ;
        RECT 25.675 238.515 26.005 238.845 ;
        RECT 25.675 237.155 26.005 237.485 ;
        RECT 25.68 237.155 26 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 244.04 27.365 245.17 ;
        RECT 27.035 239.875 27.365 240.205 ;
        RECT 27.035 238.515 27.365 238.845 ;
        RECT 27.035 237.155 27.365 237.485 ;
        RECT 27.04 237.155 27.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.035 -0.845 27.365 -0.515 ;
        RECT 27.035 -2.205 27.365 -1.875 ;
        RECT 27.035 -3.565 27.365 -3.235 ;
        RECT 27.04 -3.565 27.36 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 244.04 28.725 245.17 ;
        RECT 28.395 239.875 28.725 240.205 ;
        RECT 28.395 238.515 28.725 238.845 ;
        RECT 28.395 237.155 28.725 237.485 ;
        RECT 28.4 237.155 28.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 -0.845 28.725 -0.515 ;
        RECT 28.395 -2.205 28.725 -1.875 ;
        RECT 28.395 -3.565 28.725 -3.235 ;
        RECT 28.4 -3.565 28.72 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 28.395 -96.045 28.725 -95.715 ;
        RECT 28.395 -97.405 28.725 -97.075 ;
        RECT 28.395 -98.765 28.725 -98.435 ;
        RECT 28.395 -100.125 28.725 -99.795 ;
        RECT 28.395 -101.485 28.725 -101.155 ;
        RECT 28.395 -102.845 28.725 -102.515 ;
        RECT 28.395 -104.205 28.725 -103.875 ;
        RECT 28.395 -105.565 28.725 -105.235 ;
        RECT 28.395 -106.925 28.725 -106.595 ;
        RECT 28.395 -108.285 28.725 -107.955 ;
        RECT 28.395 -109.645 28.725 -109.315 ;
        RECT 28.395 -111.005 28.725 -110.675 ;
        RECT 28.395 -112.365 28.725 -112.035 ;
        RECT 28.395 -113.725 28.725 -113.395 ;
        RECT 28.395 -115.085 28.725 -114.755 ;
        RECT 28.395 -116.445 28.725 -116.115 ;
        RECT 28.395 -117.805 28.725 -117.475 ;
        RECT 28.395 -119.165 28.725 -118.835 ;
        RECT 28.395 -120.525 28.725 -120.195 ;
        RECT 28.395 -121.885 28.725 -121.555 ;
        RECT 28.395 -123.245 28.725 -122.915 ;
        RECT 28.395 -124.605 28.725 -124.275 ;
        RECT 28.395 -125.965 28.725 -125.635 ;
        RECT 28.395 -127.325 28.725 -126.995 ;
        RECT 28.395 -128.685 28.725 -128.355 ;
        RECT 28.395 -130.045 28.725 -129.715 ;
        RECT 28.395 -131.405 28.725 -131.075 ;
        RECT 28.395 -132.765 28.725 -132.435 ;
        RECT 28.395 -134.125 28.725 -133.795 ;
        RECT 28.395 -135.485 28.725 -135.155 ;
        RECT 28.395 -136.845 28.725 -136.515 ;
        RECT 28.395 -138.205 28.725 -137.875 ;
        RECT 28.395 -139.565 28.725 -139.235 ;
        RECT 28.395 -140.925 28.725 -140.595 ;
        RECT 28.395 -142.285 28.725 -141.955 ;
        RECT 28.395 -143.645 28.725 -143.315 ;
        RECT 28.395 -145.005 28.725 -144.675 ;
        RECT 28.395 -146.365 28.725 -146.035 ;
        RECT 28.395 -147.725 28.725 -147.395 ;
        RECT 28.395 -149.085 28.725 -148.755 ;
        RECT 28.395 -150.445 28.725 -150.115 ;
        RECT 28.395 -151.805 28.725 -151.475 ;
        RECT 28.395 -153.165 28.725 -152.835 ;
        RECT 28.395 -154.525 28.725 -154.195 ;
        RECT 28.395 -155.885 28.725 -155.555 ;
        RECT 28.395 -157.245 28.725 -156.915 ;
        RECT 28.395 -158.605 28.725 -158.275 ;
        RECT 28.395 -159.965 28.725 -159.635 ;
        RECT 28.395 -161.325 28.725 -160.995 ;
        RECT 28.395 -162.685 28.725 -162.355 ;
        RECT 28.395 -164.045 28.725 -163.715 ;
        RECT 28.395 -165.405 28.725 -165.075 ;
        RECT 28.395 -166.765 28.725 -166.435 ;
        RECT 28.395 -168.125 28.725 -167.795 ;
        RECT 28.395 -169.485 28.725 -169.155 ;
        RECT 28.395 -170.845 28.725 -170.515 ;
        RECT 28.395 -172.205 28.725 -171.875 ;
        RECT 28.395 -173.565 28.725 -173.235 ;
        RECT 28.395 -174.925 28.725 -174.595 ;
        RECT 28.395 -176.285 28.725 -175.955 ;
        RECT 28.395 -177.645 28.725 -177.315 ;
        RECT 28.395 -179.005 28.725 -178.675 ;
        RECT 28.395 -184.65 28.725 -183.52 ;
        RECT 28.4 -184.765 28.72 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 244.04 30.085 245.17 ;
        RECT 29.755 239.875 30.085 240.205 ;
        RECT 29.755 238.515 30.085 238.845 ;
        RECT 29.755 237.155 30.085 237.485 ;
        RECT 29.76 237.155 30.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 -0.845 30.085 -0.515 ;
        RECT 29.755 -2.205 30.085 -1.875 ;
        RECT 29.755 -3.565 30.085 -3.235 ;
        RECT 29.76 -3.565 30.08 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.755 -96.045 30.085 -95.715 ;
        RECT 29.755 -97.405 30.085 -97.075 ;
        RECT 29.755 -98.765 30.085 -98.435 ;
        RECT 29.755 -100.125 30.085 -99.795 ;
        RECT 29.755 -101.485 30.085 -101.155 ;
        RECT 29.755 -102.845 30.085 -102.515 ;
        RECT 29.755 -104.205 30.085 -103.875 ;
        RECT 29.755 -105.565 30.085 -105.235 ;
        RECT 29.755 -106.925 30.085 -106.595 ;
        RECT 29.755 -108.285 30.085 -107.955 ;
        RECT 29.755 -109.645 30.085 -109.315 ;
        RECT 29.755 -111.005 30.085 -110.675 ;
        RECT 29.755 -112.365 30.085 -112.035 ;
        RECT 29.755 -113.725 30.085 -113.395 ;
        RECT 29.755 -115.085 30.085 -114.755 ;
        RECT 29.755 -116.445 30.085 -116.115 ;
        RECT 29.755 -117.805 30.085 -117.475 ;
        RECT 29.755 -119.165 30.085 -118.835 ;
        RECT 29.755 -120.525 30.085 -120.195 ;
        RECT 29.755 -121.885 30.085 -121.555 ;
        RECT 29.755 -123.245 30.085 -122.915 ;
        RECT 29.755 -124.605 30.085 -124.275 ;
        RECT 29.755 -125.965 30.085 -125.635 ;
        RECT 29.755 -127.325 30.085 -126.995 ;
        RECT 29.755 -128.685 30.085 -128.355 ;
        RECT 29.755 -130.045 30.085 -129.715 ;
        RECT 29.755 -131.405 30.085 -131.075 ;
        RECT 29.755 -132.765 30.085 -132.435 ;
        RECT 29.755 -134.125 30.085 -133.795 ;
        RECT 29.755 -135.485 30.085 -135.155 ;
        RECT 29.755 -136.845 30.085 -136.515 ;
        RECT 29.755 -138.205 30.085 -137.875 ;
        RECT 29.755 -139.565 30.085 -139.235 ;
        RECT 29.755 -140.925 30.085 -140.595 ;
        RECT 29.755 -142.285 30.085 -141.955 ;
        RECT 29.755 -143.645 30.085 -143.315 ;
        RECT 29.755 -145.005 30.085 -144.675 ;
        RECT 29.755 -146.365 30.085 -146.035 ;
        RECT 29.755 -147.725 30.085 -147.395 ;
        RECT 29.755 -149.085 30.085 -148.755 ;
        RECT 29.755 -150.445 30.085 -150.115 ;
        RECT 29.755 -151.805 30.085 -151.475 ;
        RECT 29.755 -153.165 30.085 -152.835 ;
        RECT 29.755 -154.525 30.085 -154.195 ;
        RECT 29.755 -155.885 30.085 -155.555 ;
        RECT 29.755 -157.245 30.085 -156.915 ;
        RECT 29.755 -158.605 30.085 -158.275 ;
        RECT 29.755 -159.965 30.085 -159.635 ;
        RECT 29.755 -161.325 30.085 -160.995 ;
        RECT 29.755 -162.685 30.085 -162.355 ;
        RECT 29.755 -164.045 30.085 -163.715 ;
        RECT 29.755 -165.405 30.085 -165.075 ;
        RECT 29.755 -166.765 30.085 -166.435 ;
        RECT 29.755 -168.125 30.085 -167.795 ;
        RECT 29.755 -169.485 30.085 -169.155 ;
        RECT 29.755 -170.845 30.085 -170.515 ;
        RECT 29.755 -172.205 30.085 -171.875 ;
        RECT 29.755 -173.565 30.085 -173.235 ;
        RECT 29.755 -174.925 30.085 -174.595 ;
        RECT 29.755 -176.285 30.085 -175.955 ;
        RECT 29.755 -177.645 30.085 -177.315 ;
        RECT 29.755 -179.005 30.085 -178.675 ;
        RECT 29.755 -184.65 30.085 -183.52 ;
        RECT 29.76 -184.765 30.08 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 244.04 31.445 245.17 ;
        RECT 31.115 239.875 31.445 240.205 ;
        RECT 31.115 238.515 31.445 238.845 ;
        RECT 31.115 237.155 31.445 237.485 ;
        RECT 31.12 237.155 31.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 -0.845 31.445 -0.515 ;
        RECT 31.115 -2.205 31.445 -1.875 ;
        RECT 31.115 -3.565 31.445 -3.235 ;
        RECT 31.12 -3.565 31.44 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.115 -96.045 31.445 -95.715 ;
        RECT 31.115 -97.405 31.445 -97.075 ;
        RECT 31.115 -98.765 31.445 -98.435 ;
        RECT 31.115 -100.125 31.445 -99.795 ;
        RECT 31.115 -101.485 31.445 -101.155 ;
        RECT 31.115 -102.845 31.445 -102.515 ;
        RECT 31.115 -104.205 31.445 -103.875 ;
        RECT 31.115 -105.565 31.445 -105.235 ;
        RECT 31.115 -106.925 31.445 -106.595 ;
        RECT 31.115 -108.285 31.445 -107.955 ;
        RECT 31.115 -109.645 31.445 -109.315 ;
        RECT 31.115 -111.005 31.445 -110.675 ;
        RECT 31.115 -112.365 31.445 -112.035 ;
        RECT 31.115 -113.725 31.445 -113.395 ;
        RECT 31.115 -115.085 31.445 -114.755 ;
        RECT 31.115 -116.445 31.445 -116.115 ;
        RECT 31.115 -117.805 31.445 -117.475 ;
        RECT 31.115 -119.165 31.445 -118.835 ;
        RECT 31.115 -120.525 31.445 -120.195 ;
        RECT 31.115 -121.885 31.445 -121.555 ;
        RECT 31.115 -123.245 31.445 -122.915 ;
        RECT 31.115 -124.605 31.445 -124.275 ;
        RECT 31.115 -125.965 31.445 -125.635 ;
        RECT 31.115 -127.325 31.445 -126.995 ;
        RECT 31.115 -128.685 31.445 -128.355 ;
        RECT 31.115 -130.045 31.445 -129.715 ;
        RECT 31.115 -131.405 31.445 -131.075 ;
        RECT 31.115 -132.765 31.445 -132.435 ;
        RECT 31.115 -134.125 31.445 -133.795 ;
        RECT 31.115 -135.485 31.445 -135.155 ;
        RECT 31.115 -136.845 31.445 -136.515 ;
        RECT 31.115 -138.205 31.445 -137.875 ;
        RECT 31.115 -139.565 31.445 -139.235 ;
        RECT 31.115 -140.925 31.445 -140.595 ;
        RECT 31.115 -142.285 31.445 -141.955 ;
        RECT 31.115 -143.645 31.445 -143.315 ;
        RECT 31.115 -145.005 31.445 -144.675 ;
        RECT 31.115 -146.365 31.445 -146.035 ;
        RECT 31.115 -147.725 31.445 -147.395 ;
        RECT 31.115 -149.085 31.445 -148.755 ;
        RECT 31.115 -150.445 31.445 -150.115 ;
        RECT 31.115 -151.805 31.445 -151.475 ;
        RECT 31.115 -153.165 31.445 -152.835 ;
        RECT 31.115 -154.525 31.445 -154.195 ;
        RECT 31.115 -155.885 31.445 -155.555 ;
        RECT 31.115 -157.245 31.445 -156.915 ;
        RECT 31.115 -158.605 31.445 -158.275 ;
        RECT 31.115 -159.965 31.445 -159.635 ;
        RECT 31.115 -161.325 31.445 -160.995 ;
        RECT 31.115 -162.685 31.445 -162.355 ;
        RECT 31.115 -164.045 31.445 -163.715 ;
        RECT 31.115 -165.405 31.445 -165.075 ;
        RECT 31.115 -166.765 31.445 -166.435 ;
        RECT 31.115 -168.125 31.445 -167.795 ;
        RECT 31.115 -169.485 31.445 -169.155 ;
        RECT 31.115 -170.845 31.445 -170.515 ;
        RECT 31.115 -172.205 31.445 -171.875 ;
        RECT 31.115 -173.565 31.445 -173.235 ;
        RECT 31.115 -174.925 31.445 -174.595 ;
        RECT 31.115 -176.285 31.445 -175.955 ;
        RECT 31.115 -177.645 31.445 -177.315 ;
        RECT 31.115 -179.005 31.445 -178.675 ;
        RECT 31.115 -184.65 31.445 -183.52 ;
        RECT 31.12 -184.765 31.44 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 244.04 32.805 245.17 ;
        RECT 32.475 239.875 32.805 240.205 ;
        RECT 32.475 238.515 32.805 238.845 ;
        RECT 32.475 237.155 32.805 237.485 ;
        RECT 32.48 237.155 32.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 -0.845 32.805 -0.515 ;
        RECT 32.475 -2.205 32.805 -1.875 ;
        RECT 32.475 -3.565 32.805 -3.235 ;
        RECT 32.48 -3.565 32.8 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 32.475 -96.045 32.805 -95.715 ;
        RECT 32.475 -97.405 32.805 -97.075 ;
        RECT 32.475 -98.765 32.805 -98.435 ;
        RECT 32.475 -100.125 32.805 -99.795 ;
        RECT 32.475 -101.485 32.805 -101.155 ;
        RECT 32.475 -102.845 32.805 -102.515 ;
        RECT 32.475 -104.205 32.805 -103.875 ;
        RECT 32.475 -105.565 32.805 -105.235 ;
        RECT 32.475 -106.925 32.805 -106.595 ;
        RECT 32.475 -108.285 32.805 -107.955 ;
        RECT 32.475 -109.645 32.805 -109.315 ;
        RECT 32.475 -111.005 32.805 -110.675 ;
        RECT 32.475 -112.365 32.805 -112.035 ;
        RECT 32.475 -113.725 32.805 -113.395 ;
        RECT 32.475 -115.085 32.805 -114.755 ;
        RECT 32.475 -116.445 32.805 -116.115 ;
        RECT 32.475 -117.805 32.805 -117.475 ;
        RECT 32.475 -119.165 32.805 -118.835 ;
        RECT 32.475 -120.525 32.805 -120.195 ;
        RECT 32.475 -121.885 32.805 -121.555 ;
        RECT 32.475 -123.245 32.805 -122.915 ;
        RECT 32.475 -124.605 32.805 -124.275 ;
        RECT 32.475 -125.965 32.805 -125.635 ;
        RECT 32.475 -127.325 32.805 -126.995 ;
        RECT 32.475 -128.685 32.805 -128.355 ;
        RECT 32.475 -130.045 32.805 -129.715 ;
        RECT 32.475 -131.405 32.805 -131.075 ;
        RECT 32.475 -132.765 32.805 -132.435 ;
        RECT 32.475 -134.125 32.805 -133.795 ;
        RECT 32.475 -135.485 32.805 -135.155 ;
        RECT 32.475 -136.845 32.805 -136.515 ;
        RECT 32.475 -138.205 32.805 -137.875 ;
        RECT 32.475 -139.565 32.805 -139.235 ;
        RECT 32.475 -140.925 32.805 -140.595 ;
        RECT 32.475 -142.285 32.805 -141.955 ;
        RECT 32.475 -143.645 32.805 -143.315 ;
        RECT 32.475 -145.005 32.805 -144.675 ;
        RECT 32.475 -146.365 32.805 -146.035 ;
        RECT 32.475 -147.725 32.805 -147.395 ;
        RECT 32.475 -149.085 32.805 -148.755 ;
        RECT 32.475 -150.445 32.805 -150.115 ;
        RECT 32.475 -151.805 32.805 -151.475 ;
        RECT 32.475 -153.165 32.805 -152.835 ;
        RECT 32.475 -154.525 32.805 -154.195 ;
        RECT 32.475 -155.885 32.805 -155.555 ;
        RECT 32.475 -157.245 32.805 -156.915 ;
        RECT 32.475 -158.605 32.805 -158.275 ;
        RECT 32.475 -159.965 32.805 -159.635 ;
        RECT 32.475 -161.325 32.805 -160.995 ;
        RECT 32.475 -162.685 32.805 -162.355 ;
        RECT 32.475 -164.045 32.805 -163.715 ;
        RECT 32.475 -165.405 32.805 -165.075 ;
        RECT 32.475 -166.765 32.805 -166.435 ;
        RECT 32.475 -168.125 32.805 -167.795 ;
        RECT 32.475 -169.485 32.805 -169.155 ;
        RECT 32.475 -170.845 32.805 -170.515 ;
        RECT 32.475 -172.205 32.805 -171.875 ;
        RECT 32.475 -173.565 32.805 -173.235 ;
        RECT 32.475 -174.925 32.805 -174.595 ;
        RECT 32.475 -176.285 32.805 -175.955 ;
        RECT 32.475 -177.645 32.805 -177.315 ;
        RECT 32.475 -179.005 32.805 -178.675 ;
        RECT 32.475 -184.65 32.805 -183.52 ;
        RECT 32.48 -184.765 32.8 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 244.04 34.165 245.17 ;
        RECT 33.835 239.875 34.165 240.205 ;
        RECT 33.835 238.515 34.165 238.845 ;
        RECT 33.835 237.155 34.165 237.485 ;
        RECT 33.84 237.155 34.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 -0.845 34.165 -0.515 ;
        RECT 33.835 -2.205 34.165 -1.875 ;
        RECT 33.835 -3.565 34.165 -3.235 ;
        RECT 33.84 -3.565 34.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.835 -96.045 34.165 -95.715 ;
        RECT 33.835 -97.405 34.165 -97.075 ;
        RECT 33.835 -98.765 34.165 -98.435 ;
        RECT 33.835 -100.125 34.165 -99.795 ;
        RECT 33.835 -101.485 34.165 -101.155 ;
        RECT 33.835 -102.845 34.165 -102.515 ;
        RECT 33.835 -104.205 34.165 -103.875 ;
        RECT 33.835 -105.565 34.165 -105.235 ;
        RECT 33.835 -106.925 34.165 -106.595 ;
        RECT 33.835 -108.285 34.165 -107.955 ;
        RECT 33.835 -109.645 34.165 -109.315 ;
        RECT 33.835 -111.005 34.165 -110.675 ;
        RECT 33.835 -112.365 34.165 -112.035 ;
        RECT 33.835 -113.725 34.165 -113.395 ;
        RECT 33.835 -115.085 34.165 -114.755 ;
        RECT 33.835 -116.445 34.165 -116.115 ;
        RECT 33.835 -117.805 34.165 -117.475 ;
        RECT 33.835 -119.165 34.165 -118.835 ;
        RECT 33.835 -120.525 34.165 -120.195 ;
        RECT 33.835 -121.885 34.165 -121.555 ;
        RECT 33.835 -123.245 34.165 -122.915 ;
        RECT 33.835 -124.605 34.165 -124.275 ;
        RECT 33.835 -125.965 34.165 -125.635 ;
        RECT 33.835 -127.325 34.165 -126.995 ;
        RECT 33.835 -128.685 34.165 -128.355 ;
        RECT 33.835 -130.045 34.165 -129.715 ;
        RECT 33.835 -131.405 34.165 -131.075 ;
        RECT 33.835 -132.765 34.165 -132.435 ;
        RECT 33.835 -134.125 34.165 -133.795 ;
        RECT 33.835 -135.485 34.165 -135.155 ;
        RECT 33.835 -136.845 34.165 -136.515 ;
        RECT 33.835 -138.205 34.165 -137.875 ;
        RECT 33.835 -139.565 34.165 -139.235 ;
        RECT 33.835 -140.925 34.165 -140.595 ;
        RECT 33.835 -142.285 34.165 -141.955 ;
        RECT 33.835 -143.645 34.165 -143.315 ;
        RECT 33.835 -145.005 34.165 -144.675 ;
        RECT 33.835 -146.365 34.165 -146.035 ;
        RECT 33.835 -147.725 34.165 -147.395 ;
        RECT 33.835 -149.085 34.165 -148.755 ;
        RECT 33.835 -150.445 34.165 -150.115 ;
        RECT 33.835 -151.805 34.165 -151.475 ;
        RECT 33.835 -153.165 34.165 -152.835 ;
        RECT 33.835 -154.525 34.165 -154.195 ;
        RECT 33.835 -155.885 34.165 -155.555 ;
        RECT 33.835 -157.245 34.165 -156.915 ;
        RECT 33.835 -158.605 34.165 -158.275 ;
        RECT 33.835 -159.965 34.165 -159.635 ;
        RECT 33.835 -161.325 34.165 -160.995 ;
        RECT 33.835 -162.685 34.165 -162.355 ;
        RECT 33.835 -164.045 34.165 -163.715 ;
        RECT 33.835 -165.405 34.165 -165.075 ;
        RECT 33.835 -166.765 34.165 -166.435 ;
        RECT 33.835 -168.125 34.165 -167.795 ;
        RECT 33.835 -169.485 34.165 -169.155 ;
        RECT 33.835 -170.845 34.165 -170.515 ;
        RECT 33.835 -172.205 34.165 -171.875 ;
        RECT 33.835 -173.565 34.165 -173.235 ;
        RECT 33.835 -174.925 34.165 -174.595 ;
        RECT 33.835 -176.285 34.165 -175.955 ;
        RECT 33.835 -177.645 34.165 -177.315 ;
        RECT 33.835 -179.005 34.165 -178.675 ;
        RECT 33.835 -184.65 34.165 -183.52 ;
        RECT 33.84 -184.765 34.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 244.04 35.525 245.17 ;
        RECT 35.195 239.875 35.525 240.205 ;
        RECT 35.195 238.515 35.525 238.845 ;
        RECT 35.195 237.155 35.525 237.485 ;
        RECT 35.2 237.155 35.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.195 -151.805 35.525 -151.475 ;
        RECT 35.195 -153.165 35.525 -152.835 ;
        RECT 35.195 -154.525 35.525 -154.195 ;
        RECT 35.195 -155.885 35.525 -155.555 ;
        RECT 35.195 -157.245 35.525 -156.915 ;
        RECT 35.195 -158.605 35.525 -158.275 ;
        RECT 35.195 -159.965 35.525 -159.635 ;
        RECT 35.195 -161.325 35.525 -160.995 ;
        RECT 35.195 -162.685 35.525 -162.355 ;
        RECT 35.195 -164.045 35.525 -163.715 ;
        RECT 35.195 -165.405 35.525 -165.075 ;
        RECT 35.195 -166.765 35.525 -166.435 ;
        RECT 35.195 -168.125 35.525 -167.795 ;
        RECT 35.195 -169.485 35.525 -169.155 ;
        RECT 35.195 -170.845 35.525 -170.515 ;
        RECT 35.195 -172.205 35.525 -171.875 ;
        RECT 35.195 -173.565 35.525 -173.235 ;
        RECT 35.195 -174.925 35.525 -174.595 ;
        RECT 35.195 -176.285 35.525 -175.955 ;
        RECT 35.195 -177.645 35.525 -177.315 ;
        RECT 35.195 -179.005 35.525 -178.675 ;
        RECT 35.195 -184.65 35.525 -183.52 ;
        RECT 35.2 -184.765 35.52 -98.435 ;
        RECT 35.195 -98.765 35.525 -98.435 ;
        RECT 35.195 -100.125 35.525 -99.795 ;
        RECT 35.195 -101.485 35.525 -101.155 ;
        RECT 35.195 -102.845 35.525 -102.515 ;
        RECT 35.195 -104.205 35.525 -103.875 ;
        RECT 35.195 -105.565 35.525 -105.235 ;
        RECT 35.195 -106.925 35.525 -106.595 ;
        RECT 35.195 -108.285 35.525 -107.955 ;
        RECT 35.195 -109.645 35.525 -109.315 ;
        RECT 35.195 -111.005 35.525 -110.675 ;
        RECT 35.195 -112.365 35.525 -112.035 ;
        RECT 35.195 -113.725 35.525 -113.395 ;
        RECT 35.195 -115.085 35.525 -114.755 ;
        RECT 35.195 -116.445 35.525 -116.115 ;
        RECT 35.195 -117.805 35.525 -117.475 ;
        RECT 35.195 -119.165 35.525 -118.835 ;
        RECT 35.195 -120.525 35.525 -120.195 ;
        RECT 35.195 -121.885 35.525 -121.555 ;
        RECT 35.195 -123.245 35.525 -122.915 ;
        RECT 35.195 -124.605 35.525 -124.275 ;
        RECT 35.195 -125.965 35.525 -125.635 ;
        RECT 35.195 -127.325 35.525 -126.995 ;
        RECT 35.195 -128.685 35.525 -128.355 ;
        RECT 35.195 -130.045 35.525 -129.715 ;
        RECT 35.195 -131.405 35.525 -131.075 ;
        RECT 35.195 -132.765 35.525 -132.435 ;
        RECT 35.195 -134.125 35.525 -133.795 ;
        RECT 35.195 -135.485 35.525 -135.155 ;
        RECT 35.195 -136.845 35.525 -136.515 ;
        RECT 35.195 -138.205 35.525 -137.875 ;
        RECT 35.195 -139.565 35.525 -139.235 ;
        RECT 35.195 -140.925 35.525 -140.595 ;
        RECT 35.195 -142.285 35.525 -141.955 ;
        RECT 35.195 -143.645 35.525 -143.315 ;
        RECT 35.195 -145.005 35.525 -144.675 ;
        RECT 35.195 -146.365 35.525 -146.035 ;
        RECT 35.195 -147.725 35.525 -147.395 ;
        RECT 35.195 -149.085 35.525 -148.755 ;
        RECT 35.195 -150.445 35.525 -150.115 ;
    END
    PORT
      LAYER met3 ;
        RECT -1.525 244.04 -1.195 245.17 ;
        RECT -1.525 239.875 -1.195 240.205 ;
        RECT -1.525 238.515 -1.195 238.845 ;
        RECT -1.525 237.155 -1.195 237.485 ;
        RECT -1.525 235.17 -1.195 235.5 ;
        RECT -1.525 232.995 -1.195 233.325 ;
        RECT -1.525 231.415 -1.195 231.745 ;
        RECT -1.525 230.565 -1.195 230.895 ;
        RECT -1.525 228.255 -1.195 228.585 ;
        RECT -1.525 227.405 -1.195 227.735 ;
        RECT -1.525 225.095 -1.195 225.425 ;
        RECT -1.525 224.245 -1.195 224.575 ;
        RECT -1.525 221.935 -1.195 222.265 ;
        RECT -1.525 221.085 -1.195 221.415 ;
        RECT -1.525 218.775 -1.195 219.105 ;
        RECT -1.525 217.195 -1.195 217.525 ;
        RECT -1.525 216.345 -1.195 216.675 ;
        RECT -1.525 214.035 -1.195 214.365 ;
        RECT -1.525 213.185 -1.195 213.515 ;
        RECT -1.525 210.875 -1.195 211.205 ;
        RECT -1.525 210.025 -1.195 210.355 ;
        RECT -1.525 207.715 -1.195 208.045 ;
        RECT -1.525 206.865 -1.195 207.195 ;
        RECT -1.525 204.555 -1.195 204.885 ;
        RECT -1.525 202.975 -1.195 203.305 ;
        RECT -1.525 202.125 -1.195 202.455 ;
        RECT -1.525 199.815 -1.195 200.145 ;
        RECT -1.525 198.965 -1.195 199.295 ;
        RECT -1.525 196.655 -1.195 196.985 ;
        RECT -1.525 195.805 -1.195 196.135 ;
        RECT -1.525 193.495 -1.195 193.825 ;
        RECT -1.525 192.645 -1.195 192.975 ;
        RECT -1.525 190.335 -1.195 190.665 ;
        RECT -1.525 188.755 -1.195 189.085 ;
        RECT -1.525 187.905 -1.195 188.235 ;
        RECT -1.525 185.595 -1.195 185.925 ;
        RECT -1.525 184.745 -1.195 185.075 ;
        RECT -1.525 182.435 -1.195 182.765 ;
        RECT -1.525 181.585 -1.195 181.915 ;
        RECT -1.525 179.275 -1.195 179.605 ;
        RECT -1.525 178.425 -1.195 178.755 ;
        RECT -1.525 176.115 -1.195 176.445 ;
        RECT -1.525 174.535 -1.195 174.865 ;
        RECT -1.525 173.685 -1.195 174.015 ;
        RECT -1.525 171.375 -1.195 171.705 ;
        RECT -1.525 170.525 -1.195 170.855 ;
        RECT -1.525 168.215 -1.195 168.545 ;
        RECT -1.525 167.365 -1.195 167.695 ;
        RECT -1.525 165.055 -1.195 165.385 ;
        RECT -1.525 164.205 -1.195 164.535 ;
        RECT -1.525 161.895 -1.195 162.225 ;
        RECT -1.525 160.315 -1.195 160.645 ;
        RECT -1.525 159.465 -1.195 159.795 ;
        RECT -1.525 157.155 -1.195 157.485 ;
        RECT -1.525 156.305 -1.195 156.635 ;
        RECT -1.525 153.995 -1.195 154.325 ;
        RECT -1.525 153.145 -1.195 153.475 ;
        RECT -1.525 150.835 -1.195 151.165 ;
        RECT -1.525 149.985 -1.195 150.315 ;
        RECT -1.525 147.675 -1.195 148.005 ;
        RECT -1.525 146.095 -1.195 146.425 ;
        RECT -1.525 145.245 -1.195 145.575 ;
        RECT -1.525 142.935 -1.195 143.265 ;
        RECT -1.525 142.085 -1.195 142.415 ;
        RECT -1.525 139.775 -1.195 140.105 ;
        RECT -1.525 138.925 -1.195 139.255 ;
        RECT -1.525 136.615 -1.195 136.945 ;
        RECT -1.525 135.765 -1.195 136.095 ;
        RECT -1.525 133.455 -1.195 133.785 ;
        RECT -1.525 131.875 -1.195 132.205 ;
        RECT -1.525 131.025 -1.195 131.355 ;
        RECT -1.525 128.715 -1.195 129.045 ;
        RECT -1.525 127.865 -1.195 128.195 ;
        RECT -1.525 125.555 -1.195 125.885 ;
        RECT -1.525 124.705 -1.195 125.035 ;
        RECT -1.525 122.395 -1.195 122.725 ;
        RECT -1.525 121.545 -1.195 121.875 ;
        RECT -1.525 119.235 -1.195 119.565 ;
        RECT -1.525 117.655 -1.195 117.985 ;
        RECT -1.525 116.805 -1.195 117.135 ;
        RECT -1.525 114.495 -1.195 114.825 ;
        RECT -1.525 113.645 -1.195 113.975 ;
        RECT -1.525 111.335 -1.195 111.665 ;
        RECT -1.525 110.485 -1.195 110.815 ;
        RECT -1.525 108.175 -1.195 108.505 ;
        RECT -1.525 107.325 -1.195 107.655 ;
        RECT -1.525 105.015 -1.195 105.345 ;
        RECT -1.525 103.435 -1.195 103.765 ;
        RECT -1.525 102.585 -1.195 102.915 ;
        RECT -1.525 100.275 -1.195 100.605 ;
        RECT -1.525 99.425 -1.195 99.755 ;
        RECT -1.525 97.115 -1.195 97.445 ;
        RECT -1.525 96.265 -1.195 96.595 ;
        RECT -1.525 93.955 -1.195 94.285 ;
        RECT -1.525 93.105 -1.195 93.435 ;
        RECT -1.525 90.795 -1.195 91.125 ;
        RECT -1.525 89.215 -1.195 89.545 ;
        RECT -1.525 88.365 -1.195 88.695 ;
        RECT -1.525 86.055 -1.195 86.385 ;
        RECT -1.525 85.205 -1.195 85.535 ;
        RECT -1.525 82.895 -1.195 83.225 ;
        RECT -1.525 82.045 -1.195 82.375 ;
        RECT -1.525 79.735 -1.195 80.065 ;
        RECT -1.525 78.885 -1.195 79.215 ;
        RECT -1.525 76.575 -1.195 76.905 ;
        RECT -1.525 74.995 -1.195 75.325 ;
        RECT -1.525 74.145 -1.195 74.475 ;
        RECT -1.525 71.835 -1.195 72.165 ;
        RECT -1.525 70.985 -1.195 71.315 ;
        RECT -1.525 68.675 -1.195 69.005 ;
        RECT -1.525 67.825 -1.195 68.155 ;
        RECT -1.525 65.515 -1.195 65.845 ;
        RECT -1.525 64.665 -1.195 64.995 ;
        RECT -1.525 62.355 -1.195 62.685 ;
        RECT -1.525 60.775 -1.195 61.105 ;
        RECT -1.525 59.925 -1.195 60.255 ;
        RECT -1.525 57.615 -1.195 57.945 ;
        RECT -1.525 56.765 -1.195 57.095 ;
        RECT -1.525 54.455 -1.195 54.785 ;
        RECT -1.525 53.605 -1.195 53.935 ;
        RECT -1.525 51.295 -1.195 51.625 ;
        RECT -1.525 50.445 -1.195 50.775 ;
        RECT -1.525 48.135 -1.195 48.465 ;
        RECT -1.525 46.555 -1.195 46.885 ;
        RECT -1.525 45.705 -1.195 46.035 ;
        RECT -1.525 43.395 -1.195 43.725 ;
        RECT -1.525 42.545 -1.195 42.875 ;
        RECT -1.525 40.235 -1.195 40.565 ;
        RECT -1.525 39.385 -1.195 39.715 ;
        RECT -1.525 37.075 -1.195 37.405 ;
        RECT -1.525 36.225 -1.195 36.555 ;
        RECT -1.525 33.915 -1.195 34.245 ;
        RECT -1.525 32.335 -1.195 32.665 ;
        RECT -1.525 31.485 -1.195 31.815 ;
        RECT -1.525 29.175 -1.195 29.505 ;
        RECT -1.525 28.325 -1.195 28.655 ;
        RECT -1.525 26.015 -1.195 26.345 ;
        RECT -1.525 25.165 -1.195 25.495 ;
        RECT -1.525 22.855 -1.195 23.185 ;
        RECT -1.525 22.005 -1.195 22.335 ;
        RECT -1.525 19.695 -1.195 20.025 ;
        RECT -1.525 18.115 -1.195 18.445 ;
        RECT -1.525 17.265 -1.195 17.595 ;
        RECT -1.525 14.955 -1.195 15.285 ;
        RECT -1.525 14.105 -1.195 14.435 ;
        RECT -1.525 11.795 -1.195 12.125 ;
        RECT -1.525 10.945 -1.195 11.275 ;
        RECT -1.525 8.635 -1.195 8.965 ;
        RECT -1.525 7.785 -1.195 8.115 ;
        RECT -1.525 5.475 -1.195 5.805 ;
        RECT -1.525 3.895 -1.195 4.225 ;
        RECT -1.525 3.045 -1.195 3.375 ;
        RECT -1.525 0.87 -1.195 1.2 ;
        RECT -1.525 -0.845 -1.195 -0.515 ;
        RECT -1.525 -2.205 -1.195 -1.875 ;
        RECT -1.525 -3.565 -1.195 -3.235 ;
        RECT -1.525 -4.925 -1.195 -4.595 ;
        RECT -1.525 -6.285 -1.195 -5.955 ;
        RECT -1.525 -7.645 -1.195 -7.315 ;
        RECT -1.525 -9.005 -1.195 -8.675 ;
        RECT -1.525 -10.365 -1.195 -10.035 ;
        RECT -1.525 -11.725 -1.195 -11.395 ;
        RECT -1.525 -13.085 -1.195 -12.755 ;
        RECT -1.525 -14.445 -1.195 -14.115 ;
        RECT -1.525 -15.805 -1.195 -15.475 ;
        RECT -1.525 -17.165 -1.195 -16.835 ;
        RECT -1.525 -23.965 -1.195 -23.635 ;
        RECT -1.525 -25.325 -1.195 -24.995 ;
        RECT -1.525 -26.685 -1.195 -26.355 ;
        RECT -1.525 -28.045 -1.195 -27.715 ;
        RECT -1.525 -29.405 -1.195 -29.075 ;
        RECT -1.525 -30.765 -1.195 -30.435 ;
        RECT -1.525 -32.125 -1.195 -31.795 ;
        RECT -1.525 -33.485 -1.195 -33.155 ;
        RECT -1.525 -37.565 -1.195 -37.235 ;
        RECT -1.525 -40.285 -1.195 -39.955 ;
        RECT -1.525 -41.645 -1.195 -41.315 ;
        RECT -1.525 -43.005 -1.195 -42.675 ;
        RECT -1.525 -44.365 -1.195 -44.035 ;
        RECT -1.525 -45.725 -1.195 -45.395 ;
        RECT -1.525 -47.085 -1.195 -46.755 ;
        RECT -1.525 -48.445 -1.195 -48.115 ;
        RECT -1.525 -52.525 -1.195 -52.195 ;
        RECT -1.525 -53.885 -1.195 -53.555 ;
        RECT -1.525 -55.245 -1.195 -54.915 ;
        RECT -1.525 -56.605 -1.195 -56.275 ;
        RECT -1.525 -57.965 -1.195 -57.635 ;
        RECT -1.525 -59.325 -1.195 -58.995 ;
        RECT -1.525 -60.685 -1.195 -60.355 ;
        RECT -1.525 -62.045 -1.195 -61.715 ;
        RECT -1.525 -63.405 -1.195 -63.075 ;
        RECT -1.525 -64.765 -1.195 -64.435 ;
        RECT -1.525 -66.125 -1.195 -65.795 ;
        RECT -1.525 -68.845 -1.195 -68.515 ;
        RECT -1.525 -70.205 -1.195 -69.875 ;
        RECT -1.525 -71.565 -1.195 -71.235 ;
        RECT -1.525 -72.925 -1.195 -72.595 ;
        RECT -1.525 -74.285 -1.195 -73.955 ;
        RECT -1.525 -75.645 -1.195 -75.315 ;
        RECT -1.525 -77.005 -1.195 -76.675 ;
        RECT -1.525 -78.365 -1.195 -78.035 ;
        RECT -1.525 -79.725 -1.195 -79.395 ;
        RECT -1.525 -81.085 -1.195 -80.755 ;
        RECT -1.525 -82.445 -1.195 -82.115 ;
        RECT -1.525 -83.805 -1.195 -83.475 ;
        RECT -1.525 -85.165 -1.195 -84.835 ;
        RECT -1.525 -86.525 -1.195 -86.195 ;
        RECT -1.525 -87.885 -1.195 -87.555 ;
        RECT -1.525 -89.245 -1.195 -88.915 ;
        RECT -1.525 -90.605 -1.195 -90.275 ;
        RECT -1.525 -91.965 -1.195 -91.635 ;
        RECT -1.525 -93.325 -1.195 -92.995 ;
        RECT -1.525 -94.685 -1.195 -94.355 ;
        RECT -1.525 -96.045 -1.195 -95.715 ;
        RECT -1.525 -97.405 -1.195 -97.075 ;
        RECT -1.525 -98.765 -1.195 -98.435 ;
        RECT -1.525 -100.125 -1.195 -99.795 ;
        RECT -1.525 -101.485 -1.195 -101.155 ;
        RECT -1.525 -102.845 -1.195 -102.515 ;
        RECT -1.525 -104.205 -1.195 -103.875 ;
        RECT -1.525 -105.565 -1.195 -105.235 ;
        RECT -1.525 -106.925 -1.195 -106.595 ;
        RECT -1.525 -108.285 -1.195 -107.955 ;
        RECT -1.525 -109.645 -1.195 -109.315 ;
        RECT -1.525 -111.005 -1.195 -110.675 ;
        RECT -1.525 -112.365 -1.195 -112.035 ;
        RECT -1.525 -113.725 -1.195 -113.395 ;
        RECT -1.525 -115.085 -1.195 -114.755 ;
        RECT -1.525 -116.445 -1.195 -116.115 ;
        RECT -1.525 -117.805 -1.195 -117.475 ;
        RECT -1.525 -119.165 -1.195 -118.835 ;
        RECT -1.525 -120.525 -1.195 -120.195 ;
        RECT -1.525 -121.885 -1.195 -121.555 ;
        RECT -1.525 -123.245 -1.195 -122.915 ;
        RECT -1.525 -124.605 -1.195 -124.275 ;
        RECT -1.525 -125.965 -1.195 -125.635 ;
        RECT -1.525 -127.325 -1.195 -126.995 ;
        RECT -1.525 -128.685 -1.195 -128.355 ;
        RECT -1.525 -130.045 -1.195 -129.715 ;
        RECT -1.525 -131.405 -1.195 -131.075 ;
        RECT -1.525 -132.765 -1.195 -132.435 ;
        RECT -1.525 -134.125 -1.195 -133.795 ;
        RECT -1.525 -135.485 -1.195 -135.155 ;
        RECT -1.525 -136.845 -1.195 -136.515 ;
        RECT -1.525 -138.205 -1.195 -137.875 ;
        RECT -1.525 -139.565 -1.195 -139.235 ;
        RECT -1.525 -140.925 -1.195 -140.595 ;
        RECT -1.525 -142.285 -1.195 -141.955 ;
        RECT -1.525 -143.645 -1.195 -143.315 ;
        RECT -1.525 -145.005 -1.195 -144.675 ;
        RECT -1.525 -146.365 -1.195 -146.035 ;
        RECT -1.525 -147.725 -1.195 -147.395 ;
        RECT -1.525 -149.085 -1.195 -148.755 ;
        RECT -1.525 -150.445 -1.195 -150.115 ;
        RECT -1.525 -151.805 -1.195 -151.475 ;
        RECT -1.525 -153.165 -1.195 -152.835 ;
        RECT -1.525 -154.525 -1.195 -154.195 ;
        RECT -1.525 -155.885 -1.195 -155.555 ;
        RECT -1.525 -157.245 -1.195 -156.915 ;
        RECT -1.525 -158.605 -1.195 -158.275 ;
        RECT -1.525 -159.965 -1.195 -159.635 ;
        RECT -1.525 -161.325 -1.195 -160.995 ;
        RECT -1.525 -162.685 -1.195 -162.355 ;
        RECT -1.525 -164.045 -1.195 -163.715 ;
        RECT -1.525 -165.405 -1.195 -165.075 ;
        RECT -1.525 -166.765 -1.195 -166.435 ;
        RECT -1.525 -168.125 -1.195 -167.795 ;
        RECT -1.525 -169.485 -1.195 -169.155 ;
        RECT -1.525 -170.845 -1.195 -170.515 ;
        RECT -1.525 -172.205 -1.195 -171.875 ;
        RECT -1.525 -173.565 -1.195 -173.235 ;
        RECT -1.525 -174.925 -1.195 -174.595 ;
        RECT -1.525 -176.285 -1.195 -175.955 ;
        RECT -1.525 -177.645 -1.195 -177.315 ;
        RECT -1.525 -179.005 -1.195 -178.675 ;
        RECT -1.525 -184.65 -1.195 -183.52 ;
        RECT -1.52 -184.765 -1.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 244.04 0.165 245.17 ;
        RECT -0.165 239.875 0.165 240.205 ;
        RECT -0.165 238.515 0.165 238.845 ;
        RECT -0.165 237.155 0.165 237.485 ;
        RECT -0.16 237.155 0.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 -0.845 0.165 -0.515 ;
        RECT -0.165 -2.205 0.165 -1.875 ;
        RECT -0.165 -3.565 0.165 -3.235 ;
        RECT -0.16 -3.565 0.16 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.165 -96.045 0.165 -95.715 ;
        RECT -0.165 -97.405 0.165 -97.075 ;
        RECT -0.165 -98.765 0.165 -98.435 ;
        RECT -0.165 -100.125 0.165 -99.795 ;
        RECT -0.165 -101.485 0.165 -101.155 ;
        RECT -0.165 -102.845 0.165 -102.515 ;
        RECT -0.165 -104.205 0.165 -103.875 ;
        RECT -0.165 -105.565 0.165 -105.235 ;
        RECT -0.165 -106.925 0.165 -106.595 ;
        RECT -0.165 -108.285 0.165 -107.955 ;
        RECT -0.165 -109.645 0.165 -109.315 ;
        RECT -0.165 -111.005 0.165 -110.675 ;
        RECT -0.165 -112.365 0.165 -112.035 ;
        RECT -0.165 -113.725 0.165 -113.395 ;
        RECT -0.165 -115.085 0.165 -114.755 ;
        RECT -0.165 -116.445 0.165 -116.115 ;
        RECT -0.165 -117.805 0.165 -117.475 ;
        RECT -0.165 -119.165 0.165 -118.835 ;
        RECT -0.165 -120.525 0.165 -120.195 ;
        RECT -0.165 -121.885 0.165 -121.555 ;
        RECT -0.165 -123.245 0.165 -122.915 ;
        RECT -0.165 -124.605 0.165 -124.275 ;
        RECT -0.165 -125.965 0.165 -125.635 ;
        RECT -0.165 -127.325 0.165 -126.995 ;
        RECT -0.165 -128.685 0.165 -128.355 ;
        RECT -0.165 -130.045 0.165 -129.715 ;
        RECT -0.165 -131.405 0.165 -131.075 ;
        RECT -0.165 -132.765 0.165 -132.435 ;
        RECT -0.165 -134.125 0.165 -133.795 ;
        RECT -0.165 -135.485 0.165 -135.155 ;
        RECT -0.165 -136.845 0.165 -136.515 ;
        RECT -0.165 -138.205 0.165 -137.875 ;
        RECT -0.165 -139.565 0.165 -139.235 ;
        RECT -0.165 -140.925 0.165 -140.595 ;
        RECT -0.165 -142.285 0.165 -141.955 ;
        RECT -0.165 -143.645 0.165 -143.315 ;
        RECT -0.165 -145.005 0.165 -144.675 ;
        RECT -0.165 -146.365 0.165 -146.035 ;
        RECT -0.165 -147.725 0.165 -147.395 ;
        RECT -0.165 -149.085 0.165 -148.755 ;
        RECT -0.165 -150.445 0.165 -150.115 ;
        RECT -0.165 -151.805 0.165 -151.475 ;
        RECT -0.165 -153.165 0.165 -152.835 ;
        RECT -0.165 -154.525 0.165 -154.195 ;
        RECT -0.165 -155.885 0.165 -155.555 ;
        RECT -0.165 -157.245 0.165 -156.915 ;
        RECT -0.165 -158.605 0.165 -158.275 ;
        RECT -0.165 -159.965 0.165 -159.635 ;
        RECT -0.165 -161.325 0.165 -160.995 ;
        RECT -0.165 -162.685 0.165 -162.355 ;
        RECT -0.165 -164.045 0.165 -163.715 ;
        RECT -0.165 -165.405 0.165 -165.075 ;
        RECT -0.165 -166.765 0.165 -166.435 ;
        RECT -0.165 -168.125 0.165 -167.795 ;
        RECT -0.165 -169.485 0.165 -169.155 ;
        RECT -0.165 -170.845 0.165 -170.515 ;
        RECT -0.165 -172.205 0.165 -171.875 ;
        RECT -0.165 -173.565 0.165 -173.235 ;
        RECT -0.165 -174.925 0.165 -174.595 ;
        RECT -0.165 -176.285 0.165 -175.955 ;
        RECT -0.165 -177.645 0.165 -177.315 ;
        RECT -0.165 -179.005 0.165 -178.675 ;
        RECT -0.165 -184.65 0.165 -183.52 ;
        RECT -0.16 -184.765 0.16 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 244.04 1.525 245.17 ;
        RECT 1.195 239.875 1.525 240.205 ;
        RECT 1.195 238.515 1.525 238.845 ;
        RECT 1.195 237.155 1.525 237.485 ;
        RECT 1.2 237.155 1.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 -0.845 1.525 -0.515 ;
        RECT 1.195 -2.205 1.525 -1.875 ;
        RECT 1.195 -3.565 1.525 -3.235 ;
        RECT 1.2 -3.565 1.52 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.195 -96.045 1.525 -95.715 ;
        RECT 1.195 -97.405 1.525 -97.075 ;
        RECT 1.195 -98.765 1.525 -98.435 ;
        RECT 1.195 -100.125 1.525 -99.795 ;
        RECT 1.195 -101.485 1.525 -101.155 ;
        RECT 1.195 -102.845 1.525 -102.515 ;
        RECT 1.195 -104.205 1.525 -103.875 ;
        RECT 1.195 -105.565 1.525 -105.235 ;
        RECT 1.195 -106.925 1.525 -106.595 ;
        RECT 1.195 -108.285 1.525 -107.955 ;
        RECT 1.195 -109.645 1.525 -109.315 ;
        RECT 1.195 -111.005 1.525 -110.675 ;
        RECT 1.195 -112.365 1.525 -112.035 ;
        RECT 1.195 -113.725 1.525 -113.395 ;
        RECT 1.195 -115.085 1.525 -114.755 ;
        RECT 1.195 -116.445 1.525 -116.115 ;
        RECT 1.195 -117.805 1.525 -117.475 ;
        RECT 1.195 -119.165 1.525 -118.835 ;
        RECT 1.195 -120.525 1.525 -120.195 ;
        RECT 1.195 -121.885 1.525 -121.555 ;
        RECT 1.195 -123.245 1.525 -122.915 ;
        RECT 1.195 -124.605 1.525 -124.275 ;
        RECT 1.195 -125.965 1.525 -125.635 ;
        RECT 1.195 -127.325 1.525 -126.995 ;
        RECT 1.195 -128.685 1.525 -128.355 ;
        RECT 1.195 -130.045 1.525 -129.715 ;
        RECT 1.195 -131.405 1.525 -131.075 ;
        RECT 1.195 -132.765 1.525 -132.435 ;
        RECT 1.195 -134.125 1.525 -133.795 ;
        RECT 1.195 -135.485 1.525 -135.155 ;
        RECT 1.195 -136.845 1.525 -136.515 ;
        RECT 1.195 -138.205 1.525 -137.875 ;
        RECT 1.195 -139.565 1.525 -139.235 ;
        RECT 1.195 -140.925 1.525 -140.595 ;
        RECT 1.195 -142.285 1.525 -141.955 ;
        RECT 1.195 -143.645 1.525 -143.315 ;
        RECT 1.195 -145.005 1.525 -144.675 ;
        RECT 1.195 -146.365 1.525 -146.035 ;
        RECT 1.195 -147.725 1.525 -147.395 ;
        RECT 1.195 -149.085 1.525 -148.755 ;
        RECT 1.195 -150.445 1.525 -150.115 ;
        RECT 1.195 -151.805 1.525 -151.475 ;
        RECT 1.195 -153.165 1.525 -152.835 ;
        RECT 1.195 -154.525 1.525 -154.195 ;
        RECT 1.195 -155.885 1.525 -155.555 ;
        RECT 1.195 -157.245 1.525 -156.915 ;
        RECT 1.195 -158.605 1.525 -158.275 ;
        RECT 1.195 -159.965 1.525 -159.635 ;
        RECT 1.195 -161.325 1.525 -160.995 ;
        RECT 1.195 -162.685 1.525 -162.355 ;
        RECT 1.195 -164.045 1.525 -163.715 ;
        RECT 1.195 -165.405 1.525 -165.075 ;
        RECT 1.195 -166.765 1.525 -166.435 ;
        RECT 1.195 -168.125 1.525 -167.795 ;
        RECT 1.195 -169.485 1.525 -169.155 ;
        RECT 1.195 -170.845 1.525 -170.515 ;
        RECT 1.195 -172.205 1.525 -171.875 ;
        RECT 1.195 -173.565 1.525 -173.235 ;
        RECT 1.195 -174.925 1.525 -174.595 ;
        RECT 1.195 -176.285 1.525 -175.955 ;
        RECT 1.195 -177.645 1.525 -177.315 ;
        RECT 1.195 -179.005 1.525 -178.675 ;
        RECT 1.195 -184.65 1.525 -183.52 ;
        RECT 1.2 -184.765 1.52 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 244.04 2.885 245.17 ;
        RECT 2.555 239.875 2.885 240.205 ;
        RECT 2.555 238.515 2.885 238.845 ;
        RECT 2.555 237.155 2.885 237.485 ;
        RECT 2.56 237.155 2.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.555 -98.765 2.885 -98.435 ;
        RECT 2.555 -100.125 2.885 -99.795 ;
        RECT 2.555 -101.485 2.885 -101.155 ;
        RECT 2.555 -102.845 2.885 -102.515 ;
        RECT 2.555 -104.205 2.885 -103.875 ;
        RECT 2.555 -105.565 2.885 -105.235 ;
        RECT 2.555 -106.925 2.885 -106.595 ;
        RECT 2.555 -108.285 2.885 -107.955 ;
        RECT 2.555 -109.645 2.885 -109.315 ;
        RECT 2.555 -111.005 2.885 -110.675 ;
        RECT 2.555 -112.365 2.885 -112.035 ;
        RECT 2.555 -113.725 2.885 -113.395 ;
        RECT 2.555 -115.085 2.885 -114.755 ;
        RECT 2.555 -116.445 2.885 -116.115 ;
        RECT 2.555 -117.805 2.885 -117.475 ;
        RECT 2.555 -119.165 2.885 -118.835 ;
        RECT 2.555 -120.525 2.885 -120.195 ;
        RECT 2.555 -121.885 2.885 -121.555 ;
        RECT 2.555 -123.245 2.885 -122.915 ;
        RECT 2.555 -124.605 2.885 -124.275 ;
        RECT 2.555 -125.965 2.885 -125.635 ;
        RECT 2.555 -127.325 2.885 -126.995 ;
        RECT 2.555 -128.685 2.885 -128.355 ;
        RECT 2.555 -130.045 2.885 -129.715 ;
        RECT 2.555 -131.405 2.885 -131.075 ;
        RECT 2.555 -132.765 2.885 -132.435 ;
        RECT 2.555 -134.125 2.885 -133.795 ;
        RECT 2.555 -135.485 2.885 -135.155 ;
        RECT 2.555 -136.845 2.885 -136.515 ;
        RECT 2.555 -138.205 2.885 -137.875 ;
        RECT 2.555 -139.565 2.885 -139.235 ;
        RECT 2.555 -140.925 2.885 -140.595 ;
        RECT 2.555 -142.285 2.885 -141.955 ;
        RECT 2.555 -143.645 2.885 -143.315 ;
        RECT 2.555 -145.005 2.885 -144.675 ;
        RECT 2.555 -146.365 2.885 -146.035 ;
        RECT 2.555 -147.725 2.885 -147.395 ;
        RECT 2.555 -149.085 2.885 -148.755 ;
        RECT 2.555 -150.445 2.885 -150.115 ;
        RECT 2.555 -151.805 2.885 -151.475 ;
        RECT 2.555 -153.165 2.885 -152.835 ;
        RECT 2.555 -154.525 2.885 -154.195 ;
        RECT 2.555 -155.885 2.885 -155.555 ;
        RECT 2.555 -157.245 2.885 -156.915 ;
        RECT 2.555 -158.605 2.885 -158.275 ;
        RECT 2.555 -159.965 2.885 -159.635 ;
        RECT 2.555 -161.325 2.885 -160.995 ;
        RECT 2.555 -162.685 2.885 -162.355 ;
        RECT 2.555 -164.045 2.885 -163.715 ;
        RECT 2.555 -165.405 2.885 -165.075 ;
        RECT 2.555 -166.765 2.885 -166.435 ;
        RECT 2.555 -168.125 2.885 -167.795 ;
        RECT 2.555 -169.485 2.885 -169.155 ;
        RECT 2.555 -170.845 2.885 -170.515 ;
        RECT 2.555 -172.205 2.885 -171.875 ;
        RECT 2.555 -173.565 2.885 -173.235 ;
        RECT 2.555 -174.925 2.885 -174.595 ;
        RECT 2.555 -176.285 2.885 -175.955 ;
        RECT 2.555 -177.645 2.885 -177.315 ;
        RECT 2.555 -179.005 2.885 -178.675 ;
        RECT 2.555 -184.65 2.885 -183.52 ;
        RECT 2.56 -184.765 2.88 -98.435 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.66 -98.075 2.99 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.915 244.04 4.245 245.17 ;
        RECT 3.915 239.875 4.245 240.205 ;
        RECT 3.915 238.515 4.245 238.845 ;
        RECT 3.915 237.155 4.245 237.485 ;
        RECT 3.92 237.155 4.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 244.04 5.605 245.17 ;
        RECT 5.275 239.875 5.605 240.205 ;
        RECT 5.275 238.515 5.605 238.845 ;
        RECT 5.275 237.155 5.605 237.485 ;
        RECT 5.28 237.155 5.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.275 -0.845 5.605 -0.515 ;
        RECT 5.275 -2.205 5.605 -1.875 ;
        RECT 5.275 -3.565 5.605 -3.235 ;
        RECT 5.28 -3.565 5.6 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 244.04 6.965 245.17 ;
        RECT 6.635 239.875 6.965 240.205 ;
        RECT 6.635 238.515 6.965 238.845 ;
        RECT 6.635 237.155 6.965 237.485 ;
        RECT 6.64 237.155 6.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 6.635 -0.845 6.965 -0.515 ;
        RECT 6.635 -2.205 6.965 -1.875 ;
        RECT 6.635 -3.565 6.965 -3.235 ;
        RECT 6.64 -3.565 6.96 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 244.04 8.325 245.17 ;
        RECT 7.995 239.875 8.325 240.205 ;
        RECT 7.995 238.515 8.325 238.845 ;
        RECT 7.995 237.155 8.325 237.485 ;
        RECT 8 237.155 8.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 -0.845 8.325 -0.515 ;
        RECT 7.995 -2.205 8.325 -1.875 ;
        RECT 7.995 -3.565 8.325 -3.235 ;
        RECT 8 -3.565 8.32 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.995 -96.045 8.325 -95.715 ;
        RECT 7.995 -97.405 8.325 -97.075 ;
        RECT 7.995 -98.765 8.325 -98.435 ;
        RECT 7.995 -100.125 8.325 -99.795 ;
        RECT 7.995 -101.485 8.325 -101.155 ;
        RECT 7.995 -102.845 8.325 -102.515 ;
        RECT 7.995 -104.205 8.325 -103.875 ;
        RECT 7.995 -105.565 8.325 -105.235 ;
        RECT 7.995 -106.925 8.325 -106.595 ;
        RECT 7.995 -108.285 8.325 -107.955 ;
        RECT 7.995 -109.645 8.325 -109.315 ;
        RECT 7.995 -111.005 8.325 -110.675 ;
        RECT 7.995 -112.365 8.325 -112.035 ;
        RECT 7.995 -113.725 8.325 -113.395 ;
        RECT 7.995 -115.085 8.325 -114.755 ;
        RECT 7.995 -116.445 8.325 -116.115 ;
        RECT 7.995 -117.805 8.325 -117.475 ;
        RECT 7.995 -119.165 8.325 -118.835 ;
        RECT 7.995 -120.525 8.325 -120.195 ;
        RECT 7.995 -121.885 8.325 -121.555 ;
        RECT 7.995 -123.245 8.325 -122.915 ;
        RECT 7.995 -124.605 8.325 -124.275 ;
        RECT 7.995 -125.965 8.325 -125.635 ;
        RECT 7.995 -127.325 8.325 -126.995 ;
        RECT 7.995 -128.685 8.325 -128.355 ;
        RECT 7.995 -130.045 8.325 -129.715 ;
        RECT 7.995 -131.405 8.325 -131.075 ;
        RECT 7.995 -132.765 8.325 -132.435 ;
        RECT 7.995 -134.125 8.325 -133.795 ;
        RECT 7.995 -135.485 8.325 -135.155 ;
        RECT 7.995 -136.845 8.325 -136.515 ;
        RECT 7.995 -138.205 8.325 -137.875 ;
        RECT 7.995 -139.565 8.325 -139.235 ;
        RECT 7.995 -140.925 8.325 -140.595 ;
        RECT 7.995 -142.285 8.325 -141.955 ;
        RECT 7.995 -143.645 8.325 -143.315 ;
        RECT 7.995 -145.005 8.325 -144.675 ;
        RECT 7.995 -146.365 8.325 -146.035 ;
        RECT 7.995 -147.725 8.325 -147.395 ;
        RECT 7.995 -149.085 8.325 -148.755 ;
        RECT 7.995 -150.445 8.325 -150.115 ;
        RECT 7.995 -151.805 8.325 -151.475 ;
        RECT 7.995 -153.165 8.325 -152.835 ;
        RECT 7.995 -154.525 8.325 -154.195 ;
        RECT 7.995 -155.885 8.325 -155.555 ;
        RECT 7.995 -157.245 8.325 -156.915 ;
        RECT 7.995 -158.605 8.325 -158.275 ;
        RECT 7.995 -159.965 8.325 -159.635 ;
        RECT 7.995 -161.325 8.325 -160.995 ;
        RECT 7.995 -162.685 8.325 -162.355 ;
        RECT 7.995 -164.045 8.325 -163.715 ;
        RECT 7.995 -165.405 8.325 -165.075 ;
        RECT 7.995 -166.765 8.325 -166.435 ;
        RECT 7.995 -168.125 8.325 -167.795 ;
        RECT 7.995 -169.485 8.325 -169.155 ;
        RECT 7.995 -170.845 8.325 -170.515 ;
        RECT 7.995 -172.205 8.325 -171.875 ;
        RECT 7.995 -173.565 8.325 -173.235 ;
        RECT 7.995 -174.925 8.325 -174.595 ;
        RECT 7.995 -176.285 8.325 -175.955 ;
        RECT 7.995 -177.645 8.325 -177.315 ;
        RECT 7.995 -179.005 8.325 -178.675 ;
        RECT 7.995 -184.65 8.325 -183.52 ;
        RECT 8 -184.765 8.32 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 244.04 9.685 245.17 ;
        RECT 9.355 239.875 9.685 240.205 ;
        RECT 9.355 238.515 9.685 238.845 ;
        RECT 9.355 237.155 9.685 237.485 ;
        RECT 9.36 237.155 9.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 -0.845 9.685 -0.515 ;
        RECT 9.355 -2.205 9.685 -1.875 ;
        RECT 9.355 -3.565 9.685 -3.235 ;
        RECT 9.36 -3.565 9.68 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 9.355 -96.045 9.685 -95.715 ;
        RECT 9.355 -97.405 9.685 -97.075 ;
        RECT 9.355 -98.765 9.685 -98.435 ;
        RECT 9.355 -100.125 9.685 -99.795 ;
        RECT 9.355 -101.485 9.685 -101.155 ;
        RECT 9.355 -102.845 9.685 -102.515 ;
        RECT 9.355 -104.205 9.685 -103.875 ;
        RECT 9.355 -105.565 9.685 -105.235 ;
        RECT 9.355 -106.925 9.685 -106.595 ;
        RECT 9.355 -108.285 9.685 -107.955 ;
        RECT 9.355 -109.645 9.685 -109.315 ;
        RECT 9.355 -111.005 9.685 -110.675 ;
        RECT 9.355 -112.365 9.685 -112.035 ;
        RECT 9.355 -113.725 9.685 -113.395 ;
        RECT 9.355 -115.085 9.685 -114.755 ;
        RECT 9.355 -116.445 9.685 -116.115 ;
        RECT 9.355 -117.805 9.685 -117.475 ;
        RECT 9.355 -119.165 9.685 -118.835 ;
        RECT 9.355 -120.525 9.685 -120.195 ;
        RECT 9.355 -121.885 9.685 -121.555 ;
        RECT 9.355 -123.245 9.685 -122.915 ;
        RECT 9.355 -124.605 9.685 -124.275 ;
        RECT 9.355 -125.965 9.685 -125.635 ;
        RECT 9.355 -127.325 9.685 -126.995 ;
        RECT 9.355 -128.685 9.685 -128.355 ;
        RECT 9.355 -130.045 9.685 -129.715 ;
        RECT 9.355 -131.405 9.685 -131.075 ;
        RECT 9.355 -132.765 9.685 -132.435 ;
        RECT 9.355 -134.125 9.685 -133.795 ;
        RECT 9.355 -135.485 9.685 -135.155 ;
        RECT 9.355 -136.845 9.685 -136.515 ;
        RECT 9.355 -138.205 9.685 -137.875 ;
        RECT 9.355 -139.565 9.685 -139.235 ;
        RECT 9.355 -140.925 9.685 -140.595 ;
        RECT 9.355 -142.285 9.685 -141.955 ;
        RECT 9.355 -143.645 9.685 -143.315 ;
        RECT 9.355 -145.005 9.685 -144.675 ;
        RECT 9.355 -146.365 9.685 -146.035 ;
        RECT 9.355 -147.725 9.685 -147.395 ;
        RECT 9.355 -149.085 9.685 -148.755 ;
        RECT 9.355 -150.445 9.685 -150.115 ;
        RECT 9.355 -151.805 9.685 -151.475 ;
        RECT 9.355 -153.165 9.685 -152.835 ;
        RECT 9.355 -154.525 9.685 -154.195 ;
        RECT 9.355 -155.885 9.685 -155.555 ;
        RECT 9.355 -157.245 9.685 -156.915 ;
        RECT 9.355 -158.605 9.685 -158.275 ;
        RECT 9.355 -159.965 9.685 -159.635 ;
        RECT 9.355 -161.325 9.685 -160.995 ;
        RECT 9.355 -162.685 9.685 -162.355 ;
        RECT 9.355 -164.045 9.685 -163.715 ;
        RECT 9.355 -165.405 9.685 -165.075 ;
        RECT 9.355 -166.765 9.685 -166.435 ;
        RECT 9.355 -168.125 9.685 -167.795 ;
        RECT 9.355 -169.485 9.685 -169.155 ;
        RECT 9.355 -170.845 9.685 -170.515 ;
        RECT 9.355 -172.205 9.685 -171.875 ;
        RECT 9.355 -173.565 9.685 -173.235 ;
        RECT 9.355 -174.925 9.685 -174.595 ;
        RECT 9.355 -176.285 9.685 -175.955 ;
        RECT 9.355 -177.645 9.685 -177.315 ;
        RECT 9.355 -179.005 9.685 -178.675 ;
        RECT 9.355 -184.65 9.685 -183.52 ;
        RECT 9.36 -184.765 9.68 -95.04 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 244.04 11.045 245.17 ;
        RECT 10.715 239.875 11.045 240.205 ;
        RECT 10.715 238.515 11.045 238.845 ;
        RECT 10.715 237.155 11.045 237.485 ;
        RECT 10.72 237.155 11.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 -0.845 11.045 -0.515 ;
        RECT 10.715 -2.205 11.045 -1.875 ;
        RECT 10.715 -3.565 11.045 -3.235 ;
        RECT 10.72 -3.565 11.04 -0.515 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.715 -102.845 11.045 -102.515 ;
        RECT 10.715 -104.205 11.045 -103.875 ;
        RECT 10.715 -105.565 11.045 -105.235 ;
        RECT 10.715 -106.925 11.045 -106.595 ;
        RECT 10.715 -108.285 11.045 -107.955 ;
        RECT 10.715 -109.645 11.045 -109.315 ;
        RECT 10.715 -111.005 11.045 -110.675 ;
        RECT 10.715 -112.365 11.045 -112.035 ;
        RECT 10.715 -113.725 11.045 -113.395 ;
        RECT 10.715 -115.085 11.045 -114.755 ;
        RECT 10.715 -116.445 11.045 -116.115 ;
        RECT 10.715 -117.805 11.045 -117.475 ;
        RECT 10.715 -119.165 11.045 -118.835 ;
        RECT 10.715 -120.525 11.045 -120.195 ;
        RECT 10.715 -121.885 11.045 -121.555 ;
        RECT 10.715 -123.245 11.045 -122.915 ;
        RECT 10.715 -124.605 11.045 -124.275 ;
        RECT 10.715 -125.965 11.045 -125.635 ;
        RECT 10.715 -127.325 11.045 -126.995 ;
        RECT 10.715 -128.685 11.045 -128.355 ;
        RECT 10.715 -130.045 11.045 -129.715 ;
        RECT 10.715 -131.405 11.045 -131.075 ;
        RECT 10.715 -132.765 11.045 -132.435 ;
        RECT 10.715 -134.125 11.045 -133.795 ;
        RECT 10.715 -135.485 11.045 -135.155 ;
        RECT 10.715 -136.845 11.045 -136.515 ;
        RECT 10.715 -138.205 11.045 -137.875 ;
        RECT 10.715 -139.565 11.045 -139.235 ;
        RECT 10.715 -140.925 11.045 -140.595 ;
        RECT 10.715 -142.285 11.045 -141.955 ;
        RECT 10.715 -143.645 11.045 -143.315 ;
        RECT 10.715 -145.005 11.045 -144.675 ;
        RECT 10.715 -146.365 11.045 -146.035 ;
        RECT 10.715 -147.725 11.045 -147.395 ;
        RECT 10.715 -149.085 11.045 -148.755 ;
        RECT 10.715 -150.445 11.045 -150.115 ;
        RECT 10.715 -151.805 11.045 -151.475 ;
        RECT 10.715 -153.165 11.045 -152.835 ;
        RECT 10.715 -154.525 11.045 -154.195 ;
        RECT 10.715 -155.885 11.045 -155.555 ;
        RECT 10.715 -157.245 11.045 -156.915 ;
        RECT 10.715 -158.605 11.045 -158.275 ;
        RECT 10.715 -159.965 11.045 -159.635 ;
        RECT 10.715 -161.325 11.045 -160.995 ;
        RECT 10.715 -162.685 11.045 -162.355 ;
        RECT 10.715 -164.045 11.045 -163.715 ;
        RECT 10.715 -165.405 11.045 -165.075 ;
        RECT 10.715 -166.765 11.045 -166.435 ;
        RECT 10.715 -168.125 11.045 -167.795 ;
        RECT 10.715 -169.485 11.045 -169.155 ;
        RECT 10.715 -170.845 11.045 -170.515 ;
        RECT 10.715 -172.205 11.045 -171.875 ;
        RECT 10.715 -173.565 11.045 -173.235 ;
        RECT 10.715 -174.925 11.045 -174.595 ;
        RECT 10.715 -176.285 11.045 -175.955 ;
        RECT 10.715 -177.645 11.045 -177.315 ;
        RECT 10.715 -179.005 11.045 -178.675 ;
        RECT 10.715 -184.65 11.045 -183.52 ;
        RECT 10.72 -184.765 11.04 -95.04 ;
        RECT 10.715 -96.045 11.045 -95.715 ;
        RECT 10.715 -97.405 11.045 -97.075 ;
        RECT 10.715 -98.765 11.045 -98.435 ;
        RECT 10.715 -100.125 11.045 -99.795 ;
        RECT 10.715 -101.485 11.045 -101.155 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.325 244.04 -7.995 245.17 ;
        RECT -8.325 239.875 -7.995 240.205 ;
        RECT -8.325 238.515 -7.995 238.845 ;
        RECT -8.325 237.155 -7.995 237.485 ;
        RECT -8.325 235.795 -7.995 236.125 ;
        RECT -8.325 234.435 -7.995 234.765 ;
        RECT -8.325 233.075 -7.995 233.405 ;
        RECT -8.325 231.715 -7.995 232.045 ;
        RECT -8.325 227.635 -7.995 227.965 ;
        RECT -8.325 224.915 -7.995 225.245 ;
        RECT -8.325 218.115 -7.995 218.445 ;
        RECT -8.325 216.755 -7.995 217.085 ;
        RECT -8.325 207.235 -7.995 207.565 ;
        RECT -8.325 204.515 -7.995 204.845 ;
        RECT -8.325 203.155 -7.995 203.485 ;
        RECT -8.325 199.075 -7.995 199.405 ;
        RECT -8.325 196.355 -7.995 196.685 ;
        RECT -8.325 189.555 -7.995 189.885 ;
        RECT -8.325 188.195 -7.995 188.525 ;
        RECT -8.325 185.475 -7.995 185.805 ;
        RECT -8.325 178.675 -7.995 179.005 ;
        RECT -8.325 175.955 -7.995 176.285 ;
        RECT -8.325 174.595 -7.995 174.925 ;
        RECT -8.325 167.795 -7.995 168.125 ;
        RECT -8.325 160.995 -7.995 161.325 ;
        RECT -8.325 159.635 -7.995 159.965 ;
        RECT -8.325 156.915 -7.995 157.245 ;
        RECT -8.325 150.115 -7.995 150.445 ;
        RECT -8.325 147.395 -7.995 147.725 ;
        RECT -8.325 146.035 -7.995 146.365 ;
        RECT -8.325 139.235 -7.995 139.565 ;
        RECT -8.325 136.515 -7.995 136.845 ;
        RECT -8.325 132.435 -7.995 132.765 ;
        RECT -8.325 131.075 -7.995 131.405 ;
        RECT -8.325 128.355 -7.995 128.685 ;
        RECT -8.325 118.835 -7.995 119.165 ;
        RECT -8.325 117.475 -7.995 117.805 ;
        RECT -8.325 110.675 -7.995 111.005 ;
        RECT -8.325 107.955 -7.995 108.285 ;
        RECT -8.325 103.875 -7.995 104.205 ;
        RECT -8.325 99.795 -7.995 100.125 ;
        RECT -8.325 97.075 -7.995 97.405 ;
        RECT -8.325 90.275 -7.995 90.605 ;
        RECT -8.325 88.915 -7.995 89.245 ;
        RECT -8.325 82.115 -7.995 82.445 ;
        RECT -8.325 79.395 -7.995 79.725 ;
        RECT -8.325 75.315 -7.995 75.645 ;
        RECT -8.325 71.235 -7.995 71.565 ;
        RECT -8.325 68.515 -7.995 68.845 ;
        RECT -8.325 61.715 -7.995 62.045 ;
        RECT -8.325 60.355 -7.995 60.685 ;
        RECT -8.325 50.835 -7.995 51.165 ;
        RECT -8.325 46.755 -7.995 47.085 ;
        RECT -8.325 42.675 -7.995 43.005 ;
        RECT -8.325 39.955 -7.995 40.285 ;
        RECT -8.325 33.155 -7.995 33.485 ;
        RECT -8.325 31.795 -7.995 32.125 ;
        RECT -8.325 29.075 -7.995 29.405 ;
        RECT -8.325 22.275 -7.995 22.605 ;
        RECT -8.325 19.555 -7.995 19.885 ;
        RECT -8.325 18.195 -7.995 18.525 ;
        RECT -8.325 11.395 -7.995 11.725 ;
        RECT -8.325 4.595 -7.995 4.925 ;
        RECT -8.325 3.235 -7.995 3.565 ;
        RECT -8.325 1.875 -7.995 2.205 ;
        RECT -8.325 0.515 -7.995 0.845 ;
        RECT -8.325 -0.845 -7.995 -0.515 ;
        RECT -8.325 -2.205 -7.995 -1.875 ;
        RECT -8.325 -3.565 -7.995 -3.235 ;
        RECT -8.325 -4.925 -7.995 -4.595 ;
        RECT -8.325 -6.285 -7.995 -5.955 ;
        RECT -8.325 -7.645 -7.995 -7.315 ;
        RECT -8.325 -9.005 -7.995 -8.675 ;
        RECT -8.325 -10.365 -7.995 -10.035 ;
        RECT -8.325 -11.725 -7.995 -11.395 ;
        RECT -8.325 -13.085 -7.995 -12.755 ;
        RECT -8.325 -14.445 -7.995 -14.115 ;
        RECT -8.325 -15.805 -7.995 -15.475 ;
        RECT -8.325 -17.165 -7.995 -16.835 ;
        RECT -8.32 -21.24 -8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -8.325 -106.925 -7.995 -106.595 ;
        RECT -8.325 -108.285 -7.995 -107.955 ;
        RECT -8.325 -109.645 -7.995 -109.315 ;
        RECT -8.325 -111.005 -7.995 -110.675 ;
        RECT -8.325 -112.365 -7.995 -112.035 ;
        RECT -8.325 -113.725 -7.995 -113.395 ;
        RECT -8.325 -115.085 -7.995 -114.755 ;
        RECT -8.325 -116.445 -7.995 -116.115 ;
        RECT -8.325 -117.805 -7.995 -117.475 ;
        RECT -8.325 -119.165 -7.995 -118.835 ;
        RECT -8.325 -120.525 -7.995 -120.195 ;
        RECT -8.325 -121.885 -7.995 -121.555 ;
        RECT -8.325 -123.245 -7.995 -122.915 ;
        RECT -8.325 -124.605 -7.995 -124.275 ;
        RECT -8.325 -125.965 -7.995 -125.635 ;
        RECT -8.325 -127.325 -7.995 -126.995 ;
        RECT -8.325 -128.685 -7.995 -128.355 ;
        RECT -8.325 -130.045 -7.995 -129.715 ;
        RECT -8.325 -131.405 -7.995 -131.075 ;
        RECT -8.325 -132.765 -7.995 -132.435 ;
        RECT -8.325 -134.125 -7.995 -133.795 ;
        RECT -8.325 -135.485 -7.995 -135.155 ;
        RECT -8.325 -136.845 -7.995 -136.515 ;
        RECT -8.325 -138.205 -7.995 -137.875 ;
        RECT -8.325 -139.565 -7.995 -139.235 ;
        RECT -8.325 -140.925 -7.995 -140.595 ;
        RECT -8.325 -142.285 -7.995 -141.955 ;
        RECT -8.325 -143.645 -7.995 -143.315 ;
        RECT -8.325 -145.005 -7.995 -144.675 ;
        RECT -8.325 -146.365 -7.995 -146.035 ;
        RECT -8.325 -147.725 -7.995 -147.395 ;
        RECT -8.325 -149.085 -7.995 -148.755 ;
        RECT -8.325 -150.445 -7.995 -150.115 ;
        RECT -8.325 -151.805 -7.995 -151.475 ;
        RECT -8.325 -153.165 -7.995 -152.835 ;
        RECT -8.325 -154.525 -7.995 -154.195 ;
        RECT -8.325 -155.885 -7.995 -155.555 ;
        RECT -8.325 -157.245 -7.995 -156.915 ;
        RECT -8.325 -158.605 -7.995 -158.275 ;
        RECT -8.325 -159.965 -7.995 -159.635 ;
        RECT -8.325 -161.325 -7.995 -160.995 ;
        RECT -8.325 -162.685 -7.995 -162.355 ;
        RECT -8.325 -164.045 -7.995 -163.715 ;
        RECT -8.325 -165.405 -7.995 -165.075 ;
        RECT -8.32 -166.08 -8 -106.595 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.965 244.04 -6.635 245.17 ;
        RECT -6.965 239.875 -6.635 240.205 ;
        RECT -6.965 238.515 -6.635 238.845 ;
        RECT -6.965 237.155 -6.635 237.485 ;
        RECT -6.965 235.795 -6.635 236.125 ;
        RECT -6.965 234.435 -6.635 234.765 ;
        RECT -6.965 233.075 -6.635 233.405 ;
        RECT -6.965 231.715 -6.635 232.045 ;
        RECT -6.965 227.635 -6.635 227.965 ;
        RECT -6.965 224.915 -6.635 225.245 ;
        RECT -6.965 218.115 -6.635 218.445 ;
        RECT -6.965 216.755 -6.635 217.085 ;
        RECT -6.965 207.235 -6.635 207.565 ;
        RECT -6.965 204.515 -6.635 204.845 ;
        RECT -6.965 203.155 -6.635 203.485 ;
        RECT -6.965 199.075 -6.635 199.405 ;
        RECT -6.965 196.355 -6.635 196.685 ;
        RECT -6.965 189.555 -6.635 189.885 ;
        RECT -6.965 188.195 -6.635 188.525 ;
        RECT -6.965 185.475 -6.635 185.805 ;
        RECT -6.965 178.675 -6.635 179.005 ;
        RECT -6.965 175.955 -6.635 176.285 ;
        RECT -6.965 174.595 -6.635 174.925 ;
        RECT -6.965 167.795 -6.635 168.125 ;
        RECT -6.965 160.995 -6.635 161.325 ;
        RECT -6.965 159.635 -6.635 159.965 ;
        RECT -6.965 156.915 -6.635 157.245 ;
        RECT -6.965 150.115 -6.635 150.445 ;
        RECT -6.965 147.395 -6.635 147.725 ;
        RECT -6.965 146.035 -6.635 146.365 ;
        RECT -6.965 139.235 -6.635 139.565 ;
        RECT -6.965 136.515 -6.635 136.845 ;
        RECT -6.965 132.435 -6.635 132.765 ;
        RECT -6.965 131.075 -6.635 131.405 ;
        RECT -6.965 128.355 -6.635 128.685 ;
        RECT -6.965 118.835 -6.635 119.165 ;
        RECT -6.965 117.475 -6.635 117.805 ;
        RECT -6.965 110.675 -6.635 111.005 ;
        RECT -6.965 107.955 -6.635 108.285 ;
        RECT -6.965 103.875 -6.635 104.205 ;
        RECT -6.965 99.795 -6.635 100.125 ;
        RECT -6.965 97.075 -6.635 97.405 ;
        RECT -6.965 90.275 -6.635 90.605 ;
        RECT -6.965 88.915 -6.635 89.245 ;
        RECT -6.965 82.115 -6.635 82.445 ;
        RECT -6.965 79.395 -6.635 79.725 ;
        RECT -6.965 75.315 -6.635 75.645 ;
        RECT -6.965 71.235 -6.635 71.565 ;
        RECT -6.965 68.515 -6.635 68.845 ;
        RECT -6.965 61.715 -6.635 62.045 ;
        RECT -6.965 60.355 -6.635 60.685 ;
        RECT -6.965 50.835 -6.635 51.165 ;
        RECT -6.965 46.755 -6.635 47.085 ;
        RECT -6.965 42.675 -6.635 43.005 ;
        RECT -6.965 39.955 -6.635 40.285 ;
        RECT -6.965 33.155 -6.635 33.485 ;
        RECT -6.965 31.795 -6.635 32.125 ;
        RECT -6.965 29.075 -6.635 29.405 ;
        RECT -6.965 22.275 -6.635 22.605 ;
        RECT -6.965 19.555 -6.635 19.885 ;
        RECT -6.965 18.195 -6.635 18.525 ;
        RECT -6.965 11.395 -6.635 11.725 ;
        RECT -6.965 4.595 -6.635 4.925 ;
        RECT -6.965 3.235 -6.635 3.565 ;
        RECT -6.965 1.875 -6.635 2.205 ;
        RECT -6.965 0.515 -6.635 0.845 ;
        RECT -6.965 -0.845 -6.635 -0.515 ;
        RECT -6.965 -2.205 -6.635 -1.875 ;
        RECT -6.965 -3.565 -6.635 -3.235 ;
        RECT -6.965 -4.925 -6.635 -4.595 ;
        RECT -6.965 -6.285 -6.635 -5.955 ;
        RECT -6.965 -7.645 -6.635 -7.315 ;
        RECT -6.965 -9.005 -6.635 -8.675 ;
        RECT -6.965 -10.365 -6.635 -10.035 ;
        RECT -6.965 -11.725 -6.635 -11.395 ;
        RECT -6.965 -13.085 -6.635 -12.755 ;
        RECT -6.965 -14.445 -6.635 -14.115 ;
        RECT -6.965 -15.805 -6.635 -15.475 ;
        RECT -6.965 -17.165 -6.635 -16.835 ;
        RECT -6.965 -23.965 -6.635 -23.635 ;
        RECT -6.965 -25.325 -6.635 -24.995 ;
        RECT -6.965 -26.685 -6.635 -26.355 ;
        RECT -6.965 -28.045 -6.635 -27.715 ;
        RECT -6.965 -29.405 -6.635 -29.075 ;
        RECT -6.965 -30.765 -6.635 -30.435 ;
        RECT -6.965 -32.125 -6.635 -31.795 ;
        RECT -6.965 -33.485 -6.635 -33.155 ;
        RECT -6.965 -37.565 -6.635 -37.235 ;
        RECT -6.965 -40.285 -6.635 -39.955 ;
        RECT -6.965 -41.645 -6.635 -41.315 ;
        RECT -6.965 -43.005 -6.635 -42.675 ;
        RECT -6.965 -44.365 -6.635 -44.035 ;
        RECT -6.965 -45.725 -6.635 -45.395 ;
        RECT -6.965 -47.085 -6.635 -46.755 ;
        RECT -6.965 -48.445 -6.635 -48.115 ;
        RECT -6.965 -52.525 -6.635 -52.195 ;
        RECT -6.965 -53.885 -6.635 -53.555 ;
        RECT -6.965 -55.245 -6.635 -54.915 ;
        RECT -6.965 -56.605 -6.635 -56.275 ;
        RECT -6.965 -57.965 -6.635 -57.635 ;
        RECT -6.965 -59.325 -6.635 -58.995 ;
        RECT -6.965 -60.685 -6.635 -60.355 ;
        RECT -6.965 -62.045 -6.635 -61.715 ;
        RECT -6.965 -63.405 -6.635 -63.075 ;
        RECT -6.965 -64.765 -6.635 -64.435 ;
        RECT -6.965 -66.125 -6.635 -65.795 ;
        RECT -6.965 -68.845 -6.635 -68.515 ;
        RECT -6.965 -70.205 -6.635 -69.875 ;
        RECT -6.965 -71.565 -6.635 -71.235 ;
        RECT -6.965 -72.925 -6.635 -72.595 ;
        RECT -6.965 -74.285 -6.635 -73.955 ;
        RECT -6.965 -75.645 -6.635 -75.315 ;
        RECT -6.965 -77.005 -6.635 -76.675 ;
        RECT -6.965 -78.365 -6.635 -78.035 ;
        RECT -6.965 -79.725 -6.635 -79.395 ;
        RECT -6.965 -81.085 -6.635 -80.755 ;
        RECT -6.965 -82.445 -6.635 -82.115 ;
        RECT -6.965 -83.805 -6.635 -83.475 ;
        RECT -6.965 -85.165 -6.635 -84.835 ;
        RECT -6.965 -86.525 -6.635 -86.195 ;
        RECT -6.965 -87.885 -6.635 -87.555 ;
        RECT -6.965 -89.245 -6.635 -88.915 ;
        RECT -6.965 -90.605 -6.635 -90.275 ;
        RECT -6.965 -91.965 -6.635 -91.635 ;
        RECT -6.965 -93.325 -6.635 -92.995 ;
        RECT -6.965 -94.685 -6.635 -94.355 ;
        RECT -6.965 -96.045 -6.635 -95.715 ;
        RECT -6.965 -97.405 -6.635 -97.075 ;
        RECT -6.965 -98.765 -6.635 -98.435 ;
        RECT -6.965 -100.125 -6.635 -99.795 ;
        RECT -6.965 -101.485 -6.635 -101.155 ;
        RECT -6.965 -102.845 -6.635 -102.515 ;
        RECT -6.965 -104.205 -6.635 -103.875 ;
        RECT -6.965 -105.565 -6.635 -105.235 ;
        RECT -6.965 -106.925 -6.635 -106.595 ;
        RECT -6.965 -108.285 -6.635 -107.955 ;
        RECT -6.965 -109.645 -6.635 -109.315 ;
        RECT -6.965 -111.005 -6.635 -110.675 ;
        RECT -6.965 -112.365 -6.635 -112.035 ;
        RECT -6.965 -113.725 -6.635 -113.395 ;
        RECT -6.965 -115.085 -6.635 -114.755 ;
        RECT -6.965 -116.445 -6.635 -116.115 ;
        RECT -6.965 -117.805 -6.635 -117.475 ;
        RECT -6.965 -119.165 -6.635 -118.835 ;
        RECT -6.965 -120.525 -6.635 -120.195 ;
        RECT -6.965 -121.885 -6.635 -121.555 ;
        RECT -6.965 -123.245 -6.635 -122.915 ;
        RECT -6.965 -124.605 -6.635 -124.275 ;
        RECT -6.965 -125.965 -6.635 -125.635 ;
        RECT -6.965 -127.325 -6.635 -126.995 ;
        RECT -6.965 -128.685 -6.635 -128.355 ;
        RECT -6.965 -130.045 -6.635 -129.715 ;
        RECT -6.965 -131.405 -6.635 -131.075 ;
        RECT -6.965 -132.765 -6.635 -132.435 ;
        RECT -6.965 -134.125 -6.635 -133.795 ;
        RECT -6.965 -135.485 -6.635 -135.155 ;
        RECT -6.965 -136.845 -6.635 -136.515 ;
        RECT -6.965 -138.205 -6.635 -137.875 ;
        RECT -6.965 -139.565 -6.635 -139.235 ;
        RECT -6.965 -140.925 -6.635 -140.595 ;
        RECT -6.965 -142.285 -6.635 -141.955 ;
        RECT -6.965 -143.645 -6.635 -143.315 ;
        RECT -6.965 -145.005 -6.635 -144.675 ;
        RECT -6.965 -146.365 -6.635 -146.035 ;
        RECT -6.965 -147.725 -6.635 -147.395 ;
        RECT -6.965 -149.085 -6.635 -148.755 ;
        RECT -6.965 -150.445 -6.635 -150.115 ;
        RECT -6.965 -151.805 -6.635 -151.475 ;
        RECT -6.965 -153.165 -6.635 -152.835 ;
        RECT -6.965 -154.525 -6.635 -154.195 ;
        RECT -6.965 -155.885 -6.635 -155.555 ;
        RECT -6.965 -157.245 -6.635 -156.915 ;
        RECT -6.965 -158.605 -6.635 -158.275 ;
        RECT -6.965 -159.965 -6.635 -159.635 ;
        RECT -6.965 -161.325 -6.635 -160.995 ;
        RECT -6.965 -162.685 -6.635 -162.355 ;
        RECT -6.965 -164.045 -6.635 -163.715 ;
        RECT -6.965 -165.405 -6.635 -165.075 ;
        RECT -6.965 -166.765 -6.635 -166.435 ;
        RECT -6.965 -168.125 -6.635 -167.795 ;
        RECT -6.965 -169.485 -6.635 -169.155 ;
        RECT -6.965 -170.845 -6.635 -170.515 ;
        RECT -6.965 -172.205 -6.635 -171.875 ;
        RECT -6.965 -173.565 -6.635 -173.235 ;
        RECT -6.965 -174.925 -6.635 -174.595 ;
        RECT -6.965 -176.285 -6.635 -175.955 ;
        RECT -6.965 -177.645 -6.635 -177.315 ;
        RECT -6.965 -179.005 -6.635 -178.675 ;
        RECT -6.965 -184.65 -6.635 -183.52 ;
        RECT -6.96 -184.765 -6.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.605 244.04 -5.275 245.17 ;
        RECT -5.605 239.875 -5.275 240.205 ;
        RECT -5.605 238.515 -5.275 238.845 ;
        RECT -5.605 237.155 -5.275 237.485 ;
        RECT -5.605 235.17 -5.275 235.5 ;
        RECT -5.605 232.995 -5.275 233.325 ;
        RECT -5.605 231.415 -5.275 231.745 ;
        RECT -5.605 230.565 -5.275 230.895 ;
        RECT -5.605 228.255 -5.275 228.585 ;
        RECT -5.605 227.405 -5.275 227.735 ;
        RECT -5.605 225.095 -5.275 225.425 ;
        RECT -5.605 224.245 -5.275 224.575 ;
        RECT -5.605 221.935 -5.275 222.265 ;
        RECT -5.605 221.085 -5.275 221.415 ;
        RECT -5.605 218.775 -5.275 219.105 ;
        RECT -5.605 217.195 -5.275 217.525 ;
        RECT -5.605 216.345 -5.275 216.675 ;
        RECT -5.605 214.035 -5.275 214.365 ;
        RECT -5.605 213.185 -5.275 213.515 ;
        RECT -5.605 210.875 -5.275 211.205 ;
        RECT -5.605 210.025 -5.275 210.355 ;
        RECT -5.605 207.715 -5.275 208.045 ;
        RECT -5.605 206.865 -5.275 207.195 ;
        RECT -5.605 204.555 -5.275 204.885 ;
        RECT -5.605 202.975 -5.275 203.305 ;
        RECT -5.605 202.125 -5.275 202.455 ;
        RECT -5.605 199.815 -5.275 200.145 ;
        RECT -5.605 198.965 -5.275 199.295 ;
        RECT -5.605 196.655 -5.275 196.985 ;
        RECT -5.605 195.805 -5.275 196.135 ;
        RECT -5.605 193.495 -5.275 193.825 ;
        RECT -5.605 192.645 -5.275 192.975 ;
        RECT -5.605 190.335 -5.275 190.665 ;
        RECT -5.605 188.755 -5.275 189.085 ;
        RECT -5.605 187.905 -5.275 188.235 ;
        RECT -5.605 185.595 -5.275 185.925 ;
        RECT -5.605 184.745 -5.275 185.075 ;
        RECT -5.605 182.435 -5.275 182.765 ;
        RECT -5.605 181.585 -5.275 181.915 ;
        RECT -5.605 179.275 -5.275 179.605 ;
        RECT -5.605 178.425 -5.275 178.755 ;
        RECT -5.605 176.115 -5.275 176.445 ;
        RECT -5.605 174.535 -5.275 174.865 ;
        RECT -5.605 173.685 -5.275 174.015 ;
        RECT -5.605 171.375 -5.275 171.705 ;
        RECT -5.605 170.525 -5.275 170.855 ;
        RECT -5.605 168.215 -5.275 168.545 ;
        RECT -5.605 167.365 -5.275 167.695 ;
        RECT -5.605 165.055 -5.275 165.385 ;
        RECT -5.605 164.205 -5.275 164.535 ;
        RECT -5.605 161.895 -5.275 162.225 ;
        RECT -5.605 160.315 -5.275 160.645 ;
        RECT -5.605 159.465 -5.275 159.795 ;
        RECT -5.605 157.155 -5.275 157.485 ;
        RECT -5.605 156.305 -5.275 156.635 ;
        RECT -5.605 153.995 -5.275 154.325 ;
        RECT -5.605 153.145 -5.275 153.475 ;
        RECT -5.605 150.835 -5.275 151.165 ;
        RECT -5.605 149.985 -5.275 150.315 ;
        RECT -5.605 147.675 -5.275 148.005 ;
        RECT -5.605 146.095 -5.275 146.425 ;
        RECT -5.605 145.245 -5.275 145.575 ;
        RECT -5.605 142.935 -5.275 143.265 ;
        RECT -5.605 142.085 -5.275 142.415 ;
        RECT -5.605 139.775 -5.275 140.105 ;
        RECT -5.605 138.925 -5.275 139.255 ;
        RECT -5.605 136.615 -5.275 136.945 ;
        RECT -5.605 135.765 -5.275 136.095 ;
        RECT -5.605 133.455 -5.275 133.785 ;
        RECT -5.605 131.875 -5.275 132.205 ;
        RECT -5.605 131.025 -5.275 131.355 ;
        RECT -5.605 128.715 -5.275 129.045 ;
        RECT -5.605 127.865 -5.275 128.195 ;
        RECT -5.605 125.555 -5.275 125.885 ;
        RECT -5.605 124.705 -5.275 125.035 ;
        RECT -5.605 122.395 -5.275 122.725 ;
        RECT -5.605 121.545 -5.275 121.875 ;
        RECT -5.605 119.235 -5.275 119.565 ;
        RECT -5.605 117.655 -5.275 117.985 ;
        RECT -5.605 116.805 -5.275 117.135 ;
        RECT -5.605 114.495 -5.275 114.825 ;
        RECT -5.605 113.645 -5.275 113.975 ;
        RECT -5.605 111.335 -5.275 111.665 ;
        RECT -5.605 110.485 -5.275 110.815 ;
        RECT -5.605 108.175 -5.275 108.505 ;
        RECT -5.605 107.325 -5.275 107.655 ;
        RECT -5.605 105.015 -5.275 105.345 ;
        RECT -5.605 103.435 -5.275 103.765 ;
        RECT -5.605 102.585 -5.275 102.915 ;
        RECT -5.605 100.275 -5.275 100.605 ;
        RECT -5.605 99.425 -5.275 99.755 ;
        RECT -5.605 97.115 -5.275 97.445 ;
        RECT -5.605 96.265 -5.275 96.595 ;
        RECT -5.605 93.955 -5.275 94.285 ;
        RECT -5.605 93.105 -5.275 93.435 ;
        RECT -5.605 90.795 -5.275 91.125 ;
        RECT -5.605 89.215 -5.275 89.545 ;
        RECT -5.605 88.365 -5.275 88.695 ;
        RECT -5.605 86.055 -5.275 86.385 ;
        RECT -5.605 85.205 -5.275 85.535 ;
        RECT -5.605 82.895 -5.275 83.225 ;
        RECT -5.605 82.045 -5.275 82.375 ;
        RECT -5.605 79.735 -5.275 80.065 ;
        RECT -5.605 78.885 -5.275 79.215 ;
        RECT -5.605 76.575 -5.275 76.905 ;
        RECT -5.605 74.995 -5.275 75.325 ;
        RECT -5.605 74.145 -5.275 74.475 ;
        RECT -5.605 71.835 -5.275 72.165 ;
        RECT -5.605 70.985 -5.275 71.315 ;
        RECT -5.605 68.675 -5.275 69.005 ;
        RECT -5.605 67.825 -5.275 68.155 ;
        RECT -5.605 65.515 -5.275 65.845 ;
        RECT -5.605 64.665 -5.275 64.995 ;
        RECT -5.605 62.355 -5.275 62.685 ;
        RECT -5.605 60.775 -5.275 61.105 ;
        RECT -5.605 59.925 -5.275 60.255 ;
        RECT -5.605 57.615 -5.275 57.945 ;
        RECT -5.605 56.765 -5.275 57.095 ;
        RECT -5.605 54.455 -5.275 54.785 ;
        RECT -5.605 53.605 -5.275 53.935 ;
        RECT -5.605 51.295 -5.275 51.625 ;
        RECT -5.605 50.445 -5.275 50.775 ;
        RECT -5.605 48.135 -5.275 48.465 ;
        RECT -5.605 46.555 -5.275 46.885 ;
        RECT -5.605 45.705 -5.275 46.035 ;
        RECT -5.605 43.395 -5.275 43.725 ;
        RECT -5.605 42.545 -5.275 42.875 ;
        RECT -5.605 40.235 -5.275 40.565 ;
        RECT -5.605 39.385 -5.275 39.715 ;
        RECT -5.605 37.075 -5.275 37.405 ;
        RECT -5.605 36.225 -5.275 36.555 ;
        RECT -5.605 33.915 -5.275 34.245 ;
        RECT -5.605 32.335 -5.275 32.665 ;
        RECT -5.605 31.485 -5.275 31.815 ;
        RECT -5.605 29.175 -5.275 29.505 ;
        RECT -5.605 28.325 -5.275 28.655 ;
        RECT -5.605 26.015 -5.275 26.345 ;
        RECT -5.605 25.165 -5.275 25.495 ;
        RECT -5.605 22.855 -5.275 23.185 ;
        RECT -5.605 22.005 -5.275 22.335 ;
        RECT -5.605 19.695 -5.275 20.025 ;
        RECT -5.605 18.115 -5.275 18.445 ;
        RECT -5.605 17.265 -5.275 17.595 ;
        RECT -5.605 14.955 -5.275 15.285 ;
        RECT -5.605 14.105 -5.275 14.435 ;
        RECT -5.605 11.795 -5.275 12.125 ;
        RECT -5.605 10.945 -5.275 11.275 ;
        RECT -5.605 8.635 -5.275 8.965 ;
        RECT -5.605 7.785 -5.275 8.115 ;
        RECT -5.605 5.475 -5.275 5.805 ;
        RECT -5.605 3.895 -5.275 4.225 ;
        RECT -5.605 3.045 -5.275 3.375 ;
        RECT -5.605 0.87 -5.275 1.2 ;
        RECT -5.605 -0.845 -5.275 -0.515 ;
        RECT -5.605 -2.205 -5.275 -1.875 ;
        RECT -5.605 -3.565 -5.275 -3.235 ;
        RECT -5.605 -4.925 -5.275 -4.595 ;
        RECT -5.605 -6.285 -5.275 -5.955 ;
        RECT -5.605 -7.645 -5.275 -7.315 ;
        RECT -5.605 -9.005 -5.275 -8.675 ;
        RECT -5.605 -10.365 -5.275 -10.035 ;
        RECT -5.605 -11.725 -5.275 -11.395 ;
        RECT -5.605 -13.085 -5.275 -12.755 ;
        RECT -5.605 -14.445 -5.275 -14.115 ;
        RECT -5.605 -15.805 -5.275 -15.475 ;
        RECT -5.605 -17.165 -5.275 -16.835 ;
        RECT -5.605 -23.965 -5.275 -23.635 ;
        RECT -5.605 -25.325 -5.275 -24.995 ;
        RECT -5.605 -26.685 -5.275 -26.355 ;
        RECT -5.605 -28.045 -5.275 -27.715 ;
        RECT -5.605 -29.405 -5.275 -29.075 ;
        RECT -5.605 -30.765 -5.275 -30.435 ;
        RECT -5.605 -32.125 -5.275 -31.795 ;
        RECT -5.605 -33.485 -5.275 -33.155 ;
        RECT -5.605 -37.565 -5.275 -37.235 ;
        RECT -5.605 -40.285 -5.275 -39.955 ;
        RECT -5.605 -41.645 -5.275 -41.315 ;
        RECT -5.605 -43.005 -5.275 -42.675 ;
        RECT -5.605 -44.365 -5.275 -44.035 ;
        RECT -5.605 -45.725 -5.275 -45.395 ;
        RECT -5.605 -47.085 -5.275 -46.755 ;
        RECT -5.605 -48.445 -5.275 -48.115 ;
        RECT -5.605 -52.525 -5.275 -52.195 ;
        RECT -5.605 -53.885 -5.275 -53.555 ;
        RECT -5.605 -55.245 -5.275 -54.915 ;
        RECT -5.605 -56.605 -5.275 -56.275 ;
        RECT -5.605 -57.965 -5.275 -57.635 ;
        RECT -5.605 -59.325 -5.275 -58.995 ;
        RECT -5.605 -60.685 -5.275 -60.355 ;
        RECT -5.605 -62.045 -5.275 -61.715 ;
        RECT -5.605 -63.405 -5.275 -63.075 ;
        RECT -5.605 -64.765 -5.275 -64.435 ;
        RECT -5.605 -66.125 -5.275 -65.795 ;
        RECT -5.605 -68.845 -5.275 -68.515 ;
        RECT -5.605 -70.205 -5.275 -69.875 ;
        RECT -5.605 -71.565 -5.275 -71.235 ;
        RECT -5.605 -72.925 -5.275 -72.595 ;
        RECT -5.605 -74.285 -5.275 -73.955 ;
        RECT -5.605 -75.645 -5.275 -75.315 ;
        RECT -5.605 -77.005 -5.275 -76.675 ;
        RECT -5.605 -78.365 -5.275 -78.035 ;
        RECT -5.605 -79.725 -5.275 -79.395 ;
        RECT -5.605 -81.085 -5.275 -80.755 ;
        RECT -5.605 -82.445 -5.275 -82.115 ;
        RECT -5.605 -83.805 -5.275 -83.475 ;
        RECT -5.605 -85.165 -5.275 -84.835 ;
        RECT -5.605 -86.525 -5.275 -86.195 ;
        RECT -5.605 -87.885 -5.275 -87.555 ;
        RECT -5.605 -89.245 -5.275 -88.915 ;
        RECT -5.605 -90.605 -5.275 -90.275 ;
        RECT -5.605 -91.965 -5.275 -91.635 ;
        RECT -5.605 -93.325 -5.275 -92.995 ;
        RECT -5.605 -94.685 -5.275 -94.355 ;
        RECT -5.605 -96.045 -5.275 -95.715 ;
        RECT -5.605 -97.405 -5.275 -97.075 ;
        RECT -5.605 -98.765 -5.275 -98.435 ;
        RECT -5.605 -100.125 -5.275 -99.795 ;
        RECT -5.605 -101.485 -5.275 -101.155 ;
        RECT -5.605 -102.845 -5.275 -102.515 ;
        RECT -5.605 -104.205 -5.275 -103.875 ;
        RECT -5.605 -105.565 -5.275 -105.235 ;
        RECT -5.605 -106.925 -5.275 -106.595 ;
        RECT -5.605 -108.285 -5.275 -107.955 ;
        RECT -5.605 -109.645 -5.275 -109.315 ;
        RECT -5.605 -111.005 -5.275 -110.675 ;
        RECT -5.605 -112.365 -5.275 -112.035 ;
        RECT -5.605 -113.725 -5.275 -113.395 ;
        RECT -5.605 -115.085 -5.275 -114.755 ;
        RECT -5.605 -116.445 -5.275 -116.115 ;
        RECT -5.605 -117.805 -5.275 -117.475 ;
        RECT -5.605 -119.165 -5.275 -118.835 ;
        RECT -5.605 -120.525 -5.275 -120.195 ;
        RECT -5.605 -121.885 -5.275 -121.555 ;
        RECT -5.605 -123.245 -5.275 -122.915 ;
        RECT -5.605 -124.605 -5.275 -124.275 ;
        RECT -5.605 -125.965 -5.275 -125.635 ;
        RECT -5.605 -127.325 -5.275 -126.995 ;
        RECT -5.605 -128.685 -5.275 -128.355 ;
        RECT -5.605 -130.045 -5.275 -129.715 ;
        RECT -5.605 -131.405 -5.275 -131.075 ;
        RECT -5.605 -132.765 -5.275 -132.435 ;
        RECT -5.605 -134.125 -5.275 -133.795 ;
        RECT -5.605 -135.485 -5.275 -135.155 ;
        RECT -5.605 -136.845 -5.275 -136.515 ;
        RECT -5.605 -138.205 -5.275 -137.875 ;
        RECT -5.605 -139.565 -5.275 -139.235 ;
        RECT -5.605 -140.925 -5.275 -140.595 ;
        RECT -5.605 -142.285 -5.275 -141.955 ;
        RECT -5.605 -143.645 -5.275 -143.315 ;
        RECT -5.605 -145.005 -5.275 -144.675 ;
        RECT -5.605 -146.365 -5.275 -146.035 ;
        RECT -5.605 -147.725 -5.275 -147.395 ;
        RECT -5.605 -149.085 -5.275 -148.755 ;
        RECT -5.605 -150.445 -5.275 -150.115 ;
        RECT -5.605 -151.805 -5.275 -151.475 ;
        RECT -5.605 -153.165 -5.275 -152.835 ;
        RECT -5.605 -154.525 -5.275 -154.195 ;
        RECT -5.605 -155.885 -5.275 -155.555 ;
        RECT -5.605 -157.245 -5.275 -156.915 ;
        RECT -5.605 -158.605 -5.275 -158.275 ;
        RECT -5.605 -159.965 -5.275 -159.635 ;
        RECT -5.605 -161.325 -5.275 -160.995 ;
        RECT -5.605 -162.685 -5.275 -162.355 ;
        RECT -5.605 -164.045 -5.275 -163.715 ;
        RECT -5.605 -165.405 -5.275 -165.075 ;
        RECT -5.605 -166.765 -5.275 -166.435 ;
        RECT -5.605 -168.125 -5.275 -167.795 ;
        RECT -5.605 -169.485 -5.275 -169.155 ;
        RECT -5.605 -170.845 -5.275 -170.515 ;
        RECT -5.605 -172.205 -5.275 -171.875 ;
        RECT -5.605 -173.565 -5.275 -173.235 ;
        RECT -5.605 -174.925 -5.275 -174.595 ;
        RECT -5.605 -176.285 -5.275 -175.955 ;
        RECT -5.605 -177.645 -5.275 -177.315 ;
        RECT -5.605 -179.005 -5.275 -178.675 ;
        RECT -5.605 -184.65 -5.275 -183.52 ;
        RECT -5.6 -184.765 -5.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.245 244.04 -3.915 245.17 ;
        RECT -4.245 239.875 -3.915 240.205 ;
        RECT -4.245 238.515 -3.915 238.845 ;
        RECT -4.245 237.155 -3.915 237.485 ;
        RECT -4.245 235.17 -3.915 235.5 ;
        RECT -4.245 232.995 -3.915 233.325 ;
        RECT -4.245 231.415 -3.915 231.745 ;
        RECT -4.245 230.565 -3.915 230.895 ;
        RECT -4.245 228.255 -3.915 228.585 ;
        RECT -4.245 227.405 -3.915 227.735 ;
        RECT -4.245 225.095 -3.915 225.425 ;
        RECT -4.245 224.245 -3.915 224.575 ;
        RECT -4.245 221.935 -3.915 222.265 ;
        RECT -4.245 221.085 -3.915 221.415 ;
        RECT -4.245 218.775 -3.915 219.105 ;
        RECT -4.245 217.195 -3.915 217.525 ;
        RECT -4.245 216.345 -3.915 216.675 ;
        RECT -4.245 214.035 -3.915 214.365 ;
        RECT -4.245 213.185 -3.915 213.515 ;
        RECT -4.245 210.875 -3.915 211.205 ;
        RECT -4.245 210.025 -3.915 210.355 ;
        RECT -4.245 207.715 -3.915 208.045 ;
        RECT -4.245 206.865 -3.915 207.195 ;
        RECT -4.245 204.555 -3.915 204.885 ;
        RECT -4.245 202.975 -3.915 203.305 ;
        RECT -4.245 202.125 -3.915 202.455 ;
        RECT -4.245 199.815 -3.915 200.145 ;
        RECT -4.245 198.965 -3.915 199.295 ;
        RECT -4.245 196.655 -3.915 196.985 ;
        RECT -4.245 195.805 -3.915 196.135 ;
        RECT -4.245 193.495 -3.915 193.825 ;
        RECT -4.245 192.645 -3.915 192.975 ;
        RECT -4.245 190.335 -3.915 190.665 ;
        RECT -4.245 188.755 -3.915 189.085 ;
        RECT -4.245 187.905 -3.915 188.235 ;
        RECT -4.245 185.595 -3.915 185.925 ;
        RECT -4.245 184.745 -3.915 185.075 ;
        RECT -4.245 182.435 -3.915 182.765 ;
        RECT -4.245 181.585 -3.915 181.915 ;
        RECT -4.245 179.275 -3.915 179.605 ;
        RECT -4.245 178.425 -3.915 178.755 ;
        RECT -4.245 176.115 -3.915 176.445 ;
        RECT -4.245 174.535 -3.915 174.865 ;
        RECT -4.245 173.685 -3.915 174.015 ;
        RECT -4.245 171.375 -3.915 171.705 ;
        RECT -4.245 170.525 -3.915 170.855 ;
        RECT -4.245 168.215 -3.915 168.545 ;
        RECT -4.245 167.365 -3.915 167.695 ;
        RECT -4.245 165.055 -3.915 165.385 ;
        RECT -4.245 164.205 -3.915 164.535 ;
        RECT -4.245 161.895 -3.915 162.225 ;
        RECT -4.245 160.315 -3.915 160.645 ;
        RECT -4.245 159.465 -3.915 159.795 ;
        RECT -4.245 157.155 -3.915 157.485 ;
        RECT -4.245 156.305 -3.915 156.635 ;
        RECT -4.245 153.995 -3.915 154.325 ;
        RECT -4.245 153.145 -3.915 153.475 ;
        RECT -4.245 150.835 -3.915 151.165 ;
        RECT -4.245 149.985 -3.915 150.315 ;
        RECT -4.245 147.675 -3.915 148.005 ;
        RECT -4.245 146.095 -3.915 146.425 ;
        RECT -4.245 145.245 -3.915 145.575 ;
        RECT -4.245 142.935 -3.915 143.265 ;
        RECT -4.245 142.085 -3.915 142.415 ;
        RECT -4.245 139.775 -3.915 140.105 ;
        RECT -4.245 138.925 -3.915 139.255 ;
        RECT -4.245 136.615 -3.915 136.945 ;
        RECT -4.245 135.765 -3.915 136.095 ;
        RECT -4.245 133.455 -3.915 133.785 ;
        RECT -4.245 131.875 -3.915 132.205 ;
        RECT -4.245 131.025 -3.915 131.355 ;
        RECT -4.245 128.715 -3.915 129.045 ;
        RECT -4.245 127.865 -3.915 128.195 ;
        RECT -4.245 125.555 -3.915 125.885 ;
        RECT -4.245 124.705 -3.915 125.035 ;
        RECT -4.245 122.395 -3.915 122.725 ;
        RECT -4.245 121.545 -3.915 121.875 ;
        RECT -4.245 119.235 -3.915 119.565 ;
        RECT -4.245 117.655 -3.915 117.985 ;
        RECT -4.245 116.805 -3.915 117.135 ;
        RECT -4.245 114.495 -3.915 114.825 ;
        RECT -4.245 113.645 -3.915 113.975 ;
        RECT -4.245 111.335 -3.915 111.665 ;
        RECT -4.245 110.485 -3.915 110.815 ;
        RECT -4.245 108.175 -3.915 108.505 ;
        RECT -4.245 107.325 -3.915 107.655 ;
        RECT -4.245 105.015 -3.915 105.345 ;
        RECT -4.245 103.435 -3.915 103.765 ;
        RECT -4.245 102.585 -3.915 102.915 ;
        RECT -4.245 100.275 -3.915 100.605 ;
        RECT -4.245 99.425 -3.915 99.755 ;
        RECT -4.245 97.115 -3.915 97.445 ;
        RECT -4.245 96.265 -3.915 96.595 ;
        RECT -4.245 93.955 -3.915 94.285 ;
        RECT -4.245 93.105 -3.915 93.435 ;
        RECT -4.245 90.795 -3.915 91.125 ;
        RECT -4.245 89.215 -3.915 89.545 ;
        RECT -4.245 88.365 -3.915 88.695 ;
        RECT -4.245 86.055 -3.915 86.385 ;
        RECT -4.245 85.205 -3.915 85.535 ;
        RECT -4.245 82.895 -3.915 83.225 ;
        RECT -4.245 82.045 -3.915 82.375 ;
        RECT -4.245 79.735 -3.915 80.065 ;
        RECT -4.245 78.885 -3.915 79.215 ;
        RECT -4.245 76.575 -3.915 76.905 ;
        RECT -4.245 74.995 -3.915 75.325 ;
        RECT -4.245 74.145 -3.915 74.475 ;
        RECT -4.245 71.835 -3.915 72.165 ;
        RECT -4.245 70.985 -3.915 71.315 ;
        RECT -4.245 68.675 -3.915 69.005 ;
        RECT -4.245 67.825 -3.915 68.155 ;
        RECT -4.245 65.515 -3.915 65.845 ;
        RECT -4.245 64.665 -3.915 64.995 ;
        RECT -4.245 62.355 -3.915 62.685 ;
        RECT -4.245 60.775 -3.915 61.105 ;
        RECT -4.245 59.925 -3.915 60.255 ;
        RECT -4.245 57.615 -3.915 57.945 ;
        RECT -4.245 56.765 -3.915 57.095 ;
        RECT -4.245 54.455 -3.915 54.785 ;
        RECT -4.245 53.605 -3.915 53.935 ;
        RECT -4.245 51.295 -3.915 51.625 ;
        RECT -4.245 50.445 -3.915 50.775 ;
        RECT -4.245 48.135 -3.915 48.465 ;
        RECT -4.245 46.555 -3.915 46.885 ;
        RECT -4.245 45.705 -3.915 46.035 ;
        RECT -4.245 43.395 -3.915 43.725 ;
        RECT -4.245 42.545 -3.915 42.875 ;
        RECT -4.245 40.235 -3.915 40.565 ;
        RECT -4.245 39.385 -3.915 39.715 ;
        RECT -4.245 37.075 -3.915 37.405 ;
        RECT -4.245 36.225 -3.915 36.555 ;
        RECT -4.245 33.915 -3.915 34.245 ;
        RECT -4.245 32.335 -3.915 32.665 ;
        RECT -4.245 31.485 -3.915 31.815 ;
        RECT -4.245 29.175 -3.915 29.505 ;
        RECT -4.245 28.325 -3.915 28.655 ;
        RECT -4.245 26.015 -3.915 26.345 ;
        RECT -4.245 25.165 -3.915 25.495 ;
        RECT -4.245 22.855 -3.915 23.185 ;
        RECT -4.245 22.005 -3.915 22.335 ;
        RECT -4.245 19.695 -3.915 20.025 ;
        RECT -4.245 18.115 -3.915 18.445 ;
        RECT -4.245 17.265 -3.915 17.595 ;
        RECT -4.245 14.955 -3.915 15.285 ;
        RECT -4.245 14.105 -3.915 14.435 ;
        RECT -4.245 11.795 -3.915 12.125 ;
        RECT -4.245 10.945 -3.915 11.275 ;
        RECT -4.245 8.635 -3.915 8.965 ;
        RECT -4.245 7.785 -3.915 8.115 ;
        RECT -4.245 5.475 -3.915 5.805 ;
        RECT -4.245 3.895 -3.915 4.225 ;
        RECT -4.245 3.045 -3.915 3.375 ;
        RECT -4.245 0.87 -3.915 1.2 ;
        RECT -4.245 -0.845 -3.915 -0.515 ;
        RECT -4.245 -2.205 -3.915 -1.875 ;
        RECT -4.245 -3.565 -3.915 -3.235 ;
        RECT -4.245 -4.925 -3.915 -4.595 ;
        RECT -4.245 -6.285 -3.915 -5.955 ;
        RECT -4.245 -7.645 -3.915 -7.315 ;
        RECT -4.245 -9.005 -3.915 -8.675 ;
        RECT -4.245 -10.365 -3.915 -10.035 ;
        RECT -4.245 -11.725 -3.915 -11.395 ;
        RECT -4.245 -13.085 -3.915 -12.755 ;
        RECT -4.245 -14.445 -3.915 -14.115 ;
        RECT -4.245 -15.805 -3.915 -15.475 ;
        RECT -4.245 -17.165 -3.915 -16.835 ;
        RECT -4.245 -23.965 -3.915 -23.635 ;
        RECT -4.245 -25.325 -3.915 -24.995 ;
        RECT -4.245 -26.685 -3.915 -26.355 ;
        RECT -4.245 -28.045 -3.915 -27.715 ;
        RECT -4.245 -29.405 -3.915 -29.075 ;
        RECT -4.245 -30.765 -3.915 -30.435 ;
        RECT -4.245 -32.125 -3.915 -31.795 ;
        RECT -4.245 -33.485 -3.915 -33.155 ;
        RECT -4.245 -37.565 -3.915 -37.235 ;
        RECT -4.245 -40.285 -3.915 -39.955 ;
        RECT -4.245 -41.645 -3.915 -41.315 ;
        RECT -4.245 -43.005 -3.915 -42.675 ;
        RECT -4.245 -44.365 -3.915 -44.035 ;
        RECT -4.245 -45.725 -3.915 -45.395 ;
        RECT -4.245 -47.085 -3.915 -46.755 ;
        RECT -4.245 -48.445 -3.915 -48.115 ;
        RECT -4.245 -52.525 -3.915 -52.195 ;
        RECT -4.245 -53.885 -3.915 -53.555 ;
        RECT -4.245 -55.245 -3.915 -54.915 ;
        RECT -4.245 -56.605 -3.915 -56.275 ;
        RECT -4.245 -57.965 -3.915 -57.635 ;
        RECT -4.245 -59.325 -3.915 -58.995 ;
        RECT -4.245 -60.685 -3.915 -60.355 ;
        RECT -4.245 -62.045 -3.915 -61.715 ;
        RECT -4.245 -63.405 -3.915 -63.075 ;
        RECT -4.245 -64.765 -3.915 -64.435 ;
        RECT -4.245 -66.125 -3.915 -65.795 ;
        RECT -4.245 -68.845 -3.915 -68.515 ;
        RECT -4.245 -70.205 -3.915 -69.875 ;
        RECT -4.245 -71.565 -3.915 -71.235 ;
        RECT -4.245 -72.925 -3.915 -72.595 ;
        RECT -4.245 -74.285 -3.915 -73.955 ;
        RECT -4.245 -75.645 -3.915 -75.315 ;
        RECT -4.245 -77.005 -3.915 -76.675 ;
        RECT -4.245 -78.365 -3.915 -78.035 ;
        RECT -4.245 -79.725 -3.915 -79.395 ;
        RECT -4.245 -81.085 -3.915 -80.755 ;
        RECT -4.245 -82.445 -3.915 -82.115 ;
        RECT -4.245 -83.805 -3.915 -83.475 ;
        RECT -4.245 -85.165 -3.915 -84.835 ;
        RECT -4.245 -86.525 -3.915 -86.195 ;
        RECT -4.245 -87.885 -3.915 -87.555 ;
        RECT -4.245 -89.245 -3.915 -88.915 ;
        RECT -4.245 -90.605 -3.915 -90.275 ;
        RECT -4.245 -91.965 -3.915 -91.635 ;
        RECT -4.245 -93.325 -3.915 -92.995 ;
        RECT -4.245 -94.685 -3.915 -94.355 ;
        RECT -4.245 -96.045 -3.915 -95.715 ;
        RECT -4.245 -97.405 -3.915 -97.075 ;
        RECT -4.245 -98.765 -3.915 -98.435 ;
        RECT -4.245 -100.125 -3.915 -99.795 ;
        RECT -4.245 -101.485 -3.915 -101.155 ;
        RECT -4.245 -102.845 -3.915 -102.515 ;
        RECT -4.245 -104.205 -3.915 -103.875 ;
        RECT -4.245 -105.565 -3.915 -105.235 ;
        RECT -4.245 -106.925 -3.915 -106.595 ;
        RECT -4.245 -108.285 -3.915 -107.955 ;
        RECT -4.245 -109.645 -3.915 -109.315 ;
        RECT -4.245 -111.005 -3.915 -110.675 ;
        RECT -4.245 -112.365 -3.915 -112.035 ;
        RECT -4.245 -113.725 -3.915 -113.395 ;
        RECT -4.245 -115.085 -3.915 -114.755 ;
        RECT -4.245 -116.445 -3.915 -116.115 ;
        RECT -4.245 -117.805 -3.915 -117.475 ;
        RECT -4.245 -119.165 -3.915 -118.835 ;
        RECT -4.245 -120.525 -3.915 -120.195 ;
        RECT -4.245 -121.885 -3.915 -121.555 ;
        RECT -4.245 -123.245 -3.915 -122.915 ;
        RECT -4.245 -124.605 -3.915 -124.275 ;
        RECT -4.245 -125.965 -3.915 -125.635 ;
        RECT -4.245 -127.325 -3.915 -126.995 ;
        RECT -4.245 -128.685 -3.915 -128.355 ;
        RECT -4.245 -130.045 -3.915 -129.715 ;
        RECT -4.245 -131.405 -3.915 -131.075 ;
        RECT -4.245 -132.765 -3.915 -132.435 ;
        RECT -4.245 -134.125 -3.915 -133.795 ;
        RECT -4.245 -135.485 -3.915 -135.155 ;
        RECT -4.245 -136.845 -3.915 -136.515 ;
        RECT -4.245 -138.205 -3.915 -137.875 ;
        RECT -4.245 -139.565 -3.915 -139.235 ;
        RECT -4.245 -140.925 -3.915 -140.595 ;
        RECT -4.245 -142.285 -3.915 -141.955 ;
        RECT -4.245 -143.645 -3.915 -143.315 ;
        RECT -4.245 -145.005 -3.915 -144.675 ;
        RECT -4.245 -146.365 -3.915 -146.035 ;
        RECT -4.245 -147.725 -3.915 -147.395 ;
        RECT -4.245 -149.085 -3.915 -148.755 ;
        RECT -4.245 -150.445 -3.915 -150.115 ;
        RECT -4.245 -151.805 -3.915 -151.475 ;
        RECT -4.245 -153.165 -3.915 -152.835 ;
        RECT -4.245 -154.525 -3.915 -154.195 ;
        RECT -4.245 -155.885 -3.915 -155.555 ;
        RECT -4.245 -157.245 -3.915 -156.915 ;
        RECT -4.245 -158.605 -3.915 -158.275 ;
        RECT -4.245 -159.965 -3.915 -159.635 ;
        RECT -4.245 -161.325 -3.915 -160.995 ;
        RECT -4.245 -162.685 -3.915 -162.355 ;
        RECT -4.245 -164.045 -3.915 -163.715 ;
        RECT -4.245 -165.405 -3.915 -165.075 ;
        RECT -4.245 -166.765 -3.915 -166.435 ;
        RECT -4.245 -168.125 -3.915 -167.795 ;
        RECT -4.245 -169.485 -3.915 -169.155 ;
        RECT -4.245 -170.845 -3.915 -170.515 ;
        RECT -4.245 -172.205 -3.915 -171.875 ;
        RECT -4.245 -173.565 -3.915 -173.235 ;
        RECT -4.245 -174.925 -3.915 -174.595 ;
        RECT -4.245 -176.285 -3.915 -175.955 ;
        RECT -4.245 -177.645 -3.915 -177.315 ;
        RECT -4.245 -179.005 -3.915 -178.675 ;
        RECT -4.245 -184.65 -3.915 -183.52 ;
        RECT -4.24 -184.765 -3.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.885 -176.285 -2.555 -175.955 ;
        RECT -2.885 -177.645 -2.555 -177.315 ;
        RECT -2.885 -179.005 -2.555 -178.675 ;
        RECT -2.885 -184.65 -2.555 -183.52 ;
        RECT -2.88 -184.765 -2.56 245.285 ;
        RECT -2.885 244.04 -2.555 245.17 ;
        RECT -2.885 239.875 -2.555 240.205 ;
        RECT -2.885 238.515 -2.555 238.845 ;
        RECT -2.885 237.155 -2.555 237.485 ;
        RECT -2.885 235.17 -2.555 235.5 ;
        RECT -2.885 232.995 -2.555 233.325 ;
        RECT -2.885 231.415 -2.555 231.745 ;
        RECT -2.885 230.565 -2.555 230.895 ;
        RECT -2.885 228.255 -2.555 228.585 ;
        RECT -2.885 227.405 -2.555 227.735 ;
        RECT -2.885 225.095 -2.555 225.425 ;
        RECT -2.885 224.245 -2.555 224.575 ;
        RECT -2.885 221.935 -2.555 222.265 ;
        RECT -2.885 221.085 -2.555 221.415 ;
        RECT -2.885 218.775 -2.555 219.105 ;
        RECT -2.885 217.195 -2.555 217.525 ;
        RECT -2.885 216.345 -2.555 216.675 ;
        RECT -2.885 214.035 -2.555 214.365 ;
        RECT -2.885 213.185 -2.555 213.515 ;
        RECT -2.885 210.875 -2.555 211.205 ;
        RECT -2.885 210.025 -2.555 210.355 ;
        RECT -2.885 207.715 -2.555 208.045 ;
        RECT -2.885 206.865 -2.555 207.195 ;
        RECT -2.885 204.555 -2.555 204.885 ;
        RECT -2.885 202.975 -2.555 203.305 ;
        RECT -2.885 202.125 -2.555 202.455 ;
        RECT -2.885 199.815 -2.555 200.145 ;
        RECT -2.885 198.965 -2.555 199.295 ;
        RECT -2.885 196.655 -2.555 196.985 ;
        RECT -2.885 195.805 -2.555 196.135 ;
        RECT -2.885 193.495 -2.555 193.825 ;
        RECT -2.885 192.645 -2.555 192.975 ;
        RECT -2.885 190.335 -2.555 190.665 ;
        RECT -2.885 188.755 -2.555 189.085 ;
        RECT -2.885 187.905 -2.555 188.235 ;
        RECT -2.885 185.595 -2.555 185.925 ;
        RECT -2.885 184.745 -2.555 185.075 ;
        RECT -2.885 182.435 -2.555 182.765 ;
        RECT -2.885 181.585 -2.555 181.915 ;
        RECT -2.885 179.275 -2.555 179.605 ;
        RECT -2.885 178.425 -2.555 178.755 ;
        RECT -2.885 176.115 -2.555 176.445 ;
        RECT -2.885 174.535 -2.555 174.865 ;
        RECT -2.885 173.685 -2.555 174.015 ;
        RECT -2.885 171.375 -2.555 171.705 ;
        RECT -2.885 170.525 -2.555 170.855 ;
        RECT -2.885 168.215 -2.555 168.545 ;
        RECT -2.885 167.365 -2.555 167.695 ;
        RECT -2.885 165.055 -2.555 165.385 ;
        RECT -2.885 164.205 -2.555 164.535 ;
        RECT -2.885 161.895 -2.555 162.225 ;
        RECT -2.885 160.315 -2.555 160.645 ;
        RECT -2.885 159.465 -2.555 159.795 ;
        RECT -2.885 157.155 -2.555 157.485 ;
        RECT -2.885 156.305 -2.555 156.635 ;
        RECT -2.885 153.995 -2.555 154.325 ;
        RECT -2.885 153.145 -2.555 153.475 ;
        RECT -2.885 150.835 -2.555 151.165 ;
        RECT -2.885 149.985 -2.555 150.315 ;
        RECT -2.885 147.675 -2.555 148.005 ;
        RECT -2.885 146.095 -2.555 146.425 ;
        RECT -2.885 145.245 -2.555 145.575 ;
        RECT -2.885 142.935 -2.555 143.265 ;
        RECT -2.885 142.085 -2.555 142.415 ;
        RECT -2.885 139.775 -2.555 140.105 ;
        RECT -2.885 138.925 -2.555 139.255 ;
        RECT -2.885 136.615 -2.555 136.945 ;
        RECT -2.885 135.765 -2.555 136.095 ;
        RECT -2.885 133.455 -2.555 133.785 ;
        RECT -2.885 131.875 -2.555 132.205 ;
        RECT -2.885 131.025 -2.555 131.355 ;
        RECT -2.885 128.715 -2.555 129.045 ;
        RECT -2.885 127.865 -2.555 128.195 ;
        RECT -2.885 125.555 -2.555 125.885 ;
        RECT -2.885 124.705 -2.555 125.035 ;
        RECT -2.885 122.395 -2.555 122.725 ;
        RECT -2.885 121.545 -2.555 121.875 ;
        RECT -2.885 119.235 -2.555 119.565 ;
        RECT -2.885 117.655 -2.555 117.985 ;
        RECT -2.885 116.805 -2.555 117.135 ;
        RECT -2.885 114.495 -2.555 114.825 ;
        RECT -2.885 113.645 -2.555 113.975 ;
        RECT -2.885 111.335 -2.555 111.665 ;
        RECT -2.885 110.485 -2.555 110.815 ;
        RECT -2.885 108.175 -2.555 108.505 ;
        RECT -2.885 107.325 -2.555 107.655 ;
        RECT -2.885 105.015 -2.555 105.345 ;
        RECT -2.885 103.435 -2.555 103.765 ;
        RECT -2.885 102.585 -2.555 102.915 ;
        RECT -2.885 100.275 -2.555 100.605 ;
        RECT -2.885 99.425 -2.555 99.755 ;
        RECT -2.885 97.115 -2.555 97.445 ;
        RECT -2.885 96.265 -2.555 96.595 ;
        RECT -2.885 93.955 -2.555 94.285 ;
        RECT -2.885 93.105 -2.555 93.435 ;
        RECT -2.885 90.795 -2.555 91.125 ;
        RECT -2.885 89.215 -2.555 89.545 ;
        RECT -2.885 88.365 -2.555 88.695 ;
        RECT -2.885 86.055 -2.555 86.385 ;
        RECT -2.885 85.205 -2.555 85.535 ;
        RECT -2.885 82.895 -2.555 83.225 ;
        RECT -2.885 82.045 -2.555 82.375 ;
        RECT -2.885 79.735 -2.555 80.065 ;
        RECT -2.885 78.885 -2.555 79.215 ;
        RECT -2.885 76.575 -2.555 76.905 ;
        RECT -2.885 74.995 -2.555 75.325 ;
        RECT -2.885 74.145 -2.555 74.475 ;
        RECT -2.885 71.835 -2.555 72.165 ;
        RECT -2.885 70.985 -2.555 71.315 ;
        RECT -2.885 68.675 -2.555 69.005 ;
        RECT -2.885 67.825 -2.555 68.155 ;
        RECT -2.885 65.515 -2.555 65.845 ;
        RECT -2.885 64.665 -2.555 64.995 ;
        RECT -2.885 62.355 -2.555 62.685 ;
        RECT -2.885 60.775 -2.555 61.105 ;
        RECT -2.885 59.925 -2.555 60.255 ;
        RECT -2.885 57.615 -2.555 57.945 ;
        RECT -2.885 56.765 -2.555 57.095 ;
        RECT -2.885 54.455 -2.555 54.785 ;
        RECT -2.885 53.605 -2.555 53.935 ;
        RECT -2.885 51.295 -2.555 51.625 ;
        RECT -2.885 50.445 -2.555 50.775 ;
        RECT -2.885 48.135 -2.555 48.465 ;
        RECT -2.885 46.555 -2.555 46.885 ;
        RECT -2.885 45.705 -2.555 46.035 ;
        RECT -2.885 43.395 -2.555 43.725 ;
        RECT -2.885 42.545 -2.555 42.875 ;
        RECT -2.885 40.235 -2.555 40.565 ;
        RECT -2.885 39.385 -2.555 39.715 ;
        RECT -2.885 37.075 -2.555 37.405 ;
        RECT -2.885 36.225 -2.555 36.555 ;
        RECT -2.885 33.915 -2.555 34.245 ;
        RECT -2.885 32.335 -2.555 32.665 ;
        RECT -2.885 31.485 -2.555 31.815 ;
        RECT -2.885 29.175 -2.555 29.505 ;
        RECT -2.885 28.325 -2.555 28.655 ;
        RECT -2.885 26.015 -2.555 26.345 ;
        RECT -2.885 25.165 -2.555 25.495 ;
        RECT -2.885 22.855 -2.555 23.185 ;
        RECT -2.885 22.005 -2.555 22.335 ;
        RECT -2.885 19.695 -2.555 20.025 ;
        RECT -2.885 18.115 -2.555 18.445 ;
        RECT -2.885 17.265 -2.555 17.595 ;
        RECT -2.885 14.955 -2.555 15.285 ;
        RECT -2.885 14.105 -2.555 14.435 ;
        RECT -2.885 11.795 -2.555 12.125 ;
        RECT -2.885 10.945 -2.555 11.275 ;
        RECT -2.885 8.635 -2.555 8.965 ;
        RECT -2.885 7.785 -2.555 8.115 ;
        RECT -2.885 5.475 -2.555 5.805 ;
        RECT -2.885 3.895 -2.555 4.225 ;
        RECT -2.885 3.045 -2.555 3.375 ;
        RECT -2.885 0.87 -2.555 1.2 ;
        RECT -2.885 -0.845 -2.555 -0.515 ;
        RECT -2.885 -2.205 -2.555 -1.875 ;
        RECT -2.885 -3.565 -2.555 -3.235 ;
        RECT -2.885 -4.925 -2.555 -4.595 ;
        RECT -2.885 -6.285 -2.555 -5.955 ;
        RECT -2.885 -7.645 -2.555 -7.315 ;
        RECT -2.885 -9.005 -2.555 -8.675 ;
        RECT -2.885 -10.365 -2.555 -10.035 ;
        RECT -2.885 -11.725 -2.555 -11.395 ;
        RECT -2.885 -13.085 -2.555 -12.755 ;
        RECT -2.885 -14.445 -2.555 -14.115 ;
        RECT -2.885 -15.805 -2.555 -15.475 ;
        RECT -2.885 -17.165 -2.555 -16.835 ;
        RECT -2.885 -23.965 -2.555 -23.635 ;
        RECT -2.885 -25.325 -2.555 -24.995 ;
        RECT -2.885 -26.685 -2.555 -26.355 ;
        RECT -2.885 -28.045 -2.555 -27.715 ;
        RECT -2.885 -29.405 -2.555 -29.075 ;
        RECT -2.885 -30.765 -2.555 -30.435 ;
        RECT -2.885 -32.125 -2.555 -31.795 ;
        RECT -2.885 -33.485 -2.555 -33.155 ;
        RECT -2.885 -37.565 -2.555 -37.235 ;
        RECT -2.885 -40.285 -2.555 -39.955 ;
        RECT -2.885 -41.645 -2.555 -41.315 ;
        RECT -2.885 -43.005 -2.555 -42.675 ;
        RECT -2.885 -44.365 -2.555 -44.035 ;
        RECT -2.885 -45.725 -2.555 -45.395 ;
        RECT -2.885 -47.085 -2.555 -46.755 ;
        RECT -2.885 -48.445 -2.555 -48.115 ;
        RECT -2.885 -52.525 -2.555 -52.195 ;
        RECT -2.885 -53.885 -2.555 -53.555 ;
        RECT -2.885 -55.245 -2.555 -54.915 ;
        RECT -2.885 -56.605 -2.555 -56.275 ;
        RECT -2.885 -57.965 -2.555 -57.635 ;
        RECT -2.885 -59.325 -2.555 -58.995 ;
        RECT -2.885 -60.685 -2.555 -60.355 ;
        RECT -2.885 -62.045 -2.555 -61.715 ;
        RECT -2.885 -63.405 -2.555 -63.075 ;
        RECT -2.885 -64.765 -2.555 -64.435 ;
        RECT -2.885 -66.125 -2.555 -65.795 ;
        RECT -2.885 -68.845 -2.555 -68.515 ;
        RECT -2.885 -70.205 -2.555 -69.875 ;
        RECT -2.885 -71.565 -2.555 -71.235 ;
        RECT -2.885 -72.925 -2.555 -72.595 ;
        RECT -2.885 -74.285 -2.555 -73.955 ;
        RECT -2.885 -75.645 -2.555 -75.315 ;
        RECT -2.885 -77.005 -2.555 -76.675 ;
        RECT -2.885 -78.365 -2.555 -78.035 ;
        RECT -2.885 -79.725 -2.555 -79.395 ;
        RECT -2.885 -81.085 -2.555 -80.755 ;
        RECT -2.885 -82.445 -2.555 -82.115 ;
        RECT -2.885 -83.805 -2.555 -83.475 ;
        RECT -2.885 -85.165 -2.555 -84.835 ;
        RECT -2.885 -86.525 -2.555 -86.195 ;
        RECT -2.885 -87.885 -2.555 -87.555 ;
        RECT -2.885 -89.245 -2.555 -88.915 ;
        RECT -2.885 -90.605 -2.555 -90.275 ;
        RECT -2.885 -91.965 -2.555 -91.635 ;
        RECT -2.885 -93.325 -2.555 -92.995 ;
        RECT -2.885 -94.685 -2.555 -94.355 ;
        RECT -2.885 -96.045 -2.555 -95.715 ;
        RECT -2.885 -97.405 -2.555 -97.075 ;
        RECT -2.885 -98.765 -2.555 -98.435 ;
        RECT -2.885 -100.125 -2.555 -99.795 ;
        RECT -2.885 -101.485 -2.555 -101.155 ;
        RECT -2.885 -102.845 -2.555 -102.515 ;
        RECT -2.885 -104.205 -2.555 -103.875 ;
        RECT -2.885 -105.565 -2.555 -105.235 ;
        RECT -2.885 -106.925 -2.555 -106.595 ;
        RECT -2.885 -108.285 -2.555 -107.955 ;
        RECT -2.885 -109.645 -2.555 -109.315 ;
        RECT -2.885 -111.005 -2.555 -110.675 ;
        RECT -2.885 -112.365 -2.555 -112.035 ;
        RECT -2.885 -113.725 -2.555 -113.395 ;
        RECT -2.885 -115.085 -2.555 -114.755 ;
        RECT -2.885 -116.445 -2.555 -116.115 ;
        RECT -2.885 -117.805 -2.555 -117.475 ;
        RECT -2.885 -119.165 -2.555 -118.835 ;
        RECT -2.885 -120.525 -2.555 -120.195 ;
        RECT -2.885 -121.885 -2.555 -121.555 ;
        RECT -2.885 -123.245 -2.555 -122.915 ;
        RECT -2.885 -124.605 -2.555 -124.275 ;
        RECT -2.885 -125.965 -2.555 -125.635 ;
        RECT -2.885 -127.325 -2.555 -126.995 ;
        RECT -2.885 -128.685 -2.555 -128.355 ;
        RECT -2.885 -130.045 -2.555 -129.715 ;
        RECT -2.885 -131.405 -2.555 -131.075 ;
        RECT -2.885 -132.765 -2.555 -132.435 ;
        RECT -2.885 -134.125 -2.555 -133.795 ;
        RECT -2.885 -135.485 -2.555 -135.155 ;
        RECT -2.885 -136.845 -2.555 -136.515 ;
        RECT -2.885 -138.205 -2.555 -137.875 ;
        RECT -2.885 -139.565 -2.555 -139.235 ;
        RECT -2.885 -140.925 -2.555 -140.595 ;
        RECT -2.885 -142.285 -2.555 -141.955 ;
        RECT -2.885 -143.645 -2.555 -143.315 ;
        RECT -2.885 -145.005 -2.555 -144.675 ;
        RECT -2.885 -146.365 -2.555 -146.035 ;
        RECT -2.885 -147.725 -2.555 -147.395 ;
        RECT -2.885 -149.085 -2.555 -148.755 ;
        RECT -2.885 -150.445 -2.555 -150.115 ;
        RECT -2.885 -151.805 -2.555 -151.475 ;
        RECT -2.885 -153.165 -2.555 -152.835 ;
        RECT -2.885 -154.525 -2.555 -154.195 ;
        RECT -2.885 -155.885 -2.555 -155.555 ;
        RECT -2.885 -157.245 -2.555 -156.915 ;
        RECT -2.885 -158.605 -2.555 -158.275 ;
        RECT -2.885 -159.965 -2.555 -159.635 ;
        RECT -2.885 -161.325 -2.555 -160.995 ;
        RECT -2.885 -162.685 -2.555 -162.355 ;
        RECT -2.885 -164.045 -2.555 -163.715 ;
        RECT -2.885 -165.405 -2.555 -165.075 ;
        RECT -2.885 -166.765 -2.555 -166.435 ;
        RECT -2.885 -168.125 -2.555 -167.795 ;
        RECT -2.885 -169.485 -2.555 -169.155 ;
        RECT -2.885 -170.845 -2.555 -170.515 ;
        RECT -2.885 -172.205 -2.555 -171.875 ;
        RECT -2.885 -173.565 -2.555 -173.235 ;
        RECT -2.885 -174.925 -2.555 -174.595 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 -26.685 -16.155 -26.355 ;
        RECT -16.485 -28.045 -16.155 -27.715 ;
        RECT -16.485 -29.405 -16.155 -29.075 ;
        RECT -16.485 -30.765 -16.155 -30.435 ;
        RECT -16.485 -32.125 -16.155 -31.795 ;
        RECT -16.485 -33.71 -16.155 -33.38 ;
        RECT -16.485 -36.205 -16.155 -35.875 ;
        RECT -16.485 -39.75 -16.155 -39.42 ;
        RECT -16.485 -41.645 -16.155 -41.315 ;
        RECT -16.48 -43 -16.16 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 -127.325 -16.155 -126.995 ;
        RECT -16.485 -139.565 -16.155 -139.235 ;
        RECT -16.485 -142.285 -16.155 -141.955 ;
        RECT -16.485 -153.165 -16.155 -152.835 ;
        RECT -16.485 -158.605 -16.155 -158.275 ;
        RECT -16.485 -159.965 -16.155 -159.635 ;
        RECT -16.485 -161.325 -16.155 -160.995 ;
        RECT -16.485 -162.685 -16.155 -162.355 ;
        RECT -16.485 -164.045 -16.155 -163.715 ;
        RECT -16.485 -165.405 -16.155 -165.075 ;
        RECT -16.485 -166.765 -16.155 -166.435 ;
        RECT -16.485 -170.845 -16.155 -170.515 ;
        RECT -16.485 -172.205 -16.155 -171.875 ;
        RECT -16.485 -174.925 -16.155 -174.595 ;
        RECT -16.485 -177.645 -16.155 -177.315 ;
        RECT -16.485 -179.005 -16.155 -178.675 ;
        RECT -16.485 -184.65 -16.155 -183.52 ;
        RECT -16.48 -184.765 -16.16 -122.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.125 244.04 -14.795 245.17 ;
        RECT -15.125 239.875 -14.795 240.205 ;
        RECT -15.125 238.515 -14.795 238.845 ;
        RECT -15.125 237.155 -14.795 237.485 ;
        RECT -15.125 235.795 -14.795 236.125 ;
        RECT -15.125 234.435 -14.795 234.765 ;
        RECT -15.125 233.075 -14.795 233.405 ;
        RECT -15.125 231.715 -14.795 232.045 ;
        RECT -15.125 230.355 -14.795 230.685 ;
        RECT -15.125 228.995 -14.795 229.325 ;
        RECT -15.125 227.635 -14.795 227.965 ;
        RECT -15.125 226.275 -14.795 226.605 ;
        RECT -15.125 224.915 -14.795 225.245 ;
        RECT -15.125 223.555 -14.795 223.885 ;
        RECT -15.125 222.195 -14.795 222.525 ;
        RECT -15.125 220.835 -14.795 221.165 ;
        RECT -15.125 219.475 -14.795 219.805 ;
        RECT -15.125 218.115 -14.795 218.445 ;
        RECT -15.125 216.755 -14.795 217.085 ;
        RECT -15.125 215.395 -14.795 215.725 ;
        RECT -15.125 214.035 -14.795 214.365 ;
        RECT -15.125 212.675 -14.795 213.005 ;
        RECT -15.125 211.315 -14.795 211.645 ;
        RECT -15.125 209.955 -14.795 210.285 ;
        RECT -15.125 208.595 -14.795 208.925 ;
        RECT -15.125 207.235 -14.795 207.565 ;
        RECT -15.125 205.875 -14.795 206.205 ;
        RECT -15.125 204.515 -14.795 204.845 ;
        RECT -15.125 203.155 -14.795 203.485 ;
        RECT -15.125 201.795 -14.795 202.125 ;
        RECT -15.125 200.435 -14.795 200.765 ;
        RECT -15.125 199.075 -14.795 199.405 ;
        RECT -15.125 197.715 -14.795 198.045 ;
        RECT -15.125 196.355 -14.795 196.685 ;
        RECT -15.125 194.995 -14.795 195.325 ;
        RECT -15.125 193.635 -14.795 193.965 ;
        RECT -15.125 192.275 -14.795 192.605 ;
        RECT -15.125 190.915 -14.795 191.245 ;
        RECT -15.125 189.555 -14.795 189.885 ;
        RECT -15.125 188.195 -14.795 188.525 ;
        RECT -15.125 186.835 -14.795 187.165 ;
        RECT -15.125 185.475 -14.795 185.805 ;
        RECT -15.125 184.115 -14.795 184.445 ;
        RECT -15.125 182.755 -14.795 183.085 ;
        RECT -15.125 181.395 -14.795 181.725 ;
        RECT -15.125 180.035 -14.795 180.365 ;
        RECT -15.125 178.675 -14.795 179.005 ;
        RECT -15.125 177.315 -14.795 177.645 ;
        RECT -15.125 175.955 -14.795 176.285 ;
        RECT -15.125 174.595 -14.795 174.925 ;
        RECT -15.125 173.235 -14.795 173.565 ;
        RECT -15.125 171.875 -14.795 172.205 ;
        RECT -15.125 170.515 -14.795 170.845 ;
        RECT -15.125 169.155 -14.795 169.485 ;
        RECT -15.125 167.795 -14.795 168.125 ;
        RECT -15.125 166.435 -14.795 166.765 ;
        RECT -15.125 165.075 -14.795 165.405 ;
        RECT -15.125 163.715 -14.795 164.045 ;
        RECT -15.125 162.355 -14.795 162.685 ;
        RECT -15.125 160.995 -14.795 161.325 ;
        RECT -15.125 159.635 -14.795 159.965 ;
        RECT -15.125 158.275 -14.795 158.605 ;
        RECT -15.125 156.915 -14.795 157.245 ;
        RECT -15.125 155.555 -14.795 155.885 ;
        RECT -15.125 154.195 -14.795 154.525 ;
        RECT -15.125 152.835 -14.795 153.165 ;
        RECT -15.125 151.475 -14.795 151.805 ;
        RECT -15.125 150.115 -14.795 150.445 ;
        RECT -15.125 148.755 -14.795 149.085 ;
        RECT -15.125 147.395 -14.795 147.725 ;
        RECT -15.125 146.035 -14.795 146.365 ;
        RECT -15.125 144.675 -14.795 145.005 ;
        RECT -15.125 143.315 -14.795 143.645 ;
        RECT -15.125 141.955 -14.795 142.285 ;
        RECT -15.125 140.595 -14.795 140.925 ;
        RECT -15.125 139.235 -14.795 139.565 ;
        RECT -15.125 137.875 -14.795 138.205 ;
        RECT -15.125 136.515 -14.795 136.845 ;
        RECT -15.125 135.155 -14.795 135.485 ;
        RECT -15.125 133.795 -14.795 134.125 ;
        RECT -15.125 132.435 -14.795 132.765 ;
        RECT -15.125 131.075 -14.795 131.405 ;
        RECT -15.125 129.715 -14.795 130.045 ;
        RECT -15.125 128.355 -14.795 128.685 ;
        RECT -15.125 126.995 -14.795 127.325 ;
        RECT -15.125 125.635 -14.795 125.965 ;
        RECT -15.125 124.275 -14.795 124.605 ;
        RECT -15.125 122.915 -14.795 123.245 ;
        RECT -15.125 121.555 -14.795 121.885 ;
        RECT -15.125 120.195 -14.795 120.525 ;
        RECT -15.125 118.835 -14.795 119.165 ;
        RECT -15.125 117.475 -14.795 117.805 ;
        RECT -15.125 116.115 -14.795 116.445 ;
        RECT -15.125 114.755 -14.795 115.085 ;
        RECT -15.125 113.395 -14.795 113.725 ;
        RECT -15.125 112.035 -14.795 112.365 ;
        RECT -15.125 110.675 -14.795 111.005 ;
        RECT -15.125 109.315 -14.795 109.645 ;
        RECT -15.125 107.955 -14.795 108.285 ;
        RECT -15.125 106.595 -14.795 106.925 ;
        RECT -15.125 105.235 -14.795 105.565 ;
        RECT -15.125 103.875 -14.795 104.205 ;
        RECT -15.125 102.515 -14.795 102.845 ;
        RECT -15.125 101.155 -14.795 101.485 ;
        RECT -15.125 99.795 -14.795 100.125 ;
        RECT -15.125 98.435 -14.795 98.765 ;
        RECT -15.125 97.075 -14.795 97.405 ;
        RECT -15.125 95.715 -14.795 96.045 ;
        RECT -15.125 94.355 -14.795 94.685 ;
        RECT -15.125 92.995 -14.795 93.325 ;
        RECT -15.125 91.635 -14.795 91.965 ;
        RECT -15.125 90.275 -14.795 90.605 ;
        RECT -15.125 88.915 -14.795 89.245 ;
        RECT -15.125 87.555 -14.795 87.885 ;
        RECT -15.125 86.195 -14.795 86.525 ;
        RECT -15.125 84.835 -14.795 85.165 ;
        RECT -15.125 83.475 -14.795 83.805 ;
        RECT -15.125 82.115 -14.795 82.445 ;
        RECT -15.125 80.755 -14.795 81.085 ;
        RECT -15.125 79.395 -14.795 79.725 ;
        RECT -15.125 78.035 -14.795 78.365 ;
        RECT -15.125 76.675 -14.795 77.005 ;
        RECT -15.125 75.315 -14.795 75.645 ;
        RECT -15.125 73.955 -14.795 74.285 ;
        RECT -15.125 72.595 -14.795 72.925 ;
        RECT -15.125 71.235 -14.795 71.565 ;
        RECT -15.125 69.875 -14.795 70.205 ;
        RECT -15.125 68.515 -14.795 68.845 ;
        RECT -15.125 67.155 -14.795 67.485 ;
        RECT -15.125 65.795 -14.795 66.125 ;
        RECT -15.125 64.435 -14.795 64.765 ;
        RECT -15.125 63.075 -14.795 63.405 ;
        RECT -15.125 61.715 -14.795 62.045 ;
        RECT -15.125 60.355 -14.795 60.685 ;
        RECT -15.125 58.995 -14.795 59.325 ;
        RECT -15.125 57.635 -14.795 57.965 ;
        RECT -15.125 56.275 -14.795 56.605 ;
        RECT -15.125 54.915 -14.795 55.245 ;
        RECT -15.125 53.555 -14.795 53.885 ;
        RECT -15.125 52.195 -14.795 52.525 ;
        RECT -15.125 50.835 -14.795 51.165 ;
        RECT -15.125 49.475 -14.795 49.805 ;
        RECT -15.125 48.115 -14.795 48.445 ;
        RECT -15.125 46.755 -14.795 47.085 ;
        RECT -15.125 45.395 -14.795 45.725 ;
        RECT -15.125 44.035 -14.795 44.365 ;
        RECT -15.125 42.675 -14.795 43.005 ;
        RECT -15.125 41.315 -14.795 41.645 ;
        RECT -15.125 39.955 -14.795 40.285 ;
        RECT -15.125 38.595 -14.795 38.925 ;
        RECT -15.125 37.235 -14.795 37.565 ;
        RECT -15.125 35.875 -14.795 36.205 ;
        RECT -15.125 34.515 -14.795 34.845 ;
        RECT -15.125 33.155 -14.795 33.485 ;
        RECT -15.125 31.795 -14.795 32.125 ;
        RECT -15.125 30.435 -14.795 30.765 ;
        RECT -15.125 29.075 -14.795 29.405 ;
        RECT -15.125 27.715 -14.795 28.045 ;
        RECT -15.125 26.355 -14.795 26.685 ;
        RECT -15.125 24.995 -14.795 25.325 ;
        RECT -15.125 23.635 -14.795 23.965 ;
        RECT -15.125 22.275 -14.795 22.605 ;
        RECT -15.125 20.915 -14.795 21.245 ;
        RECT -15.125 19.555 -14.795 19.885 ;
        RECT -15.125 18.195 -14.795 18.525 ;
        RECT -15.125 16.835 -14.795 17.165 ;
        RECT -15.125 15.475 -14.795 15.805 ;
        RECT -15.125 14.115 -14.795 14.445 ;
        RECT -15.125 12.755 -14.795 13.085 ;
        RECT -15.125 11.395 -14.795 11.725 ;
        RECT -15.125 10.035 -14.795 10.365 ;
        RECT -15.125 8.675 -14.795 9.005 ;
        RECT -15.125 7.315 -14.795 7.645 ;
        RECT -15.125 5.955 -14.795 6.285 ;
        RECT -15.125 4.595 -14.795 4.925 ;
        RECT -15.125 3.235 -14.795 3.565 ;
        RECT -15.125 1.875 -14.795 2.205 ;
        RECT -15.125 0.515 -14.795 0.845 ;
        RECT -15.125 -0.845 -14.795 -0.515 ;
        RECT -15.125 -2.205 -14.795 -1.875 ;
        RECT -15.125 -3.565 -14.795 -3.235 ;
        RECT -15.125 -4.925 -14.795 -4.595 ;
        RECT -15.125 -7.645 -14.795 -7.315 ;
        RECT -15.125 -9.005 -14.795 -8.675 ;
        RECT -15.125 -10.73 -14.795 -10.4 ;
        RECT -15.125 -11.725 -14.795 -11.395 ;
        RECT -15.125 -13.085 -14.795 -12.755 ;
        RECT -15.125 -16.77 -14.795 -16.44 ;
        RECT -15.125 -18.525 -14.795 -18.195 ;
        RECT -15.12 -19.88 -14.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.125 -105.565 -14.795 -105.235 ;
        RECT -15.125 -113.725 -14.795 -113.395 ;
        RECT -15.125 -115.085 -14.795 -114.755 ;
        RECT -15.125 -116.445 -14.795 -116.115 ;
        RECT -15.125 -117.805 -14.795 -117.475 ;
        RECT -15.125 -119.165 -14.795 -118.835 ;
        RECT -15.125 -120.525 -14.795 -120.195 ;
        RECT -15.125 -128.685 -14.795 -128.355 ;
        RECT -15.125 -134.125 -14.795 -133.795 ;
        RECT -15.125 -135.485 -14.795 -135.155 ;
        RECT -15.125 -136.845 -14.795 -136.515 ;
        RECT -15.125 -139.565 -14.795 -139.235 ;
        RECT -15.125 -142.285 -14.795 -141.955 ;
        RECT -15.125 -147.725 -14.795 -147.395 ;
        RECT -15.125 -151.805 -14.795 -151.475 ;
        RECT -15.125 -153.165 -14.795 -152.835 ;
        RECT -15.125 -155.885 -14.795 -155.555 ;
        RECT -15.125 -158.605 -14.795 -158.275 ;
        RECT -15.125 -159.965 -14.795 -159.635 ;
        RECT -15.125 -161.325 -14.795 -160.995 ;
        RECT -15.125 -162.685 -14.795 -162.355 ;
        RECT -15.125 -164.045 -14.795 -163.715 ;
        RECT -15.125 -165.405 -14.795 -165.075 ;
        RECT -15.125 -166.765 -14.795 -166.435 ;
        RECT -15.125 -169.615 -14.795 -169.285 ;
        RECT -15.125 -170.845 -14.795 -170.515 ;
        RECT -15.125 -172.205 -14.795 -171.875 ;
        RECT -15.12 -172.88 -14.8 -105.235 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.765 244.04 -13.435 245.17 ;
        RECT -13.765 239.875 -13.435 240.205 ;
        RECT -13.765 238.515 -13.435 238.845 ;
        RECT -13.765 237.155 -13.435 237.485 ;
        RECT -13.765 235.795 -13.435 236.125 ;
        RECT -13.765 234.435 -13.435 234.765 ;
        RECT -13.765 233.075 -13.435 233.405 ;
        RECT -13.765 231.715 -13.435 232.045 ;
        RECT -13.765 230.355 -13.435 230.685 ;
        RECT -13.765 228.995 -13.435 229.325 ;
        RECT -13.765 227.635 -13.435 227.965 ;
        RECT -13.765 226.275 -13.435 226.605 ;
        RECT -13.765 224.915 -13.435 225.245 ;
        RECT -13.765 223.555 -13.435 223.885 ;
        RECT -13.765 222.195 -13.435 222.525 ;
        RECT -13.765 220.835 -13.435 221.165 ;
        RECT -13.765 219.475 -13.435 219.805 ;
        RECT -13.765 218.115 -13.435 218.445 ;
        RECT -13.765 216.755 -13.435 217.085 ;
        RECT -13.765 215.395 -13.435 215.725 ;
        RECT -13.765 214.035 -13.435 214.365 ;
        RECT -13.765 212.675 -13.435 213.005 ;
        RECT -13.765 211.315 -13.435 211.645 ;
        RECT -13.765 209.955 -13.435 210.285 ;
        RECT -13.765 208.595 -13.435 208.925 ;
        RECT -13.765 207.235 -13.435 207.565 ;
        RECT -13.765 205.875 -13.435 206.205 ;
        RECT -13.765 204.515 -13.435 204.845 ;
        RECT -13.765 203.155 -13.435 203.485 ;
        RECT -13.765 201.795 -13.435 202.125 ;
        RECT -13.765 200.435 -13.435 200.765 ;
        RECT -13.765 199.075 -13.435 199.405 ;
        RECT -13.765 197.715 -13.435 198.045 ;
        RECT -13.765 196.355 -13.435 196.685 ;
        RECT -13.765 194.995 -13.435 195.325 ;
        RECT -13.765 193.635 -13.435 193.965 ;
        RECT -13.765 192.275 -13.435 192.605 ;
        RECT -13.765 190.915 -13.435 191.245 ;
        RECT -13.765 189.555 -13.435 189.885 ;
        RECT -13.765 188.195 -13.435 188.525 ;
        RECT -13.765 186.835 -13.435 187.165 ;
        RECT -13.765 185.475 -13.435 185.805 ;
        RECT -13.765 184.115 -13.435 184.445 ;
        RECT -13.765 182.755 -13.435 183.085 ;
        RECT -13.765 181.395 -13.435 181.725 ;
        RECT -13.765 180.035 -13.435 180.365 ;
        RECT -13.765 178.675 -13.435 179.005 ;
        RECT -13.765 177.315 -13.435 177.645 ;
        RECT -13.765 175.955 -13.435 176.285 ;
        RECT -13.765 174.595 -13.435 174.925 ;
        RECT -13.765 173.235 -13.435 173.565 ;
        RECT -13.765 171.875 -13.435 172.205 ;
        RECT -13.765 170.515 -13.435 170.845 ;
        RECT -13.765 169.155 -13.435 169.485 ;
        RECT -13.765 167.795 -13.435 168.125 ;
        RECT -13.765 166.435 -13.435 166.765 ;
        RECT -13.765 165.075 -13.435 165.405 ;
        RECT -13.765 163.715 -13.435 164.045 ;
        RECT -13.765 162.355 -13.435 162.685 ;
        RECT -13.765 160.995 -13.435 161.325 ;
        RECT -13.765 159.635 -13.435 159.965 ;
        RECT -13.765 158.275 -13.435 158.605 ;
        RECT -13.765 156.915 -13.435 157.245 ;
        RECT -13.765 155.555 -13.435 155.885 ;
        RECT -13.765 154.195 -13.435 154.525 ;
        RECT -13.765 152.835 -13.435 153.165 ;
        RECT -13.765 151.475 -13.435 151.805 ;
        RECT -13.765 150.115 -13.435 150.445 ;
        RECT -13.765 148.755 -13.435 149.085 ;
        RECT -13.765 147.395 -13.435 147.725 ;
        RECT -13.765 146.035 -13.435 146.365 ;
        RECT -13.765 144.675 -13.435 145.005 ;
        RECT -13.765 143.315 -13.435 143.645 ;
        RECT -13.765 141.955 -13.435 142.285 ;
        RECT -13.765 140.595 -13.435 140.925 ;
        RECT -13.765 139.235 -13.435 139.565 ;
        RECT -13.765 137.875 -13.435 138.205 ;
        RECT -13.765 136.515 -13.435 136.845 ;
        RECT -13.765 135.155 -13.435 135.485 ;
        RECT -13.765 133.795 -13.435 134.125 ;
        RECT -13.765 132.435 -13.435 132.765 ;
        RECT -13.765 131.075 -13.435 131.405 ;
        RECT -13.765 129.715 -13.435 130.045 ;
        RECT -13.765 128.355 -13.435 128.685 ;
        RECT -13.765 126.995 -13.435 127.325 ;
        RECT -13.765 125.635 -13.435 125.965 ;
        RECT -13.765 124.275 -13.435 124.605 ;
        RECT -13.765 122.915 -13.435 123.245 ;
        RECT -13.765 121.555 -13.435 121.885 ;
        RECT -13.765 120.195 -13.435 120.525 ;
        RECT -13.765 118.835 -13.435 119.165 ;
        RECT -13.765 117.475 -13.435 117.805 ;
        RECT -13.765 116.115 -13.435 116.445 ;
        RECT -13.765 114.755 -13.435 115.085 ;
        RECT -13.765 113.395 -13.435 113.725 ;
        RECT -13.765 112.035 -13.435 112.365 ;
        RECT -13.765 110.675 -13.435 111.005 ;
        RECT -13.765 109.315 -13.435 109.645 ;
        RECT -13.765 107.955 -13.435 108.285 ;
        RECT -13.765 106.595 -13.435 106.925 ;
        RECT -13.765 105.235 -13.435 105.565 ;
        RECT -13.765 103.875 -13.435 104.205 ;
        RECT -13.765 102.515 -13.435 102.845 ;
        RECT -13.765 101.155 -13.435 101.485 ;
        RECT -13.765 99.795 -13.435 100.125 ;
        RECT -13.765 98.435 -13.435 98.765 ;
        RECT -13.765 97.075 -13.435 97.405 ;
        RECT -13.765 95.715 -13.435 96.045 ;
        RECT -13.765 94.355 -13.435 94.685 ;
        RECT -13.765 92.995 -13.435 93.325 ;
        RECT -13.765 91.635 -13.435 91.965 ;
        RECT -13.765 90.275 -13.435 90.605 ;
        RECT -13.765 88.915 -13.435 89.245 ;
        RECT -13.765 87.555 -13.435 87.885 ;
        RECT -13.765 86.195 -13.435 86.525 ;
        RECT -13.765 84.835 -13.435 85.165 ;
        RECT -13.765 83.475 -13.435 83.805 ;
        RECT -13.765 82.115 -13.435 82.445 ;
        RECT -13.765 80.755 -13.435 81.085 ;
        RECT -13.765 79.395 -13.435 79.725 ;
        RECT -13.765 78.035 -13.435 78.365 ;
        RECT -13.765 76.675 -13.435 77.005 ;
        RECT -13.765 75.315 -13.435 75.645 ;
        RECT -13.765 73.955 -13.435 74.285 ;
        RECT -13.765 72.595 -13.435 72.925 ;
        RECT -13.765 71.235 -13.435 71.565 ;
        RECT -13.765 69.875 -13.435 70.205 ;
        RECT -13.765 68.515 -13.435 68.845 ;
        RECT -13.765 67.155 -13.435 67.485 ;
        RECT -13.765 65.795 -13.435 66.125 ;
        RECT -13.765 64.435 -13.435 64.765 ;
        RECT -13.765 63.075 -13.435 63.405 ;
        RECT -13.765 61.715 -13.435 62.045 ;
        RECT -13.765 60.355 -13.435 60.685 ;
        RECT -13.765 58.995 -13.435 59.325 ;
        RECT -13.765 57.635 -13.435 57.965 ;
        RECT -13.765 56.275 -13.435 56.605 ;
        RECT -13.765 54.915 -13.435 55.245 ;
        RECT -13.765 53.555 -13.435 53.885 ;
        RECT -13.765 52.195 -13.435 52.525 ;
        RECT -13.765 50.835 -13.435 51.165 ;
        RECT -13.765 49.475 -13.435 49.805 ;
        RECT -13.765 48.115 -13.435 48.445 ;
        RECT -13.765 46.755 -13.435 47.085 ;
        RECT -13.765 45.395 -13.435 45.725 ;
        RECT -13.765 44.035 -13.435 44.365 ;
        RECT -13.765 42.675 -13.435 43.005 ;
        RECT -13.765 41.315 -13.435 41.645 ;
        RECT -13.765 39.955 -13.435 40.285 ;
        RECT -13.765 38.595 -13.435 38.925 ;
        RECT -13.765 37.235 -13.435 37.565 ;
        RECT -13.765 35.875 -13.435 36.205 ;
        RECT -13.765 34.515 -13.435 34.845 ;
        RECT -13.765 33.155 -13.435 33.485 ;
        RECT -13.765 31.795 -13.435 32.125 ;
        RECT -13.765 30.435 -13.435 30.765 ;
        RECT -13.765 29.075 -13.435 29.405 ;
        RECT -13.765 27.715 -13.435 28.045 ;
        RECT -13.765 26.355 -13.435 26.685 ;
        RECT -13.765 24.995 -13.435 25.325 ;
        RECT -13.765 23.635 -13.435 23.965 ;
        RECT -13.765 22.275 -13.435 22.605 ;
        RECT -13.765 20.915 -13.435 21.245 ;
        RECT -13.765 19.555 -13.435 19.885 ;
        RECT -13.765 18.195 -13.435 18.525 ;
        RECT -13.765 16.835 -13.435 17.165 ;
        RECT -13.765 15.475 -13.435 15.805 ;
        RECT -13.765 14.115 -13.435 14.445 ;
        RECT -13.765 12.755 -13.435 13.085 ;
        RECT -13.765 11.395 -13.435 11.725 ;
        RECT -13.765 10.035 -13.435 10.365 ;
        RECT -13.765 8.675 -13.435 9.005 ;
        RECT -13.765 7.315 -13.435 7.645 ;
        RECT -13.765 5.955 -13.435 6.285 ;
        RECT -13.765 4.595 -13.435 4.925 ;
        RECT -13.765 3.235 -13.435 3.565 ;
        RECT -13.765 1.875 -13.435 2.205 ;
        RECT -13.765 0.515 -13.435 0.845 ;
        RECT -13.765 -0.845 -13.435 -0.515 ;
        RECT -13.765 -2.205 -13.435 -1.875 ;
        RECT -13.765 -3.565 -13.435 -3.235 ;
        RECT -13.765 -4.925 -13.435 -4.595 ;
        RECT -13.765 -7.645 -13.435 -7.315 ;
        RECT -13.765 -9.005 -13.435 -8.675 ;
        RECT -13.765 -10.73 -13.435 -10.4 ;
        RECT -13.765 -11.725 -13.435 -11.395 ;
        RECT -13.765 -13.085 -13.435 -12.755 ;
        RECT -13.765 -16.77 -13.435 -16.44 ;
        RECT -13.765 -18.525 -13.435 -18.195 ;
        RECT -13.765 -26.685 -13.435 -26.355 ;
        RECT -13.765 -28.045 -13.435 -27.715 ;
        RECT -13.765 -29.405 -13.435 -29.075 ;
        RECT -13.765 -30.765 -13.435 -30.435 ;
        RECT -13.765 -32.125 -13.435 -31.795 ;
        RECT -13.765 -33.71 -13.435 -33.38 ;
        RECT -13.765 -36.205 -13.435 -35.875 ;
        RECT -13.765 -39.75 -13.435 -39.42 ;
        RECT -13.765 -41.645 -13.435 -41.315 ;
        RECT -13.765 -44.365 -13.435 -44.035 ;
        RECT -13.765 -51.165 -13.435 -50.835 ;
        RECT -13.765 -52.525 -13.435 -52.195 ;
        RECT -13.765 -53.885 -13.435 -53.555 ;
        RECT -13.765 -55.245 -13.435 -54.915 ;
        RECT -13.765 -56.605 -13.435 -56.275 ;
        RECT -13.765 -57.965 -13.435 -57.635 ;
        RECT -13.765 -59.325 -13.435 -58.995 ;
        RECT -13.765 -60.685 -13.435 -60.355 ;
        RECT -13.765 -62.045 -13.435 -61.715 ;
        RECT -13.765 -63.405 -13.435 -63.075 ;
        RECT -13.765 -64.765 -13.435 -64.435 ;
        RECT -13.765 -66.125 -13.435 -65.795 ;
        RECT -13.765 -68.845 -13.435 -68.515 ;
        RECT -13.765 -70.205 -13.435 -69.875 ;
        RECT -13.765 -71.565 -13.435 -71.235 ;
        RECT -13.765 -73.19 -13.435 -72.86 ;
        RECT -13.765 -74.285 -13.435 -73.955 ;
        RECT -13.765 -75.645 -13.435 -75.315 ;
        RECT -13.765 -78.365 -13.435 -78.035 ;
        RECT -13.765 -79.725 -13.435 -79.395 ;
        RECT -13.765 -80.73 -13.435 -80.4 ;
        RECT -13.765 -82.445 -13.435 -82.115 ;
        RECT -13.765 -83.805 -13.435 -83.475 ;
        RECT -13.765 -86.525 -13.435 -86.195 ;
        RECT -13.765 -89.245 -13.435 -88.915 ;
        RECT -13.765 -90.605 -13.435 -90.275 ;
        RECT -13.765 -91.965 -13.435 -91.635 ;
        RECT -13.765 -93.325 -13.435 -92.995 ;
        RECT -13.765 -94.685 -13.435 -94.355 ;
        RECT -13.765 -95.37 -13.435 -95.04 ;
        RECT -13.765 -97.405 -13.435 -97.075 ;
        RECT -13.765 -100.125 -13.435 -99.795 ;
        RECT -13.765 -101.485 -13.435 -101.155 ;
        RECT -13.765 -102.91 -13.435 -102.58 ;
        RECT -13.765 -113.725 -13.435 -113.395 ;
        RECT -13.765 -115.085 -13.435 -114.755 ;
        RECT -13.765 -116.445 -13.435 -116.115 ;
        RECT -13.765 -117.805 -13.435 -117.475 ;
        RECT -13.765 -119.165 -13.435 -118.835 ;
        RECT -13.765 -120.525 -13.435 -120.195 ;
        RECT -13.765 -121.885 -13.435 -121.555 ;
        RECT -13.765 -130.045 -13.435 -129.715 ;
        RECT -13.765 -134.125 -13.435 -133.795 ;
        RECT -13.765 -135.485 -13.435 -135.155 ;
        RECT -13.765 -136.845 -13.435 -136.515 ;
        RECT -13.765 -142.285 -13.435 -141.955 ;
        RECT -13.765 -147.725 -13.435 -147.395 ;
        RECT -13.765 -150.445 -13.435 -150.115 ;
        RECT -13.765 -151.805 -13.435 -151.475 ;
        RECT -13.765 -153.165 -13.435 -152.835 ;
        RECT -13.765 -155.885 -13.435 -155.555 ;
        RECT -13.765 -159.965 -13.435 -159.635 ;
        RECT -13.765 -161.325 -13.435 -160.995 ;
        RECT -13.765 -162.685 -13.435 -162.355 ;
        RECT -13.765 -164.045 -13.435 -163.715 ;
        RECT -13.765 -165.405 -13.435 -165.075 ;
        RECT -13.765 -166.765 -13.435 -166.435 ;
        RECT -13.765 -169.615 -13.435 -169.285 ;
        RECT -13.765 -170.845 -13.435 -170.515 ;
        RECT -13.765 -172.205 -13.435 -171.875 ;
        RECT -13.765 -174.925 -13.435 -174.595 ;
        RECT -13.765 -177.645 -13.435 -177.315 ;
        RECT -13.765 -179.005 -13.435 -178.675 ;
        RECT -13.765 -184.65 -13.435 -183.52 ;
        RECT -13.76 -184.765 -13.44 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.405 244.04 -12.075 245.17 ;
        RECT -12.405 239.875 -12.075 240.205 ;
        RECT -12.405 238.515 -12.075 238.845 ;
        RECT -12.405 237.155 -12.075 237.485 ;
        RECT -12.405 235.795 -12.075 236.125 ;
        RECT -12.405 234.435 -12.075 234.765 ;
        RECT -12.405 233.075 -12.075 233.405 ;
        RECT -12.405 231.715 -12.075 232.045 ;
        RECT -12.405 230.355 -12.075 230.685 ;
        RECT -12.405 228.995 -12.075 229.325 ;
        RECT -12.405 227.635 -12.075 227.965 ;
        RECT -12.405 226.275 -12.075 226.605 ;
        RECT -12.405 224.915 -12.075 225.245 ;
        RECT -12.405 223.555 -12.075 223.885 ;
        RECT -12.405 222.195 -12.075 222.525 ;
        RECT -12.405 220.835 -12.075 221.165 ;
        RECT -12.405 219.475 -12.075 219.805 ;
        RECT -12.405 218.115 -12.075 218.445 ;
        RECT -12.405 216.755 -12.075 217.085 ;
        RECT -12.405 215.395 -12.075 215.725 ;
        RECT -12.405 214.035 -12.075 214.365 ;
        RECT -12.405 212.675 -12.075 213.005 ;
        RECT -12.405 211.315 -12.075 211.645 ;
        RECT -12.405 209.955 -12.075 210.285 ;
        RECT -12.405 208.595 -12.075 208.925 ;
        RECT -12.405 207.235 -12.075 207.565 ;
        RECT -12.405 205.875 -12.075 206.205 ;
        RECT -12.405 204.515 -12.075 204.845 ;
        RECT -12.405 203.155 -12.075 203.485 ;
        RECT -12.405 201.795 -12.075 202.125 ;
        RECT -12.405 200.435 -12.075 200.765 ;
        RECT -12.405 199.075 -12.075 199.405 ;
        RECT -12.405 197.715 -12.075 198.045 ;
        RECT -12.405 196.355 -12.075 196.685 ;
        RECT -12.405 194.995 -12.075 195.325 ;
        RECT -12.405 193.635 -12.075 193.965 ;
        RECT -12.405 192.275 -12.075 192.605 ;
        RECT -12.405 190.915 -12.075 191.245 ;
        RECT -12.405 189.555 -12.075 189.885 ;
        RECT -12.405 188.195 -12.075 188.525 ;
        RECT -12.405 186.835 -12.075 187.165 ;
        RECT -12.405 185.475 -12.075 185.805 ;
        RECT -12.405 184.115 -12.075 184.445 ;
        RECT -12.405 182.755 -12.075 183.085 ;
        RECT -12.405 181.395 -12.075 181.725 ;
        RECT -12.405 180.035 -12.075 180.365 ;
        RECT -12.405 178.675 -12.075 179.005 ;
        RECT -12.405 177.315 -12.075 177.645 ;
        RECT -12.405 175.955 -12.075 176.285 ;
        RECT -12.405 174.595 -12.075 174.925 ;
        RECT -12.405 173.235 -12.075 173.565 ;
        RECT -12.405 171.875 -12.075 172.205 ;
        RECT -12.405 170.515 -12.075 170.845 ;
        RECT -12.405 169.155 -12.075 169.485 ;
        RECT -12.405 167.795 -12.075 168.125 ;
        RECT -12.405 166.435 -12.075 166.765 ;
        RECT -12.405 165.075 -12.075 165.405 ;
        RECT -12.405 163.715 -12.075 164.045 ;
        RECT -12.405 162.355 -12.075 162.685 ;
        RECT -12.405 160.995 -12.075 161.325 ;
        RECT -12.405 159.635 -12.075 159.965 ;
        RECT -12.405 158.275 -12.075 158.605 ;
        RECT -12.405 156.915 -12.075 157.245 ;
        RECT -12.405 155.555 -12.075 155.885 ;
        RECT -12.405 154.195 -12.075 154.525 ;
        RECT -12.405 152.835 -12.075 153.165 ;
        RECT -12.405 151.475 -12.075 151.805 ;
        RECT -12.405 150.115 -12.075 150.445 ;
        RECT -12.405 148.755 -12.075 149.085 ;
        RECT -12.405 147.395 -12.075 147.725 ;
        RECT -12.405 146.035 -12.075 146.365 ;
        RECT -12.405 144.675 -12.075 145.005 ;
        RECT -12.405 143.315 -12.075 143.645 ;
        RECT -12.405 141.955 -12.075 142.285 ;
        RECT -12.405 140.595 -12.075 140.925 ;
        RECT -12.405 139.235 -12.075 139.565 ;
        RECT -12.405 137.875 -12.075 138.205 ;
        RECT -12.405 136.515 -12.075 136.845 ;
        RECT -12.405 135.155 -12.075 135.485 ;
        RECT -12.405 133.795 -12.075 134.125 ;
        RECT -12.405 132.435 -12.075 132.765 ;
        RECT -12.405 131.075 -12.075 131.405 ;
        RECT -12.405 129.715 -12.075 130.045 ;
        RECT -12.405 128.355 -12.075 128.685 ;
        RECT -12.405 126.995 -12.075 127.325 ;
        RECT -12.405 125.635 -12.075 125.965 ;
        RECT -12.405 124.275 -12.075 124.605 ;
        RECT -12.405 122.915 -12.075 123.245 ;
        RECT -12.405 121.555 -12.075 121.885 ;
        RECT -12.405 120.195 -12.075 120.525 ;
        RECT -12.405 118.835 -12.075 119.165 ;
        RECT -12.405 117.475 -12.075 117.805 ;
        RECT -12.405 116.115 -12.075 116.445 ;
        RECT -12.405 114.755 -12.075 115.085 ;
        RECT -12.405 113.395 -12.075 113.725 ;
        RECT -12.405 112.035 -12.075 112.365 ;
        RECT -12.405 110.675 -12.075 111.005 ;
        RECT -12.405 109.315 -12.075 109.645 ;
        RECT -12.405 107.955 -12.075 108.285 ;
        RECT -12.405 106.595 -12.075 106.925 ;
        RECT -12.405 105.235 -12.075 105.565 ;
        RECT -12.405 103.875 -12.075 104.205 ;
        RECT -12.405 102.515 -12.075 102.845 ;
        RECT -12.405 101.155 -12.075 101.485 ;
        RECT -12.405 99.795 -12.075 100.125 ;
        RECT -12.405 98.435 -12.075 98.765 ;
        RECT -12.405 97.075 -12.075 97.405 ;
        RECT -12.405 95.715 -12.075 96.045 ;
        RECT -12.405 94.355 -12.075 94.685 ;
        RECT -12.405 92.995 -12.075 93.325 ;
        RECT -12.405 91.635 -12.075 91.965 ;
        RECT -12.405 90.275 -12.075 90.605 ;
        RECT -12.405 88.915 -12.075 89.245 ;
        RECT -12.405 87.555 -12.075 87.885 ;
        RECT -12.405 86.195 -12.075 86.525 ;
        RECT -12.405 84.835 -12.075 85.165 ;
        RECT -12.405 83.475 -12.075 83.805 ;
        RECT -12.405 82.115 -12.075 82.445 ;
        RECT -12.405 80.755 -12.075 81.085 ;
        RECT -12.405 79.395 -12.075 79.725 ;
        RECT -12.405 78.035 -12.075 78.365 ;
        RECT -12.405 76.675 -12.075 77.005 ;
        RECT -12.405 75.315 -12.075 75.645 ;
        RECT -12.405 73.955 -12.075 74.285 ;
        RECT -12.405 72.595 -12.075 72.925 ;
        RECT -12.405 71.235 -12.075 71.565 ;
        RECT -12.405 69.875 -12.075 70.205 ;
        RECT -12.405 68.515 -12.075 68.845 ;
        RECT -12.405 67.155 -12.075 67.485 ;
        RECT -12.405 65.795 -12.075 66.125 ;
        RECT -12.405 64.435 -12.075 64.765 ;
        RECT -12.405 63.075 -12.075 63.405 ;
        RECT -12.405 61.715 -12.075 62.045 ;
        RECT -12.405 60.355 -12.075 60.685 ;
        RECT -12.405 58.995 -12.075 59.325 ;
        RECT -12.405 57.635 -12.075 57.965 ;
        RECT -12.405 56.275 -12.075 56.605 ;
        RECT -12.405 54.915 -12.075 55.245 ;
        RECT -12.405 53.555 -12.075 53.885 ;
        RECT -12.405 52.195 -12.075 52.525 ;
        RECT -12.405 50.835 -12.075 51.165 ;
        RECT -12.405 49.475 -12.075 49.805 ;
        RECT -12.405 48.115 -12.075 48.445 ;
        RECT -12.405 46.755 -12.075 47.085 ;
        RECT -12.405 45.395 -12.075 45.725 ;
        RECT -12.405 44.035 -12.075 44.365 ;
        RECT -12.405 42.675 -12.075 43.005 ;
        RECT -12.405 41.315 -12.075 41.645 ;
        RECT -12.405 39.955 -12.075 40.285 ;
        RECT -12.405 38.595 -12.075 38.925 ;
        RECT -12.405 37.235 -12.075 37.565 ;
        RECT -12.405 35.875 -12.075 36.205 ;
        RECT -12.405 34.515 -12.075 34.845 ;
        RECT -12.405 33.155 -12.075 33.485 ;
        RECT -12.405 31.795 -12.075 32.125 ;
        RECT -12.405 30.435 -12.075 30.765 ;
        RECT -12.405 29.075 -12.075 29.405 ;
        RECT -12.405 27.715 -12.075 28.045 ;
        RECT -12.405 26.355 -12.075 26.685 ;
        RECT -12.405 24.995 -12.075 25.325 ;
        RECT -12.405 23.635 -12.075 23.965 ;
        RECT -12.405 22.275 -12.075 22.605 ;
        RECT -12.405 20.915 -12.075 21.245 ;
        RECT -12.405 19.555 -12.075 19.885 ;
        RECT -12.405 18.195 -12.075 18.525 ;
        RECT -12.405 16.835 -12.075 17.165 ;
        RECT -12.405 15.475 -12.075 15.805 ;
        RECT -12.405 14.115 -12.075 14.445 ;
        RECT -12.405 12.755 -12.075 13.085 ;
        RECT -12.405 11.395 -12.075 11.725 ;
        RECT -12.405 10.035 -12.075 10.365 ;
        RECT -12.405 8.675 -12.075 9.005 ;
        RECT -12.405 7.315 -12.075 7.645 ;
        RECT -12.405 5.955 -12.075 6.285 ;
        RECT -12.405 4.595 -12.075 4.925 ;
        RECT -12.405 3.235 -12.075 3.565 ;
        RECT -12.405 1.875 -12.075 2.205 ;
        RECT -12.405 0.515 -12.075 0.845 ;
        RECT -12.405 -0.845 -12.075 -0.515 ;
        RECT -12.405 -2.205 -12.075 -1.875 ;
        RECT -12.405 -3.565 -12.075 -3.235 ;
        RECT -12.405 -4.925 -12.075 -4.595 ;
        RECT -12.405 -6.285 -12.075 -5.955 ;
        RECT -12.405 -7.645 -12.075 -7.315 ;
        RECT -12.405 -9.005 -12.075 -8.675 ;
        RECT -12.405 -10.73 -12.075 -10.4 ;
        RECT -12.405 -11.725 -12.075 -11.395 ;
        RECT -12.405 -13.085 -12.075 -12.755 ;
        RECT -12.4 -15.12 -12.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -12.405 -26.685 -12.075 -26.355 ;
        RECT -12.405 -28.045 -12.075 -27.715 ;
        RECT -12.405 -29.405 -12.075 -29.075 ;
        RECT -12.405 -30.765 -12.075 -30.435 ;
        RECT -12.405 -32.125 -12.075 -31.795 ;
        RECT -12.405 -33.71 -12.075 -33.38 ;
        RECT -12.405 -39.75 -12.075 -39.42 ;
        RECT -12.405 -41.645 -12.075 -41.315 ;
        RECT -12.405 -44.365 -12.075 -44.035 ;
        RECT -12.405 -52.525 -12.075 -52.195 ;
        RECT -12.405 -53.885 -12.075 -53.555 ;
        RECT -12.405 -55.245 -12.075 -54.915 ;
        RECT -12.405 -56.605 -12.075 -56.275 ;
        RECT -12.405 -57.965 -12.075 -57.635 ;
        RECT -12.405 -59.325 -12.075 -58.995 ;
        RECT -12.405 -60.685 -12.075 -60.355 ;
        RECT -12.405 -62.045 -12.075 -61.715 ;
        RECT -12.405 -63.405 -12.075 -63.075 ;
        RECT -12.405 -64.765 -12.075 -64.435 ;
        RECT -12.405 -66.125 -12.075 -65.795 ;
        RECT -12.405 -68.845 -12.075 -68.515 ;
        RECT -12.405 -70.205 -12.075 -69.875 ;
        RECT -12.405 -71.565 -12.075 -71.235 ;
        RECT -12.405 -73.19 -12.075 -72.86 ;
        RECT -12.405 -74.285 -12.075 -73.955 ;
        RECT -12.405 -75.645 -12.075 -75.315 ;
        RECT -12.405 -78.365 -12.075 -78.035 ;
        RECT -12.405 -79.725 -12.075 -79.395 ;
        RECT -12.405 -80.73 -12.075 -80.4 ;
        RECT -12.405 -82.445 -12.075 -82.115 ;
        RECT -12.405 -83.805 -12.075 -83.475 ;
        RECT -12.405 -86.525 -12.075 -86.195 ;
        RECT -12.405 -89.245 -12.075 -88.915 ;
        RECT -12.405 -90.605 -12.075 -90.275 ;
        RECT -12.405 -91.965 -12.075 -91.635 ;
        RECT -12.405 -93.325 -12.075 -92.995 ;
        RECT -12.405 -94.685 -12.075 -94.355 ;
        RECT -12.405 -95.37 -12.075 -95.04 ;
        RECT -12.405 -97.405 -12.075 -97.075 ;
        RECT -12.405 -100.125 -12.075 -99.795 ;
        RECT -12.405 -101.485 -12.075 -101.155 ;
        RECT -12.405 -102.91 -12.075 -102.58 ;
        RECT -12.405 -113.725 -12.075 -113.395 ;
        RECT -12.405 -115.085 -12.075 -114.755 ;
        RECT -12.405 -116.445 -12.075 -116.115 ;
        RECT -12.405 -117.805 -12.075 -117.475 ;
        RECT -12.405 -119.165 -12.075 -118.835 ;
        RECT -12.405 -120.525 -12.075 -120.195 ;
        RECT -12.405 -121.885 -12.075 -121.555 ;
        RECT -12.405 -123.245 -12.075 -122.915 ;
        RECT -12.405 -130.045 -12.075 -129.715 ;
        RECT -12.405 -134.125 -12.075 -133.795 ;
        RECT -12.405 -135.485 -12.075 -135.155 ;
        RECT -12.405 -136.845 -12.075 -136.515 ;
        RECT -12.405 -138.205 -12.075 -137.875 ;
        RECT -12.405 -139.565 -12.075 -139.235 ;
        RECT -12.405 -140.925 -12.075 -140.595 ;
        RECT -12.405 -142.285 -12.075 -141.955 ;
        RECT -12.405 -145.005 -12.075 -144.675 ;
        RECT -12.405 -147.725 -12.075 -147.395 ;
        RECT -12.405 -150.445 -12.075 -150.115 ;
        RECT -12.405 -151.805 -12.075 -151.475 ;
        RECT -12.405 -153.165 -12.075 -152.835 ;
        RECT -12.405 -155.885 -12.075 -155.555 ;
        RECT -12.405 -159.965 -12.075 -159.635 ;
        RECT -12.405 -161.325 -12.075 -160.995 ;
        RECT -12.405 -162.685 -12.075 -162.355 ;
        RECT -12.405 -164.045 -12.075 -163.715 ;
        RECT -12.405 -165.405 -12.075 -165.075 ;
        RECT -12.405 -169.615 -12.075 -169.285 ;
        RECT -12.405 -170.845 -12.075 -170.515 ;
        RECT -12.405 -172.205 -12.075 -171.875 ;
        RECT -12.405 -173.565 -12.075 -173.235 ;
        RECT -12.405 -174.925 -12.075 -174.595 ;
        RECT -12.405 -177.645 -12.075 -177.315 ;
        RECT -12.405 -179.005 -12.075 -178.675 ;
        RECT -12.405 -184.65 -12.075 -183.52 ;
        RECT -12.4 -184.765 -12.08 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.045 244.04 -10.715 245.17 ;
        RECT -11.045 239.875 -10.715 240.205 ;
        RECT -11.045 238.515 -10.715 238.845 ;
        RECT -11.045 237.155 -10.715 237.485 ;
        RECT -11.045 235.795 -10.715 236.125 ;
        RECT -11.045 234.435 -10.715 234.765 ;
        RECT -11.045 233.075 -10.715 233.405 ;
        RECT -11.045 231.715 -10.715 232.045 ;
        RECT -11.045 227.635 -10.715 227.965 ;
        RECT -11.045 224.915 -10.715 225.245 ;
        RECT -11.045 218.115 -10.715 218.445 ;
        RECT -11.045 216.755 -10.715 217.085 ;
        RECT -11.045 207.235 -10.715 207.565 ;
        RECT -11.045 204.515 -10.715 204.845 ;
        RECT -11.045 203.155 -10.715 203.485 ;
        RECT -11.045 199.075 -10.715 199.405 ;
        RECT -11.045 196.355 -10.715 196.685 ;
        RECT -11.045 189.555 -10.715 189.885 ;
        RECT -11.045 188.195 -10.715 188.525 ;
        RECT -11.045 185.475 -10.715 185.805 ;
        RECT -11.045 178.675 -10.715 179.005 ;
        RECT -11.045 175.955 -10.715 176.285 ;
        RECT -11.045 174.595 -10.715 174.925 ;
        RECT -11.045 167.795 -10.715 168.125 ;
        RECT -11.045 160.995 -10.715 161.325 ;
        RECT -11.045 159.635 -10.715 159.965 ;
        RECT -11.045 156.915 -10.715 157.245 ;
        RECT -11.045 150.115 -10.715 150.445 ;
        RECT -11.045 147.395 -10.715 147.725 ;
        RECT -11.045 146.035 -10.715 146.365 ;
        RECT -11.045 139.235 -10.715 139.565 ;
        RECT -11.045 136.515 -10.715 136.845 ;
        RECT -11.045 132.435 -10.715 132.765 ;
        RECT -11.045 131.075 -10.715 131.405 ;
        RECT -11.045 128.355 -10.715 128.685 ;
        RECT -11.045 118.835 -10.715 119.165 ;
        RECT -11.045 117.475 -10.715 117.805 ;
        RECT -11.045 110.675 -10.715 111.005 ;
        RECT -11.045 107.955 -10.715 108.285 ;
        RECT -11.045 103.875 -10.715 104.205 ;
        RECT -11.045 99.795 -10.715 100.125 ;
        RECT -11.045 97.075 -10.715 97.405 ;
        RECT -11.045 90.275 -10.715 90.605 ;
        RECT -11.045 88.915 -10.715 89.245 ;
        RECT -11.045 82.115 -10.715 82.445 ;
        RECT -11.045 79.395 -10.715 79.725 ;
        RECT -11.045 75.315 -10.715 75.645 ;
        RECT -11.045 71.235 -10.715 71.565 ;
        RECT -11.045 68.515 -10.715 68.845 ;
        RECT -11.045 61.715 -10.715 62.045 ;
        RECT -11.045 60.355 -10.715 60.685 ;
        RECT -11.045 50.835 -10.715 51.165 ;
        RECT -11.045 46.755 -10.715 47.085 ;
        RECT -11.045 42.675 -10.715 43.005 ;
        RECT -11.045 39.955 -10.715 40.285 ;
        RECT -11.045 33.155 -10.715 33.485 ;
        RECT -11.045 31.795 -10.715 32.125 ;
        RECT -11.045 29.075 -10.715 29.405 ;
        RECT -11.045 22.275 -10.715 22.605 ;
        RECT -11.045 19.555 -10.715 19.885 ;
        RECT -11.045 18.195 -10.715 18.525 ;
        RECT -11.045 11.395 -10.715 11.725 ;
        RECT -11.045 4.595 -10.715 4.925 ;
        RECT -11.045 3.235 -10.715 3.565 ;
        RECT -11.045 1.875 -10.715 2.205 ;
        RECT -11.045 0.515 -10.715 0.845 ;
        RECT -11.045 -0.845 -10.715 -0.515 ;
        RECT -11.045 -2.205 -10.715 -1.875 ;
        RECT -11.045 -3.565 -10.715 -3.235 ;
        RECT -11.045 -4.925 -10.715 -4.595 ;
        RECT -11.045 -6.285 -10.715 -5.955 ;
        RECT -11.045 -7.645 -10.715 -7.315 ;
        RECT -11.045 -9.005 -10.715 -8.675 ;
        RECT -11.045 -10.73 -10.715 -10.4 ;
        RECT -11.045 -11.725 -10.715 -11.395 ;
        RECT -11.045 -13.085 -10.715 -12.755 ;
        RECT -11.045 -15.805 -10.715 -15.475 ;
        RECT -11.045 -16.77 -10.715 -16.44 ;
        RECT -11.045 -26.685 -10.715 -26.355 ;
        RECT -11.045 -28.045 -10.715 -27.715 ;
        RECT -11.045 -29.405 -10.715 -29.075 ;
        RECT -11.045 -30.765 -10.715 -30.435 ;
        RECT -11.045 -32.125 -10.715 -31.795 ;
        RECT -11.045 -33.71 -10.715 -33.38 ;
        RECT -11.045 -39.75 -10.715 -39.42 ;
        RECT -11.045 -41.645 -10.715 -41.315 ;
        RECT -11.045 -44.365 -10.715 -44.035 ;
        RECT -11.045 -52.525 -10.715 -52.195 ;
        RECT -11.045 -53.885 -10.715 -53.555 ;
        RECT -11.045 -55.245 -10.715 -54.915 ;
        RECT -11.045 -56.605 -10.715 -56.275 ;
        RECT -11.045 -57.965 -10.715 -57.635 ;
        RECT -11.045 -59.325 -10.715 -58.995 ;
        RECT -11.045 -60.685 -10.715 -60.355 ;
        RECT -11.045 -62.045 -10.715 -61.715 ;
        RECT -11.045 -63.405 -10.715 -63.075 ;
        RECT -11.045 -64.765 -10.715 -64.435 ;
        RECT -11.045 -66.125 -10.715 -65.795 ;
        RECT -11.045 -68.845 -10.715 -68.515 ;
        RECT -11.045 -70.205 -10.715 -69.875 ;
        RECT -11.045 -71.565 -10.715 -71.235 ;
        RECT -11.045 -73.19 -10.715 -72.86 ;
        RECT -11.045 -74.285 -10.715 -73.955 ;
        RECT -11.045 -75.645 -10.715 -75.315 ;
        RECT -11.045 -78.365 -10.715 -78.035 ;
        RECT -11.045 -79.725 -10.715 -79.395 ;
        RECT -11.045 -80.73 -10.715 -80.4 ;
        RECT -11.045 -82.445 -10.715 -82.115 ;
        RECT -11.045 -83.805 -10.715 -83.475 ;
        RECT -11.045 -86.525 -10.715 -86.195 ;
        RECT -11.045 -89.245 -10.715 -88.915 ;
        RECT -11.045 -90.605 -10.715 -90.275 ;
        RECT -11.045 -91.965 -10.715 -91.635 ;
        RECT -11.045 -93.325 -10.715 -92.995 ;
        RECT -11.045 -94.685 -10.715 -94.355 ;
        RECT -11.045 -95.37 -10.715 -95.04 ;
        RECT -11.045 -97.405 -10.715 -97.075 ;
        RECT -11.045 -100.125 -10.715 -99.795 ;
        RECT -11.045 -101.485 -10.715 -101.155 ;
        RECT -11.045 -102.91 -10.715 -102.58 ;
        RECT -11.045 -113.725 -10.715 -113.395 ;
        RECT -11.045 -115.085 -10.715 -114.755 ;
        RECT -11.045 -116.445 -10.715 -116.115 ;
        RECT -11.045 -117.805 -10.715 -117.475 ;
        RECT -11.045 -119.165 -10.715 -118.835 ;
        RECT -11.045 -120.525 -10.715 -120.195 ;
        RECT -11.045 -121.885 -10.715 -121.555 ;
        RECT -11.045 -123.245 -10.715 -122.915 ;
        RECT -11.045 -127.325 -10.715 -126.995 ;
        RECT -11.045 -130.045 -10.715 -129.715 ;
        RECT -11.045 -131.405 -10.715 -131.075 ;
        RECT -11.045 -134.125 -10.715 -133.795 ;
        RECT -11.045 -135.485 -10.715 -135.155 ;
        RECT -11.045 -136.845 -10.715 -136.515 ;
        RECT -11.045 -138.205 -10.715 -137.875 ;
        RECT -11.045 -139.565 -10.715 -139.235 ;
        RECT -11.045 -140.925 -10.715 -140.595 ;
        RECT -11.045 -142.285 -10.715 -141.955 ;
        RECT -11.045 -143.645 -10.715 -143.315 ;
        RECT -11.045 -145.005 -10.715 -144.675 ;
        RECT -11.045 -147.725 -10.715 -147.395 ;
        RECT -11.045 -150.445 -10.715 -150.115 ;
        RECT -11.045 -151.805 -10.715 -151.475 ;
        RECT -11.045 -153.165 -10.715 -152.835 ;
        RECT -11.045 -155.885 -10.715 -155.555 ;
        RECT -11.045 -158.605 -10.715 -158.275 ;
        RECT -11.045 -159.965 -10.715 -159.635 ;
        RECT -11.045 -161.325 -10.715 -160.995 ;
        RECT -11.045 -162.685 -10.715 -162.355 ;
        RECT -11.045 -164.045 -10.715 -163.715 ;
        RECT -11.045 -165.405 -10.715 -165.075 ;
        RECT -11.045 -169.615 -10.715 -169.285 ;
        RECT -11.045 -170.845 -10.715 -170.515 ;
        RECT -11.045 -172.205 -10.715 -171.875 ;
        RECT -11.045 -174.925 -10.715 -174.595 ;
        RECT -11.045 -177.645 -10.715 -177.315 ;
        RECT -11.045 -179.005 -10.715 -178.675 ;
        RECT -11.045 -184.65 -10.715 -183.52 ;
        RECT -11.04 -184.765 -10.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.685 -135.485 -9.355 -135.155 ;
        RECT -9.685 -136.845 -9.355 -136.515 ;
        RECT -9.685 -138.205 -9.355 -137.875 ;
        RECT -9.685 -139.565 -9.355 -139.235 ;
        RECT -9.685 -140.925 -9.355 -140.595 ;
        RECT -9.685 -142.285 -9.355 -141.955 ;
        RECT -9.685 -143.645 -9.355 -143.315 ;
        RECT -9.685 -145.005 -9.355 -144.675 ;
        RECT -9.685 -146.365 -9.355 -146.035 ;
        RECT -9.685 -147.725 -9.355 -147.395 ;
        RECT -9.685 -149.085 -9.355 -148.755 ;
        RECT -9.685 -150.445 -9.355 -150.115 ;
        RECT -9.685 -151.805 -9.355 -151.475 ;
        RECT -9.685 -153.165 -9.355 -152.835 ;
        RECT -9.685 -154.525 -9.355 -154.195 ;
        RECT -9.685 -155.885 -9.355 -155.555 ;
        RECT -9.685 -157.245 -9.355 -156.915 ;
        RECT -9.685 -158.605 -9.355 -158.275 ;
        RECT -9.685 -159.965 -9.355 -159.635 ;
        RECT -9.685 -161.325 -9.355 -160.995 ;
        RECT -9.685 -162.685 -9.355 -162.355 ;
        RECT -9.685 -164.045 -9.355 -163.715 ;
        RECT -9.685 -165.405 -9.355 -165.075 ;
        RECT -9.68 -167.44 -9.36 245.285 ;
        RECT -9.685 244.04 -9.355 245.17 ;
        RECT -9.685 239.875 -9.355 240.205 ;
        RECT -9.685 238.515 -9.355 238.845 ;
        RECT -9.685 237.155 -9.355 237.485 ;
        RECT -9.685 235.795 -9.355 236.125 ;
        RECT -9.685 234.435 -9.355 234.765 ;
        RECT -9.685 233.075 -9.355 233.405 ;
        RECT -9.685 231.715 -9.355 232.045 ;
        RECT -9.685 227.635 -9.355 227.965 ;
        RECT -9.685 224.915 -9.355 225.245 ;
        RECT -9.685 218.115 -9.355 218.445 ;
        RECT -9.685 216.755 -9.355 217.085 ;
        RECT -9.685 207.235 -9.355 207.565 ;
        RECT -9.685 204.515 -9.355 204.845 ;
        RECT -9.685 203.155 -9.355 203.485 ;
        RECT -9.685 199.075 -9.355 199.405 ;
        RECT -9.685 196.355 -9.355 196.685 ;
        RECT -9.685 189.555 -9.355 189.885 ;
        RECT -9.685 188.195 -9.355 188.525 ;
        RECT -9.685 185.475 -9.355 185.805 ;
        RECT -9.685 178.675 -9.355 179.005 ;
        RECT -9.685 175.955 -9.355 176.285 ;
        RECT -9.685 174.595 -9.355 174.925 ;
        RECT -9.685 167.795 -9.355 168.125 ;
        RECT -9.685 160.995 -9.355 161.325 ;
        RECT -9.685 159.635 -9.355 159.965 ;
        RECT -9.685 156.915 -9.355 157.245 ;
        RECT -9.685 150.115 -9.355 150.445 ;
        RECT -9.685 147.395 -9.355 147.725 ;
        RECT -9.685 146.035 -9.355 146.365 ;
        RECT -9.685 139.235 -9.355 139.565 ;
        RECT -9.685 136.515 -9.355 136.845 ;
        RECT -9.685 132.435 -9.355 132.765 ;
        RECT -9.685 131.075 -9.355 131.405 ;
        RECT -9.685 128.355 -9.355 128.685 ;
        RECT -9.685 118.835 -9.355 119.165 ;
        RECT -9.685 117.475 -9.355 117.805 ;
        RECT -9.685 110.675 -9.355 111.005 ;
        RECT -9.685 107.955 -9.355 108.285 ;
        RECT -9.685 103.875 -9.355 104.205 ;
        RECT -9.685 99.795 -9.355 100.125 ;
        RECT -9.685 97.075 -9.355 97.405 ;
        RECT -9.685 90.275 -9.355 90.605 ;
        RECT -9.685 88.915 -9.355 89.245 ;
        RECT -9.685 82.115 -9.355 82.445 ;
        RECT -9.685 79.395 -9.355 79.725 ;
        RECT -9.685 75.315 -9.355 75.645 ;
        RECT -9.685 71.235 -9.355 71.565 ;
        RECT -9.685 68.515 -9.355 68.845 ;
        RECT -9.685 61.715 -9.355 62.045 ;
        RECT -9.685 60.355 -9.355 60.685 ;
        RECT -9.685 50.835 -9.355 51.165 ;
        RECT -9.685 46.755 -9.355 47.085 ;
        RECT -9.685 42.675 -9.355 43.005 ;
        RECT -9.685 39.955 -9.355 40.285 ;
        RECT -9.685 33.155 -9.355 33.485 ;
        RECT -9.685 31.795 -9.355 32.125 ;
        RECT -9.685 29.075 -9.355 29.405 ;
        RECT -9.685 22.275 -9.355 22.605 ;
        RECT -9.685 19.555 -9.355 19.885 ;
        RECT -9.685 18.195 -9.355 18.525 ;
        RECT -9.685 11.395 -9.355 11.725 ;
        RECT -9.685 4.595 -9.355 4.925 ;
        RECT -9.685 3.235 -9.355 3.565 ;
        RECT -9.685 1.875 -9.355 2.205 ;
        RECT -9.685 0.515 -9.355 0.845 ;
        RECT -9.685 -0.845 -9.355 -0.515 ;
        RECT -9.685 -2.205 -9.355 -1.875 ;
        RECT -9.685 -3.565 -9.355 -3.235 ;
        RECT -9.685 -4.925 -9.355 -4.595 ;
        RECT -9.685 -6.285 -9.355 -5.955 ;
        RECT -9.685 -7.645 -9.355 -7.315 ;
        RECT -9.685 -9.005 -9.355 -8.675 ;
        RECT -9.685 -11.725 -9.355 -11.395 ;
        RECT -9.685 -13.085 -9.355 -12.755 ;
        RECT -9.685 -15.805 -9.355 -15.475 ;
        RECT -9.685 -26.685 -9.355 -26.355 ;
        RECT -9.685 -28.045 -9.355 -27.715 ;
        RECT -9.685 -29.405 -9.355 -29.075 ;
        RECT -9.685 -30.765 -9.355 -30.435 ;
        RECT -9.685 -32.125 -9.355 -31.795 ;
        RECT -9.685 -41.645 -9.355 -41.315 ;
        RECT -9.685 -44.365 -9.355 -44.035 ;
        RECT -9.685 -52.525 -9.355 -52.195 ;
        RECT -9.685 -53.885 -9.355 -53.555 ;
        RECT -9.685 -55.245 -9.355 -54.915 ;
        RECT -9.685 -56.605 -9.355 -56.275 ;
        RECT -9.685 -57.965 -9.355 -57.635 ;
        RECT -9.685 -59.325 -9.355 -58.995 ;
        RECT -9.685 -60.685 -9.355 -60.355 ;
        RECT -9.685 -62.045 -9.355 -61.715 ;
        RECT -9.685 -63.405 -9.355 -63.075 ;
        RECT -9.685 -64.765 -9.355 -64.435 ;
        RECT -9.685 -66.125 -9.355 -65.795 ;
        RECT -9.685 -68.845 -9.355 -68.515 ;
        RECT -9.685 -70.205 -9.355 -69.875 ;
        RECT -9.685 -71.565 -9.355 -71.235 ;
        RECT -9.685 -74.285 -9.355 -73.955 ;
        RECT -9.685 -75.645 -9.355 -75.315 ;
        RECT -9.685 -78.365 -9.355 -78.035 ;
        RECT -9.685 -79.725 -9.355 -79.395 ;
        RECT -9.685 -82.445 -9.355 -82.115 ;
        RECT -9.685 -83.805 -9.355 -83.475 ;
        RECT -9.685 -86.525 -9.355 -86.195 ;
        RECT -9.685 -89.245 -9.355 -88.915 ;
        RECT -9.685 -90.605 -9.355 -90.275 ;
        RECT -9.685 -91.965 -9.355 -91.635 ;
        RECT -9.685 -93.325 -9.355 -92.995 ;
        RECT -9.685 -94.685 -9.355 -94.355 ;
        RECT -9.685 -97.405 -9.355 -97.075 ;
        RECT -9.685 -100.125 -9.355 -99.795 ;
        RECT -9.685 -101.485 -9.355 -101.155 ;
        RECT -9.685 -113.725 -9.355 -113.395 ;
        RECT -9.685 -115.085 -9.355 -114.755 ;
        RECT -9.685 -116.445 -9.355 -116.115 ;
        RECT -9.685 -117.805 -9.355 -117.475 ;
        RECT -9.685 -119.165 -9.355 -118.835 ;
        RECT -9.685 -120.525 -9.355 -120.195 ;
        RECT -9.685 -121.885 -9.355 -121.555 ;
        RECT -9.685 -123.245 -9.355 -122.915 ;
        RECT -9.685 -124.605 -9.355 -124.275 ;
        RECT -9.685 -127.325 -9.355 -126.995 ;
        RECT -9.685 -128.685 -9.355 -128.355 ;
        RECT -9.685 -130.045 -9.355 -129.715 ;
        RECT -9.685 -131.405 -9.355 -131.075 ;
        RECT -9.685 -134.125 -9.355 -133.795 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 -30.765 -21.595 -30.435 ;
        RECT -21.925 -32.125 -21.595 -31.795 ;
        RECT -21.925 -33.71 -21.595 -33.38 ;
        RECT -21.925 -34.845 -21.595 -34.515 ;
        RECT -21.925 -36.205 -21.595 -35.875 ;
        RECT -21.925 -39.75 -21.595 -39.42 ;
        RECT -21.925 -41.645 -21.595 -41.315 ;
        RECT -21.925 -44.365 -21.595 -44.035 ;
        RECT -21.925 -51.165 -21.595 -50.835 ;
        RECT -21.925 -52.525 -21.595 -52.195 ;
        RECT -21.925 -53.885 -21.595 -53.555 ;
        RECT -21.925 -55.245 -21.595 -54.915 ;
        RECT -21.925 -56.605 -21.595 -56.275 ;
        RECT -21.925 -57.965 -21.595 -57.635 ;
        RECT -21.925 -59.325 -21.595 -58.995 ;
        RECT -21.925 -60.685 -21.595 -60.355 ;
        RECT -21.925 -62.045 -21.595 -61.715 ;
        RECT -21.925 -63.405 -21.595 -63.075 ;
        RECT -21.925 -64.765 -21.595 -64.435 ;
        RECT -21.925 -66.125 -21.595 -65.795 ;
        RECT -21.925 -68.845 -21.595 -68.515 ;
        RECT -21.925 -70.205 -21.595 -69.875 ;
        RECT -21.925 -71.565 -21.595 -71.235 ;
        RECT -21.925 -73.19 -21.595 -72.86 ;
        RECT -21.925 -74.285 -21.595 -73.955 ;
        RECT -21.925 -75.645 -21.595 -75.315 ;
        RECT -21.925 -78.365 -21.595 -78.035 ;
        RECT -21.925 -79.725 -21.595 -79.395 ;
        RECT -21.925 -80.73 -21.595 -80.4 ;
        RECT -21.925 -82.445 -21.595 -82.115 ;
        RECT -21.925 -83.805 -21.595 -83.475 ;
        RECT -21.925 -86.525 -21.595 -86.195 ;
        RECT -21.925 -89.245 -21.595 -88.915 ;
        RECT -21.925 -90.605 -21.595 -90.275 ;
        RECT -21.925 -91.965 -21.595 -91.635 ;
        RECT -21.925 -93.325 -21.595 -92.995 ;
        RECT -21.925 -94.685 -21.595 -94.355 ;
        RECT -21.925 -95.37 -21.595 -95.04 ;
        RECT -21.925 -97.405 -21.595 -97.075 ;
        RECT -21.925 -100.125 -21.595 -99.795 ;
        RECT -21.925 -101.485 -21.595 -101.155 ;
        RECT -21.925 -102.91 -21.595 -102.58 ;
        RECT -21.925 -104.205 -21.595 -103.875 ;
        RECT -21.92 -111.68 -21.6 -29.76 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 -117.805 -21.595 -117.475 ;
        RECT -21.925 -119.165 -21.595 -118.835 ;
        RECT -21.925 -120.525 -21.595 -120.195 ;
        RECT -21.925 -123.245 -21.595 -122.915 ;
        RECT -21.925 -124.605 -21.595 -124.275 ;
        RECT -21.925 -125.965 -21.595 -125.635 ;
        RECT -21.925 -127.325 -21.595 -126.995 ;
        RECT -21.925 -128.685 -21.595 -128.355 ;
        RECT -21.925 -135.485 -21.595 -135.155 ;
        RECT -21.925 -139.565 -21.595 -139.235 ;
        RECT -21.925 -142.285 -21.595 -141.955 ;
        RECT -21.925 -143.645 -21.595 -143.315 ;
        RECT -21.925 -147.725 -21.595 -147.395 ;
        RECT -21.925 -149.085 -21.595 -148.755 ;
        RECT -21.925 -151.805 -21.595 -151.475 ;
        RECT -21.925 -153.165 -21.595 -152.835 ;
        RECT -21.925 -158.605 -21.595 -158.275 ;
        RECT -21.925 -159.965 -21.595 -159.635 ;
        RECT -21.925 -161.325 -21.595 -160.995 ;
        RECT -21.925 -162.685 -21.595 -162.355 ;
        RECT -21.925 -164.045 -21.595 -163.715 ;
        RECT -21.925 -165.405 -21.595 -165.075 ;
        RECT -21.925 -166.765 -21.595 -166.435 ;
        RECT -21.925 -169.615 -21.595 -169.285 ;
        RECT -21.925 -170.845 -21.595 -170.515 ;
        RECT -21.925 -172.205 -21.595 -171.875 ;
        RECT -21.925 -177.645 -21.595 -177.315 ;
        RECT -21.925 -179.005 -21.595 -178.675 ;
        RECT -21.925 -184.65 -21.595 -183.52 ;
        RECT -21.92 -184.765 -21.6 -116.8 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 244.04 -20.235 245.17 ;
        RECT -20.565 239.875 -20.235 240.205 ;
        RECT -20.565 238.515 -20.235 238.845 ;
        RECT -20.565 237.155 -20.235 237.485 ;
        RECT -20.565 235.795 -20.235 236.125 ;
        RECT -20.565 234.435 -20.235 234.765 ;
        RECT -20.565 233.075 -20.235 233.405 ;
        RECT -20.565 231.715 -20.235 232.045 ;
        RECT -20.565 230.355 -20.235 230.685 ;
        RECT -20.565 228.995 -20.235 229.325 ;
        RECT -20.565 227.635 -20.235 227.965 ;
        RECT -20.565 226.275 -20.235 226.605 ;
        RECT -20.565 224.915 -20.235 225.245 ;
        RECT -20.565 223.555 -20.235 223.885 ;
        RECT -20.565 222.195 -20.235 222.525 ;
        RECT -20.565 220.835 -20.235 221.165 ;
        RECT -20.565 219.475 -20.235 219.805 ;
        RECT -20.565 218.115 -20.235 218.445 ;
        RECT -20.565 216.755 -20.235 217.085 ;
        RECT -20.565 215.395 -20.235 215.725 ;
        RECT -20.565 214.035 -20.235 214.365 ;
        RECT -20.565 212.675 -20.235 213.005 ;
        RECT -20.565 211.315 -20.235 211.645 ;
        RECT -20.565 209.955 -20.235 210.285 ;
        RECT -20.565 208.595 -20.235 208.925 ;
        RECT -20.565 207.235 -20.235 207.565 ;
        RECT -20.565 205.875 -20.235 206.205 ;
        RECT -20.565 204.515 -20.235 204.845 ;
        RECT -20.565 203.155 -20.235 203.485 ;
        RECT -20.565 201.795 -20.235 202.125 ;
        RECT -20.565 200.435 -20.235 200.765 ;
        RECT -20.565 199.075 -20.235 199.405 ;
        RECT -20.565 197.715 -20.235 198.045 ;
        RECT -20.565 196.355 -20.235 196.685 ;
        RECT -20.565 194.995 -20.235 195.325 ;
        RECT -20.565 193.635 -20.235 193.965 ;
        RECT -20.565 192.275 -20.235 192.605 ;
        RECT -20.565 190.915 -20.235 191.245 ;
        RECT -20.565 189.555 -20.235 189.885 ;
        RECT -20.565 188.195 -20.235 188.525 ;
        RECT -20.565 186.835 -20.235 187.165 ;
        RECT -20.565 185.475 -20.235 185.805 ;
        RECT -20.565 184.115 -20.235 184.445 ;
        RECT -20.565 182.755 -20.235 183.085 ;
        RECT -20.565 181.395 -20.235 181.725 ;
        RECT -20.565 180.035 -20.235 180.365 ;
        RECT -20.565 178.675 -20.235 179.005 ;
        RECT -20.565 177.315 -20.235 177.645 ;
        RECT -20.565 175.955 -20.235 176.285 ;
        RECT -20.565 174.595 -20.235 174.925 ;
        RECT -20.565 173.235 -20.235 173.565 ;
        RECT -20.565 171.875 -20.235 172.205 ;
        RECT -20.565 170.515 -20.235 170.845 ;
        RECT -20.565 169.155 -20.235 169.485 ;
        RECT -20.565 167.795 -20.235 168.125 ;
        RECT -20.565 166.435 -20.235 166.765 ;
        RECT -20.565 165.075 -20.235 165.405 ;
        RECT -20.565 163.715 -20.235 164.045 ;
        RECT -20.565 162.355 -20.235 162.685 ;
        RECT -20.565 160.995 -20.235 161.325 ;
        RECT -20.565 159.635 -20.235 159.965 ;
        RECT -20.565 158.275 -20.235 158.605 ;
        RECT -20.565 156.915 -20.235 157.245 ;
        RECT -20.565 155.555 -20.235 155.885 ;
        RECT -20.565 154.195 -20.235 154.525 ;
        RECT -20.565 152.835 -20.235 153.165 ;
        RECT -20.565 151.475 -20.235 151.805 ;
        RECT -20.565 150.115 -20.235 150.445 ;
        RECT -20.565 148.755 -20.235 149.085 ;
        RECT -20.565 147.395 -20.235 147.725 ;
        RECT -20.565 146.035 -20.235 146.365 ;
        RECT -20.565 144.675 -20.235 145.005 ;
        RECT -20.565 143.315 -20.235 143.645 ;
        RECT -20.565 141.955 -20.235 142.285 ;
        RECT -20.565 140.595 -20.235 140.925 ;
        RECT -20.565 139.235 -20.235 139.565 ;
        RECT -20.565 137.875 -20.235 138.205 ;
        RECT -20.565 136.515 -20.235 136.845 ;
        RECT -20.565 135.155 -20.235 135.485 ;
        RECT -20.565 133.795 -20.235 134.125 ;
        RECT -20.565 132.435 -20.235 132.765 ;
        RECT -20.565 131.075 -20.235 131.405 ;
        RECT -20.565 129.715 -20.235 130.045 ;
        RECT -20.565 128.355 -20.235 128.685 ;
        RECT -20.565 126.995 -20.235 127.325 ;
        RECT -20.565 125.635 -20.235 125.965 ;
        RECT -20.565 124.275 -20.235 124.605 ;
        RECT -20.565 122.915 -20.235 123.245 ;
        RECT -20.565 121.555 -20.235 121.885 ;
        RECT -20.565 120.195 -20.235 120.525 ;
        RECT -20.565 118.835 -20.235 119.165 ;
        RECT -20.565 117.475 -20.235 117.805 ;
        RECT -20.565 116.115 -20.235 116.445 ;
        RECT -20.565 114.755 -20.235 115.085 ;
        RECT -20.565 113.395 -20.235 113.725 ;
        RECT -20.565 112.035 -20.235 112.365 ;
        RECT -20.565 110.675 -20.235 111.005 ;
        RECT -20.565 109.315 -20.235 109.645 ;
        RECT -20.565 107.955 -20.235 108.285 ;
        RECT -20.565 106.595 -20.235 106.925 ;
        RECT -20.565 105.235 -20.235 105.565 ;
        RECT -20.565 103.875 -20.235 104.205 ;
        RECT -20.565 102.515 -20.235 102.845 ;
        RECT -20.565 101.155 -20.235 101.485 ;
        RECT -20.565 99.795 -20.235 100.125 ;
        RECT -20.565 98.435 -20.235 98.765 ;
        RECT -20.565 97.075 -20.235 97.405 ;
        RECT -20.565 95.715 -20.235 96.045 ;
        RECT -20.565 94.355 -20.235 94.685 ;
        RECT -20.565 92.995 -20.235 93.325 ;
        RECT -20.565 91.635 -20.235 91.965 ;
        RECT -20.565 90.275 -20.235 90.605 ;
        RECT -20.565 88.915 -20.235 89.245 ;
        RECT -20.565 87.555 -20.235 87.885 ;
        RECT -20.565 86.195 -20.235 86.525 ;
        RECT -20.565 84.835 -20.235 85.165 ;
        RECT -20.565 83.475 -20.235 83.805 ;
        RECT -20.565 82.115 -20.235 82.445 ;
        RECT -20.565 80.755 -20.235 81.085 ;
        RECT -20.565 79.395 -20.235 79.725 ;
        RECT -20.565 78.035 -20.235 78.365 ;
        RECT -20.565 76.675 -20.235 77.005 ;
        RECT -20.565 75.315 -20.235 75.645 ;
        RECT -20.565 73.955 -20.235 74.285 ;
        RECT -20.565 72.595 -20.235 72.925 ;
        RECT -20.565 71.235 -20.235 71.565 ;
        RECT -20.565 69.875 -20.235 70.205 ;
        RECT -20.565 68.515 -20.235 68.845 ;
        RECT -20.565 67.155 -20.235 67.485 ;
        RECT -20.565 65.795 -20.235 66.125 ;
        RECT -20.565 64.435 -20.235 64.765 ;
        RECT -20.565 63.075 -20.235 63.405 ;
        RECT -20.565 61.715 -20.235 62.045 ;
        RECT -20.565 60.355 -20.235 60.685 ;
        RECT -20.565 58.995 -20.235 59.325 ;
        RECT -20.565 57.635 -20.235 57.965 ;
        RECT -20.565 56.275 -20.235 56.605 ;
        RECT -20.565 54.915 -20.235 55.245 ;
        RECT -20.565 53.555 -20.235 53.885 ;
        RECT -20.565 52.195 -20.235 52.525 ;
        RECT -20.565 50.835 -20.235 51.165 ;
        RECT -20.565 49.475 -20.235 49.805 ;
        RECT -20.565 48.115 -20.235 48.445 ;
        RECT -20.565 46.755 -20.235 47.085 ;
        RECT -20.565 45.395 -20.235 45.725 ;
        RECT -20.565 44.035 -20.235 44.365 ;
        RECT -20.565 42.675 -20.235 43.005 ;
        RECT -20.565 41.315 -20.235 41.645 ;
        RECT -20.565 39.955 -20.235 40.285 ;
        RECT -20.565 38.595 -20.235 38.925 ;
        RECT -20.565 37.235 -20.235 37.565 ;
        RECT -20.565 35.875 -20.235 36.205 ;
        RECT -20.565 34.515 -20.235 34.845 ;
        RECT -20.565 33.155 -20.235 33.485 ;
        RECT -20.565 31.795 -20.235 32.125 ;
        RECT -20.565 30.435 -20.235 30.765 ;
        RECT -20.565 29.075 -20.235 29.405 ;
        RECT -20.565 27.715 -20.235 28.045 ;
        RECT -20.565 26.355 -20.235 26.685 ;
        RECT -20.565 24.995 -20.235 25.325 ;
        RECT -20.565 23.635 -20.235 23.965 ;
        RECT -20.565 22.275 -20.235 22.605 ;
        RECT -20.565 20.915 -20.235 21.245 ;
        RECT -20.565 19.555 -20.235 19.885 ;
        RECT -20.565 18.195 -20.235 18.525 ;
        RECT -20.565 16.835 -20.235 17.165 ;
        RECT -20.565 15.475 -20.235 15.805 ;
        RECT -20.565 14.115 -20.235 14.445 ;
        RECT -20.565 12.755 -20.235 13.085 ;
        RECT -20.565 11.395 -20.235 11.725 ;
        RECT -20.565 10.035 -20.235 10.365 ;
        RECT -20.565 8.675 -20.235 9.005 ;
        RECT -20.565 7.315 -20.235 7.645 ;
        RECT -20.565 5.955 -20.235 6.285 ;
        RECT -20.565 4.595 -20.235 4.925 ;
        RECT -20.565 3.235 -20.235 3.565 ;
        RECT -20.565 1.875 -20.235 2.205 ;
        RECT -20.565 0.515 -20.235 0.845 ;
        RECT -20.565 -0.845 -20.235 -0.515 ;
        RECT -20.565 -2.205 -20.235 -1.875 ;
        RECT -20.565 -3.565 -20.235 -3.235 ;
        RECT -20.565 -7.645 -20.235 -7.315 ;
        RECT -20.565 -9.005 -20.235 -8.675 ;
        RECT -20.565 -10.73 -20.235 -10.4 ;
        RECT -20.565 -11.725 -20.235 -11.395 ;
        RECT -20.565 -16.77 -20.235 -16.44 ;
        RECT -20.565 -18.525 -20.235 -18.195 ;
        RECT -20.565 -21.245 -20.235 -20.915 ;
        RECT -20.56 -22.6 -20.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 -29.405 -20.235 -29.075 ;
        RECT -20.565 -30.765 -20.235 -30.435 ;
        RECT -20.565 -32.125 -20.235 -31.795 ;
        RECT -20.565 -33.71 -20.235 -33.38 ;
        RECT -20.565 -34.845 -20.235 -34.515 ;
        RECT -20.565 -36.205 -20.235 -35.875 ;
        RECT -20.565 -39.75 -20.235 -39.42 ;
        RECT -20.565 -41.645 -20.235 -41.315 ;
        RECT -20.565 -44.365 -20.235 -44.035 ;
        RECT -20.565 -51.165 -20.235 -50.835 ;
        RECT -20.565 -52.525 -20.235 -52.195 ;
        RECT -20.565 -53.885 -20.235 -53.555 ;
        RECT -20.565 -55.245 -20.235 -54.915 ;
        RECT -20.565 -56.605 -20.235 -56.275 ;
        RECT -20.565 -57.965 -20.235 -57.635 ;
        RECT -20.565 -59.325 -20.235 -58.995 ;
        RECT -20.565 -60.685 -20.235 -60.355 ;
        RECT -20.565 -62.045 -20.235 -61.715 ;
        RECT -20.565 -63.405 -20.235 -63.075 ;
        RECT -20.565 -64.765 -20.235 -64.435 ;
        RECT -20.565 -66.125 -20.235 -65.795 ;
        RECT -20.565 -68.845 -20.235 -68.515 ;
        RECT -20.565 -70.205 -20.235 -69.875 ;
        RECT -20.565 -71.565 -20.235 -71.235 ;
        RECT -20.565 -73.19 -20.235 -72.86 ;
        RECT -20.565 -74.285 -20.235 -73.955 ;
        RECT -20.565 -75.645 -20.235 -75.315 ;
        RECT -20.565 -78.365 -20.235 -78.035 ;
        RECT -20.565 -79.725 -20.235 -79.395 ;
        RECT -20.565 -80.73 -20.235 -80.4 ;
        RECT -20.565 -82.445 -20.235 -82.115 ;
        RECT -20.565 -83.805 -20.235 -83.475 ;
        RECT -20.565 -86.525 -20.235 -86.195 ;
        RECT -20.565 -89.245 -20.235 -88.915 ;
        RECT -20.565 -90.605 -20.235 -90.275 ;
        RECT -20.565 -91.965 -20.235 -91.635 ;
        RECT -20.565 -93.325 -20.235 -92.995 ;
        RECT -20.565 -94.685 -20.235 -94.355 ;
        RECT -20.565 -95.37 -20.235 -95.04 ;
        RECT -20.565 -97.405 -20.235 -97.075 ;
        RECT -20.565 -100.125 -20.235 -99.795 ;
        RECT -20.565 -101.485 -20.235 -101.155 ;
        RECT -20.565 -102.91 -20.235 -102.58 ;
        RECT -20.565 -104.205 -20.235 -103.875 ;
        RECT -20.56 -110.32 -20.24 -28.4 ;
    END
    PORT
      LAYER met3 ;
        RECT -20.565 -177.645 -20.235 -177.315 ;
        RECT -20.565 -179.005 -20.235 -178.675 ;
        RECT -20.565 -184.65 -20.235 -183.52 ;
        RECT -20.56 -184.765 -20.24 -175.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 244.04 -18.875 245.17 ;
        RECT -19.205 239.875 -18.875 240.205 ;
        RECT -19.205 238.515 -18.875 238.845 ;
        RECT -19.205 237.155 -18.875 237.485 ;
        RECT -19.205 235.795 -18.875 236.125 ;
        RECT -19.205 234.435 -18.875 234.765 ;
        RECT -19.205 233.075 -18.875 233.405 ;
        RECT -19.205 231.715 -18.875 232.045 ;
        RECT -19.205 230.355 -18.875 230.685 ;
        RECT -19.205 228.995 -18.875 229.325 ;
        RECT -19.205 227.635 -18.875 227.965 ;
        RECT -19.205 226.275 -18.875 226.605 ;
        RECT -19.205 224.915 -18.875 225.245 ;
        RECT -19.205 223.555 -18.875 223.885 ;
        RECT -19.205 222.195 -18.875 222.525 ;
        RECT -19.205 220.835 -18.875 221.165 ;
        RECT -19.205 219.475 -18.875 219.805 ;
        RECT -19.205 218.115 -18.875 218.445 ;
        RECT -19.205 216.755 -18.875 217.085 ;
        RECT -19.205 215.395 -18.875 215.725 ;
        RECT -19.205 214.035 -18.875 214.365 ;
        RECT -19.205 212.675 -18.875 213.005 ;
        RECT -19.205 211.315 -18.875 211.645 ;
        RECT -19.205 209.955 -18.875 210.285 ;
        RECT -19.205 208.595 -18.875 208.925 ;
        RECT -19.205 207.235 -18.875 207.565 ;
        RECT -19.205 205.875 -18.875 206.205 ;
        RECT -19.205 204.515 -18.875 204.845 ;
        RECT -19.205 203.155 -18.875 203.485 ;
        RECT -19.205 201.795 -18.875 202.125 ;
        RECT -19.205 200.435 -18.875 200.765 ;
        RECT -19.205 199.075 -18.875 199.405 ;
        RECT -19.205 197.715 -18.875 198.045 ;
        RECT -19.205 196.355 -18.875 196.685 ;
        RECT -19.205 194.995 -18.875 195.325 ;
        RECT -19.205 193.635 -18.875 193.965 ;
        RECT -19.205 192.275 -18.875 192.605 ;
        RECT -19.205 190.915 -18.875 191.245 ;
        RECT -19.205 189.555 -18.875 189.885 ;
        RECT -19.205 188.195 -18.875 188.525 ;
        RECT -19.205 186.835 -18.875 187.165 ;
        RECT -19.205 185.475 -18.875 185.805 ;
        RECT -19.205 184.115 -18.875 184.445 ;
        RECT -19.205 182.755 -18.875 183.085 ;
        RECT -19.205 181.395 -18.875 181.725 ;
        RECT -19.205 180.035 -18.875 180.365 ;
        RECT -19.205 178.675 -18.875 179.005 ;
        RECT -19.205 177.315 -18.875 177.645 ;
        RECT -19.205 175.955 -18.875 176.285 ;
        RECT -19.205 174.595 -18.875 174.925 ;
        RECT -19.205 173.235 -18.875 173.565 ;
        RECT -19.205 171.875 -18.875 172.205 ;
        RECT -19.205 170.515 -18.875 170.845 ;
        RECT -19.205 169.155 -18.875 169.485 ;
        RECT -19.205 167.795 -18.875 168.125 ;
        RECT -19.205 166.435 -18.875 166.765 ;
        RECT -19.205 165.075 -18.875 165.405 ;
        RECT -19.205 163.715 -18.875 164.045 ;
        RECT -19.205 162.355 -18.875 162.685 ;
        RECT -19.205 160.995 -18.875 161.325 ;
        RECT -19.205 159.635 -18.875 159.965 ;
        RECT -19.205 158.275 -18.875 158.605 ;
        RECT -19.205 156.915 -18.875 157.245 ;
        RECT -19.205 155.555 -18.875 155.885 ;
        RECT -19.205 154.195 -18.875 154.525 ;
        RECT -19.205 152.835 -18.875 153.165 ;
        RECT -19.205 151.475 -18.875 151.805 ;
        RECT -19.205 150.115 -18.875 150.445 ;
        RECT -19.205 148.755 -18.875 149.085 ;
        RECT -19.205 147.395 -18.875 147.725 ;
        RECT -19.205 146.035 -18.875 146.365 ;
        RECT -19.205 144.675 -18.875 145.005 ;
        RECT -19.205 143.315 -18.875 143.645 ;
        RECT -19.205 141.955 -18.875 142.285 ;
        RECT -19.205 140.595 -18.875 140.925 ;
        RECT -19.205 139.235 -18.875 139.565 ;
        RECT -19.205 137.875 -18.875 138.205 ;
        RECT -19.205 136.515 -18.875 136.845 ;
        RECT -19.205 135.155 -18.875 135.485 ;
        RECT -19.205 133.795 -18.875 134.125 ;
        RECT -19.205 132.435 -18.875 132.765 ;
        RECT -19.205 131.075 -18.875 131.405 ;
        RECT -19.205 129.715 -18.875 130.045 ;
        RECT -19.205 128.355 -18.875 128.685 ;
        RECT -19.205 126.995 -18.875 127.325 ;
        RECT -19.205 125.635 -18.875 125.965 ;
        RECT -19.205 124.275 -18.875 124.605 ;
        RECT -19.205 122.915 -18.875 123.245 ;
        RECT -19.205 121.555 -18.875 121.885 ;
        RECT -19.205 120.195 -18.875 120.525 ;
        RECT -19.205 118.835 -18.875 119.165 ;
        RECT -19.205 117.475 -18.875 117.805 ;
        RECT -19.205 116.115 -18.875 116.445 ;
        RECT -19.205 114.755 -18.875 115.085 ;
        RECT -19.205 113.395 -18.875 113.725 ;
        RECT -19.205 112.035 -18.875 112.365 ;
        RECT -19.205 110.675 -18.875 111.005 ;
        RECT -19.205 109.315 -18.875 109.645 ;
        RECT -19.205 107.955 -18.875 108.285 ;
        RECT -19.205 106.595 -18.875 106.925 ;
        RECT -19.205 105.235 -18.875 105.565 ;
        RECT -19.205 103.875 -18.875 104.205 ;
        RECT -19.205 102.515 -18.875 102.845 ;
        RECT -19.205 101.155 -18.875 101.485 ;
        RECT -19.205 99.795 -18.875 100.125 ;
        RECT -19.205 98.435 -18.875 98.765 ;
        RECT -19.205 97.075 -18.875 97.405 ;
        RECT -19.205 95.715 -18.875 96.045 ;
        RECT -19.205 94.355 -18.875 94.685 ;
        RECT -19.205 92.995 -18.875 93.325 ;
        RECT -19.205 91.635 -18.875 91.965 ;
        RECT -19.205 90.275 -18.875 90.605 ;
        RECT -19.205 88.915 -18.875 89.245 ;
        RECT -19.205 87.555 -18.875 87.885 ;
        RECT -19.205 86.195 -18.875 86.525 ;
        RECT -19.205 84.835 -18.875 85.165 ;
        RECT -19.205 83.475 -18.875 83.805 ;
        RECT -19.205 82.115 -18.875 82.445 ;
        RECT -19.205 80.755 -18.875 81.085 ;
        RECT -19.205 79.395 -18.875 79.725 ;
        RECT -19.205 78.035 -18.875 78.365 ;
        RECT -19.205 76.675 -18.875 77.005 ;
        RECT -19.205 75.315 -18.875 75.645 ;
        RECT -19.205 73.955 -18.875 74.285 ;
        RECT -19.205 72.595 -18.875 72.925 ;
        RECT -19.205 71.235 -18.875 71.565 ;
        RECT -19.205 69.875 -18.875 70.205 ;
        RECT -19.205 68.515 -18.875 68.845 ;
        RECT -19.205 67.155 -18.875 67.485 ;
        RECT -19.205 65.795 -18.875 66.125 ;
        RECT -19.205 64.435 -18.875 64.765 ;
        RECT -19.205 63.075 -18.875 63.405 ;
        RECT -19.205 61.715 -18.875 62.045 ;
        RECT -19.205 60.355 -18.875 60.685 ;
        RECT -19.205 58.995 -18.875 59.325 ;
        RECT -19.205 57.635 -18.875 57.965 ;
        RECT -19.205 56.275 -18.875 56.605 ;
        RECT -19.205 54.915 -18.875 55.245 ;
        RECT -19.205 53.555 -18.875 53.885 ;
        RECT -19.205 52.195 -18.875 52.525 ;
        RECT -19.205 50.835 -18.875 51.165 ;
        RECT -19.205 49.475 -18.875 49.805 ;
        RECT -19.205 48.115 -18.875 48.445 ;
        RECT -19.205 46.755 -18.875 47.085 ;
        RECT -19.205 45.395 -18.875 45.725 ;
        RECT -19.205 44.035 -18.875 44.365 ;
        RECT -19.205 42.675 -18.875 43.005 ;
        RECT -19.205 41.315 -18.875 41.645 ;
        RECT -19.205 39.955 -18.875 40.285 ;
        RECT -19.205 38.595 -18.875 38.925 ;
        RECT -19.205 37.235 -18.875 37.565 ;
        RECT -19.205 35.875 -18.875 36.205 ;
        RECT -19.205 34.515 -18.875 34.845 ;
        RECT -19.205 33.155 -18.875 33.485 ;
        RECT -19.205 31.795 -18.875 32.125 ;
        RECT -19.205 30.435 -18.875 30.765 ;
        RECT -19.205 29.075 -18.875 29.405 ;
        RECT -19.205 27.715 -18.875 28.045 ;
        RECT -19.205 26.355 -18.875 26.685 ;
        RECT -19.205 24.995 -18.875 25.325 ;
        RECT -19.205 23.635 -18.875 23.965 ;
        RECT -19.205 22.275 -18.875 22.605 ;
        RECT -19.205 20.915 -18.875 21.245 ;
        RECT -19.205 19.555 -18.875 19.885 ;
        RECT -19.205 18.195 -18.875 18.525 ;
        RECT -19.205 16.835 -18.875 17.165 ;
        RECT -19.205 15.475 -18.875 15.805 ;
        RECT -19.205 14.115 -18.875 14.445 ;
        RECT -19.205 12.755 -18.875 13.085 ;
        RECT -19.205 11.395 -18.875 11.725 ;
        RECT -19.205 10.035 -18.875 10.365 ;
        RECT -19.205 8.675 -18.875 9.005 ;
        RECT -19.205 7.315 -18.875 7.645 ;
        RECT -19.205 5.955 -18.875 6.285 ;
        RECT -19.205 4.595 -18.875 4.925 ;
        RECT -19.205 3.235 -18.875 3.565 ;
        RECT -19.205 1.875 -18.875 2.205 ;
        RECT -19.205 0.515 -18.875 0.845 ;
        RECT -19.205 -0.845 -18.875 -0.515 ;
        RECT -19.205 -2.205 -18.875 -1.875 ;
        RECT -19.205 -3.565 -18.875 -3.235 ;
        RECT -19.205 -7.645 -18.875 -7.315 ;
        RECT -19.205 -9.005 -18.875 -8.675 ;
        RECT -19.205 -10.73 -18.875 -10.4 ;
        RECT -19.205 -11.725 -18.875 -11.395 ;
        RECT -19.205 -16.77 -18.875 -16.44 ;
        RECT -19.205 -18.525 -18.875 -18.195 ;
        RECT -19.205 -21.245 -18.875 -20.915 ;
        RECT -19.2 -21.92 -18.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 -28.045 -18.875 -27.715 ;
        RECT -19.205 -29.405 -18.875 -29.075 ;
        RECT -19.205 -30.765 -18.875 -30.435 ;
        RECT -19.205 -32.125 -18.875 -31.795 ;
        RECT -19.205 -33.71 -18.875 -33.38 ;
        RECT -19.205 -34.845 -18.875 -34.515 ;
        RECT -19.205 -36.205 -18.875 -35.875 ;
        RECT -19.205 -39.75 -18.875 -39.42 ;
        RECT -19.205 -41.645 -18.875 -41.315 ;
        RECT -19.205 -44.365 -18.875 -44.035 ;
        RECT -19.205 -51.165 -18.875 -50.835 ;
        RECT -19.205 -52.525 -18.875 -52.195 ;
        RECT -19.205 -53.885 -18.875 -53.555 ;
        RECT -19.205 -55.245 -18.875 -54.915 ;
        RECT -19.205 -56.605 -18.875 -56.275 ;
        RECT -19.205 -57.965 -18.875 -57.635 ;
        RECT -19.205 -59.325 -18.875 -58.995 ;
        RECT -19.205 -60.685 -18.875 -60.355 ;
        RECT -19.205 -62.045 -18.875 -61.715 ;
        RECT -19.205 -63.405 -18.875 -63.075 ;
        RECT -19.205 -64.765 -18.875 -64.435 ;
        RECT -19.205 -66.125 -18.875 -65.795 ;
        RECT -19.205 -68.845 -18.875 -68.515 ;
        RECT -19.205 -70.205 -18.875 -69.875 ;
        RECT -19.205 -71.565 -18.875 -71.235 ;
        RECT -19.205 -73.19 -18.875 -72.86 ;
        RECT -19.205 -74.285 -18.875 -73.955 ;
        RECT -19.205 -75.645 -18.875 -75.315 ;
        RECT -19.205 -78.365 -18.875 -78.035 ;
        RECT -19.205 -79.725 -18.875 -79.395 ;
        RECT -19.205 -80.73 -18.875 -80.4 ;
        RECT -19.205 -82.445 -18.875 -82.115 ;
        RECT -19.205 -83.805 -18.875 -83.475 ;
        RECT -19.205 -86.525 -18.875 -86.195 ;
        RECT -19.205 -89.245 -18.875 -88.915 ;
        RECT -19.205 -90.605 -18.875 -90.275 ;
        RECT -19.205 -91.965 -18.875 -91.635 ;
        RECT -19.205 -93.325 -18.875 -92.995 ;
        RECT -19.205 -94.685 -18.875 -94.355 ;
        RECT -19.205 -95.37 -18.875 -95.04 ;
        RECT -19.205 -97.405 -18.875 -97.075 ;
        RECT -19.205 -100.125 -18.875 -99.795 ;
        RECT -19.205 -101.485 -18.875 -101.155 ;
        RECT -19.205 -102.91 -18.875 -102.58 ;
        RECT -19.205 -104.205 -18.875 -103.875 ;
        RECT -19.2 -109.64 -18.88 -27.04 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.205 -173.565 -18.875 -173.235 ;
        RECT -19.205 -174.925 -18.875 -174.595 ;
        RECT -19.205 -177.645 -18.875 -177.315 ;
        RECT -19.205 -179.005 -18.875 -178.675 ;
        RECT -19.205 -184.65 -18.875 -183.52 ;
        RECT -19.2 -184.765 -18.88 -173.235 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.845 244.04 -17.515 245.17 ;
        RECT -17.845 239.875 -17.515 240.205 ;
        RECT -17.845 238.515 -17.515 238.845 ;
        RECT -17.845 237.155 -17.515 237.485 ;
        RECT -17.845 235.795 -17.515 236.125 ;
        RECT -17.845 234.435 -17.515 234.765 ;
        RECT -17.845 233.075 -17.515 233.405 ;
        RECT -17.845 231.715 -17.515 232.045 ;
        RECT -17.845 230.355 -17.515 230.685 ;
        RECT -17.845 228.995 -17.515 229.325 ;
        RECT -17.845 227.635 -17.515 227.965 ;
        RECT -17.845 226.275 -17.515 226.605 ;
        RECT -17.845 224.915 -17.515 225.245 ;
        RECT -17.845 223.555 -17.515 223.885 ;
        RECT -17.845 222.195 -17.515 222.525 ;
        RECT -17.845 220.835 -17.515 221.165 ;
        RECT -17.845 219.475 -17.515 219.805 ;
        RECT -17.845 218.115 -17.515 218.445 ;
        RECT -17.845 216.755 -17.515 217.085 ;
        RECT -17.845 215.395 -17.515 215.725 ;
        RECT -17.845 214.035 -17.515 214.365 ;
        RECT -17.845 212.675 -17.515 213.005 ;
        RECT -17.845 211.315 -17.515 211.645 ;
        RECT -17.845 209.955 -17.515 210.285 ;
        RECT -17.845 208.595 -17.515 208.925 ;
        RECT -17.845 207.235 -17.515 207.565 ;
        RECT -17.845 205.875 -17.515 206.205 ;
        RECT -17.845 204.515 -17.515 204.845 ;
        RECT -17.845 203.155 -17.515 203.485 ;
        RECT -17.845 201.795 -17.515 202.125 ;
        RECT -17.845 200.435 -17.515 200.765 ;
        RECT -17.845 199.075 -17.515 199.405 ;
        RECT -17.845 197.715 -17.515 198.045 ;
        RECT -17.845 196.355 -17.515 196.685 ;
        RECT -17.845 194.995 -17.515 195.325 ;
        RECT -17.845 193.635 -17.515 193.965 ;
        RECT -17.845 192.275 -17.515 192.605 ;
        RECT -17.845 190.915 -17.515 191.245 ;
        RECT -17.845 189.555 -17.515 189.885 ;
        RECT -17.845 188.195 -17.515 188.525 ;
        RECT -17.845 186.835 -17.515 187.165 ;
        RECT -17.845 185.475 -17.515 185.805 ;
        RECT -17.845 184.115 -17.515 184.445 ;
        RECT -17.845 182.755 -17.515 183.085 ;
        RECT -17.845 181.395 -17.515 181.725 ;
        RECT -17.845 180.035 -17.515 180.365 ;
        RECT -17.845 178.675 -17.515 179.005 ;
        RECT -17.845 177.315 -17.515 177.645 ;
        RECT -17.845 175.955 -17.515 176.285 ;
        RECT -17.845 174.595 -17.515 174.925 ;
        RECT -17.845 173.235 -17.515 173.565 ;
        RECT -17.845 171.875 -17.515 172.205 ;
        RECT -17.845 170.515 -17.515 170.845 ;
        RECT -17.845 169.155 -17.515 169.485 ;
        RECT -17.845 167.795 -17.515 168.125 ;
        RECT -17.845 166.435 -17.515 166.765 ;
        RECT -17.845 165.075 -17.515 165.405 ;
        RECT -17.845 163.715 -17.515 164.045 ;
        RECT -17.845 162.355 -17.515 162.685 ;
        RECT -17.845 160.995 -17.515 161.325 ;
        RECT -17.845 159.635 -17.515 159.965 ;
        RECT -17.845 158.275 -17.515 158.605 ;
        RECT -17.845 156.915 -17.515 157.245 ;
        RECT -17.845 155.555 -17.515 155.885 ;
        RECT -17.845 154.195 -17.515 154.525 ;
        RECT -17.845 152.835 -17.515 153.165 ;
        RECT -17.845 151.475 -17.515 151.805 ;
        RECT -17.845 150.115 -17.515 150.445 ;
        RECT -17.845 148.755 -17.515 149.085 ;
        RECT -17.845 147.395 -17.515 147.725 ;
        RECT -17.845 146.035 -17.515 146.365 ;
        RECT -17.845 144.675 -17.515 145.005 ;
        RECT -17.845 143.315 -17.515 143.645 ;
        RECT -17.845 141.955 -17.515 142.285 ;
        RECT -17.845 140.595 -17.515 140.925 ;
        RECT -17.845 139.235 -17.515 139.565 ;
        RECT -17.845 137.875 -17.515 138.205 ;
        RECT -17.845 136.515 -17.515 136.845 ;
        RECT -17.845 135.155 -17.515 135.485 ;
        RECT -17.845 133.795 -17.515 134.125 ;
        RECT -17.845 132.435 -17.515 132.765 ;
        RECT -17.845 131.075 -17.515 131.405 ;
        RECT -17.845 129.715 -17.515 130.045 ;
        RECT -17.845 128.355 -17.515 128.685 ;
        RECT -17.845 126.995 -17.515 127.325 ;
        RECT -17.845 125.635 -17.515 125.965 ;
        RECT -17.845 124.275 -17.515 124.605 ;
        RECT -17.845 122.915 -17.515 123.245 ;
        RECT -17.845 121.555 -17.515 121.885 ;
        RECT -17.845 120.195 -17.515 120.525 ;
        RECT -17.845 118.835 -17.515 119.165 ;
        RECT -17.845 117.475 -17.515 117.805 ;
        RECT -17.845 116.115 -17.515 116.445 ;
        RECT -17.845 114.755 -17.515 115.085 ;
        RECT -17.845 113.395 -17.515 113.725 ;
        RECT -17.845 112.035 -17.515 112.365 ;
        RECT -17.845 110.675 -17.515 111.005 ;
        RECT -17.845 109.315 -17.515 109.645 ;
        RECT -17.845 107.955 -17.515 108.285 ;
        RECT -17.845 106.595 -17.515 106.925 ;
        RECT -17.845 105.235 -17.515 105.565 ;
        RECT -17.845 103.875 -17.515 104.205 ;
        RECT -17.845 102.515 -17.515 102.845 ;
        RECT -17.845 101.155 -17.515 101.485 ;
        RECT -17.845 99.795 -17.515 100.125 ;
        RECT -17.845 98.435 -17.515 98.765 ;
        RECT -17.845 97.075 -17.515 97.405 ;
        RECT -17.845 95.715 -17.515 96.045 ;
        RECT -17.845 94.355 -17.515 94.685 ;
        RECT -17.845 92.995 -17.515 93.325 ;
        RECT -17.845 91.635 -17.515 91.965 ;
        RECT -17.845 90.275 -17.515 90.605 ;
        RECT -17.845 88.915 -17.515 89.245 ;
        RECT -17.845 87.555 -17.515 87.885 ;
        RECT -17.845 86.195 -17.515 86.525 ;
        RECT -17.845 84.835 -17.515 85.165 ;
        RECT -17.845 83.475 -17.515 83.805 ;
        RECT -17.845 82.115 -17.515 82.445 ;
        RECT -17.845 80.755 -17.515 81.085 ;
        RECT -17.845 79.395 -17.515 79.725 ;
        RECT -17.845 78.035 -17.515 78.365 ;
        RECT -17.845 76.675 -17.515 77.005 ;
        RECT -17.845 75.315 -17.515 75.645 ;
        RECT -17.845 73.955 -17.515 74.285 ;
        RECT -17.845 72.595 -17.515 72.925 ;
        RECT -17.845 71.235 -17.515 71.565 ;
        RECT -17.845 69.875 -17.515 70.205 ;
        RECT -17.845 68.515 -17.515 68.845 ;
        RECT -17.845 67.155 -17.515 67.485 ;
        RECT -17.845 65.795 -17.515 66.125 ;
        RECT -17.845 64.435 -17.515 64.765 ;
        RECT -17.845 63.075 -17.515 63.405 ;
        RECT -17.845 61.715 -17.515 62.045 ;
        RECT -17.845 60.355 -17.515 60.685 ;
        RECT -17.845 58.995 -17.515 59.325 ;
        RECT -17.845 57.635 -17.515 57.965 ;
        RECT -17.845 56.275 -17.515 56.605 ;
        RECT -17.845 54.915 -17.515 55.245 ;
        RECT -17.845 53.555 -17.515 53.885 ;
        RECT -17.845 52.195 -17.515 52.525 ;
        RECT -17.845 50.835 -17.515 51.165 ;
        RECT -17.845 49.475 -17.515 49.805 ;
        RECT -17.845 48.115 -17.515 48.445 ;
        RECT -17.845 46.755 -17.515 47.085 ;
        RECT -17.845 45.395 -17.515 45.725 ;
        RECT -17.845 44.035 -17.515 44.365 ;
        RECT -17.845 42.675 -17.515 43.005 ;
        RECT -17.845 41.315 -17.515 41.645 ;
        RECT -17.845 39.955 -17.515 40.285 ;
        RECT -17.845 38.595 -17.515 38.925 ;
        RECT -17.845 37.235 -17.515 37.565 ;
        RECT -17.845 35.875 -17.515 36.205 ;
        RECT -17.845 34.515 -17.515 34.845 ;
        RECT -17.845 33.155 -17.515 33.485 ;
        RECT -17.845 31.795 -17.515 32.125 ;
        RECT -17.845 30.435 -17.515 30.765 ;
        RECT -17.845 29.075 -17.515 29.405 ;
        RECT -17.845 27.715 -17.515 28.045 ;
        RECT -17.845 26.355 -17.515 26.685 ;
        RECT -17.845 24.995 -17.515 25.325 ;
        RECT -17.845 23.635 -17.515 23.965 ;
        RECT -17.845 22.275 -17.515 22.605 ;
        RECT -17.845 20.915 -17.515 21.245 ;
        RECT -17.845 19.555 -17.515 19.885 ;
        RECT -17.845 18.195 -17.515 18.525 ;
        RECT -17.845 16.835 -17.515 17.165 ;
        RECT -17.845 15.475 -17.515 15.805 ;
        RECT -17.845 14.115 -17.515 14.445 ;
        RECT -17.845 12.755 -17.515 13.085 ;
        RECT -17.845 11.395 -17.515 11.725 ;
        RECT -17.845 10.035 -17.515 10.365 ;
        RECT -17.845 8.675 -17.515 9.005 ;
        RECT -17.845 7.315 -17.515 7.645 ;
        RECT -17.845 5.955 -17.515 6.285 ;
        RECT -17.845 4.595 -17.515 4.925 ;
        RECT -17.845 3.235 -17.515 3.565 ;
        RECT -17.845 1.875 -17.515 2.205 ;
        RECT -17.845 0.515 -17.515 0.845 ;
        RECT -17.845 -0.845 -17.515 -0.515 ;
        RECT -17.845 -2.205 -17.515 -1.875 ;
        RECT -17.845 -3.565 -17.515 -3.235 ;
        RECT -17.845 -7.645 -17.515 -7.315 ;
        RECT -17.845 -9.005 -17.515 -8.675 ;
        RECT -17.845 -10.73 -17.515 -10.4 ;
        RECT -17.845 -11.725 -17.515 -11.395 ;
        RECT -17.84 -11.725 -17.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.845 -26.685 -17.515 -26.355 ;
        RECT -17.845 -28.045 -17.515 -27.715 ;
        RECT -17.845 -29.405 -17.515 -29.075 ;
        RECT -17.845 -30.765 -17.515 -30.435 ;
        RECT -17.845 -32.125 -17.515 -31.795 ;
        RECT -17.845 -33.71 -17.515 -33.38 ;
        RECT -17.84 -34.16 -17.52 -26.355 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.845 -127.325 -17.515 -126.995 ;
        RECT -17.845 -139.565 -17.515 -139.235 ;
        RECT -17.845 -143.645 -17.515 -143.315 ;
        RECT -17.845 -145.005 -17.515 -144.675 ;
        RECT -17.845 -149.085 -17.515 -148.755 ;
        RECT -17.845 -153.165 -17.515 -152.835 ;
        RECT -17.845 -158.605 -17.515 -158.275 ;
        RECT -17.845 -159.965 -17.515 -159.635 ;
        RECT -17.845 -161.325 -17.515 -160.995 ;
        RECT -17.845 -162.685 -17.515 -162.355 ;
        RECT -17.845 -164.045 -17.515 -163.715 ;
        RECT -17.845 -165.405 -17.515 -165.075 ;
        RECT -17.845 -166.765 -17.515 -166.435 ;
        RECT -17.845 -169.615 -17.515 -169.285 ;
        RECT -17.845 -170.845 -17.515 -170.515 ;
        RECT -17.845 -172.205 -17.515 -171.875 ;
        RECT -17.845 -173.565 -17.515 -173.235 ;
        RECT -17.845 -177.645 -17.515 -177.315 ;
        RECT -17.845 -179.005 -17.515 -178.675 ;
        RECT -17.845 -184.65 -17.515 -183.52 ;
        RECT -17.84 -184.765 -17.52 -120.88 ;
    END
    PORT
      LAYER met3 ;
        RECT -16.485 186.835 -16.155 187.165 ;
        RECT -16.485 185.475 -16.155 185.805 ;
        RECT -16.485 184.115 -16.155 184.445 ;
        RECT -16.485 182.755 -16.155 183.085 ;
        RECT -16.485 181.395 -16.155 181.725 ;
        RECT -16.485 180.035 -16.155 180.365 ;
        RECT -16.485 178.675 -16.155 179.005 ;
        RECT -16.485 177.315 -16.155 177.645 ;
        RECT -16.485 175.955 -16.155 176.285 ;
        RECT -16.485 174.595 -16.155 174.925 ;
        RECT -16.485 173.235 -16.155 173.565 ;
        RECT -16.485 171.875 -16.155 172.205 ;
        RECT -16.485 170.515 -16.155 170.845 ;
        RECT -16.485 169.155 -16.155 169.485 ;
        RECT -16.485 167.795 -16.155 168.125 ;
        RECT -16.485 166.435 -16.155 166.765 ;
        RECT -16.485 165.075 -16.155 165.405 ;
        RECT -16.485 163.715 -16.155 164.045 ;
        RECT -16.485 162.355 -16.155 162.685 ;
        RECT -16.485 160.995 -16.155 161.325 ;
        RECT -16.485 159.635 -16.155 159.965 ;
        RECT -16.485 158.275 -16.155 158.605 ;
        RECT -16.485 156.915 -16.155 157.245 ;
        RECT -16.485 155.555 -16.155 155.885 ;
        RECT -16.485 154.195 -16.155 154.525 ;
        RECT -16.485 152.835 -16.155 153.165 ;
        RECT -16.485 151.475 -16.155 151.805 ;
        RECT -16.485 150.115 -16.155 150.445 ;
        RECT -16.485 148.755 -16.155 149.085 ;
        RECT -16.485 147.395 -16.155 147.725 ;
        RECT -16.485 146.035 -16.155 146.365 ;
        RECT -16.485 144.675 -16.155 145.005 ;
        RECT -16.485 143.315 -16.155 143.645 ;
        RECT -16.485 141.955 -16.155 142.285 ;
        RECT -16.485 140.595 -16.155 140.925 ;
        RECT -16.485 139.235 -16.155 139.565 ;
        RECT -16.485 137.875 -16.155 138.205 ;
        RECT -16.485 136.515 -16.155 136.845 ;
        RECT -16.485 135.155 -16.155 135.485 ;
        RECT -16.485 133.795 -16.155 134.125 ;
        RECT -16.485 132.435 -16.155 132.765 ;
        RECT -16.485 131.075 -16.155 131.405 ;
        RECT -16.485 129.715 -16.155 130.045 ;
        RECT -16.485 128.355 -16.155 128.685 ;
        RECT -16.485 126.995 -16.155 127.325 ;
        RECT -16.485 125.635 -16.155 125.965 ;
        RECT -16.485 124.275 -16.155 124.605 ;
        RECT -16.485 122.915 -16.155 123.245 ;
        RECT -16.485 121.555 -16.155 121.885 ;
        RECT -16.485 120.195 -16.155 120.525 ;
        RECT -16.485 118.835 -16.155 119.165 ;
        RECT -16.485 117.475 -16.155 117.805 ;
        RECT -16.485 116.115 -16.155 116.445 ;
        RECT -16.485 114.755 -16.155 115.085 ;
        RECT -16.485 113.395 -16.155 113.725 ;
        RECT -16.485 112.035 -16.155 112.365 ;
        RECT -16.485 110.675 -16.155 111.005 ;
        RECT -16.485 109.315 -16.155 109.645 ;
        RECT -16.485 107.955 -16.155 108.285 ;
        RECT -16.485 106.595 -16.155 106.925 ;
        RECT -16.485 105.235 -16.155 105.565 ;
        RECT -16.485 103.875 -16.155 104.205 ;
        RECT -16.485 102.515 -16.155 102.845 ;
        RECT -16.485 101.155 -16.155 101.485 ;
        RECT -16.485 99.795 -16.155 100.125 ;
        RECT -16.485 98.435 -16.155 98.765 ;
        RECT -16.485 97.075 -16.155 97.405 ;
        RECT -16.485 95.715 -16.155 96.045 ;
        RECT -16.485 94.355 -16.155 94.685 ;
        RECT -16.485 92.995 -16.155 93.325 ;
        RECT -16.485 91.635 -16.155 91.965 ;
        RECT -16.485 90.275 -16.155 90.605 ;
        RECT -16.485 88.915 -16.155 89.245 ;
        RECT -16.485 87.555 -16.155 87.885 ;
        RECT -16.485 86.195 -16.155 86.525 ;
        RECT -16.485 84.835 -16.155 85.165 ;
        RECT -16.485 83.475 -16.155 83.805 ;
        RECT -16.485 82.115 -16.155 82.445 ;
        RECT -16.485 80.755 -16.155 81.085 ;
        RECT -16.485 79.395 -16.155 79.725 ;
        RECT -16.485 78.035 -16.155 78.365 ;
        RECT -16.485 76.675 -16.155 77.005 ;
        RECT -16.485 75.315 -16.155 75.645 ;
        RECT -16.485 73.955 -16.155 74.285 ;
        RECT -16.485 72.595 -16.155 72.925 ;
        RECT -16.485 71.235 -16.155 71.565 ;
        RECT -16.485 69.875 -16.155 70.205 ;
        RECT -16.485 68.515 -16.155 68.845 ;
        RECT -16.485 67.155 -16.155 67.485 ;
        RECT -16.485 65.795 -16.155 66.125 ;
        RECT -16.485 64.435 -16.155 64.765 ;
        RECT -16.485 63.075 -16.155 63.405 ;
        RECT -16.485 61.715 -16.155 62.045 ;
        RECT -16.485 60.355 -16.155 60.685 ;
        RECT -16.485 58.995 -16.155 59.325 ;
        RECT -16.485 57.635 -16.155 57.965 ;
        RECT -16.485 56.275 -16.155 56.605 ;
        RECT -16.485 54.915 -16.155 55.245 ;
        RECT -16.485 53.555 -16.155 53.885 ;
        RECT -16.485 52.195 -16.155 52.525 ;
        RECT -16.485 50.835 -16.155 51.165 ;
        RECT -16.485 49.475 -16.155 49.805 ;
        RECT -16.485 48.115 -16.155 48.445 ;
        RECT -16.485 46.755 -16.155 47.085 ;
        RECT -16.485 45.395 -16.155 45.725 ;
        RECT -16.485 44.035 -16.155 44.365 ;
        RECT -16.485 42.675 -16.155 43.005 ;
        RECT -16.485 41.315 -16.155 41.645 ;
        RECT -16.485 39.955 -16.155 40.285 ;
        RECT -16.485 38.595 -16.155 38.925 ;
        RECT -16.485 37.235 -16.155 37.565 ;
        RECT -16.485 35.875 -16.155 36.205 ;
        RECT -16.485 34.515 -16.155 34.845 ;
        RECT -16.485 33.155 -16.155 33.485 ;
        RECT -16.485 31.795 -16.155 32.125 ;
        RECT -16.485 30.435 -16.155 30.765 ;
        RECT -16.485 29.075 -16.155 29.405 ;
        RECT -16.485 27.715 -16.155 28.045 ;
        RECT -16.485 26.355 -16.155 26.685 ;
        RECT -16.485 24.995 -16.155 25.325 ;
        RECT -16.485 23.635 -16.155 23.965 ;
        RECT -16.485 22.275 -16.155 22.605 ;
        RECT -16.485 20.915 -16.155 21.245 ;
        RECT -16.485 19.555 -16.155 19.885 ;
        RECT -16.485 18.195 -16.155 18.525 ;
        RECT -16.485 16.835 -16.155 17.165 ;
        RECT -16.485 15.475 -16.155 15.805 ;
        RECT -16.485 14.115 -16.155 14.445 ;
        RECT -16.485 12.755 -16.155 13.085 ;
        RECT -16.485 11.395 -16.155 11.725 ;
        RECT -16.485 10.035 -16.155 10.365 ;
        RECT -16.485 8.675 -16.155 9.005 ;
        RECT -16.485 7.315 -16.155 7.645 ;
        RECT -16.485 5.955 -16.155 6.285 ;
        RECT -16.485 4.595 -16.155 4.925 ;
        RECT -16.485 3.235 -16.155 3.565 ;
        RECT -16.485 1.875 -16.155 2.205 ;
        RECT -16.485 0.515 -16.155 0.845 ;
        RECT -16.485 -0.845 -16.155 -0.515 ;
        RECT -16.485 -2.205 -16.155 -1.875 ;
        RECT -16.485 -3.565 -16.155 -3.235 ;
        RECT -16.485 -4.925 -16.155 -4.595 ;
        RECT -16.485 -7.645 -16.155 -7.315 ;
        RECT -16.485 -9.005 -16.155 -8.675 ;
        RECT -16.485 -10.73 -16.155 -10.4 ;
        RECT -16.485 -11.725 -16.155 -11.395 ;
        RECT -16.485 -13.085 -16.155 -12.755 ;
        RECT -16.48 -13.085 -16.16 245.285 ;
        RECT -16.485 244.04 -16.155 245.17 ;
        RECT -16.485 239.875 -16.155 240.205 ;
        RECT -16.485 238.515 -16.155 238.845 ;
        RECT -16.485 237.155 -16.155 237.485 ;
        RECT -16.485 235.795 -16.155 236.125 ;
        RECT -16.485 234.435 -16.155 234.765 ;
        RECT -16.485 233.075 -16.155 233.405 ;
        RECT -16.485 231.715 -16.155 232.045 ;
        RECT -16.485 230.355 -16.155 230.685 ;
        RECT -16.485 228.995 -16.155 229.325 ;
        RECT -16.485 227.635 -16.155 227.965 ;
        RECT -16.485 226.275 -16.155 226.605 ;
        RECT -16.485 224.915 -16.155 225.245 ;
        RECT -16.485 223.555 -16.155 223.885 ;
        RECT -16.485 222.195 -16.155 222.525 ;
        RECT -16.485 220.835 -16.155 221.165 ;
        RECT -16.485 219.475 -16.155 219.805 ;
        RECT -16.485 218.115 -16.155 218.445 ;
        RECT -16.485 216.755 -16.155 217.085 ;
        RECT -16.485 215.395 -16.155 215.725 ;
        RECT -16.485 214.035 -16.155 214.365 ;
        RECT -16.485 212.675 -16.155 213.005 ;
        RECT -16.485 211.315 -16.155 211.645 ;
        RECT -16.485 209.955 -16.155 210.285 ;
        RECT -16.485 208.595 -16.155 208.925 ;
        RECT -16.485 207.235 -16.155 207.565 ;
        RECT -16.485 205.875 -16.155 206.205 ;
        RECT -16.485 204.515 -16.155 204.845 ;
        RECT -16.485 203.155 -16.155 203.485 ;
        RECT -16.485 201.795 -16.155 202.125 ;
        RECT -16.485 200.435 -16.155 200.765 ;
        RECT -16.485 199.075 -16.155 199.405 ;
        RECT -16.485 197.715 -16.155 198.045 ;
        RECT -16.485 196.355 -16.155 196.685 ;
        RECT -16.485 194.995 -16.155 195.325 ;
        RECT -16.485 193.635 -16.155 193.965 ;
        RECT -16.485 192.275 -16.155 192.605 ;
        RECT -16.485 190.915 -16.155 191.245 ;
        RECT -16.485 189.555 -16.155 189.885 ;
        RECT -16.485 188.195 -16.155 188.525 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.365 -32.125 -27.035 -31.795 ;
        RECT -27.365 -33.71 -27.035 -33.38 ;
        RECT -27.365 -34.845 -27.035 -34.515 ;
        RECT -27.365 -36.205 -27.035 -35.875 ;
        RECT -27.365 -38.925 -27.035 -38.595 ;
        RECT -27.365 -39.75 -27.035 -39.42 ;
        RECT -27.365 -41.645 -27.035 -41.315 ;
        RECT -27.365 -44.365 -27.035 -44.035 ;
        RECT -27.365 -49.805 -27.035 -49.475 ;
        RECT -27.365 -51.165 -27.035 -50.835 ;
        RECT -27.365 -53.885 -27.035 -53.555 ;
        RECT -27.365 -55.245 -27.035 -54.915 ;
        RECT -27.365 -59.325 -27.035 -58.995 ;
        RECT -27.365 -60.685 -27.035 -60.355 ;
        RECT -27.365 -63.405 -27.035 -63.075 ;
        RECT -27.365 -67.485 -27.035 -67.155 ;
        RECT -27.365 -68.845 -27.035 -68.515 ;
        RECT -27.365 -70.205 -27.035 -69.875 ;
        RECT -27.365 -71.565 -27.035 -71.235 ;
        RECT -27.365 -73.19 -27.035 -72.86 ;
        RECT -27.365 -74.285 -27.035 -73.955 ;
        RECT -27.365 -75.645 -27.035 -75.315 ;
        RECT -27.365 -78.365 -27.035 -78.035 ;
        RECT -27.365 -79.725 -27.035 -79.395 ;
        RECT -27.365 -80.73 -27.035 -80.4 ;
        RECT -27.365 -82.445 -27.035 -82.115 ;
        RECT -27.365 -83.805 -27.035 -83.475 ;
        RECT -27.365 -86.525 -27.035 -86.195 ;
        RECT -27.365 -89.245 -27.035 -88.915 ;
        RECT -27.365 -90.605 -27.035 -90.275 ;
        RECT -27.365 -91.965 -27.035 -91.635 ;
        RECT -27.365 -93.325 -27.035 -92.995 ;
        RECT -27.365 -94.685 -27.035 -94.355 ;
        RECT -27.365 -95.37 -27.035 -95.04 ;
        RECT -27.365 -97.405 -27.035 -97.075 ;
        RECT -27.365 -100.125 -27.035 -99.795 ;
        RECT -27.365 -101.485 -27.035 -101.155 ;
        RECT -27.365 -102.91 -27.035 -102.58 ;
        RECT -27.365 -104.205 -27.035 -103.875 ;
        RECT -27.365 -105.565 -27.035 -105.235 ;
        RECT -27.365 -108.285 -27.035 -107.955 ;
        RECT -27.365 -115.085 -27.035 -114.755 ;
        RECT -27.365 -116.445 -27.035 -116.115 ;
        RECT -27.365 -117.805 -27.035 -117.475 ;
        RECT -27.365 -119.165 -27.035 -118.835 ;
        RECT -27.365 -120.525 -27.035 -120.195 ;
        RECT -27.365 -123.245 -27.035 -122.915 ;
        RECT -27.365 -125.965 -27.035 -125.635 ;
        RECT -27.365 -127.325 -27.035 -126.995 ;
        RECT -27.365 -128.685 -27.035 -128.355 ;
        RECT -27.365 -130.045 -27.035 -129.715 ;
        RECT -27.365 -134.125 -27.035 -133.795 ;
        RECT -27.365 -135.485 -27.035 -135.155 ;
        RECT -27.365 -136.845 -27.035 -136.515 ;
        RECT -27.365 -139.565 -27.035 -139.235 ;
        RECT -27.365 -142.285 -27.035 -141.955 ;
        RECT -27.365 -143.645 -27.035 -143.315 ;
        RECT -27.365 -145.005 -27.035 -144.675 ;
        RECT -27.365 -146.365 -27.035 -146.035 ;
        RECT -27.365 -147.725 -27.035 -147.395 ;
        RECT -27.365 -149.085 -27.035 -148.755 ;
        RECT -27.365 -151.805 -27.035 -151.475 ;
        RECT -27.365 -153.165 -27.035 -152.835 ;
        RECT -27.365 -157.245 -27.035 -156.915 ;
        RECT -27.365 -158.605 -27.035 -158.275 ;
        RECT -27.365 -159.965 -27.035 -159.635 ;
        RECT -27.365 -161.325 -27.035 -160.995 ;
        RECT -27.365 -162.685 -27.035 -162.355 ;
        RECT -27.365 -164.045 -27.035 -163.715 ;
        RECT -27.365 -165.405 -27.035 -165.075 ;
        RECT -27.365 -166.765 -27.035 -166.435 ;
        RECT -27.365 -169.615 -27.035 -169.285 ;
        RECT -27.365 -170.845 -27.035 -170.515 ;
        RECT -27.365 -172.205 -27.035 -171.875 ;
        RECT -27.365 -177.645 -27.035 -177.315 ;
        RECT -27.365 -179.005 -27.035 -178.675 ;
        RECT -27.365 -184.65 -27.035 -183.52 ;
        RECT -27.36 -184.765 -27.04 -30.44 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.005 244.04 -25.675 245.17 ;
        RECT -26.005 239.875 -25.675 240.205 ;
        RECT -26.005 238.515 -25.675 238.845 ;
        RECT -26.005 237.155 -25.675 237.485 ;
        RECT -26.005 235.795 -25.675 236.125 ;
        RECT -26.005 234.435 -25.675 234.765 ;
        RECT -26.005 233.075 -25.675 233.405 ;
        RECT -26.005 231.715 -25.675 232.045 ;
        RECT -26.005 230.355 -25.675 230.685 ;
        RECT -26.005 228.995 -25.675 229.325 ;
        RECT -26.005 227.635 -25.675 227.965 ;
        RECT -26.005 226.275 -25.675 226.605 ;
        RECT -26.005 224.915 -25.675 225.245 ;
        RECT -26.005 223.555 -25.675 223.885 ;
        RECT -26.005 222.195 -25.675 222.525 ;
        RECT -26.005 220.835 -25.675 221.165 ;
        RECT -26.005 219.475 -25.675 219.805 ;
        RECT -26.005 218.115 -25.675 218.445 ;
        RECT -26.005 216.755 -25.675 217.085 ;
        RECT -26.005 215.395 -25.675 215.725 ;
        RECT -26.005 214.035 -25.675 214.365 ;
        RECT -26.005 212.675 -25.675 213.005 ;
        RECT -26.005 211.315 -25.675 211.645 ;
        RECT -26.005 209.955 -25.675 210.285 ;
        RECT -26.005 208.595 -25.675 208.925 ;
        RECT -26.005 207.235 -25.675 207.565 ;
        RECT -26.005 205.875 -25.675 206.205 ;
        RECT -26.005 204.515 -25.675 204.845 ;
        RECT -26.005 203.155 -25.675 203.485 ;
        RECT -26.005 201.795 -25.675 202.125 ;
        RECT -26.005 200.435 -25.675 200.765 ;
        RECT -26.005 199.075 -25.675 199.405 ;
        RECT -26.005 197.715 -25.675 198.045 ;
        RECT -26.005 196.355 -25.675 196.685 ;
        RECT -26.005 194.995 -25.675 195.325 ;
        RECT -26.005 193.635 -25.675 193.965 ;
        RECT -26.005 192.275 -25.675 192.605 ;
        RECT -26.005 190.915 -25.675 191.245 ;
        RECT -26.005 189.555 -25.675 189.885 ;
        RECT -26.005 188.195 -25.675 188.525 ;
        RECT -26.005 186.835 -25.675 187.165 ;
        RECT -26.005 185.475 -25.675 185.805 ;
        RECT -26.005 184.115 -25.675 184.445 ;
        RECT -26.005 182.755 -25.675 183.085 ;
        RECT -26.005 181.395 -25.675 181.725 ;
        RECT -26.005 180.035 -25.675 180.365 ;
        RECT -26.005 178.675 -25.675 179.005 ;
        RECT -26.005 177.315 -25.675 177.645 ;
        RECT -26.005 175.955 -25.675 176.285 ;
        RECT -26.005 174.595 -25.675 174.925 ;
        RECT -26.005 173.235 -25.675 173.565 ;
        RECT -26.005 171.875 -25.675 172.205 ;
        RECT -26.005 170.515 -25.675 170.845 ;
        RECT -26.005 169.155 -25.675 169.485 ;
        RECT -26.005 167.795 -25.675 168.125 ;
        RECT -26.005 166.435 -25.675 166.765 ;
        RECT -26.005 165.075 -25.675 165.405 ;
        RECT -26.005 163.715 -25.675 164.045 ;
        RECT -26.005 162.355 -25.675 162.685 ;
        RECT -26.005 160.995 -25.675 161.325 ;
        RECT -26.005 159.635 -25.675 159.965 ;
        RECT -26.005 158.275 -25.675 158.605 ;
        RECT -26.005 156.915 -25.675 157.245 ;
        RECT -26.005 155.555 -25.675 155.885 ;
        RECT -26.005 154.195 -25.675 154.525 ;
        RECT -26.005 152.835 -25.675 153.165 ;
        RECT -26.005 151.475 -25.675 151.805 ;
        RECT -26.005 150.115 -25.675 150.445 ;
        RECT -26.005 148.755 -25.675 149.085 ;
        RECT -26.005 147.395 -25.675 147.725 ;
        RECT -26.005 146.035 -25.675 146.365 ;
        RECT -26.005 144.675 -25.675 145.005 ;
        RECT -26.005 143.315 -25.675 143.645 ;
        RECT -26.005 141.955 -25.675 142.285 ;
        RECT -26.005 140.595 -25.675 140.925 ;
        RECT -26.005 139.235 -25.675 139.565 ;
        RECT -26.005 137.875 -25.675 138.205 ;
        RECT -26.005 136.515 -25.675 136.845 ;
        RECT -26.005 135.155 -25.675 135.485 ;
        RECT -26.005 133.795 -25.675 134.125 ;
        RECT -26.005 132.435 -25.675 132.765 ;
        RECT -26.005 131.075 -25.675 131.405 ;
        RECT -26.005 129.715 -25.675 130.045 ;
        RECT -26.005 128.355 -25.675 128.685 ;
        RECT -26.005 126.995 -25.675 127.325 ;
        RECT -26.005 125.635 -25.675 125.965 ;
        RECT -26.005 124.275 -25.675 124.605 ;
        RECT -26.005 122.915 -25.675 123.245 ;
        RECT -26.005 121.555 -25.675 121.885 ;
        RECT -26.005 120.195 -25.675 120.525 ;
        RECT -26.005 118.835 -25.675 119.165 ;
        RECT -26.005 117.475 -25.675 117.805 ;
        RECT -26.005 116.115 -25.675 116.445 ;
        RECT -26.005 114.755 -25.675 115.085 ;
        RECT -26.005 113.395 -25.675 113.725 ;
        RECT -26.005 112.035 -25.675 112.365 ;
        RECT -26.005 110.675 -25.675 111.005 ;
        RECT -26.005 109.315 -25.675 109.645 ;
        RECT -26.005 107.955 -25.675 108.285 ;
        RECT -26.005 106.595 -25.675 106.925 ;
        RECT -26.005 105.235 -25.675 105.565 ;
        RECT -26.005 103.875 -25.675 104.205 ;
        RECT -26.005 102.515 -25.675 102.845 ;
        RECT -26.005 101.155 -25.675 101.485 ;
        RECT -26.005 99.795 -25.675 100.125 ;
        RECT -26.005 98.435 -25.675 98.765 ;
        RECT -26.005 97.075 -25.675 97.405 ;
        RECT -26.005 95.715 -25.675 96.045 ;
        RECT -26.005 94.355 -25.675 94.685 ;
        RECT -26.005 92.995 -25.675 93.325 ;
        RECT -26.005 91.635 -25.675 91.965 ;
        RECT -26.005 90.275 -25.675 90.605 ;
        RECT -26.005 88.915 -25.675 89.245 ;
        RECT -26.005 87.555 -25.675 87.885 ;
        RECT -26.005 86.195 -25.675 86.525 ;
        RECT -26.005 84.835 -25.675 85.165 ;
        RECT -26.005 83.475 -25.675 83.805 ;
        RECT -26.005 82.115 -25.675 82.445 ;
        RECT -26.005 80.755 -25.675 81.085 ;
        RECT -26.005 79.395 -25.675 79.725 ;
        RECT -26.005 78.035 -25.675 78.365 ;
        RECT -26.005 76.675 -25.675 77.005 ;
        RECT -26.005 75.315 -25.675 75.645 ;
        RECT -26.005 73.955 -25.675 74.285 ;
        RECT -26.005 72.595 -25.675 72.925 ;
        RECT -26.005 71.235 -25.675 71.565 ;
        RECT -26.005 69.875 -25.675 70.205 ;
        RECT -26.005 68.515 -25.675 68.845 ;
        RECT -26.005 67.155 -25.675 67.485 ;
        RECT -26.005 65.795 -25.675 66.125 ;
        RECT -26.005 64.435 -25.675 64.765 ;
        RECT -26.005 63.075 -25.675 63.405 ;
        RECT -26.005 61.715 -25.675 62.045 ;
        RECT -26.005 60.355 -25.675 60.685 ;
        RECT -26.005 58.995 -25.675 59.325 ;
        RECT -26.005 57.635 -25.675 57.965 ;
        RECT -26.005 56.275 -25.675 56.605 ;
        RECT -26.005 54.915 -25.675 55.245 ;
        RECT -26.005 53.555 -25.675 53.885 ;
        RECT -26.005 52.195 -25.675 52.525 ;
        RECT -26.005 50.835 -25.675 51.165 ;
        RECT -26.005 49.475 -25.675 49.805 ;
        RECT -26.005 48.115 -25.675 48.445 ;
        RECT -26.005 46.755 -25.675 47.085 ;
        RECT -26.005 45.395 -25.675 45.725 ;
        RECT -26.005 44.035 -25.675 44.365 ;
        RECT -26.005 42.675 -25.675 43.005 ;
        RECT -26.005 41.315 -25.675 41.645 ;
        RECT -26.005 39.955 -25.675 40.285 ;
        RECT -26.005 38.595 -25.675 38.925 ;
        RECT -26.005 37.235 -25.675 37.565 ;
        RECT -26.005 35.875 -25.675 36.205 ;
        RECT -26.005 34.515 -25.675 34.845 ;
        RECT -26.005 33.155 -25.675 33.485 ;
        RECT -26.005 31.795 -25.675 32.125 ;
        RECT -26.005 30.435 -25.675 30.765 ;
        RECT -26.005 29.075 -25.675 29.405 ;
        RECT -26.005 27.715 -25.675 28.045 ;
        RECT -26.005 26.355 -25.675 26.685 ;
        RECT -26.005 24.995 -25.675 25.325 ;
        RECT -26.005 23.635 -25.675 23.965 ;
        RECT -26.005 22.275 -25.675 22.605 ;
        RECT -26.005 20.915 -25.675 21.245 ;
        RECT -26.005 19.555 -25.675 19.885 ;
        RECT -26.005 18.195 -25.675 18.525 ;
        RECT -26.005 16.835 -25.675 17.165 ;
        RECT -26.005 15.475 -25.675 15.805 ;
        RECT -26.005 14.115 -25.675 14.445 ;
        RECT -26.005 12.755 -25.675 13.085 ;
        RECT -26.005 11.395 -25.675 11.725 ;
        RECT -26.005 10.035 -25.675 10.365 ;
        RECT -26.005 8.675 -25.675 9.005 ;
        RECT -26.005 7.315 -25.675 7.645 ;
        RECT -26.005 5.955 -25.675 6.285 ;
        RECT -26.005 4.595 -25.675 4.925 ;
        RECT -26.005 3.235 -25.675 3.565 ;
        RECT -26.005 1.875 -25.675 2.205 ;
        RECT -26.005 0.515 -25.675 0.845 ;
        RECT -26.005 -0.845 -25.675 -0.515 ;
        RECT -26.005 -2.205 -25.675 -1.875 ;
        RECT -26.005 -7.645 -25.675 -7.315 ;
        RECT -26.005 -9.005 -25.675 -8.675 ;
        RECT -26.005 -10.73 -25.675 -10.4 ;
        RECT -26.005 -11.725 -25.675 -11.395 ;
        RECT -26.005 -16.77 -25.675 -16.44 ;
        RECT -26.005 -18.525 -25.675 -18.195 ;
        RECT -26.005 -21.245 -25.675 -20.915 ;
        RECT -26.005 -30.765 -25.675 -30.435 ;
        RECT -26.005 -32.125 -25.675 -31.795 ;
        RECT -26.005 -33.71 -25.675 -33.38 ;
        RECT -26.005 -34.845 -25.675 -34.515 ;
        RECT -26.005 -36.205 -25.675 -35.875 ;
        RECT -26.005 -38.925 -25.675 -38.595 ;
        RECT -26.005 -39.75 -25.675 -39.42 ;
        RECT -26.005 -41.645 -25.675 -41.315 ;
        RECT -26.005 -44.365 -25.675 -44.035 ;
        RECT -26.005 -49.805 -25.675 -49.475 ;
        RECT -26.005 -51.165 -25.675 -50.835 ;
        RECT -26.005 -53.885 -25.675 -53.555 ;
        RECT -26.005 -55.245 -25.675 -54.915 ;
        RECT -26.005 -59.325 -25.675 -58.995 ;
        RECT -26.005 -60.685 -25.675 -60.355 ;
        RECT -26.005 -63.405 -25.675 -63.075 ;
        RECT -26.005 -68.845 -25.675 -68.515 ;
        RECT -26.005 -70.205 -25.675 -69.875 ;
        RECT -26.005 -71.565 -25.675 -71.235 ;
        RECT -26.005 -73.19 -25.675 -72.86 ;
        RECT -26.005 -74.285 -25.675 -73.955 ;
        RECT -26.005 -75.645 -25.675 -75.315 ;
        RECT -26.005 -78.365 -25.675 -78.035 ;
        RECT -26.005 -79.725 -25.675 -79.395 ;
        RECT -26.005 -80.73 -25.675 -80.4 ;
        RECT -26.005 -82.445 -25.675 -82.115 ;
        RECT -26.005 -83.805 -25.675 -83.475 ;
        RECT -26.005 -86.525 -25.675 -86.195 ;
        RECT -26.005 -89.245 -25.675 -88.915 ;
        RECT -26.005 -90.605 -25.675 -90.275 ;
        RECT -26.005 -91.965 -25.675 -91.635 ;
        RECT -26.005 -93.325 -25.675 -92.995 ;
        RECT -26.005 -94.685 -25.675 -94.355 ;
        RECT -26.005 -95.37 -25.675 -95.04 ;
        RECT -26.005 -97.405 -25.675 -97.075 ;
        RECT -26.005 -100.125 -25.675 -99.795 ;
        RECT -26.005 -101.485 -25.675 -101.155 ;
        RECT -26.005 -102.91 -25.675 -102.58 ;
        RECT -26.005 -104.205 -25.675 -103.875 ;
        RECT -26.005 -105.565 -25.675 -105.235 ;
        RECT -26.005 -115.085 -25.675 -114.755 ;
        RECT -26.005 -116.445 -25.675 -116.115 ;
        RECT -26.005 -117.805 -25.675 -117.475 ;
        RECT -26.005 -119.165 -25.675 -118.835 ;
        RECT -26.005 -120.525 -25.675 -120.195 ;
        RECT -26.005 -123.245 -25.675 -122.915 ;
        RECT -26.005 -124.605 -25.675 -124.275 ;
        RECT -26.005 -125.965 -25.675 -125.635 ;
        RECT -26.005 -127.325 -25.675 -126.995 ;
        RECT -26.005 -128.685 -25.675 -128.355 ;
        RECT -26.005 -130.045 -25.675 -129.715 ;
        RECT -26.005 -135.485 -25.675 -135.155 ;
        RECT -26.005 -136.845 -25.675 -136.515 ;
        RECT -26.005 -139.565 -25.675 -139.235 ;
        RECT -26.005 -142.285 -25.675 -141.955 ;
        RECT -26.005 -143.645 -25.675 -143.315 ;
        RECT -26.005 -145.005 -25.675 -144.675 ;
        RECT -26.005 -147.725 -25.675 -147.395 ;
        RECT -26.005 -149.085 -25.675 -148.755 ;
        RECT -26.005 -151.805 -25.675 -151.475 ;
        RECT -26.005 -153.165 -25.675 -152.835 ;
        RECT -26.005 -157.245 -25.675 -156.915 ;
        RECT -26.005 -158.605 -25.675 -158.275 ;
        RECT -26.005 -159.965 -25.675 -159.635 ;
        RECT -26.005 -161.325 -25.675 -160.995 ;
        RECT -26.005 -162.685 -25.675 -162.355 ;
        RECT -26.005 -164.045 -25.675 -163.715 ;
        RECT -26.005 -165.405 -25.675 -165.075 ;
        RECT -26.005 -166.765 -25.675 -166.435 ;
        RECT -26.005 -169.615 -25.675 -169.285 ;
        RECT -26.005 -170.845 -25.675 -170.515 ;
        RECT -26.005 -172.205 -25.675 -171.875 ;
        RECT -26.005 -177.645 -25.675 -177.315 ;
        RECT -26.005 -179.005 -25.675 -178.675 ;
        RECT -26.005 -184.65 -25.675 -183.52 ;
        RECT -26 -184.765 -25.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.645 244.04 -24.315 245.17 ;
        RECT -24.645 239.875 -24.315 240.205 ;
        RECT -24.645 238.515 -24.315 238.845 ;
        RECT -24.645 237.155 -24.315 237.485 ;
        RECT -24.645 235.795 -24.315 236.125 ;
        RECT -24.645 234.435 -24.315 234.765 ;
        RECT -24.645 233.075 -24.315 233.405 ;
        RECT -24.645 231.715 -24.315 232.045 ;
        RECT -24.645 230.355 -24.315 230.685 ;
        RECT -24.645 228.995 -24.315 229.325 ;
        RECT -24.645 227.635 -24.315 227.965 ;
        RECT -24.645 226.275 -24.315 226.605 ;
        RECT -24.645 224.915 -24.315 225.245 ;
        RECT -24.645 223.555 -24.315 223.885 ;
        RECT -24.645 222.195 -24.315 222.525 ;
        RECT -24.645 220.835 -24.315 221.165 ;
        RECT -24.645 219.475 -24.315 219.805 ;
        RECT -24.645 218.115 -24.315 218.445 ;
        RECT -24.645 216.755 -24.315 217.085 ;
        RECT -24.645 215.395 -24.315 215.725 ;
        RECT -24.645 214.035 -24.315 214.365 ;
        RECT -24.645 212.675 -24.315 213.005 ;
        RECT -24.645 211.315 -24.315 211.645 ;
        RECT -24.645 209.955 -24.315 210.285 ;
        RECT -24.645 208.595 -24.315 208.925 ;
        RECT -24.645 207.235 -24.315 207.565 ;
        RECT -24.645 205.875 -24.315 206.205 ;
        RECT -24.645 204.515 -24.315 204.845 ;
        RECT -24.645 203.155 -24.315 203.485 ;
        RECT -24.645 201.795 -24.315 202.125 ;
        RECT -24.645 200.435 -24.315 200.765 ;
        RECT -24.645 199.075 -24.315 199.405 ;
        RECT -24.645 197.715 -24.315 198.045 ;
        RECT -24.645 196.355 -24.315 196.685 ;
        RECT -24.645 194.995 -24.315 195.325 ;
        RECT -24.645 193.635 -24.315 193.965 ;
        RECT -24.645 192.275 -24.315 192.605 ;
        RECT -24.645 190.915 -24.315 191.245 ;
        RECT -24.645 189.555 -24.315 189.885 ;
        RECT -24.645 188.195 -24.315 188.525 ;
        RECT -24.645 186.835 -24.315 187.165 ;
        RECT -24.645 185.475 -24.315 185.805 ;
        RECT -24.645 184.115 -24.315 184.445 ;
        RECT -24.645 182.755 -24.315 183.085 ;
        RECT -24.645 181.395 -24.315 181.725 ;
        RECT -24.645 180.035 -24.315 180.365 ;
        RECT -24.645 178.675 -24.315 179.005 ;
        RECT -24.645 177.315 -24.315 177.645 ;
        RECT -24.645 175.955 -24.315 176.285 ;
        RECT -24.645 174.595 -24.315 174.925 ;
        RECT -24.645 173.235 -24.315 173.565 ;
        RECT -24.645 171.875 -24.315 172.205 ;
        RECT -24.645 170.515 -24.315 170.845 ;
        RECT -24.645 169.155 -24.315 169.485 ;
        RECT -24.645 167.795 -24.315 168.125 ;
        RECT -24.645 166.435 -24.315 166.765 ;
        RECT -24.645 165.075 -24.315 165.405 ;
        RECT -24.645 163.715 -24.315 164.045 ;
        RECT -24.645 162.355 -24.315 162.685 ;
        RECT -24.645 160.995 -24.315 161.325 ;
        RECT -24.645 159.635 -24.315 159.965 ;
        RECT -24.645 158.275 -24.315 158.605 ;
        RECT -24.645 156.915 -24.315 157.245 ;
        RECT -24.645 155.555 -24.315 155.885 ;
        RECT -24.645 154.195 -24.315 154.525 ;
        RECT -24.645 152.835 -24.315 153.165 ;
        RECT -24.645 151.475 -24.315 151.805 ;
        RECT -24.645 150.115 -24.315 150.445 ;
        RECT -24.645 148.755 -24.315 149.085 ;
        RECT -24.645 147.395 -24.315 147.725 ;
        RECT -24.645 146.035 -24.315 146.365 ;
        RECT -24.645 144.675 -24.315 145.005 ;
        RECT -24.645 143.315 -24.315 143.645 ;
        RECT -24.645 141.955 -24.315 142.285 ;
        RECT -24.645 140.595 -24.315 140.925 ;
        RECT -24.645 139.235 -24.315 139.565 ;
        RECT -24.645 137.875 -24.315 138.205 ;
        RECT -24.645 136.515 -24.315 136.845 ;
        RECT -24.645 135.155 -24.315 135.485 ;
        RECT -24.645 133.795 -24.315 134.125 ;
        RECT -24.645 132.435 -24.315 132.765 ;
        RECT -24.645 131.075 -24.315 131.405 ;
        RECT -24.645 129.715 -24.315 130.045 ;
        RECT -24.645 128.355 -24.315 128.685 ;
        RECT -24.645 126.995 -24.315 127.325 ;
        RECT -24.645 125.635 -24.315 125.965 ;
        RECT -24.645 124.275 -24.315 124.605 ;
        RECT -24.645 122.915 -24.315 123.245 ;
        RECT -24.645 121.555 -24.315 121.885 ;
        RECT -24.645 120.195 -24.315 120.525 ;
        RECT -24.645 118.835 -24.315 119.165 ;
        RECT -24.645 117.475 -24.315 117.805 ;
        RECT -24.645 116.115 -24.315 116.445 ;
        RECT -24.645 114.755 -24.315 115.085 ;
        RECT -24.645 113.395 -24.315 113.725 ;
        RECT -24.645 112.035 -24.315 112.365 ;
        RECT -24.645 110.675 -24.315 111.005 ;
        RECT -24.645 109.315 -24.315 109.645 ;
        RECT -24.645 107.955 -24.315 108.285 ;
        RECT -24.645 106.595 -24.315 106.925 ;
        RECT -24.645 105.235 -24.315 105.565 ;
        RECT -24.645 103.875 -24.315 104.205 ;
        RECT -24.645 102.515 -24.315 102.845 ;
        RECT -24.645 101.155 -24.315 101.485 ;
        RECT -24.645 99.795 -24.315 100.125 ;
        RECT -24.645 98.435 -24.315 98.765 ;
        RECT -24.645 97.075 -24.315 97.405 ;
        RECT -24.645 95.715 -24.315 96.045 ;
        RECT -24.645 94.355 -24.315 94.685 ;
        RECT -24.645 92.995 -24.315 93.325 ;
        RECT -24.645 91.635 -24.315 91.965 ;
        RECT -24.645 90.275 -24.315 90.605 ;
        RECT -24.645 88.915 -24.315 89.245 ;
        RECT -24.645 87.555 -24.315 87.885 ;
        RECT -24.645 86.195 -24.315 86.525 ;
        RECT -24.645 84.835 -24.315 85.165 ;
        RECT -24.645 83.475 -24.315 83.805 ;
        RECT -24.645 82.115 -24.315 82.445 ;
        RECT -24.645 80.755 -24.315 81.085 ;
        RECT -24.645 79.395 -24.315 79.725 ;
        RECT -24.645 78.035 -24.315 78.365 ;
        RECT -24.645 76.675 -24.315 77.005 ;
        RECT -24.645 75.315 -24.315 75.645 ;
        RECT -24.645 73.955 -24.315 74.285 ;
        RECT -24.645 72.595 -24.315 72.925 ;
        RECT -24.645 71.235 -24.315 71.565 ;
        RECT -24.645 69.875 -24.315 70.205 ;
        RECT -24.645 68.515 -24.315 68.845 ;
        RECT -24.645 67.155 -24.315 67.485 ;
        RECT -24.645 65.795 -24.315 66.125 ;
        RECT -24.645 64.435 -24.315 64.765 ;
        RECT -24.645 63.075 -24.315 63.405 ;
        RECT -24.645 61.715 -24.315 62.045 ;
        RECT -24.645 60.355 -24.315 60.685 ;
        RECT -24.645 58.995 -24.315 59.325 ;
        RECT -24.645 57.635 -24.315 57.965 ;
        RECT -24.645 56.275 -24.315 56.605 ;
        RECT -24.645 54.915 -24.315 55.245 ;
        RECT -24.645 53.555 -24.315 53.885 ;
        RECT -24.645 52.195 -24.315 52.525 ;
        RECT -24.645 50.835 -24.315 51.165 ;
        RECT -24.645 49.475 -24.315 49.805 ;
        RECT -24.645 48.115 -24.315 48.445 ;
        RECT -24.645 46.755 -24.315 47.085 ;
        RECT -24.645 45.395 -24.315 45.725 ;
        RECT -24.645 44.035 -24.315 44.365 ;
        RECT -24.645 42.675 -24.315 43.005 ;
        RECT -24.645 41.315 -24.315 41.645 ;
        RECT -24.645 39.955 -24.315 40.285 ;
        RECT -24.645 38.595 -24.315 38.925 ;
        RECT -24.645 37.235 -24.315 37.565 ;
        RECT -24.645 35.875 -24.315 36.205 ;
        RECT -24.645 34.515 -24.315 34.845 ;
        RECT -24.645 33.155 -24.315 33.485 ;
        RECT -24.645 31.795 -24.315 32.125 ;
        RECT -24.645 30.435 -24.315 30.765 ;
        RECT -24.645 29.075 -24.315 29.405 ;
        RECT -24.645 27.715 -24.315 28.045 ;
        RECT -24.645 26.355 -24.315 26.685 ;
        RECT -24.645 24.995 -24.315 25.325 ;
        RECT -24.645 23.635 -24.315 23.965 ;
        RECT -24.645 22.275 -24.315 22.605 ;
        RECT -24.645 20.915 -24.315 21.245 ;
        RECT -24.645 19.555 -24.315 19.885 ;
        RECT -24.645 18.195 -24.315 18.525 ;
        RECT -24.645 16.835 -24.315 17.165 ;
        RECT -24.645 15.475 -24.315 15.805 ;
        RECT -24.645 14.115 -24.315 14.445 ;
        RECT -24.645 12.755 -24.315 13.085 ;
        RECT -24.645 11.395 -24.315 11.725 ;
        RECT -24.645 10.035 -24.315 10.365 ;
        RECT -24.645 8.675 -24.315 9.005 ;
        RECT -24.645 7.315 -24.315 7.645 ;
        RECT -24.645 5.955 -24.315 6.285 ;
        RECT -24.645 4.595 -24.315 4.925 ;
        RECT -24.645 3.235 -24.315 3.565 ;
        RECT -24.645 1.875 -24.315 2.205 ;
        RECT -24.645 0.515 -24.315 0.845 ;
        RECT -24.645 -0.845 -24.315 -0.515 ;
        RECT -24.645 -2.205 -24.315 -1.875 ;
        RECT -24.645 -7.645 -24.315 -7.315 ;
        RECT -24.645 -9.005 -24.315 -8.675 ;
        RECT -24.645 -10.73 -24.315 -10.4 ;
        RECT -24.645 -11.725 -24.315 -11.395 ;
        RECT -24.645 -16.77 -24.315 -16.44 ;
        RECT -24.645 -18.525 -24.315 -18.195 ;
        RECT -24.645 -21.245 -24.315 -20.915 ;
        RECT -24.645 -30.765 -24.315 -30.435 ;
        RECT -24.645 -32.125 -24.315 -31.795 ;
        RECT -24.645 -33.71 -24.315 -33.38 ;
        RECT -24.645 -34.845 -24.315 -34.515 ;
        RECT -24.645 -36.205 -24.315 -35.875 ;
        RECT -24.645 -38.925 -24.315 -38.595 ;
        RECT -24.645 -39.75 -24.315 -39.42 ;
        RECT -24.645 -41.645 -24.315 -41.315 ;
        RECT -24.645 -44.365 -24.315 -44.035 ;
        RECT -24.645 -49.805 -24.315 -49.475 ;
        RECT -24.645 -51.165 -24.315 -50.835 ;
        RECT -24.645 -53.885 -24.315 -53.555 ;
        RECT -24.645 -55.245 -24.315 -54.915 ;
        RECT -24.645 -59.325 -24.315 -58.995 ;
        RECT -24.645 -60.685 -24.315 -60.355 ;
        RECT -24.645 -63.405 -24.315 -63.075 ;
        RECT -24.645 -68.845 -24.315 -68.515 ;
        RECT -24.645 -70.205 -24.315 -69.875 ;
        RECT -24.645 -71.565 -24.315 -71.235 ;
        RECT -24.645 -73.19 -24.315 -72.86 ;
        RECT -24.645 -74.285 -24.315 -73.955 ;
        RECT -24.645 -75.645 -24.315 -75.315 ;
        RECT -24.645 -78.365 -24.315 -78.035 ;
        RECT -24.645 -79.725 -24.315 -79.395 ;
        RECT -24.645 -80.73 -24.315 -80.4 ;
        RECT -24.645 -82.445 -24.315 -82.115 ;
        RECT -24.645 -83.805 -24.315 -83.475 ;
        RECT -24.645 -86.525 -24.315 -86.195 ;
        RECT -24.645 -89.245 -24.315 -88.915 ;
        RECT -24.645 -90.605 -24.315 -90.275 ;
        RECT -24.645 -91.965 -24.315 -91.635 ;
        RECT -24.645 -93.325 -24.315 -92.995 ;
        RECT -24.645 -94.685 -24.315 -94.355 ;
        RECT -24.645 -95.37 -24.315 -95.04 ;
        RECT -24.645 -97.405 -24.315 -97.075 ;
        RECT -24.645 -100.125 -24.315 -99.795 ;
        RECT -24.645 -101.485 -24.315 -101.155 ;
        RECT -24.645 -102.91 -24.315 -102.58 ;
        RECT -24.645 -104.205 -24.315 -103.875 ;
        RECT -24.645 -105.565 -24.315 -105.235 ;
        RECT -24.64 -113.72 -24.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -24.645 -177.645 -24.315 -177.315 ;
        RECT -24.645 -179.005 -24.315 -178.675 ;
        RECT -24.645 -184.65 -24.315 -183.52 ;
        RECT -24.64 -184.765 -24.32 -175.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.285 244.04 -22.955 245.17 ;
        RECT -23.285 239.875 -22.955 240.205 ;
        RECT -23.285 238.515 -22.955 238.845 ;
        RECT -23.285 237.155 -22.955 237.485 ;
        RECT -23.285 235.795 -22.955 236.125 ;
        RECT -23.285 234.435 -22.955 234.765 ;
        RECT -23.285 233.075 -22.955 233.405 ;
        RECT -23.285 231.715 -22.955 232.045 ;
        RECT -23.285 230.355 -22.955 230.685 ;
        RECT -23.285 228.995 -22.955 229.325 ;
        RECT -23.285 227.635 -22.955 227.965 ;
        RECT -23.285 226.275 -22.955 226.605 ;
        RECT -23.285 224.915 -22.955 225.245 ;
        RECT -23.285 223.555 -22.955 223.885 ;
        RECT -23.285 222.195 -22.955 222.525 ;
        RECT -23.285 220.835 -22.955 221.165 ;
        RECT -23.285 219.475 -22.955 219.805 ;
        RECT -23.285 218.115 -22.955 218.445 ;
        RECT -23.285 216.755 -22.955 217.085 ;
        RECT -23.285 215.395 -22.955 215.725 ;
        RECT -23.285 214.035 -22.955 214.365 ;
        RECT -23.285 212.675 -22.955 213.005 ;
        RECT -23.285 211.315 -22.955 211.645 ;
        RECT -23.285 209.955 -22.955 210.285 ;
        RECT -23.285 208.595 -22.955 208.925 ;
        RECT -23.285 207.235 -22.955 207.565 ;
        RECT -23.285 205.875 -22.955 206.205 ;
        RECT -23.285 204.515 -22.955 204.845 ;
        RECT -23.285 203.155 -22.955 203.485 ;
        RECT -23.285 201.795 -22.955 202.125 ;
        RECT -23.285 200.435 -22.955 200.765 ;
        RECT -23.285 199.075 -22.955 199.405 ;
        RECT -23.285 197.715 -22.955 198.045 ;
        RECT -23.285 196.355 -22.955 196.685 ;
        RECT -23.285 194.995 -22.955 195.325 ;
        RECT -23.285 193.635 -22.955 193.965 ;
        RECT -23.285 192.275 -22.955 192.605 ;
        RECT -23.285 190.915 -22.955 191.245 ;
        RECT -23.285 189.555 -22.955 189.885 ;
        RECT -23.285 188.195 -22.955 188.525 ;
        RECT -23.285 186.835 -22.955 187.165 ;
        RECT -23.285 185.475 -22.955 185.805 ;
        RECT -23.285 184.115 -22.955 184.445 ;
        RECT -23.285 182.755 -22.955 183.085 ;
        RECT -23.285 181.395 -22.955 181.725 ;
        RECT -23.285 180.035 -22.955 180.365 ;
        RECT -23.285 178.675 -22.955 179.005 ;
        RECT -23.285 177.315 -22.955 177.645 ;
        RECT -23.285 175.955 -22.955 176.285 ;
        RECT -23.285 174.595 -22.955 174.925 ;
        RECT -23.285 173.235 -22.955 173.565 ;
        RECT -23.285 171.875 -22.955 172.205 ;
        RECT -23.285 170.515 -22.955 170.845 ;
        RECT -23.285 169.155 -22.955 169.485 ;
        RECT -23.285 167.795 -22.955 168.125 ;
        RECT -23.285 166.435 -22.955 166.765 ;
        RECT -23.285 165.075 -22.955 165.405 ;
        RECT -23.285 163.715 -22.955 164.045 ;
        RECT -23.285 162.355 -22.955 162.685 ;
        RECT -23.285 160.995 -22.955 161.325 ;
        RECT -23.285 159.635 -22.955 159.965 ;
        RECT -23.285 158.275 -22.955 158.605 ;
        RECT -23.285 156.915 -22.955 157.245 ;
        RECT -23.285 155.555 -22.955 155.885 ;
        RECT -23.285 154.195 -22.955 154.525 ;
        RECT -23.285 152.835 -22.955 153.165 ;
        RECT -23.285 151.475 -22.955 151.805 ;
        RECT -23.285 150.115 -22.955 150.445 ;
        RECT -23.285 148.755 -22.955 149.085 ;
        RECT -23.285 147.395 -22.955 147.725 ;
        RECT -23.285 146.035 -22.955 146.365 ;
        RECT -23.285 144.675 -22.955 145.005 ;
        RECT -23.285 143.315 -22.955 143.645 ;
        RECT -23.285 141.955 -22.955 142.285 ;
        RECT -23.285 140.595 -22.955 140.925 ;
        RECT -23.285 139.235 -22.955 139.565 ;
        RECT -23.285 137.875 -22.955 138.205 ;
        RECT -23.285 136.515 -22.955 136.845 ;
        RECT -23.285 135.155 -22.955 135.485 ;
        RECT -23.285 133.795 -22.955 134.125 ;
        RECT -23.285 132.435 -22.955 132.765 ;
        RECT -23.285 131.075 -22.955 131.405 ;
        RECT -23.285 129.715 -22.955 130.045 ;
        RECT -23.285 128.355 -22.955 128.685 ;
        RECT -23.285 126.995 -22.955 127.325 ;
        RECT -23.285 125.635 -22.955 125.965 ;
        RECT -23.285 124.275 -22.955 124.605 ;
        RECT -23.285 122.915 -22.955 123.245 ;
        RECT -23.285 121.555 -22.955 121.885 ;
        RECT -23.285 120.195 -22.955 120.525 ;
        RECT -23.285 118.835 -22.955 119.165 ;
        RECT -23.285 117.475 -22.955 117.805 ;
        RECT -23.285 116.115 -22.955 116.445 ;
        RECT -23.285 114.755 -22.955 115.085 ;
        RECT -23.285 113.395 -22.955 113.725 ;
        RECT -23.285 112.035 -22.955 112.365 ;
        RECT -23.285 110.675 -22.955 111.005 ;
        RECT -23.285 109.315 -22.955 109.645 ;
        RECT -23.285 107.955 -22.955 108.285 ;
        RECT -23.285 106.595 -22.955 106.925 ;
        RECT -23.285 105.235 -22.955 105.565 ;
        RECT -23.285 103.875 -22.955 104.205 ;
        RECT -23.285 102.515 -22.955 102.845 ;
        RECT -23.285 101.155 -22.955 101.485 ;
        RECT -23.285 99.795 -22.955 100.125 ;
        RECT -23.285 98.435 -22.955 98.765 ;
        RECT -23.285 97.075 -22.955 97.405 ;
        RECT -23.285 95.715 -22.955 96.045 ;
        RECT -23.285 94.355 -22.955 94.685 ;
        RECT -23.285 92.995 -22.955 93.325 ;
        RECT -23.285 91.635 -22.955 91.965 ;
        RECT -23.285 90.275 -22.955 90.605 ;
        RECT -23.285 88.915 -22.955 89.245 ;
        RECT -23.285 87.555 -22.955 87.885 ;
        RECT -23.285 86.195 -22.955 86.525 ;
        RECT -23.285 84.835 -22.955 85.165 ;
        RECT -23.285 83.475 -22.955 83.805 ;
        RECT -23.285 82.115 -22.955 82.445 ;
        RECT -23.285 80.755 -22.955 81.085 ;
        RECT -23.285 79.395 -22.955 79.725 ;
        RECT -23.285 78.035 -22.955 78.365 ;
        RECT -23.285 76.675 -22.955 77.005 ;
        RECT -23.285 75.315 -22.955 75.645 ;
        RECT -23.285 73.955 -22.955 74.285 ;
        RECT -23.285 72.595 -22.955 72.925 ;
        RECT -23.285 71.235 -22.955 71.565 ;
        RECT -23.285 69.875 -22.955 70.205 ;
        RECT -23.285 68.515 -22.955 68.845 ;
        RECT -23.285 67.155 -22.955 67.485 ;
        RECT -23.285 65.795 -22.955 66.125 ;
        RECT -23.285 64.435 -22.955 64.765 ;
        RECT -23.285 63.075 -22.955 63.405 ;
        RECT -23.285 61.715 -22.955 62.045 ;
        RECT -23.285 60.355 -22.955 60.685 ;
        RECT -23.285 58.995 -22.955 59.325 ;
        RECT -23.285 57.635 -22.955 57.965 ;
        RECT -23.285 56.275 -22.955 56.605 ;
        RECT -23.285 54.915 -22.955 55.245 ;
        RECT -23.285 53.555 -22.955 53.885 ;
        RECT -23.285 52.195 -22.955 52.525 ;
        RECT -23.285 50.835 -22.955 51.165 ;
        RECT -23.285 49.475 -22.955 49.805 ;
        RECT -23.285 48.115 -22.955 48.445 ;
        RECT -23.285 46.755 -22.955 47.085 ;
        RECT -23.285 45.395 -22.955 45.725 ;
        RECT -23.285 44.035 -22.955 44.365 ;
        RECT -23.285 42.675 -22.955 43.005 ;
        RECT -23.285 41.315 -22.955 41.645 ;
        RECT -23.285 39.955 -22.955 40.285 ;
        RECT -23.285 38.595 -22.955 38.925 ;
        RECT -23.285 37.235 -22.955 37.565 ;
        RECT -23.285 35.875 -22.955 36.205 ;
        RECT -23.285 34.515 -22.955 34.845 ;
        RECT -23.285 33.155 -22.955 33.485 ;
        RECT -23.285 31.795 -22.955 32.125 ;
        RECT -23.285 30.435 -22.955 30.765 ;
        RECT -23.285 29.075 -22.955 29.405 ;
        RECT -23.285 27.715 -22.955 28.045 ;
        RECT -23.285 26.355 -22.955 26.685 ;
        RECT -23.285 24.995 -22.955 25.325 ;
        RECT -23.285 23.635 -22.955 23.965 ;
        RECT -23.285 22.275 -22.955 22.605 ;
        RECT -23.285 20.915 -22.955 21.245 ;
        RECT -23.285 19.555 -22.955 19.885 ;
        RECT -23.285 18.195 -22.955 18.525 ;
        RECT -23.285 16.835 -22.955 17.165 ;
        RECT -23.285 15.475 -22.955 15.805 ;
        RECT -23.285 14.115 -22.955 14.445 ;
        RECT -23.285 12.755 -22.955 13.085 ;
        RECT -23.285 11.395 -22.955 11.725 ;
        RECT -23.285 10.035 -22.955 10.365 ;
        RECT -23.285 8.675 -22.955 9.005 ;
        RECT -23.285 7.315 -22.955 7.645 ;
        RECT -23.285 5.955 -22.955 6.285 ;
        RECT -23.285 4.595 -22.955 4.925 ;
        RECT -23.285 3.235 -22.955 3.565 ;
        RECT -23.285 1.875 -22.955 2.205 ;
        RECT -23.285 0.515 -22.955 0.845 ;
        RECT -23.285 -0.845 -22.955 -0.515 ;
        RECT -23.285 -2.205 -22.955 -1.875 ;
        RECT -23.285 -7.645 -22.955 -7.315 ;
        RECT -23.285 -9.005 -22.955 -8.675 ;
        RECT -23.285 -10.73 -22.955 -10.4 ;
        RECT -23.285 -11.725 -22.955 -11.395 ;
        RECT -23.285 -16.77 -22.955 -16.44 ;
        RECT -23.285 -18.525 -22.955 -18.195 ;
        RECT -23.285 -21.245 -22.955 -20.915 ;
        RECT -23.285 -30.765 -22.955 -30.435 ;
        RECT -23.285 -32.125 -22.955 -31.795 ;
        RECT -23.285 -33.71 -22.955 -33.38 ;
        RECT -23.285 -34.845 -22.955 -34.515 ;
        RECT -23.285 -36.205 -22.955 -35.875 ;
        RECT -23.285 -38.925 -22.955 -38.595 ;
        RECT -23.285 -39.75 -22.955 -39.42 ;
        RECT -23.285 -41.645 -22.955 -41.315 ;
        RECT -23.285 -44.365 -22.955 -44.035 ;
        RECT -23.285 -49.805 -22.955 -49.475 ;
        RECT -23.285 -51.165 -22.955 -50.835 ;
        RECT -23.285 -52.525 -22.955 -52.195 ;
        RECT -23.285 -53.885 -22.955 -53.555 ;
        RECT -23.285 -55.245 -22.955 -54.915 ;
        RECT -23.285 -56.605 -22.955 -56.275 ;
        RECT -23.285 -57.965 -22.955 -57.635 ;
        RECT -23.285 -59.325 -22.955 -58.995 ;
        RECT -23.285 -60.685 -22.955 -60.355 ;
        RECT -23.285 -62.045 -22.955 -61.715 ;
        RECT -23.285 -63.405 -22.955 -63.075 ;
        RECT -23.285 -64.765 -22.955 -64.435 ;
        RECT -23.285 -66.125 -22.955 -65.795 ;
        RECT -23.285 -68.845 -22.955 -68.515 ;
        RECT -23.285 -70.205 -22.955 -69.875 ;
        RECT -23.285 -71.565 -22.955 -71.235 ;
        RECT -23.285 -73.19 -22.955 -72.86 ;
        RECT -23.285 -74.285 -22.955 -73.955 ;
        RECT -23.285 -75.645 -22.955 -75.315 ;
        RECT -23.285 -78.365 -22.955 -78.035 ;
        RECT -23.285 -79.725 -22.955 -79.395 ;
        RECT -23.285 -80.73 -22.955 -80.4 ;
        RECT -23.285 -82.445 -22.955 -82.115 ;
        RECT -23.285 -83.805 -22.955 -83.475 ;
        RECT -23.285 -86.525 -22.955 -86.195 ;
        RECT -23.285 -89.245 -22.955 -88.915 ;
        RECT -23.285 -90.605 -22.955 -90.275 ;
        RECT -23.285 -91.965 -22.955 -91.635 ;
        RECT -23.285 -93.325 -22.955 -92.995 ;
        RECT -23.285 -94.685 -22.955 -94.355 ;
        RECT -23.285 -95.37 -22.955 -95.04 ;
        RECT -23.285 -97.405 -22.955 -97.075 ;
        RECT -23.285 -100.125 -22.955 -99.795 ;
        RECT -23.285 -101.485 -22.955 -101.155 ;
        RECT -23.285 -102.91 -22.955 -102.58 ;
        RECT -23.285 -104.205 -22.955 -103.875 ;
        RECT -23.285 -105.565 -22.955 -105.235 ;
        RECT -23.28 -114.4 -22.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.285 -177.645 -22.955 -177.315 ;
        RECT -23.285 -179.005 -22.955 -178.675 ;
        RECT -23.285 -184.65 -22.955 -183.52 ;
        RECT -23.28 -184.765 -22.96 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.925 125.635 -21.595 125.965 ;
        RECT -21.925 124.275 -21.595 124.605 ;
        RECT -21.925 122.915 -21.595 123.245 ;
        RECT -21.925 121.555 -21.595 121.885 ;
        RECT -21.925 120.195 -21.595 120.525 ;
        RECT -21.925 118.835 -21.595 119.165 ;
        RECT -21.925 117.475 -21.595 117.805 ;
        RECT -21.925 116.115 -21.595 116.445 ;
        RECT -21.925 114.755 -21.595 115.085 ;
        RECT -21.925 113.395 -21.595 113.725 ;
        RECT -21.925 112.035 -21.595 112.365 ;
        RECT -21.925 110.675 -21.595 111.005 ;
        RECT -21.925 109.315 -21.595 109.645 ;
        RECT -21.925 107.955 -21.595 108.285 ;
        RECT -21.925 106.595 -21.595 106.925 ;
        RECT -21.925 105.235 -21.595 105.565 ;
        RECT -21.925 103.875 -21.595 104.205 ;
        RECT -21.925 102.515 -21.595 102.845 ;
        RECT -21.925 101.155 -21.595 101.485 ;
        RECT -21.925 99.795 -21.595 100.125 ;
        RECT -21.925 98.435 -21.595 98.765 ;
        RECT -21.925 97.075 -21.595 97.405 ;
        RECT -21.925 95.715 -21.595 96.045 ;
        RECT -21.925 94.355 -21.595 94.685 ;
        RECT -21.925 92.995 -21.595 93.325 ;
        RECT -21.925 91.635 -21.595 91.965 ;
        RECT -21.925 90.275 -21.595 90.605 ;
        RECT -21.925 88.915 -21.595 89.245 ;
        RECT -21.925 87.555 -21.595 87.885 ;
        RECT -21.925 86.195 -21.595 86.525 ;
        RECT -21.925 84.835 -21.595 85.165 ;
        RECT -21.925 83.475 -21.595 83.805 ;
        RECT -21.925 82.115 -21.595 82.445 ;
        RECT -21.925 80.755 -21.595 81.085 ;
        RECT -21.925 79.395 -21.595 79.725 ;
        RECT -21.925 78.035 -21.595 78.365 ;
        RECT -21.925 76.675 -21.595 77.005 ;
        RECT -21.925 75.315 -21.595 75.645 ;
        RECT -21.925 73.955 -21.595 74.285 ;
        RECT -21.925 72.595 -21.595 72.925 ;
        RECT -21.925 71.235 -21.595 71.565 ;
        RECT -21.925 69.875 -21.595 70.205 ;
        RECT -21.925 68.515 -21.595 68.845 ;
        RECT -21.925 67.155 -21.595 67.485 ;
        RECT -21.925 65.795 -21.595 66.125 ;
        RECT -21.925 64.435 -21.595 64.765 ;
        RECT -21.925 63.075 -21.595 63.405 ;
        RECT -21.925 61.715 -21.595 62.045 ;
        RECT -21.925 60.355 -21.595 60.685 ;
        RECT -21.925 58.995 -21.595 59.325 ;
        RECT -21.925 57.635 -21.595 57.965 ;
        RECT -21.925 56.275 -21.595 56.605 ;
        RECT -21.925 54.915 -21.595 55.245 ;
        RECT -21.925 53.555 -21.595 53.885 ;
        RECT -21.925 52.195 -21.595 52.525 ;
        RECT -21.925 50.835 -21.595 51.165 ;
        RECT -21.925 49.475 -21.595 49.805 ;
        RECT -21.925 48.115 -21.595 48.445 ;
        RECT -21.925 46.755 -21.595 47.085 ;
        RECT -21.925 45.395 -21.595 45.725 ;
        RECT -21.925 44.035 -21.595 44.365 ;
        RECT -21.925 42.675 -21.595 43.005 ;
        RECT -21.925 41.315 -21.595 41.645 ;
        RECT -21.925 39.955 -21.595 40.285 ;
        RECT -21.925 38.595 -21.595 38.925 ;
        RECT -21.925 37.235 -21.595 37.565 ;
        RECT -21.925 35.875 -21.595 36.205 ;
        RECT -21.925 34.515 -21.595 34.845 ;
        RECT -21.925 33.155 -21.595 33.485 ;
        RECT -21.925 31.795 -21.595 32.125 ;
        RECT -21.925 30.435 -21.595 30.765 ;
        RECT -21.925 29.075 -21.595 29.405 ;
        RECT -21.925 27.715 -21.595 28.045 ;
        RECT -21.925 26.355 -21.595 26.685 ;
        RECT -21.925 24.995 -21.595 25.325 ;
        RECT -21.925 23.635 -21.595 23.965 ;
        RECT -21.925 22.275 -21.595 22.605 ;
        RECT -21.925 20.915 -21.595 21.245 ;
        RECT -21.925 19.555 -21.595 19.885 ;
        RECT -21.925 18.195 -21.595 18.525 ;
        RECT -21.925 16.835 -21.595 17.165 ;
        RECT -21.925 15.475 -21.595 15.805 ;
        RECT -21.925 14.115 -21.595 14.445 ;
        RECT -21.925 12.755 -21.595 13.085 ;
        RECT -21.925 11.395 -21.595 11.725 ;
        RECT -21.925 10.035 -21.595 10.365 ;
        RECT -21.925 8.675 -21.595 9.005 ;
        RECT -21.925 7.315 -21.595 7.645 ;
        RECT -21.925 5.955 -21.595 6.285 ;
        RECT -21.925 4.595 -21.595 4.925 ;
        RECT -21.925 3.235 -21.595 3.565 ;
        RECT -21.925 1.875 -21.595 2.205 ;
        RECT -21.925 0.515 -21.595 0.845 ;
        RECT -21.925 -0.845 -21.595 -0.515 ;
        RECT -21.925 -2.205 -21.595 -1.875 ;
        RECT -21.925 -3.565 -21.595 -3.235 ;
        RECT -21.925 -7.645 -21.595 -7.315 ;
        RECT -21.925 -9.005 -21.595 -8.675 ;
        RECT -21.925 -10.73 -21.595 -10.4 ;
        RECT -21.925 -11.725 -21.595 -11.395 ;
        RECT -21.925 -16.77 -21.595 -16.44 ;
        RECT -21.925 -18.525 -21.595 -18.195 ;
        RECT -21.925 -21.245 -21.595 -20.915 ;
        RECT -21.92 -23.96 -21.6 245.285 ;
        RECT -21.925 244.04 -21.595 245.17 ;
        RECT -21.925 239.875 -21.595 240.205 ;
        RECT -21.925 238.515 -21.595 238.845 ;
        RECT -21.925 237.155 -21.595 237.485 ;
        RECT -21.925 235.795 -21.595 236.125 ;
        RECT -21.925 234.435 -21.595 234.765 ;
        RECT -21.925 233.075 -21.595 233.405 ;
        RECT -21.925 231.715 -21.595 232.045 ;
        RECT -21.925 230.355 -21.595 230.685 ;
        RECT -21.925 228.995 -21.595 229.325 ;
        RECT -21.925 227.635 -21.595 227.965 ;
        RECT -21.925 226.275 -21.595 226.605 ;
        RECT -21.925 224.915 -21.595 225.245 ;
        RECT -21.925 223.555 -21.595 223.885 ;
        RECT -21.925 222.195 -21.595 222.525 ;
        RECT -21.925 220.835 -21.595 221.165 ;
        RECT -21.925 219.475 -21.595 219.805 ;
        RECT -21.925 218.115 -21.595 218.445 ;
        RECT -21.925 216.755 -21.595 217.085 ;
        RECT -21.925 215.395 -21.595 215.725 ;
        RECT -21.925 214.035 -21.595 214.365 ;
        RECT -21.925 212.675 -21.595 213.005 ;
        RECT -21.925 211.315 -21.595 211.645 ;
        RECT -21.925 209.955 -21.595 210.285 ;
        RECT -21.925 208.595 -21.595 208.925 ;
        RECT -21.925 207.235 -21.595 207.565 ;
        RECT -21.925 205.875 -21.595 206.205 ;
        RECT -21.925 204.515 -21.595 204.845 ;
        RECT -21.925 203.155 -21.595 203.485 ;
        RECT -21.925 201.795 -21.595 202.125 ;
        RECT -21.925 200.435 -21.595 200.765 ;
        RECT -21.925 199.075 -21.595 199.405 ;
        RECT -21.925 197.715 -21.595 198.045 ;
        RECT -21.925 196.355 -21.595 196.685 ;
        RECT -21.925 194.995 -21.595 195.325 ;
        RECT -21.925 193.635 -21.595 193.965 ;
        RECT -21.925 192.275 -21.595 192.605 ;
        RECT -21.925 190.915 -21.595 191.245 ;
        RECT -21.925 189.555 -21.595 189.885 ;
        RECT -21.925 188.195 -21.595 188.525 ;
        RECT -21.925 186.835 -21.595 187.165 ;
        RECT -21.925 185.475 -21.595 185.805 ;
        RECT -21.925 184.115 -21.595 184.445 ;
        RECT -21.925 182.755 -21.595 183.085 ;
        RECT -21.925 181.395 -21.595 181.725 ;
        RECT -21.925 180.035 -21.595 180.365 ;
        RECT -21.925 178.675 -21.595 179.005 ;
        RECT -21.925 177.315 -21.595 177.645 ;
        RECT -21.925 175.955 -21.595 176.285 ;
        RECT -21.925 174.595 -21.595 174.925 ;
        RECT -21.925 173.235 -21.595 173.565 ;
        RECT -21.925 171.875 -21.595 172.205 ;
        RECT -21.925 170.515 -21.595 170.845 ;
        RECT -21.925 169.155 -21.595 169.485 ;
        RECT -21.925 167.795 -21.595 168.125 ;
        RECT -21.925 166.435 -21.595 166.765 ;
        RECT -21.925 165.075 -21.595 165.405 ;
        RECT -21.925 163.715 -21.595 164.045 ;
        RECT -21.925 162.355 -21.595 162.685 ;
        RECT -21.925 160.995 -21.595 161.325 ;
        RECT -21.925 159.635 -21.595 159.965 ;
        RECT -21.925 158.275 -21.595 158.605 ;
        RECT -21.925 156.915 -21.595 157.245 ;
        RECT -21.925 155.555 -21.595 155.885 ;
        RECT -21.925 154.195 -21.595 154.525 ;
        RECT -21.925 152.835 -21.595 153.165 ;
        RECT -21.925 151.475 -21.595 151.805 ;
        RECT -21.925 150.115 -21.595 150.445 ;
        RECT -21.925 148.755 -21.595 149.085 ;
        RECT -21.925 147.395 -21.595 147.725 ;
        RECT -21.925 146.035 -21.595 146.365 ;
        RECT -21.925 144.675 -21.595 145.005 ;
        RECT -21.925 143.315 -21.595 143.645 ;
        RECT -21.925 141.955 -21.595 142.285 ;
        RECT -21.925 140.595 -21.595 140.925 ;
        RECT -21.925 139.235 -21.595 139.565 ;
        RECT -21.925 137.875 -21.595 138.205 ;
        RECT -21.925 136.515 -21.595 136.845 ;
        RECT -21.925 135.155 -21.595 135.485 ;
        RECT -21.925 133.795 -21.595 134.125 ;
        RECT -21.925 132.435 -21.595 132.765 ;
        RECT -21.925 131.075 -21.595 131.405 ;
        RECT -21.925 129.715 -21.595 130.045 ;
        RECT -21.925 128.355 -21.595 128.685 ;
        RECT -21.925 126.995 -21.595 127.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.805 -174.925 -32.475 -174.595 ;
        RECT -32.805 -177.645 -32.475 -177.315 ;
        RECT -32.805 -179.005 -32.475 -178.675 ;
        RECT -32.805 -184.65 -32.475 -183.52 ;
        RECT -32.8 -184.765 -32.48 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -31.445 244.04 -31.115 245.17 ;
        RECT -31.445 239.875 -31.115 240.205 ;
        RECT -31.445 238.515 -31.115 238.845 ;
        RECT -31.445 237.155 -31.115 237.485 ;
        RECT -31.445 235.795 -31.115 236.125 ;
        RECT -31.445 234.435 -31.115 234.765 ;
        RECT -31.445 233.075 -31.115 233.405 ;
        RECT -31.445 231.715 -31.115 232.045 ;
        RECT -31.445 230.355 -31.115 230.685 ;
        RECT -31.445 228.995 -31.115 229.325 ;
        RECT -31.445 227.635 -31.115 227.965 ;
        RECT -31.445 226.275 -31.115 226.605 ;
        RECT -31.445 224.915 -31.115 225.245 ;
        RECT -31.445 223.555 -31.115 223.885 ;
        RECT -31.445 222.195 -31.115 222.525 ;
        RECT -31.445 220.835 -31.115 221.165 ;
        RECT -31.445 219.475 -31.115 219.805 ;
        RECT -31.445 218.115 -31.115 218.445 ;
        RECT -31.445 216.755 -31.115 217.085 ;
        RECT -31.445 215.395 -31.115 215.725 ;
        RECT -31.445 214.035 -31.115 214.365 ;
        RECT -31.445 212.675 -31.115 213.005 ;
        RECT -31.445 211.315 -31.115 211.645 ;
        RECT -31.445 209.955 -31.115 210.285 ;
        RECT -31.445 208.595 -31.115 208.925 ;
        RECT -31.445 207.235 -31.115 207.565 ;
        RECT -31.445 205.875 -31.115 206.205 ;
        RECT -31.445 204.515 -31.115 204.845 ;
        RECT -31.445 203.155 -31.115 203.485 ;
        RECT -31.445 201.795 -31.115 202.125 ;
        RECT -31.445 200.435 -31.115 200.765 ;
        RECT -31.445 199.075 -31.115 199.405 ;
        RECT -31.445 197.715 -31.115 198.045 ;
        RECT -31.445 196.355 -31.115 196.685 ;
        RECT -31.445 194.995 -31.115 195.325 ;
        RECT -31.445 193.635 -31.115 193.965 ;
        RECT -31.445 192.275 -31.115 192.605 ;
        RECT -31.445 190.915 -31.115 191.245 ;
        RECT -31.445 189.555 -31.115 189.885 ;
        RECT -31.445 188.195 -31.115 188.525 ;
        RECT -31.445 186.835 -31.115 187.165 ;
        RECT -31.445 185.475 -31.115 185.805 ;
        RECT -31.445 184.115 -31.115 184.445 ;
        RECT -31.445 182.755 -31.115 183.085 ;
        RECT -31.445 181.395 -31.115 181.725 ;
        RECT -31.445 180.035 -31.115 180.365 ;
        RECT -31.445 178.675 -31.115 179.005 ;
        RECT -31.445 177.315 -31.115 177.645 ;
        RECT -31.445 175.955 -31.115 176.285 ;
        RECT -31.445 174.595 -31.115 174.925 ;
        RECT -31.445 173.235 -31.115 173.565 ;
        RECT -31.445 171.875 -31.115 172.205 ;
        RECT -31.445 170.515 -31.115 170.845 ;
        RECT -31.445 169.155 -31.115 169.485 ;
        RECT -31.445 167.795 -31.115 168.125 ;
        RECT -31.445 166.435 -31.115 166.765 ;
        RECT -31.445 165.075 -31.115 165.405 ;
        RECT -31.445 163.715 -31.115 164.045 ;
        RECT -31.445 162.355 -31.115 162.685 ;
        RECT -31.445 160.995 -31.115 161.325 ;
        RECT -31.445 159.635 -31.115 159.965 ;
        RECT -31.445 158.275 -31.115 158.605 ;
        RECT -31.445 156.915 -31.115 157.245 ;
        RECT -31.445 155.555 -31.115 155.885 ;
        RECT -31.445 154.195 -31.115 154.525 ;
        RECT -31.445 152.835 -31.115 153.165 ;
        RECT -31.445 151.475 -31.115 151.805 ;
        RECT -31.445 150.115 -31.115 150.445 ;
        RECT -31.445 148.755 -31.115 149.085 ;
        RECT -31.445 147.395 -31.115 147.725 ;
        RECT -31.445 146.035 -31.115 146.365 ;
        RECT -31.445 144.675 -31.115 145.005 ;
        RECT -31.445 143.315 -31.115 143.645 ;
        RECT -31.445 141.955 -31.115 142.285 ;
        RECT -31.445 140.595 -31.115 140.925 ;
        RECT -31.445 139.235 -31.115 139.565 ;
        RECT -31.445 137.875 -31.115 138.205 ;
        RECT -31.445 136.515 -31.115 136.845 ;
        RECT -31.445 135.155 -31.115 135.485 ;
        RECT -31.445 133.795 -31.115 134.125 ;
        RECT -31.445 132.435 -31.115 132.765 ;
        RECT -31.445 131.075 -31.115 131.405 ;
        RECT -31.445 129.715 -31.115 130.045 ;
        RECT -31.445 128.355 -31.115 128.685 ;
        RECT -31.445 126.995 -31.115 127.325 ;
        RECT -31.445 125.635 -31.115 125.965 ;
        RECT -31.445 124.275 -31.115 124.605 ;
        RECT -31.445 122.915 -31.115 123.245 ;
        RECT -31.445 121.555 -31.115 121.885 ;
        RECT -31.445 120.195 -31.115 120.525 ;
        RECT -31.445 118.835 -31.115 119.165 ;
        RECT -31.445 117.475 -31.115 117.805 ;
        RECT -31.445 116.115 -31.115 116.445 ;
        RECT -31.445 114.755 -31.115 115.085 ;
        RECT -31.445 113.395 -31.115 113.725 ;
        RECT -31.445 112.035 -31.115 112.365 ;
        RECT -31.445 110.675 -31.115 111.005 ;
        RECT -31.445 109.315 -31.115 109.645 ;
        RECT -31.445 107.955 -31.115 108.285 ;
        RECT -31.445 106.595 -31.115 106.925 ;
        RECT -31.445 105.235 -31.115 105.565 ;
        RECT -31.445 103.875 -31.115 104.205 ;
        RECT -31.445 102.515 -31.115 102.845 ;
        RECT -31.445 101.155 -31.115 101.485 ;
        RECT -31.445 99.795 -31.115 100.125 ;
        RECT -31.445 98.435 -31.115 98.765 ;
        RECT -31.445 97.075 -31.115 97.405 ;
        RECT -31.445 95.715 -31.115 96.045 ;
        RECT -31.445 94.355 -31.115 94.685 ;
        RECT -31.445 92.995 -31.115 93.325 ;
        RECT -31.445 91.635 -31.115 91.965 ;
        RECT -31.445 90.275 -31.115 90.605 ;
        RECT -31.445 88.915 -31.115 89.245 ;
        RECT -31.445 87.555 -31.115 87.885 ;
        RECT -31.445 86.195 -31.115 86.525 ;
        RECT -31.445 84.835 -31.115 85.165 ;
        RECT -31.445 83.475 -31.115 83.805 ;
        RECT -31.445 82.115 -31.115 82.445 ;
        RECT -31.445 80.755 -31.115 81.085 ;
        RECT -31.445 79.395 -31.115 79.725 ;
        RECT -31.445 78.035 -31.115 78.365 ;
        RECT -31.445 76.675 -31.115 77.005 ;
        RECT -31.445 75.315 -31.115 75.645 ;
        RECT -31.445 73.955 -31.115 74.285 ;
        RECT -31.445 72.595 -31.115 72.925 ;
        RECT -31.445 71.235 -31.115 71.565 ;
        RECT -31.445 69.875 -31.115 70.205 ;
        RECT -31.445 68.515 -31.115 68.845 ;
        RECT -31.445 67.155 -31.115 67.485 ;
        RECT -31.445 65.795 -31.115 66.125 ;
        RECT -31.445 64.435 -31.115 64.765 ;
        RECT -31.445 63.075 -31.115 63.405 ;
        RECT -31.445 61.715 -31.115 62.045 ;
        RECT -31.445 60.355 -31.115 60.685 ;
        RECT -31.445 58.995 -31.115 59.325 ;
        RECT -31.445 57.635 -31.115 57.965 ;
        RECT -31.445 56.275 -31.115 56.605 ;
        RECT -31.445 54.915 -31.115 55.245 ;
        RECT -31.445 53.555 -31.115 53.885 ;
        RECT -31.445 52.195 -31.115 52.525 ;
        RECT -31.445 50.835 -31.115 51.165 ;
        RECT -31.445 49.475 -31.115 49.805 ;
        RECT -31.445 48.115 -31.115 48.445 ;
        RECT -31.445 46.755 -31.115 47.085 ;
        RECT -31.445 45.395 -31.115 45.725 ;
        RECT -31.445 44.035 -31.115 44.365 ;
        RECT -31.445 42.675 -31.115 43.005 ;
        RECT -31.445 41.315 -31.115 41.645 ;
        RECT -31.445 39.955 -31.115 40.285 ;
        RECT -31.445 38.595 -31.115 38.925 ;
        RECT -31.445 37.235 -31.115 37.565 ;
        RECT -31.445 35.875 -31.115 36.205 ;
        RECT -31.445 34.515 -31.115 34.845 ;
        RECT -31.445 33.155 -31.115 33.485 ;
        RECT -31.445 31.795 -31.115 32.125 ;
        RECT -31.445 30.435 -31.115 30.765 ;
        RECT -31.445 29.075 -31.115 29.405 ;
        RECT -31.445 27.715 -31.115 28.045 ;
        RECT -31.445 26.355 -31.115 26.685 ;
        RECT -31.445 24.995 -31.115 25.325 ;
        RECT -31.445 23.635 -31.115 23.965 ;
        RECT -31.445 22.275 -31.115 22.605 ;
        RECT -31.445 20.915 -31.115 21.245 ;
        RECT -31.445 19.555 -31.115 19.885 ;
        RECT -31.445 18.195 -31.115 18.525 ;
        RECT -31.445 16.835 -31.115 17.165 ;
        RECT -31.445 15.475 -31.115 15.805 ;
        RECT -31.445 14.115 -31.115 14.445 ;
        RECT -31.445 12.755 -31.115 13.085 ;
        RECT -31.445 11.395 -31.115 11.725 ;
        RECT -31.445 10.035 -31.115 10.365 ;
        RECT -31.445 8.675 -31.115 9.005 ;
        RECT -31.445 7.315 -31.115 7.645 ;
        RECT -31.445 5.955 -31.115 6.285 ;
        RECT -31.445 4.595 -31.115 4.925 ;
        RECT -31.445 3.235 -31.115 3.565 ;
        RECT -31.445 1.875 -31.115 2.205 ;
        RECT -31.445 0.515 -31.115 0.845 ;
        RECT -31.445 -0.845 -31.115 -0.515 ;
        RECT -31.445 -7.645 -31.115 -7.315 ;
        RECT -31.445 -9.005 -31.115 -8.675 ;
        RECT -31.445 -10.365 -31.115 -10.035 ;
        RECT -31.445 -14.445 -31.115 -14.115 ;
        RECT -31.445 -17.165 -31.115 -16.835 ;
        RECT -31.445 -18.525 -31.115 -18.195 ;
        RECT -31.445 -19.885 -31.115 -19.555 ;
        RECT -31.445 -21.245 -31.115 -20.915 ;
        RECT -31.445 -22.605 -31.115 -22.275 ;
        RECT -31.445 -23.965 -31.115 -23.635 ;
        RECT -31.445 -25.325 -31.115 -24.995 ;
        RECT -31.445 -32.125 -31.115 -31.795 ;
        RECT -31.445 -33.71 -31.115 -33.38 ;
        RECT -31.445 -34.845 -31.115 -34.515 ;
        RECT -31.445 -36.205 -31.115 -35.875 ;
        RECT -31.445 -38.925 -31.115 -38.595 ;
        RECT -31.445 -39.75 -31.115 -39.42 ;
        RECT -31.445 -41.645 -31.115 -41.315 ;
        RECT -31.445 -44.365 -31.115 -44.035 ;
        RECT -31.445 -49.805 -31.115 -49.475 ;
        RECT -31.445 -51.165 -31.115 -50.835 ;
        RECT -31.445 -53.885 -31.115 -53.555 ;
        RECT -31.445 -55.245 -31.115 -54.915 ;
        RECT -31.445 -59.325 -31.115 -58.995 ;
        RECT -31.445 -60.685 -31.115 -60.355 ;
        RECT -31.445 -63.405 -31.115 -63.075 ;
        RECT -31.445 -70.205 -31.115 -69.875 ;
        RECT -31.445 -71.565 -31.115 -71.235 ;
        RECT -31.445 -72.925 -31.115 -72.595 ;
        RECT -31.445 -74.285 -31.115 -73.955 ;
        RECT -31.445 -75.645 -31.115 -75.315 ;
        RECT -31.445 -77.005 -31.115 -76.675 ;
        RECT -31.445 -78.365 -31.115 -78.035 ;
        RECT -31.445 -79.725 -31.115 -79.395 ;
        RECT -31.445 -81.085 -31.115 -80.755 ;
        RECT -31.445 -82.445 -31.115 -82.115 ;
        RECT -31.445 -83.805 -31.115 -83.475 ;
        RECT -31.445 -85.165 -31.115 -84.835 ;
        RECT -31.445 -86.525 -31.115 -86.195 ;
        RECT -31.445 -87.885 -31.115 -87.555 ;
        RECT -31.445 -89.245 -31.115 -88.915 ;
        RECT -31.445 -90.605 -31.115 -90.275 ;
        RECT -31.445 -91.965 -31.115 -91.635 ;
        RECT -31.445 -93.325 -31.115 -92.995 ;
        RECT -31.445 -94.685 -31.115 -94.355 ;
        RECT -31.445 -96.045 -31.115 -95.715 ;
        RECT -31.445 -97.405 -31.115 -97.075 ;
        RECT -31.445 -98.765 -31.115 -98.435 ;
        RECT -31.445 -100.125 -31.115 -99.795 ;
        RECT -31.445 -101.485 -31.115 -101.155 ;
        RECT -31.445 -102.845 -31.115 -102.515 ;
        RECT -31.445 -104.205 -31.115 -103.875 ;
        RECT -31.445 -105.565 -31.115 -105.235 ;
        RECT -31.445 -106.925 -31.115 -106.595 ;
        RECT -31.445 -108.285 -31.115 -107.955 ;
        RECT -31.445 -109.645 -31.115 -109.315 ;
        RECT -31.445 -111.005 -31.115 -110.675 ;
        RECT -31.445 -112.365 -31.115 -112.035 ;
        RECT -31.445 -113.725 -31.115 -113.395 ;
        RECT -31.445 -115.085 -31.115 -114.755 ;
        RECT -31.445 -116.445 -31.115 -116.115 ;
        RECT -31.445 -117.805 -31.115 -117.475 ;
        RECT -31.445 -119.165 -31.115 -118.835 ;
        RECT -31.445 -120.525 -31.115 -120.195 ;
        RECT -31.445 -123.245 -31.115 -122.915 ;
        RECT -31.445 -124.605 -31.115 -124.275 ;
        RECT -31.445 -125.965 -31.115 -125.635 ;
        RECT -31.445 -127.325 -31.115 -126.995 ;
        RECT -31.445 -128.685 -31.115 -128.355 ;
        RECT -31.445 -130.045 -31.115 -129.715 ;
        RECT -31.445 -134.125 -31.115 -133.795 ;
        RECT -31.445 -135.485 -31.115 -135.155 ;
        RECT -31.445 -136.845 -31.115 -136.515 ;
        RECT -31.445 -139.565 -31.115 -139.235 ;
        RECT -31.445 -142.285 -31.115 -141.955 ;
        RECT -31.445 -143.645 -31.115 -143.315 ;
        RECT -31.445 -145.005 -31.115 -144.675 ;
        RECT -31.445 -146.365 -31.115 -146.035 ;
        RECT -31.445 -147.725 -31.115 -147.395 ;
        RECT -31.445 -149.085 -31.115 -148.755 ;
        RECT -31.445 -151.805 -31.115 -151.475 ;
        RECT -31.445 -153.165 -31.115 -152.835 ;
        RECT -31.445 -157.245 -31.115 -156.915 ;
        RECT -31.445 -158.605 -31.115 -158.275 ;
        RECT -31.445 -159.965 -31.115 -159.635 ;
        RECT -31.445 -161.325 -31.115 -160.995 ;
        RECT -31.445 -162.685 -31.115 -162.355 ;
        RECT -31.445 -164.045 -31.115 -163.715 ;
        RECT -31.445 -165.405 -31.115 -165.075 ;
        RECT -31.445 -166.765 -31.115 -166.435 ;
        RECT -31.445 -169.615 -31.115 -169.285 ;
        RECT -31.445 -170.845 -31.115 -170.515 ;
        RECT -31.445 -172.205 -31.115 -171.875 ;
        RECT -31.445 -173.565 -31.115 -173.235 ;
        RECT -31.445 -174.925 -31.115 -174.595 ;
        RECT -31.445 -177.645 -31.115 -177.315 ;
        RECT -31.445 -179.005 -31.115 -178.675 ;
        RECT -31.445 -184.65 -31.115 -183.52 ;
        RECT -31.44 -184.765 -31.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 244.04 -29.755 245.17 ;
        RECT -30.085 239.875 -29.755 240.205 ;
        RECT -30.085 238.515 -29.755 238.845 ;
        RECT -30.085 237.155 -29.755 237.485 ;
        RECT -30.085 235.795 -29.755 236.125 ;
        RECT -30.085 234.435 -29.755 234.765 ;
        RECT -30.085 233.075 -29.755 233.405 ;
        RECT -30.085 231.715 -29.755 232.045 ;
        RECT -30.085 230.355 -29.755 230.685 ;
        RECT -30.085 228.995 -29.755 229.325 ;
        RECT -30.085 227.635 -29.755 227.965 ;
        RECT -30.085 226.275 -29.755 226.605 ;
        RECT -30.085 224.915 -29.755 225.245 ;
        RECT -30.085 223.555 -29.755 223.885 ;
        RECT -30.085 222.195 -29.755 222.525 ;
        RECT -30.085 220.835 -29.755 221.165 ;
        RECT -30.085 219.475 -29.755 219.805 ;
        RECT -30.085 218.115 -29.755 218.445 ;
        RECT -30.085 216.755 -29.755 217.085 ;
        RECT -30.085 215.395 -29.755 215.725 ;
        RECT -30.085 214.035 -29.755 214.365 ;
        RECT -30.085 212.675 -29.755 213.005 ;
        RECT -30.085 211.315 -29.755 211.645 ;
        RECT -30.085 209.955 -29.755 210.285 ;
        RECT -30.085 208.595 -29.755 208.925 ;
        RECT -30.085 207.235 -29.755 207.565 ;
        RECT -30.085 205.875 -29.755 206.205 ;
        RECT -30.085 204.515 -29.755 204.845 ;
        RECT -30.085 203.155 -29.755 203.485 ;
        RECT -30.085 201.795 -29.755 202.125 ;
        RECT -30.085 200.435 -29.755 200.765 ;
        RECT -30.085 199.075 -29.755 199.405 ;
        RECT -30.085 197.715 -29.755 198.045 ;
        RECT -30.085 196.355 -29.755 196.685 ;
        RECT -30.085 194.995 -29.755 195.325 ;
        RECT -30.085 193.635 -29.755 193.965 ;
        RECT -30.085 192.275 -29.755 192.605 ;
        RECT -30.085 190.915 -29.755 191.245 ;
        RECT -30.085 189.555 -29.755 189.885 ;
        RECT -30.085 188.195 -29.755 188.525 ;
        RECT -30.085 186.835 -29.755 187.165 ;
        RECT -30.085 185.475 -29.755 185.805 ;
        RECT -30.085 184.115 -29.755 184.445 ;
        RECT -30.085 182.755 -29.755 183.085 ;
        RECT -30.085 181.395 -29.755 181.725 ;
        RECT -30.085 180.035 -29.755 180.365 ;
        RECT -30.085 178.675 -29.755 179.005 ;
        RECT -30.085 177.315 -29.755 177.645 ;
        RECT -30.085 175.955 -29.755 176.285 ;
        RECT -30.085 174.595 -29.755 174.925 ;
        RECT -30.085 173.235 -29.755 173.565 ;
        RECT -30.085 171.875 -29.755 172.205 ;
        RECT -30.085 170.515 -29.755 170.845 ;
        RECT -30.085 169.155 -29.755 169.485 ;
        RECT -30.085 167.795 -29.755 168.125 ;
        RECT -30.085 166.435 -29.755 166.765 ;
        RECT -30.085 165.075 -29.755 165.405 ;
        RECT -30.085 163.715 -29.755 164.045 ;
        RECT -30.085 162.355 -29.755 162.685 ;
        RECT -30.085 160.995 -29.755 161.325 ;
        RECT -30.085 159.635 -29.755 159.965 ;
        RECT -30.085 158.275 -29.755 158.605 ;
        RECT -30.085 156.915 -29.755 157.245 ;
        RECT -30.085 155.555 -29.755 155.885 ;
        RECT -30.085 154.195 -29.755 154.525 ;
        RECT -30.085 152.835 -29.755 153.165 ;
        RECT -30.085 151.475 -29.755 151.805 ;
        RECT -30.085 150.115 -29.755 150.445 ;
        RECT -30.085 148.755 -29.755 149.085 ;
        RECT -30.085 147.395 -29.755 147.725 ;
        RECT -30.085 146.035 -29.755 146.365 ;
        RECT -30.085 144.675 -29.755 145.005 ;
        RECT -30.085 143.315 -29.755 143.645 ;
        RECT -30.085 141.955 -29.755 142.285 ;
        RECT -30.085 140.595 -29.755 140.925 ;
        RECT -30.085 139.235 -29.755 139.565 ;
        RECT -30.085 137.875 -29.755 138.205 ;
        RECT -30.085 136.515 -29.755 136.845 ;
        RECT -30.085 135.155 -29.755 135.485 ;
        RECT -30.085 133.795 -29.755 134.125 ;
        RECT -30.085 132.435 -29.755 132.765 ;
        RECT -30.085 131.075 -29.755 131.405 ;
        RECT -30.085 129.715 -29.755 130.045 ;
        RECT -30.085 128.355 -29.755 128.685 ;
        RECT -30.085 126.995 -29.755 127.325 ;
        RECT -30.085 125.635 -29.755 125.965 ;
        RECT -30.085 124.275 -29.755 124.605 ;
        RECT -30.085 122.915 -29.755 123.245 ;
        RECT -30.085 121.555 -29.755 121.885 ;
        RECT -30.085 120.195 -29.755 120.525 ;
        RECT -30.085 118.835 -29.755 119.165 ;
        RECT -30.085 117.475 -29.755 117.805 ;
        RECT -30.085 116.115 -29.755 116.445 ;
        RECT -30.085 114.755 -29.755 115.085 ;
        RECT -30.085 113.395 -29.755 113.725 ;
        RECT -30.085 112.035 -29.755 112.365 ;
        RECT -30.085 110.675 -29.755 111.005 ;
        RECT -30.085 109.315 -29.755 109.645 ;
        RECT -30.085 107.955 -29.755 108.285 ;
        RECT -30.085 106.595 -29.755 106.925 ;
        RECT -30.085 105.235 -29.755 105.565 ;
        RECT -30.085 103.875 -29.755 104.205 ;
        RECT -30.085 102.515 -29.755 102.845 ;
        RECT -30.085 101.155 -29.755 101.485 ;
        RECT -30.085 99.795 -29.755 100.125 ;
        RECT -30.085 98.435 -29.755 98.765 ;
        RECT -30.085 97.075 -29.755 97.405 ;
        RECT -30.085 95.715 -29.755 96.045 ;
        RECT -30.085 94.355 -29.755 94.685 ;
        RECT -30.085 92.995 -29.755 93.325 ;
        RECT -30.085 91.635 -29.755 91.965 ;
        RECT -30.085 90.275 -29.755 90.605 ;
        RECT -30.085 88.915 -29.755 89.245 ;
        RECT -30.085 87.555 -29.755 87.885 ;
        RECT -30.085 86.195 -29.755 86.525 ;
        RECT -30.085 84.835 -29.755 85.165 ;
        RECT -30.085 83.475 -29.755 83.805 ;
        RECT -30.085 82.115 -29.755 82.445 ;
        RECT -30.085 80.755 -29.755 81.085 ;
        RECT -30.085 79.395 -29.755 79.725 ;
        RECT -30.085 78.035 -29.755 78.365 ;
        RECT -30.085 76.675 -29.755 77.005 ;
        RECT -30.085 75.315 -29.755 75.645 ;
        RECT -30.085 73.955 -29.755 74.285 ;
        RECT -30.085 72.595 -29.755 72.925 ;
        RECT -30.085 71.235 -29.755 71.565 ;
        RECT -30.085 69.875 -29.755 70.205 ;
        RECT -30.085 68.515 -29.755 68.845 ;
        RECT -30.085 67.155 -29.755 67.485 ;
        RECT -30.085 65.795 -29.755 66.125 ;
        RECT -30.085 64.435 -29.755 64.765 ;
        RECT -30.085 63.075 -29.755 63.405 ;
        RECT -30.085 61.715 -29.755 62.045 ;
        RECT -30.085 60.355 -29.755 60.685 ;
        RECT -30.085 58.995 -29.755 59.325 ;
        RECT -30.085 57.635 -29.755 57.965 ;
        RECT -30.085 56.275 -29.755 56.605 ;
        RECT -30.085 54.915 -29.755 55.245 ;
        RECT -30.085 53.555 -29.755 53.885 ;
        RECT -30.085 52.195 -29.755 52.525 ;
        RECT -30.085 50.835 -29.755 51.165 ;
        RECT -30.085 49.475 -29.755 49.805 ;
        RECT -30.085 48.115 -29.755 48.445 ;
        RECT -30.085 46.755 -29.755 47.085 ;
        RECT -30.085 45.395 -29.755 45.725 ;
        RECT -30.085 44.035 -29.755 44.365 ;
        RECT -30.085 42.675 -29.755 43.005 ;
        RECT -30.085 41.315 -29.755 41.645 ;
        RECT -30.085 39.955 -29.755 40.285 ;
        RECT -30.085 38.595 -29.755 38.925 ;
        RECT -30.085 37.235 -29.755 37.565 ;
        RECT -30.085 35.875 -29.755 36.205 ;
        RECT -30.085 34.515 -29.755 34.845 ;
        RECT -30.085 33.155 -29.755 33.485 ;
        RECT -30.085 31.795 -29.755 32.125 ;
        RECT -30.085 30.435 -29.755 30.765 ;
        RECT -30.085 29.075 -29.755 29.405 ;
        RECT -30.085 27.715 -29.755 28.045 ;
        RECT -30.085 26.355 -29.755 26.685 ;
        RECT -30.085 24.995 -29.755 25.325 ;
        RECT -30.085 23.635 -29.755 23.965 ;
        RECT -30.085 22.275 -29.755 22.605 ;
        RECT -30.085 20.915 -29.755 21.245 ;
        RECT -30.085 19.555 -29.755 19.885 ;
        RECT -30.085 18.195 -29.755 18.525 ;
        RECT -30.085 16.835 -29.755 17.165 ;
        RECT -30.085 15.475 -29.755 15.805 ;
        RECT -30.085 14.115 -29.755 14.445 ;
        RECT -30.085 12.755 -29.755 13.085 ;
        RECT -30.085 11.395 -29.755 11.725 ;
        RECT -30.085 10.035 -29.755 10.365 ;
        RECT -30.085 8.675 -29.755 9.005 ;
        RECT -30.085 7.315 -29.755 7.645 ;
        RECT -30.085 5.955 -29.755 6.285 ;
        RECT -30.085 4.595 -29.755 4.925 ;
        RECT -30.085 3.235 -29.755 3.565 ;
        RECT -30.085 1.875 -29.755 2.205 ;
        RECT -30.085 0.515 -29.755 0.845 ;
        RECT -30.085 -0.845 -29.755 -0.515 ;
        RECT -30.085 -7.645 -29.755 -7.315 ;
        RECT -30.085 -9.005 -29.755 -8.675 ;
        RECT -30.085 -18.525 -29.755 -18.195 ;
        RECT -30.085 -21.245 -29.755 -20.915 ;
        RECT -30.085 -32.125 -29.755 -31.795 ;
        RECT -30.085 -33.71 -29.755 -33.38 ;
        RECT -30.085 -34.845 -29.755 -34.515 ;
        RECT -30.085 -36.205 -29.755 -35.875 ;
        RECT -30.085 -38.925 -29.755 -38.595 ;
        RECT -30.085 -39.75 -29.755 -39.42 ;
        RECT -30.085 -41.645 -29.755 -41.315 ;
        RECT -30.085 -44.365 -29.755 -44.035 ;
        RECT -30.085 -49.805 -29.755 -49.475 ;
        RECT -30.085 -51.165 -29.755 -50.835 ;
        RECT -30.085 -53.885 -29.755 -53.555 ;
        RECT -30.085 -55.245 -29.755 -54.915 ;
        RECT -30.085 -59.325 -29.755 -58.995 ;
        RECT -30.085 -60.685 -29.755 -60.355 ;
        RECT -30.085 -63.405 -29.755 -63.075 ;
        RECT -30.08 -64.08 -29.76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.085 -67.485 -29.755 -67.155 ;
        RECT -30.085 -70.205 -29.755 -69.875 ;
        RECT -30.085 -71.565 -29.755 -71.235 ;
        RECT -30.085 -74.285 -29.755 -73.955 ;
        RECT -30.085 -75.645 -29.755 -75.315 ;
        RECT -30.085 -78.365 -29.755 -78.035 ;
        RECT -30.085 -79.725 -29.755 -79.395 ;
        RECT -30.085 -82.445 -29.755 -82.115 ;
        RECT -30.085 -83.805 -29.755 -83.475 ;
        RECT -30.085 -86.525 -29.755 -86.195 ;
        RECT -30.085 -89.245 -29.755 -88.915 ;
        RECT -30.085 -90.605 -29.755 -90.275 ;
        RECT -30.085 -91.965 -29.755 -91.635 ;
        RECT -30.085 -93.325 -29.755 -92.995 ;
        RECT -30.085 -94.685 -29.755 -94.355 ;
        RECT -30.085 -97.405 -29.755 -97.075 ;
        RECT -30.085 -100.125 -29.755 -99.795 ;
        RECT -30.085 -101.485 -29.755 -101.155 ;
        RECT -30.085 -104.205 -29.755 -103.875 ;
        RECT -30.085 -105.565 -29.755 -105.235 ;
        RECT -30.085 -108.285 -29.755 -107.955 ;
        RECT -30.085 -113.725 -29.755 -113.395 ;
        RECT -30.085 -115.085 -29.755 -114.755 ;
        RECT -30.085 -116.445 -29.755 -116.115 ;
        RECT -30.085 -117.805 -29.755 -117.475 ;
        RECT -30.085 -119.165 -29.755 -118.835 ;
        RECT -30.085 -120.525 -29.755 -120.195 ;
        RECT -30.085 -123.245 -29.755 -122.915 ;
        RECT -30.085 -125.965 -29.755 -125.635 ;
        RECT -30.085 -127.325 -29.755 -126.995 ;
        RECT -30.085 -128.685 -29.755 -128.355 ;
        RECT -30.085 -130.045 -29.755 -129.715 ;
        RECT -30.085 -134.125 -29.755 -133.795 ;
        RECT -30.085 -135.485 -29.755 -135.155 ;
        RECT -30.085 -136.845 -29.755 -136.515 ;
        RECT -30.085 -139.565 -29.755 -139.235 ;
        RECT -30.085 -142.285 -29.755 -141.955 ;
        RECT -30.085 -143.645 -29.755 -143.315 ;
        RECT -30.085 -145.005 -29.755 -144.675 ;
        RECT -30.085 -146.365 -29.755 -146.035 ;
        RECT -30.085 -147.725 -29.755 -147.395 ;
        RECT -30.085 -149.085 -29.755 -148.755 ;
        RECT -30.085 -151.805 -29.755 -151.475 ;
        RECT -30.085 -153.165 -29.755 -152.835 ;
        RECT -30.085 -157.245 -29.755 -156.915 ;
        RECT -30.085 -158.605 -29.755 -158.275 ;
        RECT -30.085 -159.965 -29.755 -159.635 ;
        RECT -30.085 -161.325 -29.755 -160.995 ;
        RECT -30.085 -162.685 -29.755 -162.355 ;
        RECT -30.085 -164.045 -29.755 -163.715 ;
        RECT -30.085 -165.405 -29.755 -165.075 ;
        RECT -30.085 -166.765 -29.755 -166.435 ;
        RECT -30.085 -169.615 -29.755 -169.285 ;
        RECT -30.085 -170.845 -29.755 -170.515 ;
        RECT -30.085 -172.205 -29.755 -171.875 ;
        RECT -30.085 -173.565 -29.755 -173.235 ;
        RECT -30.085 -177.645 -29.755 -177.315 ;
        RECT -30.085 -179.005 -29.755 -178.675 ;
        RECT -30.085 -184.65 -29.755 -183.52 ;
        RECT -30.08 -184.765 -29.76 -67.155 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.725 244.04 -28.395 245.17 ;
        RECT -28.725 239.875 -28.395 240.205 ;
        RECT -28.725 238.515 -28.395 238.845 ;
        RECT -28.725 237.155 -28.395 237.485 ;
        RECT -28.725 235.795 -28.395 236.125 ;
        RECT -28.725 234.435 -28.395 234.765 ;
        RECT -28.725 233.075 -28.395 233.405 ;
        RECT -28.725 231.715 -28.395 232.045 ;
        RECT -28.725 230.355 -28.395 230.685 ;
        RECT -28.725 228.995 -28.395 229.325 ;
        RECT -28.725 227.635 -28.395 227.965 ;
        RECT -28.725 226.275 -28.395 226.605 ;
        RECT -28.725 224.915 -28.395 225.245 ;
        RECT -28.725 223.555 -28.395 223.885 ;
        RECT -28.725 222.195 -28.395 222.525 ;
        RECT -28.725 220.835 -28.395 221.165 ;
        RECT -28.725 219.475 -28.395 219.805 ;
        RECT -28.725 218.115 -28.395 218.445 ;
        RECT -28.725 216.755 -28.395 217.085 ;
        RECT -28.725 215.395 -28.395 215.725 ;
        RECT -28.725 214.035 -28.395 214.365 ;
        RECT -28.725 212.675 -28.395 213.005 ;
        RECT -28.725 211.315 -28.395 211.645 ;
        RECT -28.725 209.955 -28.395 210.285 ;
        RECT -28.725 208.595 -28.395 208.925 ;
        RECT -28.725 207.235 -28.395 207.565 ;
        RECT -28.725 205.875 -28.395 206.205 ;
        RECT -28.725 204.515 -28.395 204.845 ;
        RECT -28.725 203.155 -28.395 203.485 ;
        RECT -28.725 201.795 -28.395 202.125 ;
        RECT -28.725 200.435 -28.395 200.765 ;
        RECT -28.725 199.075 -28.395 199.405 ;
        RECT -28.725 197.715 -28.395 198.045 ;
        RECT -28.725 196.355 -28.395 196.685 ;
        RECT -28.725 194.995 -28.395 195.325 ;
        RECT -28.725 193.635 -28.395 193.965 ;
        RECT -28.725 192.275 -28.395 192.605 ;
        RECT -28.725 190.915 -28.395 191.245 ;
        RECT -28.725 189.555 -28.395 189.885 ;
        RECT -28.725 188.195 -28.395 188.525 ;
        RECT -28.725 186.835 -28.395 187.165 ;
        RECT -28.725 185.475 -28.395 185.805 ;
        RECT -28.725 184.115 -28.395 184.445 ;
        RECT -28.725 182.755 -28.395 183.085 ;
        RECT -28.725 181.395 -28.395 181.725 ;
        RECT -28.725 180.035 -28.395 180.365 ;
        RECT -28.725 178.675 -28.395 179.005 ;
        RECT -28.725 177.315 -28.395 177.645 ;
        RECT -28.725 175.955 -28.395 176.285 ;
        RECT -28.725 174.595 -28.395 174.925 ;
        RECT -28.725 173.235 -28.395 173.565 ;
        RECT -28.725 171.875 -28.395 172.205 ;
        RECT -28.725 170.515 -28.395 170.845 ;
        RECT -28.725 169.155 -28.395 169.485 ;
        RECT -28.725 167.795 -28.395 168.125 ;
        RECT -28.725 166.435 -28.395 166.765 ;
        RECT -28.725 165.075 -28.395 165.405 ;
        RECT -28.725 163.715 -28.395 164.045 ;
        RECT -28.725 162.355 -28.395 162.685 ;
        RECT -28.725 160.995 -28.395 161.325 ;
        RECT -28.725 159.635 -28.395 159.965 ;
        RECT -28.725 158.275 -28.395 158.605 ;
        RECT -28.725 156.915 -28.395 157.245 ;
        RECT -28.725 155.555 -28.395 155.885 ;
        RECT -28.725 154.195 -28.395 154.525 ;
        RECT -28.725 152.835 -28.395 153.165 ;
        RECT -28.725 151.475 -28.395 151.805 ;
        RECT -28.725 150.115 -28.395 150.445 ;
        RECT -28.725 148.755 -28.395 149.085 ;
        RECT -28.725 147.395 -28.395 147.725 ;
        RECT -28.725 146.035 -28.395 146.365 ;
        RECT -28.725 144.675 -28.395 145.005 ;
        RECT -28.725 143.315 -28.395 143.645 ;
        RECT -28.725 141.955 -28.395 142.285 ;
        RECT -28.725 140.595 -28.395 140.925 ;
        RECT -28.725 139.235 -28.395 139.565 ;
        RECT -28.725 137.875 -28.395 138.205 ;
        RECT -28.725 136.515 -28.395 136.845 ;
        RECT -28.725 135.155 -28.395 135.485 ;
        RECT -28.725 133.795 -28.395 134.125 ;
        RECT -28.725 132.435 -28.395 132.765 ;
        RECT -28.725 131.075 -28.395 131.405 ;
        RECT -28.725 129.715 -28.395 130.045 ;
        RECT -28.725 128.355 -28.395 128.685 ;
        RECT -28.725 126.995 -28.395 127.325 ;
        RECT -28.725 125.635 -28.395 125.965 ;
        RECT -28.725 124.275 -28.395 124.605 ;
        RECT -28.725 122.915 -28.395 123.245 ;
        RECT -28.725 121.555 -28.395 121.885 ;
        RECT -28.725 120.195 -28.395 120.525 ;
        RECT -28.725 118.835 -28.395 119.165 ;
        RECT -28.725 117.475 -28.395 117.805 ;
        RECT -28.725 116.115 -28.395 116.445 ;
        RECT -28.725 114.755 -28.395 115.085 ;
        RECT -28.725 113.395 -28.395 113.725 ;
        RECT -28.725 112.035 -28.395 112.365 ;
        RECT -28.725 110.675 -28.395 111.005 ;
        RECT -28.725 109.315 -28.395 109.645 ;
        RECT -28.725 107.955 -28.395 108.285 ;
        RECT -28.725 106.595 -28.395 106.925 ;
        RECT -28.725 105.235 -28.395 105.565 ;
        RECT -28.725 103.875 -28.395 104.205 ;
        RECT -28.725 102.515 -28.395 102.845 ;
        RECT -28.725 101.155 -28.395 101.485 ;
        RECT -28.725 99.795 -28.395 100.125 ;
        RECT -28.725 98.435 -28.395 98.765 ;
        RECT -28.725 97.075 -28.395 97.405 ;
        RECT -28.725 95.715 -28.395 96.045 ;
        RECT -28.725 94.355 -28.395 94.685 ;
        RECT -28.725 92.995 -28.395 93.325 ;
        RECT -28.725 91.635 -28.395 91.965 ;
        RECT -28.725 90.275 -28.395 90.605 ;
        RECT -28.725 88.915 -28.395 89.245 ;
        RECT -28.725 87.555 -28.395 87.885 ;
        RECT -28.725 86.195 -28.395 86.525 ;
        RECT -28.725 84.835 -28.395 85.165 ;
        RECT -28.725 83.475 -28.395 83.805 ;
        RECT -28.725 82.115 -28.395 82.445 ;
        RECT -28.725 80.755 -28.395 81.085 ;
        RECT -28.725 79.395 -28.395 79.725 ;
        RECT -28.725 78.035 -28.395 78.365 ;
        RECT -28.725 76.675 -28.395 77.005 ;
        RECT -28.725 75.315 -28.395 75.645 ;
        RECT -28.725 73.955 -28.395 74.285 ;
        RECT -28.725 72.595 -28.395 72.925 ;
        RECT -28.725 71.235 -28.395 71.565 ;
        RECT -28.725 69.875 -28.395 70.205 ;
        RECT -28.725 68.515 -28.395 68.845 ;
        RECT -28.725 67.155 -28.395 67.485 ;
        RECT -28.725 65.795 -28.395 66.125 ;
        RECT -28.725 64.435 -28.395 64.765 ;
        RECT -28.725 63.075 -28.395 63.405 ;
        RECT -28.725 61.715 -28.395 62.045 ;
        RECT -28.725 60.355 -28.395 60.685 ;
        RECT -28.725 58.995 -28.395 59.325 ;
        RECT -28.725 57.635 -28.395 57.965 ;
        RECT -28.725 56.275 -28.395 56.605 ;
        RECT -28.725 54.915 -28.395 55.245 ;
        RECT -28.725 53.555 -28.395 53.885 ;
        RECT -28.725 52.195 -28.395 52.525 ;
        RECT -28.725 50.835 -28.395 51.165 ;
        RECT -28.725 49.475 -28.395 49.805 ;
        RECT -28.725 48.115 -28.395 48.445 ;
        RECT -28.725 46.755 -28.395 47.085 ;
        RECT -28.725 45.395 -28.395 45.725 ;
        RECT -28.725 44.035 -28.395 44.365 ;
        RECT -28.725 42.675 -28.395 43.005 ;
        RECT -28.725 41.315 -28.395 41.645 ;
        RECT -28.725 39.955 -28.395 40.285 ;
        RECT -28.725 38.595 -28.395 38.925 ;
        RECT -28.725 37.235 -28.395 37.565 ;
        RECT -28.725 35.875 -28.395 36.205 ;
        RECT -28.725 34.515 -28.395 34.845 ;
        RECT -28.725 33.155 -28.395 33.485 ;
        RECT -28.725 31.795 -28.395 32.125 ;
        RECT -28.725 30.435 -28.395 30.765 ;
        RECT -28.725 29.075 -28.395 29.405 ;
        RECT -28.725 27.715 -28.395 28.045 ;
        RECT -28.725 26.355 -28.395 26.685 ;
        RECT -28.725 24.995 -28.395 25.325 ;
        RECT -28.725 23.635 -28.395 23.965 ;
        RECT -28.725 22.275 -28.395 22.605 ;
        RECT -28.725 20.915 -28.395 21.245 ;
        RECT -28.725 19.555 -28.395 19.885 ;
        RECT -28.725 18.195 -28.395 18.525 ;
        RECT -28.725 16.835 -28.395 17.165 ;
        RECT -28.725 15.475 -28.395 15.805 ;
        RECT -28.725 14.115 -28.395 14.445 ;
        RECT -28.725 12.755 -28.395 13.085 ;
        RECT -28.725 11.395 -28.395 11.725 ;
        RECT -28.725 10.035 -28.395 10.365 ;
        RECT -28.725 8.675 -28.395 9.005 ;
        RECT -28.725 7.315 -28.395 7.645 ;
        RECT -28.725 5.955 -28.395 6.285 ;
        RECT -28.725 4.595 -28.395 4.925 ;
        RECT -28.725 3.235 -28.395 3.565 ;
        RECT -28.725 1.875 -28.395 2.205 ;
        RECT -28.725 0.515 -28.395 0.845 ;
        RECT -28.725 -0.845 -28.395 -0.515 ;
        RECT -28.725 -7.645 -28.395 -7.315 ;
        RECT -28.725 -9.005 -28.395 -8.675 ;
        RECT -28.725 -10.73 -28.395 -10.4 ;
        RECT -28.725 -16.77 -28.395 -16.44 ;
        RECT -28.725 -18.525 -28.395 -18.195 ;
        RECT -28.725 -21.245 -28.395 -20.915 ;
        RECT -28.725 -32.125 -28.395 -31.795 ;
        RECT -28.725 -33.71 -28.395 -33.38 ;
        RECT -28.725 -34.845 -28.395 -34.515 ;
        RECT -28.725 -36.205 -28.395 -35.875 ;
        RECT -28.725 -38.925 -28.395 -38.595 ;
        RECT -28.725 -39.75 -28.395 -39.42 ;
        RECT -28.725 -41.645 -28.395 -41.315 ;
        RECT -28.725 -44.365 -28.395 -44.035 ;
        RECT -28.725 -49.805 -28.395 -49.475 ;
        RECT -28.725 -51.165 -28.395 -50.835 ;
        RECT -28.725 -53.885 -28.395 -53.555 ;
        RECT -28.725 -55.245 -28.395 -54.915 ;
        RECT -28.725 -59.325 -28.395 -58.995 ;
        RECT -28.725 -60.685 -28.395 -60.355 ;
        RECT -28.725 -63.405 -28.395 -63.075 ;
        RECT -28.72 -63.405 -28.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.725 -70.205 -28.395 -69.875 ;
        RECT -28.725 -71.565 -28.395 -71.235 ;
        RECT -28.725 -73.19 -28.395 -72.86 ;
        RECT -28.725 -74.285 -28.395 -73.955 ;
        RECT -28.725 -75.645 -28.395 -75.315 ;
        RECT -28.725 -78.365 -28.395 -78.035 ;
        RECT -28.725 -79.725 -28.395 -79.395 ;
        RECT -28.725 -80.73 -28.395 -80.4 ;
        RECT -28.725 -82.445 -28.395 -82.115 ;
        RECT -28.725 -83.805 -28.395 -83.475 ;
        RECT -28.725 -86.525 -28.395 -86.195 ;
        RECT -28.725 -89.245 -28.395 -88.915 ;
        RECT -28.725 -90.605 -28.395 -90.275 ;
        RECT -28.725 -91.965 -28.395 -91.635 ;
        RECT -28.725 -93.325 -28.395 -92.995 ;
        RECT -28.725 -94.685 -28.395 -94.355 ;
        RECT -28.725 -95.37 -28.395 -95.04 ;
        RECT -28.725 -97.405 -28.395 -97.075 ;
        RECT -28.725 -100.125 -28.395 -99.795 ;
        RECT -28.725 -101.485 -28.395 -101.155 ;
        RECT -28.725 -102.91 -28.395 -102.58 ;
        RECT -28.725 -104.205 -28.395 -103.875 ;
        RECT -28.725 -105.565 -28.395 -105.235 ;
        RECT -28.725 -108.285 -28.395 -107.955 ;
        RECT -28.725 -115.085 -28.395 -114.755 ;
        RECT -28.725 -116.445 -28.395 -116.115 ;
        RECT -28.725 -117.805 -28.395 -117.475 ;
        RECT -28.725 -119.165 -28.395 -118.835 ;
        RECT -28.725 -120.525 -28.395 -120.195 ;
        RECT -28.725 -123.245 -28.395 -122.915 ;
        RECT -28.725 -125.965 -28.395 -125.635 ;
        RECT -28.725 -127.325 -28.395 -126.995 ;
        RECT -28.725 -128.685 -28.395 -128.355 ;
        RECT -28.725 -130.045 -28.395 -129.715 ;
        RECT -28.725 -134.125 -28.395 -133.795 ;
        RECT -28.725 -135.485 -28.395 -135.155 ;
        RECT -28.725 -136.845 -28.395 -136.515 ;
        RECT -28.725 -139.565 -28.395 -139.235 ;
        RECT -28.725 -142.285 -28.395 -141.955 ;
        RECT -28.725 -143.645 -28.395 -143.315 ;
        RECT -28.725 -145.005 -28.395 -144.675 ;
        RECT -28.725 -146.365 -28.395 -146.035 ;
        RECT -28.725 -147.725 -28.395 -147.395 ;
        RECT -28.725 -149.085 -28.395 -148.755 ;
        RECT -28.725 -151.805 -28.395 -151.475 ;
        RECT -28.725 -153.165 -28.395 -152.835 ;
        RECT -28.725 -157.245 -28.395 -156.915 ;
        RECT -28.725 -158.605 -28.395 -158.275 ;
        RECT -28.725 -159.965 -28.395 -159.635 ;
        RECT -28.725 -161.325 -28.395 -160.995 ;
        RECT -28.725 -162.685 -28.395 -162.355 ;
        RECT -28.725 -164.045 -28.395 -163.715 ;
        RECT -28.725 -165.405 -28.395 -165.075 ;
        RECT -28.725 -166.765 -28.395 -166.435 ;
        RECT -28.725 -170.845 -28.395 -170.515 ;
        RECT -28.725 -172.205 -28.395 -171.875 ;
        RECT -28.725 -177.645 -28.395 -177.315 ;
        RECT -28.725 -179.005 -28.395 -178.675 ;
        RECT -28.725 -184.65 -28.395 -183.52 ;
        RECT -28.72 -184.765 -28.4 -69.2 ;
    END
    PORT
      LAYER met3 ;
        RECT -27.365 125.635 -27.035 125.965 ;
        RECT -27.365 124.275 -27.035 124.605 ;
        RECT -27.365 122.915 -27.035 123.245 ;
        RECT -27.365 121.555 -27.035 121.885 ;
        RECT -27.365 120.195 -27.035 120.525 ;
        RECT -27.365 118.835 -27.035 119.165 ;
        RECT -27.365 117.475 -27.035 117.805 ;
        RECT -27.365 116.115 -27.035 116.445 ;
        RECT -27.365 114.755 -27.035 115.085 ;
        RECT -27.365 113.395 -27.035 113.725 ;
        RECT -27.365 112.035 -27.035 112.365 ;
        RECT -27.365 110.675 -27.035 111.005 ;
        RECT -27.365 109.315 -27.035 109.645 ;
        RECT -27.365 107.955 -27.035 108.285 ;
        RECT -27.365 106.595 -27.035 106.925 ;
        RECT -27.365 105.235 -27.035 105.565 ;
        RECT -27.365 103.875 -27.035 104.205 ;
        RECT -27.365 102.515 -27.035 102.845 ;
        RECT -27.365 101.155 -27.035 101.485 ;
        RECT -27.365 99.795 -27.035 100.125 ;
        RECT -27.365 98.435 -27.035 98.765 ;
        RECT -27.365 97.075 -27.035 97.405 ;
        RECT -27.365 95.715 -27.035 96.045 ;
        RECT -27.365 94.355 -27.035 94.685 ;
        RECT -27.365 92.995 -27.035 93.325 ;
        RECT -27.365 91.635 -27.035 91.965 ;
        RECT -27.365 90.275 -27.035 90.605 ;
        RECT -27.365 88.915 -27.035 89.245 ;
        RECT -27.365 87.555 -27.035 87.885 ;
        RECT -27.365 86.195 -27.035 86.525 ;
        RECT -27.365 84.835 -27.035 85.165 ;
        RECT -27.365 83.475 -27.035 83.805 ;
        RECT -27.365 82.115 -27.035 82.445 ;
        RECT -27.365 80.755 -27.035 81.085 ;
        RECT -27.365 79.395 -27.035 79.725 ;
        RECT -27.365 78.035 -27.035 78.365 ;
        RECT -27.365 76.675 -27.035 77.005 ;
        RECT -27.365 75.315 -27.035 75.645 ;
        RECT -27.365 73.955 -27.035 74.285 ;
        RECT -27.365 72.595 -27.035 72.925 ;
        RECT -27.365 71.235 -27.035 71.565 ;
        RECT -27.365 69.875 -27.035 70.205 ;
        RECT -27.365 68.515 -27.035 68.845 ;
        RECT -27.365 67.155 -27.035 67.485 ;
        RECT -27.365 65.795 -27.035 66.125 ;
        RECT -27.365 64.435 -27.035 64.765 ;
        RECT -27.365 63.075 -27.035 63.405 ;
        RECT -27.365 61.715 -27.035 62.045 ;
        RECT -27.365 60.355 -27.035 60.685 ;
        RECT -27.365 58.995 -27.035 59.325 ;
        RECT -27.365 57.635 -27.035 57.965 ;
        RECT -27.365 56.275 -27.035 56.605 ;
        RECT -27.365 54.915 -27.035 55.245 ;
        RECT -27.365 53.555 -27.035 53.885 ;
        RECT -27.365 52.195 -27.035 52.525 ;
        RECT -27.365 50.835 -27.035 51.165 ;
        RECT -27.365 49.475 -27.035 49.805 ;
        RECT -27.365 48.115 -27.035 48.445 ;
        RECT -27.365 46.755 -27.035 47.085 ;
        RECT -27.365 45.395 -27.035 45.725 ;
        RECT -27.365 44.035 -27.035 44.365 ;
        RECT -27.365 42.675 -27.035 43.005 ;
        RECT -27.365 41.315 -27.035 41.645 ;
        RECT -27.365 39.955 -27.035 40.285 ;
        RECT -27.365 38.595 -27.035 38.925 ;
        RECT -27.365 37.235 -27.035 37.565 ;
        RECT -27.365 35.875 -27.035 36.205 ;
        RECT -27.365 34.515 -27.035 34.845 ;
        RECT -27.365 33.155 -27.035 33.485 ;
        RECT -27.365 31.795 -27.035 32.125 ;
        RECT -27.365 30.435 -27.035 30.765 ;
        RECT -27.365 29.075 -27.035 29.405 ;
        RECT -27.365 27.715 -27.035 28.045 ;
        RECT -27.365 26.355 -27.035 26.685 ;
        RECT -27.365 24.995 -27.035 25.325 ;
        RECT -27.365 23.635 -27.035 23.965 ;
        RECT -27.365 22.275 -27.035 22.605 ;
        RECT -27.365 20.915 -27.035 21.245 ;
        RECT -27.365 19.555 -27.035 19.885 ;
        RECT -27.365 18.195 -27.035 18.525 ;
        RECT -27.365 16.835 -27.035 17.165 ;
        RECT -27.365 15.475 -27.035 15.805 ;
        RECT -27.365 14.115 -27.035 14.445 ;
        RECT -27.365 12.755 -27.035 13.085 ;
        RECT -27.365 11.395 -27.035 11.725 ;
        RECT -27.365 10.035 -27.035 10.365 ;
        RECT -27.365 8.675 -27.035 9.005 ;
        RECT -27.365 7.315 -27.035 7.645 ;
        RECT -27.365 5.955 -27.035 6.285 ;
        RECT -27.365 4.595 -27.035 4.925 ;
        RECT -27.365 3.235 -27.035 3.565 ;
        RECT -27.365 1.875 -27.035 2.205 ;
        RECT -27.365 0.515 -27.035 0.845 ;
        RECT -27.365 -0.845 -27.035 -0.515 ;
        RECT -27.365 -2.205 -27.035 -1.875 ;
        RECT -27.365 -7.645 -27.035 -7.315 ;
        RECT -27.365 -9.005 -27.035 -8.675 ;
        RECT -27.365 -10.73 -27.035 -10.4 ;
        RECT -27.36 -11.04 -27.04 245.285 ;
        RECT -27.365 244.04 -27.035 245.17 ;
        RECT -27.365 239.875 -27.035 240.205 ;
        RECT -27.365 238.515 -27.035 238.845 ;
        RECT -27.365 237.155 -27.035 237.485 ;
        RECT -27.365 235.795 -27.035 236.125 ;
        RECT -27.365 234.435 -27.035 234.765 ;
        RECT -27.365 233.075 -27.035 233.405 ;
        RECT -27.365 231.715 -27.035 232.045 ;
        RECT -27.365 230.355 -27.035 230.685 ;
        RECT -27.365 228.995 -27.035 229.325 ;
        RECT -27.365 227.635 -27.035 227.965 ;
        RECT -27.365 226.275 -27.035 226.605 ;
        RECT -27.365 224.915 -27.035 225.245 ;
        RECT -27.365 223.555 -27.035 223.885 ;
        RECT -27.365 222.195 -27.035 222.525 ;
        RECT -27.365 220.835 -27.035 221.165 ;
        RECT -27.365 219.475 -27.035 219.805 ;
        RECT -27.365 218.115 -27.035 218.445 ;
        RECT -27.365 216.755 -27.035 217.085 ;
        RECT -27.365 215.395 -27.035 215.725 ;
        RECT -27.365 214.035 -27.035 214.365 ;
        RECT -27.365 212.675 -27.035 213.005 ;
        RECT -27.365 211.315 -27.035 211.645 ;
        RECT -27.365 209.955 -27.035 210.285 ;
        RECT -27.365 208.595 -27.035 208.925 ;
        RECT -27.365 207.235 -27.035 207.565 ;
        RECT -27.365 205.875 -27.035 206.205 ;
        RECT -27.365 204.515 -27.035 204.845 ;
        RECT -27.365 203.155 -27.035 203.485 ;
        RECT -27.365 201.795 -27.035 202.125 ;
        RECT -27.365 200.435 -27.035 200.765 ;
        RECT -27.365 199.075 -27.035 199.405 ;
        RECT -27.365 197.715 -27.035 198.045 ;
        RECT -27.365 196.355 -27.035 196.685 ;
        RECT -27.365 194.995 -27.035 195.325 ;
        RECT -27.365 193.635 -27.035 193.965 ;
        RECT -27.365 192.275 -27.035 192.605 ;
        RECT -27.365 190.915 -27.035 191.245 ;
        RECT -27.365 189.555 -27.035 189.885 ;
        RECT -27.365 188.195 -27.035 188.525 ;
        RECT -27.365 186.835 -27.035 187.165 ;
        RECT -27.365 185.475 -27.035 185.805 ;
        RECT -27.365 184.115 -27.035 184.445 ;
        RECT -27.365 182.755 -27.035 183.085 ;
        RECT -27.365 181.395 -27.035 181.725 ;
        RECT -27.365 180.035 -27.035 180.365 ;
        RECT -27.365 178.675 -27.035 179.005 ;
        RECT -27.365 177.315 -27.035 177.645 ;
        RECT -27.365 175.955 -27.035 176.285 ;
        RECT -27.365 174.595 -27.035 174.925 ;
        RECT -27.365 173.235 -27.035 173.565 ;
        RECT -27.365 171.875 -27.035 172.205 ;
        RECT -27.365 170.515 -27.035 170.845 ;
        RECT -27.365 169.155 -27.035 169.485 ;
        RECT -27.365 167.795 -27.035 168.125 ;
        RECT -27.365 166.435 -27.035 166.765 ;
        RECT -27.365 165.075 -27.035 165.405 ;
        RECT -27.365 163.715 -27.035 164.045 ;
        RECT -27.365 162.355 -27.035 162.685 ;
        RECT -27.365 160.995 -27.035 161.325 ;
        RECT -27.365 159.635 -27.035 159.965 ;
        RECT -27.365 158.275 -27.035 158.605 ;
        RECT -27.365 156.915 -27.035 157.245 ;
        RECT -27.365 155.555 -27.035 155.885 ;
        RECT -27.365 154.195 -27.035 154.525 ;
        RECT -27.365 152.835 -27.035 153.165 ;
        RECT -27.365 151.475 -27.035 151.805 ;
        RECT -27.365 150.115 -27.035 150.445 ;
        RECT -27.365 148.755 -27.035 149.085 ;
        RECT -27.365 147.395 -27.035 147.725 ;
        RECT -27.365 146.035 -27.035 146.365 ;
        RECT -27.365 144.675 -27.035 145.005 ;
        RECT -27.365 143.315 -27.035 143.645 ;
        RECT -27.365 141.955 -27.035 142.285 ;
        RECT -27.365 140.595 -27.035 140.925 ;
        RECT -27.365 139.235 -27.035 139.565 ;
        RECT -27.365 137.875 -27.035 138.205 ;
        RECT -27.365 136.515 -27.035 136.845 ;
        RECT -27.365 135.155 -27.035 135.485 ;
        RECT -27.365 133.795 -27.035 134.125 ;
        RECT -27.365 132.435 -27.035 132.765 ;
        RECT -27.365 131.075 -27.035 131.405 ;
        RECT -27.365 129.715 -27.035 130.045 ;
        RECT -27.365 128.355 -27.035 128.685 ;
        RECT -27.365 126.995 -27.035 127.325 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.245 -173.565 -37.915 -173.235 ;
        RECT -38.245 -174.925 -37.915 -174.595 ;
        RECT -38.245 -177.645 -37.915 -177.315 ;
        RECT -38.245 -179.005 -37.915 -178.675 ;
        RECT -38.245 -184.65 -37.915 -183.52 ;
        RECT -38.24 -184.765 -37.92 -173.235 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.885 244.04 -36.555 245.17 ;
        RECT -36.885 239.875 -36.555 240.205 ;
        RECT -36.885 238.515 -36.555 238.845 ;
        RECT -36.885 237.155 -36.555 237.485 ;
        RECT -36.885 235.795 -36.555 236.125 ;
        RECT -36.885 234.435 -36.555 234.765 ;
        RECT -36.885 233.075 -36.555 233.405 ;
        RECT -36.885 231.715 -36.555 232.045 ;
        RECT -36.885 230.355 -36.555 230.685 ;
        RECT -36.885 228.995 -36.555 229.325 ;
        RECT -36.885 227.635 -36.555 227.965 ;
        RECT -36.885 226.275 -36.555 226.605 ;
        RECT -36.885 224.915 -36.555 225.245 ;
        RECT -36.885 223.555 -36.555 223.885 ;
        RECT -36.885 222.195 -36.555 222.525 ;
        RECT -36.885 220.835 -36.555 221.165 ;
        RECT -36.885 219.475 -36.555 219.805 ;
        RECT -36.885 218.115 -36.555 218.445 ;
        RECT -36.885 216.755 -36.555 217.085 ;
        RECT -36.885 215.395 -36.555 215.725 ;
        RECT -36.885 214.035 -36.555 214.365 ;
        RECT -36.885 212.675 -36.555 213.005 ;
        RECT -36.885 211.315 -36.555 211.645 ;
        RECT -36.885 209.955 -36.555 210.285 ;
        RECT -36.885 208.595 -36.555 208.925 ;
        RECT -36.885 207.235 -36.555 207.565 ;
        RECT -36.885 205.875 -36.555 206.205 ;
        RECT -36.885 204.515 -36.555 204.845 ;
        RECT -36.885 203.155 -36.555 203.485 ;
        RECT -36.885 201.795 -36.555 202.125 ;
        RECT -36.885 200.435 -36.555 200.765 ;
        RECT -36.885 199.075 -36.555 199.405 ;
        RECT -36.885 197.715 -36.555 198.045 ;
        RECT -36.885 196.355 -36.555 196.685 ;
        RECT -36.885 194.995 -36.555 195.325 ;
        RECT -36.885 193.635 -36.555 193.965 ;
        RECT -36.885 192.275 -36.555 192.605 ;
        RECT -36.885 190.915 -36.555 191.245 ;
        RECT -36.885 189.555 -36.555 189.885 ;
        RECT -36.885 188.195 -36.555 188.525 ;
        RECT -36.885 186.835 -36.555 187.165 ;
        RECT -36.885 185.475 -36.555 185.805 ;
        RECT -36.885 184.115 -36.555 184.445 ;
        RECT -36.885 182.755 -36.555 183.085 ;
        RECT -36.885 181.395 -36.555 181.725 ;
        RECT -36.885 180.035 -36.555 180.365 ;
        RECT -36.885 178.675 -36.555 179.005 ;
        RECT -36.885 177.315 -36.555 177.645 ;
        RECT -36.885 175.955 -36.555 176.285 ;
        RECT -36.885 174.595 -36.555 174.925 ;
        RECT -36.885 173.235 -36.555 173.565 ;
        RECT -36.885 171.875 -36.555 172.205 ;
        RECT -36.885 170.515 -36.555 170.845 ;
        RECT -36.885 169.155 -36.555 169.485 ;
        RECT -36.885 167.795 -36.555 168.125 ;
        RECT -36.885 166.435 -36.555 166.765 ;
        RECT -36.885 165.075 -36.555 165.405 ;
        RECT -36.885 163.715 -36.555 164.045 ;
        RECT -36.885 162.355 -36.555 162.685 ;
        RECT -36.885 160.995 -36.555 161.325 ;
        RECT -36.885 159.635 -36.555 159.965 ;
        RECT -36.885 158.275 -36.555 158.605 ;
        RECT -36.885 156.915 -36.555 157.245 ;
        RECT -36.885 155.555 -36.555 155.885 ;
        RECT -36.885 154.195 -36.555 154.525 ;
        RECT -36.885 152.835 -36.555 153.165 ;
        RECT -36.885 151.475 -36.555 151.805 ;
        RECT -36.885 150.115 -36.555 150.445 ;
        RECT -36.885 148.755 -36.555 149.085 ;
        RECT -36.885 147.395 -36.555 147.725 ;
        RECT -36.885 146.035 -36.555 146.365 ;
        RECT -36.885 144.675 -36.555 145.005 ;
        RECT -36.885 143.315 -36.555 143.645 ;
        RECT -36.885 141.955 -36.555 142.285 ;
        RECT -36.885 140.595 -36.555 140.925 ;
        RECT -36.885 139.235 -36.555 139.565 ;
        RECT -36.885 137.875 -36.555 138.205 ;
        RECT -36.885 136.515 -36.555 136.845 ;
        RECT -36.885 135.155 -36.555 135.485 ;
        RECT -36.885 133.795 -36.555 134.125 ;
        RECT -36.885 132.435 -36.555 132.765 ;
        RECT -36.885 131.075 -36.555 131.405 ;
        RECT -36.885 129.715 -36.555 130.045 ;
        RECT -36.885 128.355 -36.555 128.685 ;
        RECT -36.885 126.995 -36.555 127.325 ;
        RECT -36.885 125.635 -36.555 125.965 ;
        RECT -36.885 124.275 -36.555 124.605 ;
        RECT -36.885 122.915 -36.555 123.245 ;
        RECT -36.885 121.555 -36.555 121.885 ;
        RECT -36.885 120.195 -36.555 120.525 ;
        RECT -36.885 118.835 -36.555 119.165 ;
        RECT -36.885 117.475 -36.555 117.805 ;
        RECT -36.885 116.115 -36.555 116.445 ;
        RECT -36.885 114.755 -36.555 115.085 ;
        RECT -36.885 113.395 -36.555 113.725 ;
        RECT -36.885 112.035 -36.555 112.365 ;
        RECT -36.885 110.675 -36.555 111.005 ;
        RECT -36.885 109.315 -36.555 109.645 ;
        RECT -36.885 107.955 -36.555 108.285 ;
        RECT -36.885 106.595 -36.555 106.925 ;
        RECT -36.885 105.235 -36.555 105.565 ;
        RECT -36.885 103.875 -36.555 104.205 ;
        RECT -36.885 102.515 -36.555 102.845 ;
        RECT -36.885 101.155 -36.555 101.485 ;
        RECT -36.885 99.795 -36.555 100.125 ;
        RECT -36.885 98.435 -36.555 98.765 ;
        RECT -36.885 97.075 -36.555 97.405 ;
        RECT -36.885 95.715 -36.555 96.045 ;
        RECT -36.885 94.355 -36.555 94.685 ;
        RECT -36.885 92.995 -36.555 93.325 ;
        RECT -36.885 91.635 -36.555 91.965 ;
        RECT -36.885 90.275 -36.555 90.605 ;
        RECT -36.885 88.915 -36.555 89.245 ;
        RECT -36.885 87.555 -36.555 87.885 ;
        RECT -36.885 86.195 -36.555 86.525 ;
        RECT -36.885 84.835 -36.555 85.165 ;
        RECT -36.885 83.475 -36.555 83.805 ;
        RECT -36.885 82.115 -36.555 82.445 ;
        RECT -36.885 80.755 -36.555 81.085 ;
        RECT -36.885 79.395 -36.555 79.725 ;
        RECT -36.885 78.035 -36.555 78.365 ;
        RECT -36.885 76.675 -36.555 77.005 ;
        RECT -36.885 75.315 -36.555 75.645 ;
        RECT -36.885 73.955 -36.555 74.285 ;
        RECT -36.885 72.595 -36.555 72.925 ;
        RECT -36.885 71.235 -36.555 71.565 ;
        RECT -36.885 69.875 -36.555 70.205 ;
        RECT -36.885 68.515 -36.555 68.845 ;
        RECT -36.885 67.155 -36.555 67.485 ;
        RECT -36.885 65.795 -36.555 66.125 ;
        RECT -36.885 64.435 -36.555 64.765 ;
        RECT -36.885 63.075 -36.555 63.405 ;
        RECT -36.885 61.715 -36.555 62.045 ;
        RECT -36.885 60.355 -36.555 60.685 ;
        RECT -36.885 58.995 -36.555 59.325 ;
        RECT -36.885 57.635 -36.555 57.965 ;
        RECT -36.885 56.275 -36.555 56.605 ;
        RECT -36.885 54.915 -36.555 55.245 ;
        RECT -36.885 53.555 -36.555 53.885 ;
        RECT -36.885 52.195 -36.555 52.525 ;
        RECT -36.885 50.835 -36.555 51.165 ;
        RECT -36.885 49.475 -36.555 49.805 ;
        RECT -36.885 48.115 -36.555 48.445 ;
        RECT -36.885 46.755 -36.555 47.085 ;
        RECT -36.885 45.395 -36.555 45.725 ;
        RECT -36.885 44.035 -36.555 44.365 ;
        RECT -36.885 42.675 -36.555 43.005 ;
        RECT -36.885 41.315 -36.555 41.645 ;
        RECT -36.885 39.955 -36.555 40.285 ;
        RECT -36.885 38.595 -36.555 38.925 ;
        RECT -36.885 37.235 -36.555 37.565 ;
        RECT -36.885 35.875 -36.555 36.205 ;
        RECT -36.885 34.515 -36.555 34.845 ;
        RECT -36.885 33.155 -36.555 33.485 ;
        RECT -36.885 31.795 -36.555 32.125 ;
        RECT -36.885 30.435 -36.555 30.765 ;
        RECT -36.885 29.075 -36.555 29.405 ;
        RECT -36.885 27.715 -36.555 28.045 ;
        RECT -36.885 26.355 -36.555 26.685 ;
        RECT -36.885 24.995 -36.555 25.325 ;
        RECT -36.885 23.635 -36.555 23.965 ;
        RECT -36.885 22.275 -36.555 22.605 ;
        RECT -36.885 20.915 -36.555 21.245 ;
        RECT -36.885 19.555 -36.555 19.885 ;
        RECT -36.885 18.195 -36.555 18.525 ;
        RECT -36.885 16.835 -36.555 17.165 ;
        RECT -36.885 15.475 -36.555 15.805 ;
        RECT -36.885 14.115 -36.555 14.445 ;
        RECT -36.885 12.755 -36.555 13.085 ;
        RECT -36.885 11.395 -36.555 11.725 ;
        RECT -36.885 10.035 -36.555 10.365 ;
        RECT -36.885 8.675 -36.555 9.005 ;
        RECT -36.885 7.315 -36.555 7.645 ;
        RECT -36.885 5.955 -36.555 6.285 ;
        RECT -36.885 4.595 -36.555 4.925 ;
        RECT -36.885 3.235 -36.555 3.565 ;
        RECT -36.885 1.875 -36.555 2.205 ;
        RECT -36.885 0.515 -36.555 0.845 ;
        RECT -36.885 -0.845 -36.555 -0.515 ;
        RECT -36.885 -2.205 -36.555 -1.875 ;
        RECT -36.885 -7.645 -36.555 -7.315 ;
        RECT -36.885 -10.365 -36.555 -10.035 ;
        RECT -36.885 -14.445 -36.555 -14.115 ;
        RECT -36.885 -17.165 -36.555 -16.835 ;
        RECT -36.885 -18.525 -36.555 -18.195 ;
        RECT -36.885 -19.885 -36.555 -19.555 ;
        RECT -36.885 -21.245 -36.555 -20.915 ;
        RECT -36.885 -22.605 -36.555 -22.275 ;
        RECT -36.885 -23.965 -36.555 -23.635 ;
        RECT -36.885 -25.325 -36.555 -24.995 ;
        RECT -36.885 -32.125 -36.555 -31.795 ;
        RECT -36.885 -33.71 -36.555 -33.38 ;
        RECT -36.885 -34.845 -36.555 -34.515 ;
        RECT -36.885 -36.205 -36.555 -35.875 ;
        RECT -36.885 -38.925 -36.555 -38.595 ;
        RECT -36.885 -39.75 -36.555 -39.42 ;
        RECT -36.885 -41.645 -36.555 -41.315 ;
        RECT -36.885 -44.365 -36.555 -44.035 ;
        RECT -36.885 -49.805 -36.555 -49.475 ;
        RECT -36.885 -51.165 -36.555 -50.835 ;
        RECT -36.885 -52.525 -36.555 -52.195 ;
        RECT -36.885 -53.885 -36.555 -53.555 ;
        RECT -36.885 -55.245 -36.555 -54.915 ;
        RECT -36.885 -56.605 -36.555 -56.275 ;
        RECT -36.885 -57.965 -36.555 -57.635 ;
        RECT -36.885 -59.325 -36.555 -58.995 ;
        RECT -36.885 -60.685 -36.555 -60.355 ;
        RECT -36.885 -62.045 -36.555 -61.715 ;
        RECT -36.885 -63.405 -36.555 -63.075 ;
        RECT -36.885 -64.765 -36.555 -64.435 ;
        RECT -36.885 -66.125 -36.555 -65.795 ;
        RECT -36.885 -70.205 -36.555 -69.875 ;
        RECT -36.885 -71.565 -36.555 -71.235 ;
        RECT -36.885 -72.925 -36.555 -72.595 ;
        RECT -36.885 -74.285 -36.555 -73.955 ;
        RECT -36.885 -75.645 -36.555 -75.315 ;
        RECT -36.885 -77.005 -36.555 -76.675 ;
        RECT -36.885 -78.365 -36.555 -78.035 ;
        RECT -36.885 -79.725 -36.555 -79.395 ;
        RECT -36.885 -81.085 -36.555 -80.755 ;
        RECT -36.885 -82.445 -36.555 -82.115 ;
        RECT -36.885 -83.805 -36.555 -83.475 ;
        RECT -36.885 -85.165 -36.555 -84.835 ;
        RECT -36.885 -86.525 -36.555 -86.195 ;
        RECT -36.885 -87.885 -36.555 -87.555 ;
        RECT -36.885 -89.245 -36.555 -88.915 ;
        RECT -36.885 -90.605 -36.555 -90.275 ;
        RECT -36.885 -91.77 -36.555 -91.44 ;
        RECT -36.885 -93.325 -36.555 -92.995 ;
        RECT -36.885 -94.685 -36.555 -94.355 ;
        RECT -36.885 -96.045 -36.555 -95.715 ;
        RECT -36.885 -97.405 -36.555 -97.075 ;
        RECT -36.885 -98.765 -36.555 -98.435 ;
        RECT -36.885 -101.485 -36.555 -101.155 ;
        RECT -36.885 -102.31 -36.555 -101.98 ;
        RECT -36.885 -104.205 -36.555 -103.875 ;
        RECT -36.885 -105.565 -36.555 -105.235 ;
        RECT -36.885 -106.925 -36.555 -106.595 ;
        RECT -36.885 -109.645 -36.555 -109.315 ;
        RECT -36.885 -111.005 -36.555 -110.675 ;
        RECT -36.885 -113.725 -36.555 -113.395 ;
        RECT -36.885 -115.085 -36.555 -114.755 ;
        RECT -36.885 -116.445 -36.555 -116.115 ;
        RECT -36.885 -117.805 -36.555 -117.475 ;
        RECT -36.885 -119.165 -36.555 -118.835 ;
        RECT -36.885 -120.525 -36.555 -120.195 ;
        RECT -36.885 -123.245 -36.555 -122.915 ;
        RECT -36.885 -124.605 -36.555 -124.275 ;
        RECT -36.885 -125.965 -36.555 -125.635 ;
        RECT -36.885 -127.325 -36.555 -126.995 ;
        RECT -36.885 -128.685 -36.555 -128.355 ;
        RECT -36.885 -130.045 -36.555 -129.715 ;
        RECT -36.885 -134.125 -36.555 -133.795 ;
        RECT -36.885 -135.485 -36.555 -135.155 ;
        RECT -36.885 -136.845 -36.555 -136.515 ;
        RECT -36.885 -138.205 -36.555 -137.875 ;
        RECT -36.885 -139.565 -36.555 -139.235 ;
        RECT -36.885 -140.925 -36.555 -140.595 ;
        RECT -36.885 -142.285 -36.555 -141.955 ;
        RECT -36.885 -143.645 -36.555 -143.315 ;
        RECT -36.885 -145.005 -36.555 -144.675 ;
        RECT -36.885 -146.365 -36.555 -146.035 ;
        RECT -36.885 -147.725 -36.555 -147.395 ;
        RECT -36.885 -149.085 -36.555 -148.755 ;
        RECT -36.885 -151.805 -36.555 -151.475 ;
        RECT -36.885 -153.165 -36.555 -152.835 ;
        RECT -36.885 -157.245 -36.555 -156.915 ;
        RECT -36.885 -158.605 -36.555 -158.275 ;
        RECT -36.885 -159.965 -36.555 -159.635 ;
        RECT -36.885 -161.325 -36.555 -160.995 ;
        RECT -36.885 -162.685 -36.555 -162.355 ;
        RECT -36.885 -164.045 -36.555 -163.715 ;
        RECT -36.885 -165.405 -36.555 -165.075 ;
        RECT -36.885 -166.765 -36.555 -166.435 ;
        RECT -36.885 -169.615 -36.555 -169.285 ;
        RECT -36.885 -170.845 -36.555 -170.515 ;
        RECT -36.885 -172.205 -36.555 -171.875 ;
        RECT -36.885 -173.565 -36.555 -173.235 ;
        RECT -36.885 -174.925 -36.555 -174.595 ;
        RECT -36.885 -177.645 -36.555 -177.315 ;
        RECT -36.885 -179.005 -36.555 -178.675 ;
        RECT -36.885 -184.65 -36.555 -183.52 ;
        RECT -36.88 -184.765 -36.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.525 244.04 -35.195 245.17 ;
        RECT -35.525 239.875 -35.195 240.205 ;
        RECT -35.525 238.515 -35.195 238.845 ;
        RECT -35.525 237.155 -35.195 237.485 ;
        RECT -35.525 235.795 -35.195 236.125 ;
        RECT -35.525 234.435 -35.195 234.765 ;
        RECT -35.525 233.075 -35.195 233.405 ;
        RECT -35.525 231.715 -35.195 232.045 ;
        RECT -35.525 230.355 -35.195 230.685 ;
        RECT -35.525 228.995 -35.195 229.325 ;
        RECT -35.525 227.635 -35.195 227.965 ;
        RECT -35.525 226.275 -35.195 226.605 ;
        RECT -35.525 224.915 -35.195 225.245 ;
        RECT -35.525 223.555 -35.195 223.885 ;
        RECT -35.525 222.195 -35.195 222.525 ;
        RECT -35.525 220.835 -35.195 221.165 ;
        RECT -35.525 219.475 -35.195 219.805 ;
        RECT -35.525 218.115 -35.195 218.445 ;
        RECT -35.525 216.755 -35.195 217.085 ;
        RECT -35.525 215.395 -35.195 215.725 ;
        RECT -35.525 214.035 -35.195 214.365 ;
        RECT -35.525 212.675 -35.195 213.005 ;
        RECT -35.525 211.315 -35.195 211.645 ;
        RECT -35.525 209.955 -35.195 210.285 ;
        RECT -35.525 208.595 -35.195 208.925 ;
        RECT -35.525 207.235 -35.195 207.565 ;
        RECT -35.525 205.875 -35.195 206.205 ;
        RECT -35.525 204.515 -35.195 204.845 ;
        RECT -35.525 203.155 -35.195 203.485 ;
        RECT -35.525 201.795 -35.195 202.125 ;
        RECT -35.525 200.435 -35.195 200.765 ;
        RECT -35.525 199.075 -35.195 199.405 ;
        RECT -35.525 197.715 -35.195 198.045 ;
        RECT -35.525 196.355 -35.195 196.685 ;
        RECT -35.525 194.995 -35.195 195.325 ;
        RECT -35.525 193.635 -35.195 193.965 ;
        RECT -35.525 192.275 -35.195 192.605 ;
        RECT -35.525 190.915 -35.195 191.245 ;
        RECT -35.525 189.555 -35.195 189.885 ;
        RECT -35.525 188.195 -35.195 188.525 ;
        RECT -35.525 186.835 -35.195 187.165 ;
        RECT -35.525 185.475 -35.195 185.805 ;
        RECT -35.525 184.115 -35.195 184.445 ;
        RECT -35.525 182.755 -35.195 183.085 ;
        RECT -35.525 181.395 -35.195 181.725 ;
        RECT -35.525 180.035 -35.195 180.365 ;
        RECT -35.525 178.675 -35.195 179.005 ;
        RECT -35.525 177.315 -35.195 177.645 ;
        RECT -35.525 175.955 -35.195 176.285 ;
        RECT -35.525 174.595 -35.195 174.925 ;
        RECT -35.525 173.235 -35.195 173.565 ;
        RECT -35.525 171.875 -35.195 172.205 ;
        RECT -35.525 170.515 -35.195 170.845 ;
        RECT -35.525 169.155 -35.195 169.485 ;
        RECT -35.525 167.795 -35.195 168.125 ;
        RECT -35.525 166.435 -35.195 166.765 ;
        RECT -35.525 165.075 -35.195 165.405 ;
        RECT -35.525 163.715 -35.195 164.045 ;
        RECT -35.525 162.355 -35.195 162.685 ;
        RECT -35.525 160.995 -35.195 161.325 ;
        RECT -35.525 159.635 -35.195 159.965 ;
        RECT -35.525 158.275 -35.195 158.605 ;
        RECT -35.525 156.915 -35.195 157.245 ;
        RECT -35.525 155.555 -35.195 155.885 ;
        RECT -35.525 154.195 -35.195 154.525 ;
        RECT -35.525 152.835 -35.195 153.165 ;
        RECT -35.525 151.475 -35.195 151.805 ;
        RECT -35.525 150.115 -35.195 150.445 ;
        RECT -35.525 148.755 -35.195 149.085 ;
        RECT -35.525 147.395 -35.195 147.725 ;
        RECT -35.525 146.035 -35.195 146.365 ;
        RECT -35.525 144.675 -35.195 145.005 ;
        RECT -35.525 143.315 -35.195 143.645 ;
        RECT -35.525 141.955 -35.195 142.285 ;
        RECT -35.525 140.595 -35.195 140.925 ;
        RECT -35.525 139.235 -35.195 139.565 ;
        RECT -35.525 137.875 -35.195 138.205 ;
        RECT -35.525 136.515 -35.195 136.845 ;
        RECT -35.525 135.155 -35.195 135.485 ;
        RECT -35.525 133.795 -35.195 134.125 ;
        RECT -35.525 132.435 -35.195 132.765 ;
        RECT -35.525 131.075 -35.195 131.405 ;
        RECT -35.525 129.715 -35.195 130.045 ;
        RECT -35.525 128.355 -35.195 128.685 ;
        RECT -35.525 126.995 -35.195 127.325 ;
        RECT -35.525 125.635 -35.195 125.965 ;
        RECT -35.525 124.275 -35.195 124.605 ;
        RECT -35.525 122.915 -35.195 123.245 ;
        RECT -35.525 121.555 -35.195 121.885 ;
        RECT -35.525 120.195 -35.195 120.525 ;
        RECT -35.525 118.835 -35.195 119.165 ;
        RECT -35.525 117.475 -35.195 117.805 ;
        RECT -35.525 116.115 -35.195 116.445 ;
        RECT -35.525 114.755 -35.195 115.085 ;
        RECT -35.525 113.395 -35.195 113.725 ;
        RECT -35.525 112.035 -35.195 112.365 ;
        RECT -35.525 110.675 -35.195 111.005 ;
        RECT -35.525 109.315 -35.195 109.645 ;
        RECT -35.525 107.955 -35.195 108.285 ;
        RECT -35.525 106.595 -35.195 106.925 ;
        RECT -35.525 105.235 -35.195 105.565 ;
        RECT -35.525 103.875 -35.195 104.205 ;
        RECT -35.525 102.515 -35.195 102.845 ;
        RECT -35.525 101.155 -35.195 101.485 ;
        RECT -35.525 99.795 -35.195 100.125 ;
        RECT -35.525 98.435 -35.195 98.765 ;
        RECT -35.525 97.075 -35.195 97.405 ;
        RECT -35.525 95.715 -35.195 96.045 ;
        RECT -35.525 94.355 -35.195 94.685 ;
        RECT -35.525 92.995 -35.195 93.325 ;
        RECT -35.525 91.635 -35.195 91.965 ;
        RECT -35.525 90.275 -35.195 90.605 ;
        RECT -35.525 88.915 -35.195 89.245 ;
        RECT -35.525 87.555 -35.195 87.885 ;
        RECT -35.525 86.195 -35.195 86.525 ;
        RECT -35.525 84.835 -35.195 85.165 ;
        RECT -35.525 83.475 -35.195 83.805 ;
        RECT -35.525 82.115 -35.195 82.445 ;
        RECT -35.525 80.755 -35.195 81.085 ;
        RECT -35.525 79.395 -35.195 79.725 ;
        RECT -35.525 78.035 -35.195 78.365 ;
        RECT -35.525 76.675 -35.195 77.005 ;
        RECT -35.525 75.315 -35.195 75.645 ;
        RECT -35.525 73.955 -35.195 74.285 ;
        RECT -35.525 72.595 -35.195 72.925 ;
        RECT -35.525 71.235 -35.195 71.565 ;
        RECT -35.525 69.875 -35.195 70.205 ;
        RECT -35.525 68.515 -35.195 68.845 ;
        RECT -35.525 67.155 -35.195 67.485 ;
        RECT -35.525 65.795 -35.195 66.125 ;
        RECT -35.525 64.435 -35.195 64.765 ;
        RECT -35.525 63.075 -35.195 63.405 ;
        RECT -35.525 61.715 -35.195 62.045 ;
        RECT -35.525 60.355 -35.195 60.685 ;
        RECT -35.525 58.995 -35.195 59.325 ;
        RECT -35.525 57.635 -35.195 57.965 ;
        RECT -35.525 56.275 -35.195 56.605 ;
        RECT -35.525 54.915 -35.195 55.245 ;
        RECT -35.525 53.555 -35.195 53.885 ;
        RECT -35.525 52.195 -35.195 52.525 ;
        RECT -35.525 50.835 -35.195 51.165 ;
        RECT -35.525 49.475 -35.195 49.805 ;
        RECT -35.525 48.115 -35.195 48.445 ;
        RECT -35.525 46.755 -35.195 47.085 ;
        RECT -35.525 45.395 -35.195 45.725 ;
        RECT -35.525 44.035 -35.195 44.365 ;
        RECT -35.525 42.675 -35.195 43.005 ;
        RECT -35.525 41.315 -35.195 41.645 ;
        RECT -35.525 39.955 -35.195 40.285 ;
        RECT -35.525 38.595 -35.195 38.925 ;
        RECT -35.525 37.235 -35.195 37.565 ;
        RECT -35.525 35.875 -35.195 36.205 ;
        RECT -35.525 34.515 -35.195 34.845 ;
        RECT -35.525 33.155 -35.195 33.485 ;
        RECT -35.525 31.795 -35.195 32.125 ;
        RECT -35.525 30.435 -35.195 30.765 ;
        RECT -35.525 29.075 -35.195 29.405 ;
        RECT -35.525 27.715 -35.195 28.045 ;
        RECT -35.525 26.355 -35.195 26.685 ;
        RECT -35.525 24.995 -35.195 25.325 ;
        RECT -35.525 23.635 -35.195 23.965 ;
        RECT -35.525 22.275 -35.195 22.605 ;
        RECT -35.525 20.915 -35.195 21.245 ;
        RECT -35.525 19.555 -35.195 19.885 ;
        RECT -35.525 18.195 -35.195 18.525 ;
        RECT -35.525 16.835 -35.195 17.165 ;
        RECT -35.525 15.475 -35.195 15.805 ;
        RECT -35.525 14.115 -35.195 14.445 ;
        RECT -35.525 12.755 -35.195 13.085 ;
        RECT -35.525 11.395 -35.195 11.725 ;
        RECT -35.525 10.035 -35.195 10.365 ;
        RECT -35.525 8.675 -35.195 9.005 ;
        RECT -35.525 7.315 -35.195 7.645 ;
        RECT -35.525 5.955 -35.195 6.285 ;
        RECT -35.525 4.595 -35.195 4.925 ;
        RECT -35.525 3.235 -35.195 3.565 ;
        RECT -35.525 1.875 -35.195 2.205 ;
        RECT -35.525 0.515 -35.195 0.845 ;
        RECT -35.525 -0.845 -35.195 -0.515 ;
        RECT -35.525 -7.645 -35.195 -7.315 ;
        RECT -35.525 -10.365 -35.195 -10.035 ;
        RECT -35.525 -14.445 -35.195 -14.115 ;
        RECT -35.525 -17.165 -35.195 -16.835 ;
        RECT -35.525 -18.525 -35.195 -18.195 ;
        RECT -35.525 -19.885 -35.195 -19.555 ;
        RECT -35.525 -21.245 -35.195 -20.915 ;
        RECT -35.525 -22.605 -35.195 -22.275 ;
        RECT -35.525 -23.965 -35.195 -23.635 ;
        RECT -35.525 -25.325 -35.195 -24.995 ;
        RECT -35.525 -32.125 -35.195 -31.795 ;
        RECT -35.525 -33.71 -35.195 -33.38 ;
        RECT -35.525 -34.845 -35.195 -34.515 ;
        RECT -35.525 -36.205 -35.195 -35.875 ;
        RECT -35.525 -38.925 -35.195 -38.595 ;
        RECT -35.525 -39.75 -35.195 -39.42 ;
        RECT -35.525 -41.645 -35.195 -41.315 ;
        RECT -35.525 -44.365 -35.195 -44.035 ;
        RECT -35.525 -49.805 -35.195 -49.475 ;
        RECT -35.525 -51.165 -35.195 -50.835 ;
        RECT -35.525 -52.525 -35.195 -52.195 ;
        RECT -35.525 -53.885 -35.195 -53.555 ;
        RECT -35.525 -55.245 -35.195 -54.915 ;
        RECT -35.525 -56.605 -35.195 -56.275 ;
        RECT -35.525 -57.965 -35.195 -57.635 ;
        RECT -35.525 -59.325 -35.195 -58.995 ;
        RECT -35.525 -60.685 -35.195 -60.355 ;
        RECT -35.525 -62.045 -35.195 -61.715 ;
        RECT -35.525 -63.405 -35.195 -63.075 ;
        RECT -35.525 -64.765 -35.195 -64.435 ;
        RECT -35.525 -66.125 -35.195 -65.795 ;
        RECT -35.525 -70.205 -35.195 -69.875 ;
        RECT -35.525 -71.565 -35.195 -71.235 ;
        RECT -35.525 -72.925 -35.195 -72.595 ;
        RECT -35.525 -74.285 -35.195 -73.955 ;
        RECT -35.525 -75.645 -35.195 -75.315 ;
        RECT -35.525 -77.005 -35.195 -76.675 ;
        RECT -35.525 -78.365 -35.195 -78.035 ;
        RECT -35.525 -79.725 -35.195 -79.395 ;
        RECT -35.525 -81.085 -35.195 -80.755 ;
        RECT -35.525 -82.445 -35.195 -82.115 ;
        RECT -35.525 -83.805 -35.195 -83.475 ;
        RECT -35.525 -85.165 -35.195 -84.835 ;
        RECT -35.525 -86.525 -35.195 -86.195 ;
        RECT -35.525 -87.885 -35.195 -87.555 ;
        RECT -35.525 -89.245 -35.195 -88.915 ;
        RECT -35.525 -90.605 -35.195 -90.275 ;
        RECT -35.525 -91.965 -35.195 -91.635 ;
        RECT -35.525 -93.325 -35.195 -92.995 ;
        RECT -35.525 -94.685 -35.195 -94.355 ;
        RECT -35.525 -96.045 -35.195 -95.715 ;
        RECT -35.525 -97.405 -35.195 -97.075 ;
        RECT -35.525 -98.765 -35.195 -98.435 ;
        RECT -35.525 -100.125 -35.195 -99.795 ;
        RECT -35.525 -101.485 -35.195 -101.155 ;
        RECT -35.525 -102.845 -35.195 -102.515 ;
        RECT -35.525 -104.205 -35.195 -103.875 ;
        RECT -35.525 -105.565 -35.195 -105.235 ;
        RECT -35.525 -106.925 -35.195 -106.595 ;
        RECT -35.525 -108.285 -35.195 -107.955 ;
        RECT -35.525 -109.645 -35.195 -109.315 ;
        RECT -35.525 -111.005 -35.195 -110.675 ;
        RECT -35.525 -112.365 -35.195 -112.035 ;
        RECT -35.525 -113.725 -35.195 -113.395 ;
        RECT -35.52 -113.725 -35.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -35.525 -177.645 -35.195 -177.315 ;
        RECT -35.525 -179.005 -35.195 -178.675 ;
        RECT -35.525 -184.65 -35.195 -183.52 ;
        RECT -35.52 -184.765 -35.2 -175.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.165 244.04 -33.835 245.17 ;
        RECT -34.165 239.875 -33.835 240.205 ;
        RECT -34.165 238.515 -33.835 238.845 ;
        RECT -34.165 237.155 -33.835 237.485 ;
        RECT -34.165 235.795 -33.835 236.125 ;
        RECT -34.165 234.435 -33.835 234.765 ;
        RECT -34.165 233.075 -33.835 233.405 ;
        RECT -34.165 231.715 -33.835 232.045 ;
        RECT -34.165 230.355 -33.835 230.685 ;
        RECT -34.165 228.995 -33.835 229.325 ;
        RECT -34.165 227.635 -33.835 227.965 ;
        RECT -34.165 226.275 -33.835 226.605 ;
        RECT -34.165 224.915 -33.835 225.245 ;
        RECT -34.165 223.555 -33.835 223.885 ;
        RECT -34.165 222.195 -33.835 222.525 ;
        RECT -34.165 220.835 -33.835 221.165 ;
        RECT -34.165 219.475 -33.835 219.805 ;
        RECT -34.165 218.115 -33.835 218.445 ;
        RECT -34.165 216.755 -33.835 217.085 ;
        RECT -34.165 215.395 -33.835 215.725 ;
        RECT -34.165 214.035 -33.835 214.365 ;
        RECT -34.165 212.675 -33.835 213.005 ;
        RECT -34.165 211.315 -33.835 211.645 ;
        RECT -34.165 209.955 -33.835 210.285 ;
        RECT -34.165 208.595 -33.835 208.925 ;
        RECT -34.165 207.235 -33.835 207.565 ;
        RECT -34.165 205.875 -33.835 206.205 ;
        RECT -34.165 204.515 -33.835 204.845 ;
        RECT -34.165 203.155 -33.835 203.485 ;
        RECT -34.165 201.795 -33.835 202.125 ;
        RECT -34.165 200.435 -33.835 200.765 ;
        RECT -34.165 199.075 -33.835 199.405 ;
        RECT -34.165 197.715 -33.835 198.045 ;
        RECT -34.165 196.355 -33.835 196.685 ;
        RECT -34.165 194.995 -33.835 195.325 ;
        RECT -34.165 193.635 -33.835 193.965 ;
        RECT -34.165 192.275 -33.835 192.605 ;
        RECT -34.165 190.915 -33.835 191.245 ;
        RECT -34.165 189.555 -33.835 189.885 ;
        RECT -34.165 188.195 -33.835 188.525 ;
        RECT -34.165 186.835 -33.835 187.165 ;
        RECT -34.165 185.475 -33.835 185.805 ;
        RECT -34.165 184.115 -33.835 184.445 ;
        RECT -34.165 182.755 -33.835 183.085 ;
        RECT -34.165 181.395 -33.835 181.725 ;
        RECT -34.165 180.035 -33.835 180.365 ;
        RECT -34.165 178.675 -33.835 179.005 ;
        RECT -34.165 177.315 -33.835 177.645 ;
        RECT -34.165 175.955 -33.835 176.285 ;
        RECT -34.165 174.595 -33.835 174.925 ;
        RECT -34.165 173.235 -33.835 173.565 ;
        RECT -34.165 171.875 -33.835 172.205 ;
        RECT -34.165 170.515 -33.835 170.845 ;
        RECT -34.165 169.155 -33.835 169.485 ;
        RECT -34.165 167.795 -33.835 168.125 ;
        RECT -34.165 166.435 -33.835 166.765 ;
        RECT -34.165 165.075 -33.835 165.405 ;
        RECT -34.165 163.715 -33.835 164.045 ;
        RECT -34.165 162.355 -33.835 162.685 ;
        RECT -34.165 160.995 -33.835 161.325 ;
        RECT -34.165 159.635 -33.835 159.965 ;
        RECT -34.165 158.275 -33.835 158.605 ;
        RECT -34.165 156.915 -33.835 157.245 ;
        RECT -34.165 155.555 -33.835 155.885 ;
        RECT -34.165 154.195 -33.835 154.525 ;
        RECT -34.165 152.835 -33.835 153.165 ;
        RECT -34.165 151.475 -33.835 151.805 ;
        RECT -34.165 150.115 -33.835 150.445 ;
        RECT -34.165 148.755 -33.835 149.085 ;
        RECT -34.165 147.395 -33.835 147.725 ;
        RECT -34.165 146.035 -33.835 146.365 ;
        RECT -34.165 144.675 -33.835 145.005 ;
        RECT -34.165 143.315 -33.835 143.645 ;
        RECT -34.165 141.955 -33.835 142.285 ;
        RECT -34.165 140.595 -33.835 140.925 ;
        RECT -34.165 139.235 -33.835 139.565 ;
        RECT -34.165 137.875 -33.835 138.205 ;
        RECT -34.165 136.515 -33.835 136.845 ;
        RECT -34.165 135.155 -33.835 135.485 ;
        RECT -34.165 133.795 -33.835 134.125 ;
        RECT -34.165 132.435 -33.835 132.765 ;
        RECT -34.165 131.075 -33.835 131.405 ;
        RECT -34.165 129.715 -33.835 130.045 ;
        RECT -34.165 128.355 -33.835 128.685 ;
        RECT -34.165 126.995 -33.835 127.325 ;
        RECT -34.165 125.635 -33.835 125.965 ;
        RECT -34.165 124.275 -33.835 124.605 ;
        RECT -34.165 122.915 -33.835 123.245 ;
        RECT -34.165 121.555 -33.835 121.885 ;
        RECT -34.165 120.195 -33.835 120.525 ;
        RECT -34.165 118.835 -33.835 119.165 ;
        RECT -34.165 117.475 -33.835 117.805 ;
        RECT -34.165 116.115 -33.835 116.445 ;
        RECT -34.165 114.755 -33.835 115.085 ;
        RECT -34.165 113.395 -33.835 113.725 ;
        RECT -34.165 112.035 -33.835 112.365 ;
        RECT -34.165 110.675 -33.835 111.005 ;
        RECT -34.165 109.315 -33.835 109.645 ;
        RECT -34.165 107.955 -33.835 108.285 ;
        RECT -34.165 106.595 -33.835 106.925 ;
        RECT -34.165 105.235 -33.835 105.565 ;
        RECT -34.165 103.875 -33.835 104.205 ;
        RECT -34.165 102.515 -33.835 102.845 ;
        RECT -34.165 101.155 -33.835 101.485 ;
        RECT -34.165 99.795 -33.835 100.125 ;
        RECT -34.165 98.435 -33.835 98.765 ;
        RECT -34.165 97.075 -33.835 97.405 ;
        RECT -34.165 95.715 -33.835 96.045 ;
        RECT -34.165 94.355 -33.835 94.685 ;
        RECT -34.165 92.995 -33.835 93.325 ;
        RECT -34.165 91.635 -33.835 91.965 ;
        RECT -34.165 90.275 -33.835 90.605 ;
        RECT -34.165 88.915 -33.835 89.245 ;
        RECT -34.165 87.555 -33.835 87.885 ;
        RECT -34.165 86.195 -33.835 86.525 ;
        RECT -34.165 84.835 -33.835 85.165 ;
        RECT -34.165 83.475 -33.835 83.805 ;
        RECT -34.165 82.115 -33.835 82.445 ;
        RECT -34.165 80.755 -33.835 81.085 ;
        RECT -34.165 79.395 -33.835 79.725 ;
        RECT -34.165 78.035 -33.835 78.365 ;
        RECT -34.165 76.675 -33.835 77.005 ;
        RECT -34.165 75.315 -33.835 75.645 ;
        RECT -34.165 73.955 -33.835 74.285 ;
        RECT -34.165 72.595 -33.835 72.925 ;
        RECT -34.165 71.235 -33.835 71.565 ;
        RECT -34.165 69.875 -33.835 70.205 ;
        RECT -34.165 68.515 -33.835 68.845 ;
        RECT -34.165 67.155 -33.835 67.485 ;
        RECT -34.165 65.795 -33.835 66.125 ;
        RECT -34.165 64.435 -33.835 64.765 ;
        RECT -34.165 63.075 -33.835 63.405 ;
        RECT -34.165 61.715 -33.835 62.045 ;
        RECT -34.165 60.355 -33.835 60.685 ;
        RECT -34.165 58.995 -33.835 59.325 ;
        RECT -34.165 57.635 -33.835 57.965 ;
        RECT -34.165 56.275 -33.835 56.605 ;
        RECT -34.165 54.915 -33.835 55.245 ;
        RECT -34.165 53.555 -33.835 53.885 ;
        RECT -34.165 52.195 -33.835 52.525 ;
        RECT -34.165 50.835 -33.835 51.165 ;
        RECT -34.165 49.475 -33.835 49.805 ;
        RECT -34.165 48.115 -33.835 48.445 ;
        RECT -34.165 46.755 -33.835 47.085 ;
        RECT -34.165 45.395 -33.835 45.725 ;
        RECT -34.165 44.035 -33.835 44.365 ;
        RECT -34.165 42.675 -33.835 43.005 ;
        RECT -34.165 41.315 -33.835 41.645 ;
        RECT -34.165 39.955 -33.835 40.285 ;
        RECT -34.165 38.595 -33.835 38.925 ;
        RECT -34.165 37.235 -33.835 37.565 ;
        RECT -34.165 35.875 -33.835 36.205 ;
        RECT -34.165 34.515 -33.835 34.845 ;
        RECT -34.165 33.155 -33.835 33.485 ;
        RECT -34.165 31.795 -33.835 32.125 ;
        RECT -34.165 30.435 -33.835 30.765 ;
        RECT -34.165 29.075 -33.835 29.405 ;
        RECT -34.165 27.715 -33.835 28.045 ;
        RECT -34.165 26.355 -33.835 26.685 ;
        RECT -34.165 24.995 -33.835 25.325 ;
        RECT -34.165 23.635 -33.835 23.965 ;
        RECT -34.165 22.275 -33.835 22.605 ;
        RECT -34.165 20.915 -33.835 21.245 ;
        RECT -34.165 19.555 -33.835 19.885 ;
        RECT -34.165 18.195 -33.835 18.525 ;
        RECT -34.165 16.835 -33.835 17.165 ;
        RECT -34.165 15.475 -33.835 15.805 ;
        RECT -34.165 14.115 -33.835 14.445 ;
        RECT -34.165 12.755 -33.835 13.085 ;
        RECT -34.165 11.395 -33.835 11.725 ;
        RECT -34.165 10.035 -33.835 10.365 ;
        RECT -34.165 8.675 -33.835 9.005 ;
        RECT -34.165 7.315 -33.835 7.645 ;
        RECT -34.165 5.955 -33.835 6.285 ;
        RECT -34.165 4.595 -33.835 4.925 ;
        RECT -34.165 3.235 -33.835 3.565 ;
        RECT -34.165 1.875 -33.835 2.205 ;
        RECT -34.165 0.515 -33.835 0.845 ;
        RECT -34.165 -0.845 -33.835 -0.515 ;
        RECT -34.165 -7.645 -33.835 -7.315 ;
        RECT -34.165 -10.365 -33.835 -10.035 ;
        RECT -34.165 -14.445 -33.835 -14.115 ;
        RECT -34.165 -17.165 -33.835 -16.835 ;
        RECT -34.165 -18.525 -33.835 -18.195 ;
        RECT -34.165 -19.885 -33.835 -19.555 ;
        RECT -34.165 -21.245 -33.835 -20.915 ;
        RECT -34.165 -22.605 -33.835 -22.275 ;
        RECT -34.165 -23.965 -33.835 -23.635 ;
        RECT -34.165 -25.325 -33.835 -24.995 ;
        RECT -34.165 -32.125 -33.835 -31.795 ;
        RECT -34.165 -33.71 -33.835 -33.38 ;
        RECT -34.165 -34.845 -33.835 -34.515 ;
        RECT -34.165 -36.205 -33.835 -35.875 ;
        RECT -34.165 -38.925 -33.835 -38.595 ;
        RECT -34.165 -39.75 -33.835 -39.42 ;
        RECT -34.165 -41.645 -33.835 -41.315 ;
        RECT -34.165 -44.365 -33.835 -44.035 ;
        RECT -34.165 -49.805 -33.835 -49.475 ;
        RECT -34.165 -51.165 -33.835 -50.835 ;
        RECT -34.165 -53.885 -33.835 -53.555 ;
        RECT -34.165 -55.245 -33.835 -54.915 ;
        RECT -34.165 -59.325 -33.835 -58.995 ;
        RECT -34.165 -60.685 -33.835 -60.355 ;
        RECT -34.165 -63.405 -33.835 -63.075 ;
        RECT -34.165 -70.205 -33.835 -69.875 ;
        RECT -34.165 -71.565 -33.835 -71.235 ;
        RECT -34.165 -72.925 -33.835 -72.595 ;
        RECT -34.165 -74.285 -33.835 -73.955 ;
        RECT -34.165 -75.645 -33.835 -75.315 ;
        RECT -34.165 -77.005 -33.835 -76.675 ;
        RECT -34.165 -78.365 -33.835 -78.035 ;
        RECT -34.165 -79.725 -33.835 -79.395 ;
        RECT -34.165 -81.085 -33.835 -80.755 ;
        RECT -34.165 -82.445 -33.835 -82.115 ;
        RECT -34.165 -83.805 -33.835 -83.475 ;
        RECT -34.165 -85.165 -33.835 -84.835 ;
        RECT -34.165 -86.525 -33.835 -86.195 ;
        RECT -34.165 -87.885 -33.835 -87.555 ;
        RECT -34.165 -89.245 -33.835 -88.915 ;
        RECT -34.165 -90.605 -33.835 -90.275 ;
        RECT -34.165 -91.965 -33.835 -91.635 ;
        RECT -34.165 -93.325 -33.835 -92.995 ;
        RECT -34.165 -94.685 -33.835 -94.355 ;
        RECT -34.165 -96.045 -33.835 -95.715 ;
        RECT -34.165 -97.405 -33.835 -97.075 ;
        RECT -34.165 -98.765 -33.835 -98.435 ;
        RECT -34.165 -100.125 -33.835 -99.795 ;
        RECT -34.165 -101.485 -33.835 -101.155 ;
        RECT -34.165 -102.845 -33.835 -102.515 ;
        RECT -34.165 -104.205 -33.835 -103.875 ;
        RECT -34.165 -105.565 -33.835 -105.235 ;
        RECT -34.165 -106.925 -33.835 -106.595 ;
        RECT -34.165 -108.285 -33.835 -107.955 ;
        RECT -34.165 -109.645 -33.835 -109.315 ;
        RECT -34.165 -111.005 -33.835 -110.675 ;
        RECT -34.165 -112.365 -33.835 -112.035 ;
        RECT -34.165 -113.725 -33.835 -113.395 ;
        RECT -34.165 -115.085 -33.835 -114.755 ;
        RECT -34.165 -116.445 -33.835 -116.115 ;
        RECT -34.165 -117.805 -33.835 -117.475 ;
        RECT -34.165 -119.165 -33.835 -118.835 ;
        RECT -34.165 -120.525 -33.835 -120.195 ;
        RECT -34.165 -123.245 -33.835 -122.915 ;
        RECT -34.165 -125.965 -33.835 -125.635 ;
        RECT -34.165 -127.325 -33.835 -126.995 ;
        RECT -34.165 -128.685 -33.835 -128.355 ;
        RECT -34.165 -130.045 -33.835 -129.715 ;
        RECT -34.165 -134.125 -33.835 -133.795 ;
        RECT -34.165 -135.485 -33.835 -135.155 ;
        RECT -34.165 -136.845 -33.835 -136.515 ;
        RECT -34.165 -138.205 -33.835 -137.875 ;
        RECT -34.165 -139.565 -33.835 -139.235 ;
        RECT -34.165 -142.285 -33.835 -141.955 ;
        RECT -34.165 -143.645 -33.835 -143.315 ;
        RECT -34.165 -145.005 -33.835 -144.675 ;
        RECT -34.165 -146.365 -33.835 -146.035 ;
        RECT -34.165 -147.725 -33.835 -147.395 ;
        RECT -34.165 -149.085 -33.835 -148.755 ;
        RECT -34.165 -151.805 -33.835 -151.475 ;
        RECT -34.165 -153.165 -33.835 -152.835 ;
        RECT -34.165 -157.245 -33.835 -156.915 ;
        RECT -34.165 -158.605 -33.835 -158.275 ;
        RECT -34.165 -159.965 -33.835 -159.635 ;
        RECT -34.165 -161.325 -33.835 -160.995 ;
        RECT -34.165 -162.685 -33.835 -162.355 ;
        RECT -34.165 -164.045 -33.835 -163.715 ;
        RECT -34.165 -165.405 -33.835 -165.075 ;
        RECT -34.165 -166.765 -33.835 -166.435 ;
        RECT -34.165 -169.615 -33.835 -169.285 ;
        RECT -34.165 -170.845 -33.835 -170.515 ;
        RECT -34.165 -172.205 -33.835 -171.875 ;
        RECT -34.16 -172.88 -33.84 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.805 107.955 -32.475 108.285 ;
        RECT -32.805 106.595 -32.475 106.925 ;
        RECT -32.805 105.235 -32.475 105.565 ;
        RECT -32.805 103.875 -32.475 104.205 ;
        RECT -32.805 102.515 -32.475 102.845 ;
        RECT -32.805 101.155 -32.475 101.485 ;
        RECT -32.805 99.795 -32.475 100.125 ;
        RECT -32.805 98.435 -32.475 98.765 ;
        RECT -32.805 97.075 -32.475 97.405 ;
        RECT -32.805 95.715 -32.475 96.045 ;
        RECT -32.805 94.355 -32.475 94.685 ;
        RECT -32.805 92.995 -32.475 93.325 ;
        RECT -32.805 91.635 -32.475 91.965 ;
        RECT -32.805 90.275 -32.475 90.605 ;
        RECT -32.805 88.915 -32.475 89.245 ;
        RECT -32.805 87.555 -32.475 87.885 ;
        RECT -32.805 86.195 -32.475 86.525 ;
        RECT -32.805 84.835 -32.475 85.165 ;
        RECT -32.805 83.475 -32.475 83.805 ;
        RECT -32.805 82.115 -32.475 82.445 ;
        RECT -32.805 80.755 -32.475 81.085 ;
        RECT -32.805 79.395 -32.475 79.725 ;
        RECT -32.805 78.035 -32.475 78.365 ;
        RECT -32.805 76.675 -32.475 77.005 ;
        RECT -32.805 75.315 -32.475 75.645 ;
        RECT -32.805 73.955 -32.475 74.285 ;
        RECT -32.805 72.595 -32.475 72.925 ;
        RECT -32.805 71.235 -32.475 71.565 ;
        RECT -32.805 69.875 -32.475 70.205 ;
        RECT -32.805 68.515 -32.475 68.845 ;
        RECT -32.805 67.155 -32.475 67.485 ;
        RECT -32.805 65.795 -32.475 66.125 ;
        RECT -32.805 64.435 -32.475 64.765 ;
        RECT -32.805 63.075 -32.475 63.405 ;
        RECT -32.805 61.715 -32.475 62.045 ;
        RECT -32.805 60.355 -32.475 60.685 ;
        RECT -32.805 58.995 -32.475 59.325 ;
        RECT -32.805 57.635 -32.475 57.965 ;
        RECT -32.805 56.275 -32.475 56.605 ;
        RECT -32.805 54.915 -32.475 55.245 ;
        RECT -32.805 53.555 -32.475 53.885 ;
        RECT -32.805 52.195 -32.475 52.525 ;
        RECT -32.805 50.835 -32.475 51.165 ;
        RECT -32.805 49.475 -32.475 49.805 ;
        RECT -32.805 48.115 -32.475 48.445 ;
        RECT -32.805 46.755 -32.475 47.085 ;
        RECT -32.805 45.395 -32.475 45.725 ;
        RECT -32.805 44.035 -32.475 44.365 ;
        RECT -32.805 42.675 -32.475 43.005 ;
        RECT -32.805 41.315 -32.475 41.645 ;
        RECT -32.805 39.955 -32.475 40.285 ;
        RECT -32.805 38.595 -32.475 38.925 ;
        RECT -32.805 37.235 -32.475 37.565 ;
        RECT -32.805 35.875 -32.475 36.205 ;
        RECT -32.805 34.515 -32.475 34.845 ;
        RECT -32.805 33.155 -32.475 33.485 ;
        RECT -32.805 31.795 -32.475 32.125 ;
        RECT -32.805 30.435 -32.475 30.765 ;
        RECT -32.805 29.075 -32.475 29.405 ;
        RECT -32.805 27.715 -32.475 28.045 ;
        RECT -32.805 26.355 -32.475 26.685 ;
        RECT -32.805 24.995 -32.475 25.325 ;
        RECT -32.805 23.635 -32.475 23.965 ;
        RECT -32.805 22.275 -32.475 22.605 ;
        RECT -32.805 20.915 -32.475 21.245 ;
        RECT -32.805 19.555 -32.475 19.885 ;
        RECT -32.805 18.195 -32.475 18.525 ;
        RECT -32.805 16.835 -32.475 17.165 ;
        RECT -32.805 15.475 -32.475 15.805 ;
        RECT -32.805 14.115 -32.475 14.445 ;
        RECT -32.805 12.755 -32.475 13.085 ;
        RECT -32.805 11.395 -32.475 11.725 ;
        RECT -32.805 10.035 -32.475 10.365 ;
        RECT -32.805 8.675 -32.475 9.005 ;
        RECT -32.805 7.315 -32.475 7.645 ;
        RECT -32.805 5.955 -32.475 6.285 ;
        RECT -32.805 4.595 -32.475 4.925 ;
        RECT -32.805 3.235 -32.475 3.565 ;
        RECT -32.805 1.875 -32.475 2.205 ;
        RECT -32.805 0.515 -32.475 0.845 ;
        RECT -32.805 -0.845 -32.475 -0.515 ;
        RECT -32.805 -7.645 -32.475 -7.315 ;
        RECT -32.805 -10.365 -32.475 -10.035 ;
        RECT -32.805 -14.445 -32.475 -14.115 ;
        RECT -32.805 -17.165 -32.475 -16.835 ;
        RECT -32.805 -18.525 -32.475 -18.195 ;
        RECT -32.805 -19.885 -32.475 -19.555 ;
        RECT -32.805 -21.245 -32.475 -20.915 ;
        RECT -32.805 -22.605 -32.475 -22.275 ;
        RECT -32.805 -23.965 -32.475 -23.635 ;
        RECT -32.805 -25.325 -32.475 -24.995 ;
        RECT -32.805 -32.125 -32.475 -31.795 ;
        RECT -32.805 -33.71 -32.475 -33.38 ;
        RECT -32.805 -34.845 -32.475 -34.515 ;
        RECT -32.805 -36.205 -32.475 -35.875 ;
        RECT -32.805 -38.925 -32.475 -38.595 ;
        RECT -32.805 -39.75 -32.475 -39.42 ;
        RECT -32.805 -41.645 -32.475 -41.315 ;
        RECT -32.805 -44.365 -32.475 -44.035 ;
        RECT -32.805 -49.805 -32.475 -49.475 ;
        RECT -32.805 -51.165 -32.475 -50.835 ;
        RECT -32.805 -53.885 -32.475 -53.555 ;
        RECT -32.805 -55.245 -32.475 -54.915 ;
        RECT -32.805 -59.325 -32.475 -58.995 ;
        RECT -32.805 -60.685 -32.475 -60.355 ;
        RECT -32.805 -63.405 -32.475 -63.075 ;
        RECT -32.805 -70.205 -32.475 -69.875 ;
        RECT -32.805 -71.565 -32.475 -71.235 ;
        RECT -32.805 -72.925 -32.475 -72.595 ;
        RECT -32.805 -74.285 -32.475 -73.955 ;
        RECT -32.805 -75.645 -32.475 -75.315 ;
        RECT -32.805 -77.005 -32.475 -76.675 ;
        RECT -32.805 -78.365 -32.475 -78.035 ;
        RECT -32.805 -79.725 -32.475 -79.395 ;
        RECT -32.805 -81.085 -32.475 -80.755 ;
        RECT -32.805 -82.445 -32.475 -82.115 ;
        RECT -32.805 -83.805 -32.475 -83.475 ;
        RECT -32.805 -85.165 -32.475 -84.835 ;
        RECT -32.805 -86.525 -32.475 -86.195 ;
        RECT -32.805 -87.885 -32.475 -87.555 ;
        RECT -32.805 -89.245 -32.475 -88.915 ;
        RECT -32.805 -90.605 -32.475 -90.275 ;
        RECT -32.805 -91.965 -32.475 -91.635 ;
        RECT -32.805 -93.325 -32.475 -92.995 ;
        RECT -32.805 -94.685 -32.475 -94.355 ;
        RECT -32.805 -96.045 -32.475 -95.715 ;
        RECT -32.805 -97.405 -32.475 -97.075 ;
        RECT -32.805 -98.765 -32.475 -98.435 ;
        RECT -32.805 -100.125 -32.475 -99.795 ;
        RECT -32.805 -101.485 -32.475 -101.155 ;
        RECT -32.805 -102.845 -32.475 -102.515 ;
        RECT -32.805 -104.205 -32.475 -103.875 ;
        RECT -32.805 -105.565 -32.475 -105.235 ;
        RECT -32.805 -106.925 -32.475 -106.595 ;
        RECT -32.805 -108.285 -32.475 -107.955 ;
        RECT -32.805 -109.645 -32.475 -109.315 ;
        RECT -32.805 -111.005 -32.475 -110.675 ;
        RECT -32.805 -112.365 -32.475 -112.035 ;
        RECT -32.805 -113.725 -32.475 -113.395 ;
        RECT -32.805 -115.085 -32.475 -114.755 ;
        RECT -32.805 -116.445 -32.475 -116.115 ;
        RECT -32.805 -117.805 -32.475 -117.475 ;
        RECT -32.805 -119.165 -32.475 -118.835 ;
        RECT -32.805 -120.525 -32.475 -120.195 ;
        RECT -32.805 -123.245 -32.475 -122.915 ;
        RECT -32.805 -125.965 -32.475 -125.635 ;
        RECT -32.805 -127.325 -32.475 -126.995 ;
        RECT -32.805 -128.685 -32.475 -128.355 ;
        RECT -32.805 -130.045 -32.475 -129.715 ;
        RECT -32.805 -134.125 -32.475 -133.795 ;
        RECT -32.805 -135.485 -32.475 -135.155 ;
        RECT -32.805 -136.845 -32.475 -136.515 ;
        RECT -32.805 -138.205 -32.475 -137.875 ;
        RECT -32.805 -139.565 -32.475 -139.235 ;
        RECT -32.805 -142.285 -32.475 -141.955 ;
        RECT -32.805 -143.645 -32.475 -143.315 ;
        RECT -32.805 -145.005 -32.475 -144.675 ;
        RECT -32.805 -146.365 -32.475 -146.035 ;
        RECT -32.805 -147.725 -32.475 -147.395 ;
        RECT -32.805 -149.085 -32.475 -148.755 ;
        RECT -32.805 -151.805 -32.475 -151.475 ;
        RECT -32.805 -153.165 -32.475 -152.835 ;
        RECT -32.805 -157.245 -32.475 -156.915 ;
        RECT -32.805 -158.605 -32.475 -158.275 ;
        RECT -32.805 -159.965 -32.475 -159.635 ;
        RECT -32.805 -161.325 -32.475 -160.995 ;
        RECT -32.805 -162.685 -32.475 -162.355 ;
        RECT -32.805 -164.045 -32.475 -163.715 ;
        RECT -32.805 -165.405 -32.475 -165.075 ;
        RECT -32.805 -166.765 -32.475 -166.435 ;
        RECT -32.8 -167.44 -32.48 245.285 ;
        RECT -32.805 244.04 -32.475 245.17 ;
        RECT -32.805 239.875 -32.475 240.205 ;
        RECT -32.805 238.515 -32.475 238.845 ;
        RECT -32.805 237.155 -32.475 237.485 ;
        RECT -32.805 235.795 -32.475 236.125 ;
        RECT -32.805 234.435 -32.475 234.765 ;
        RECT -32.805 233.075 -32.475 233.405 ;
        RECT -32.805 231.715 -32.475 232.045 ;
        RECT -32.805 230.355 -32.475 230.685 ;
        RECT -32.805 228.995 -32.475 229.325 ;
        RECT -32.805 227.635 -32.475 227.965 ;
        RECT -32.805 226.275 -32.475 226.605 ;
        RECT -32.805 224.915 -32.475 225.245 ;
        RECT -32.805 223.555 -32.475 223.885 ;
        RECT -32.805 222.195 -32.475 222.525 ;
        RECT -32.805 220.835 -32.475 221.165 ;
        RECT -32.805 219.475 -32.475 219.805 ;
        RECT -32.805 218.115 -32.475 218.445 ;
        RECT -32.805 216.755 -32.475 217.085 ;
        RECT -32.805 215.395 -32.475 215.725 ;
        RECT -32.805 214.035 -32.475 214.365 ;
        RECT -32.805 212.675 -32.475 213.005 ;
        RECT -32.805 211.315 -32.475 211.645 ;
        RECT -32.805 209.955 -32.475 210.285 ;
        RECT -32.805 208.595 -32.475 208.925 ;
        RECT -32.805 207.235 -32.475 207.565 ;
        RECT -32.805 205.875 -32.475 206.205 ;
        RECT -32.805 204.515 -32.475 204.845 ;
        RECT -32.805 203.155 -32.475 203.485 ;
        RECT -32.805 201.795 -32.475 202.125 ;
        RECT -32.805 200.435 -32.475 200.765 ;
        RECT -32.805 199.075 -32.475 199.405 ;
        RECT -32.805 197.715 -32.475 198.045 ;
        RECT -32.805 196.355 -32.475 196.685 ;
        RECT -32.805 194.995 -32.475 195.325 ;
        RECT -32.805 193.635 -32.475 193.965 ;
        RECT -32.805 192.275 -32.475 192.605 ;
        RECT -32.805 190.915 -32.475 191.245 ;
        RECT -32.805 189.555 -32.475 189.885 ;
        RECT -32.805 188.195 -32.475 188.525 ;
        RECT -32.805 186.835 -32.475 187.165 ;
        RECT -32.805 185.475 -32.475 185.805 ;
        RECT -32.805 184.115 -32.475 184.445 ;
        RECT -32.805 182.755 -32.475 183.085 ;
        RECT -32.805 181.395 -32.475 181.725 ;
        RECT -32.805 180.035 -32.475 180.365 ;
        RECT -32.805 178.675 -32.475 179.005 ;
        RECT -32.805 177.315 -32.475 177.645 ;
        RECT -32.805 175.955 -32.475 176.285 ;
        RECT -32.805 174.595 -32.475 174.925 ;
        RECT -32.805 173.235 -32.475 173.565 ;
        RECT -32.805 171.875 -32.475 172.205 ;
        RECT -32.805 170.515 -32.475 170.845 ;
        RECT -32.805 169.155 -32.475 169.485 ;
        RECT -32.805 167.795 -32.475 168.125 ;
        RECT -32.805 166.435 -32.475 166.765 ;
        RECT -32.805 165.075 -32.475 165.405 ;
        RECT -32.805 163.715 -32.475 164.045 ;
        RECT -32.805 162.355 -32.475 162.685 ;
        RECT -32.805 160.995 -32.475 161.325 ;
        RECT -32.805 159.635 -32.475 159.965 ;
        RECT -32.805 158.275 -32.475 158.605 ;
        RECT -32.805 156.915 -32.475 157.245 ;
        RECT -32.805 155.555 -32.475 155.885 ;
        RECT -32.805 154.195 -32.475 154.525 ;
        RECT -32.805 152.835 -32.475 153.165 ;
        RECT -32.805 151.475 -32.475 151.805 ;
        RECT -32.805 150.115 -32.475 150.445 ;
        RECT -32.805 148.755 -32.475 149.085 ;
        RECT -32.805 147.395 -32.475 147.725 ;
        RECT -32.805 146.035 -32.475 146.365 ;
        RECT -32.805 144.675 -32.475 145.005 ;
        RECT -32.805 143.315 -32.475 143.645 ;
        RECT -32.805 141.955 -32.475 142.285 ;
        RECT -32.805 140.595 -32.475 140.925 ;
        RECT -32.805 139.235 -32.475 139.565 ;
        RECT -32.805 137.875 -32.475 138.205 ;
        RECT -32.805 136.515 -32.475 136.845 ;
        RECT -32.805 135.155 -32.475 135.485 ;
        RECT -32.805 133.795 -32.475 134.125 ;
        RECT -32.805 132.435 -32.475 132.765 ;
        RECT -32.805 131.075 -32.475 131.405 ;
        RECT -32.805 129.715 -32.475 130.045 ;
        RECT -32.805 128.355 -32.475 128.685 ;
        RECT -32.805 126.995 -32.475 127.325 ;
        RECT -32.805 125.635 -32.475 125.965 ;
        RECT -32.805 124.275 -32.475 124.605 ;
        RECT -32.805 122.915 -32.475 123.245 ;
        RECT -32.805 121.555 -32.475 121.885 ;
        RECT -32.805 120.195 -32.475 120.525 ;
        RECT -32.805 118.835 -32.475 119.165 ;
        RECT -32.805 117.475 -32.475 117.805 ;
        RECT -32.805 116.115 -32.475 116.445 ;
        RECT -32.805 114.755 -32.475 115.085 ;
        RECT -32.805 113.395 -32.475 113.725 ;
        RECT -32.805 112.035 -32.475 112.365 ;
        RECT -32.805 110.675 -32.475 111.005 ;
        RECT -32.805 109.315 -32.475 109.645 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.965 244.04 -40.635 245.17 ;
        RECT -40.965 239.875 -40.635 240.205 ;
        RECT -40.965 238.515 -40.635 238.845 ;
        RECT -40.965 237.155 -40.635 237.485 ;
        RECT -40.965 235.795 -40.635 236.125 ;
        RECT -40.965 234.435 -40.635 234.765 ;
        RECT -40.965 233.075 -40.635 233.405 ;
        RECT -40.965 231.715 -40.635 232.045 ;
        RECT -40.965 230.355 -40.635 230.685 ;
        RECT -40.965 228.995 -40.635 229.325 ;
        RECT -40.965 227.635 -40.635 227.965 ;
        RECT -40.965 226.275 -40.635 226.605 ;
        RECT -40.965 224.915 -40.635 225.245 ;
        RECT -40.965 223.555 -40.635 223.885 ;
        RECT -40.965 222.195 -40.635 222.525 ;
        RECT -40.965 220.835 -40.635 221.165 ;
        RECT -40.965 219.475 -40.635 219.805 ;
        RECT -40.965 218.115 -40.635 218.445 ;
        RECT -40.965 216.755 -40.635 217.085 ;
        RECT -40.965 215.395 -40.635 215.725 ;
        RECT -40.965 214.035 -40.635 214.365 ;
        RECT -40.965 212.675 -40.635 213.005 ;
        RECT -40.965 211.315 -40.635 211.645 ;
        RECT -40.965 209.955 -40.635 210.285 ;
        RECT -40.965 208.595 -40.635 208.925 ;
        RECT -40.965 207.235 -40.635 207.565 ;
        RECT -40.965 205.875 -40.635 206.205 ;
        RECT -40.965 204.515 -40.635 204.845 ;
        RECT -40.965 203.155 -40.635 203.485 ;
        RECT -40.965 201.795 -40.635 202.125 ;
        RECT -40.965 200.435 -40.635 200.765 ;
        RECT -40.965 199.075 -40.635 199.405 ;
        RECT -40.965 197.715 -40.635 198.045 ;
        RECT -40.965 196.355 -40.635 196.685 ;
        RECT -40.965 194.995 -40.635 195.325 ;
        RECT -40.965 193.635 -40.635 193.965 ;
        RECT -40.965 192.275 -40.635 192.605 ;
        RECT -40.965 190.915 -40.635 191.245 ;
        RECT -40.965 189.555 -40.635 189.885 ;
        RECT -40.965 188.195 -40.635 188.525 ;
        RECT -40.965 186.835 -40.635 187.165 ;
        RECT -40.965 185.475 -40.635 185.805 ;
        RECT -40.965 184.115 -40.635 184.445 ;
        RECT -40.965 182.755 -40.635 183.085 ;
        RECT -40.965 181.395 -40.635 181.725 ;
        RECT -40.965 180.035 -40.635 180.365 ;
        RECT -40.965 178.675 -40.635 179.005 ;
        RECT -40.965 177.315 -40.635 177.645 ;
        RECT -40.965 175.955 -40.635 176.285 ;
        RECT -40.965 174.595 -40.635 174.925 ;
        RECT -40.965 173.235 -40.635 173.565 ;
        RECT -40.965 171.875 -40.635 172.205 ;
        RECT -40.965 170.515 -40.635 170.845 ;
        RECT -40.965 169.155 -40.635 169.485 ;
        RECT -40.965 167.795 -40.635 168.125 ;
        RECT -40.965 166.435 -40.635 166.765 ;
        RECT -40.965 165.075 -40.635 165.405 ;
        RECT -40.965 163.715 -40.635 164.045 ;
        RECT -40.965 162.355 -40.635 162.685 ;
        RECT -40.965 160.995 -40.635 161.325 ;
        RECT -40.965 159.635 -40.635 159.965 ;
        RECT -40.965 158.275 -40.635 158.605 ;
        RECT -40.965 156.915 -40.635 157.245 ;
        RECT -40.965 155.555 -40.635 155.885 ;
        RECT -40.965 154.195 -40.635 154.525 ;
        RECT -40.965 152.835 -40.635 153.165 ;
        RECT -40.965 151.475 -40.635 151.805 ;
        RECT -40.965 150.115 -40.635 150.445 ;
        RECT -40.965 148.755 -40.635 149.085 ;
        RECT -40.965 147.395 -40.635 147.725 ;
        RECT -40.965 146.035 -40.635 146.365 ;
        RECT -40.965 144.675 -40.635 145.005 ;
        RECT -40.965 143.315 -40.635 143.645 ;
        RECT -40.965 141.955 -40.635 142.285 ;
        RECT -40.965 140.595 -40.635 140.925 ;
        RECT -40.965 139.235 -40.635 139.565 ;
        RECT -40.965 137.875 -40.635 138.205 ;
        RECT -40.965 136.515 -40.635 136.845 ;
        RECT -40.965 135.155 -40.635 135.485 ;
        RECT -40.965 133.795 -40.635 134.125 ;
        RECT -40.965 132.435 -40.635 132.765 ;
        RECT -40.965 131.075 -40.635 131.405 ;
        RECT -40.965 129.715 -40.635 130.045 ;
        RECT -40.965 128.355 -40.635 128.685 ;
        RECT -40.965 126.995 -40.635 127.325 ;
        RECT -40.965 125.635 -40.635 125.965 ;
        RECT -40.965 124.275 -40.635 124.605 ;
        RECT -40.965 122.915 -40.635 123.245 ;
        RECT -40.965 121.555 -40.635 121.885 ;
        RECT -40.965 120.195 -40.635 120.525 ;
        RECT -40.965 118.835 -40.635 119.165 ;
        RECT -40.965 117.475 -40.635 117.805 ;
        RECT -40.965 116.115 -40.635 116.445 ;
        RECT -40.965 114.755 -40.635 115.085 ;
        RECT -40.965 113.395 -40.635 113.725 ;
        RECT -40.965 112.035 -40.635 112.365 ;
        RECT -40.965 110.675 -40.635 111.005 ;
        RECT -40.965 109.315 -40.635 109.645 ;
        RECT -40.965 107.955 -40.635 108.285 ;
        RECT -40.965 106.595 -40.635 106.925 ;
        RECT -40.965 105.235 -40.635 105.565 ;
        RECT -40.965 103.875 -40.635 104.205 ;
        RECT -40.965 102.515 -40.635 102.845 ;
        RECT -40.965 101.155 -40.635 101.485 ;
        RECT -40.965 99.795 -40.635 100.125 ;
        RECT -40.965 98.435 -40.635 98.765 ;
        RECT -40.965 97.075 -40.635 97.405 ;
        RECT -40.965 95.715 -40.635 96.045 ;
        RECT -40.965 94.355 -40.635 94.685 ;
        RECT -40.965 92.995 -40.635 93.325 ;
        RECT -40.965 91.635 -40.635 91.965 ;
        RECT -40.965 90.275 -40.635 90.605 ;
        RECT -40.965 88.915 -40.635 89.245 ;
        RECT -40.965 87.555 -40.635 87.885 ;
        RECT -40.965 86.195 -40.635 86.525 ;
        RECT -40.965 84.835 -40.635 85.165 ;
        RECT -40.965 83.475 -40.635 83.805 ;
        RECT -40.965 82.115 -40.635 82.445 ;
        RECT -40.965 80.755 -40.635 81.085 ;
        RECT -40.965 79.395 -40.635 79.725 ;
        RECT -40.965 78.035 -40.635 78.365 ;
        RECT -40.965 76.675 -40.635 77.005 ;
        RECT -40.965 75.315 -40.635 75.645 ;
        RECT -40.965 73.955 -40.635 74.285 ;
        RECT -40.965 72.595 -40.635 72.925 ;
        RECT -40.965 71.235 -40.635 71.565 ;
        RECT -40.965 69.875 -40.635 70.205 ;
        RECT -40.965 68.515 -40.635 68.845 ;
        RECT -40.965 67.155 -40.635 67.485 ;
        RECT -40.965 65.795 -40.635 66.125 ;
        RECT -40.965 64.435 -40.635 64.765 ;
        RECT -40.965 63.075 -40.635 63.405 ;
        RECT -40.965 61.715 -40.635 62.045 ;
        RECT -40.965 60.355 -40.635 60.685 ;
        RECT -40.965 58.995 -40.635 59.325 ;
        RECT -40.965 57.635 -40.635 57.965 ;
        RECT -40.965 56.275 -40.635 56.605 ;
        RECT -40.965 54.915 -40.635 55.245 ;
        RECT -40.965 53.555 -40.635 53.885 ;
        RECT -40.965 52.195 -40.635 52.525 ;
        RECT -40.965 50.835 -40.635 51.165 ;
        RECT -40.965 49.475 -40.635 49.805 ;
        RECT -40.965 48.115 -40.635 48.445 ;
        RECT -40.965 46.755 -40.635 47.085 ;
        RECT -40.965 45.395 -40.635 45.725 ;
        RECT -40.965 44.035 -40.635 44.365 ;
        RECT -40.965 42.675 -40.635 43.005 ;
        RECT -40.965 41.315 -40.635 41.645 ;
        RECT -40.965 39.955 -40.635 40.285 ;
        RECT -40.965 38.595 -40.635 38.925 ;
        RECT -40.965 37.235 -40.635 37.565 ;
        RECT -40.965 35.875 -40.635 36.205 ;
        RECT -40.965 34.515 -40.635 34.845 ;
        RECT -40.965 33.155 -40.635 33.485 ;
        RECT -40.965 31.795 -40.635 32.125 ;
        RECT -40.965 30.435 -40.635 30.765 ;
        RECT -40.965 29.075 -40.635 29.405 ;
        RECT -40.965 27.715 -40.635 28.045 ;
        RECT -40.965 26.355 -40.635 26.685 ;
        RECT -40.965 24.995 -40.635 25.325 ;
        RECT -40.965 23.635 -40.635 23.965 ;
        RECT -40.965 22.275 -40.635 22.605 ;
        RECT -40.965 20.915 -40.635 21.245 ;
        RECT -40.965 19.555 -40.635 19.885 ;
        RECT -40.965 18.195 -40.635 18.525 ;
        RECT -40.965 16.835 -40.635 17.165 ;
        RECT -40.965 15.475 -40.635 15.805 ;
        RECT -40.965 14.115 -40.635 14.445 ;
        RECT -40.965 12.755 -40.635 13.085 ;
        RECT -40.965 11.395 -40.635 11.725 ;
        RECT -40.965 10.035 -40.635 10.365 ;
        RECT -40.965 8.675 -40.635 9.005 ;
        RECT -40.965 7.315 -40.635 7.645 ;
        RECT -40.965 5.955 -40.635 6.285 ;
        RECT -40.965 4.595 -40.635 4.925 ;
        RECT -40.965 3.235 -40.635 3.565 ;
        RECT -40.965 1.875 -40.635 2.205 ;
        RECT -40.965 0.515 -40.635 0.845 ;
        RECT -40.965 -0.845 -40.635 -0.515 ;
        RECT -40.965 -2.205 -40.635 -1.875 ;
        RECT -40.965 -3.565 -40.635 -3.235 ;
        RECT -40.965 -4.925 -40.635 -4.595 ;
        RECT -40.965 -6.285 -40.635 -5.955 ;
        RECT -40.965 -10.365 -40.635 -10.035 ;
        RECT -40.965 -14.445 -40.635 -14.115 ;
        RECT -40.965 -17.165 -40.635 -16.835 ;
        RECT -40.965 -18.525 -40.635 -18.195 ;
        RECT -40.965 -19.885 -40.635 -19.555 ;
        RECT -40.965 -21.245 -40.635 -20.915 ;
        RECT -40.965 -22.605 -40.635 -22.275 ;
        RECT -40.965 -23.965 -40.635 -23.635 ;
        RECT -40.965 -25.325 -40.635 -24.995 ;
        RECT -40.965 -32.125 -40.635 -31.795 ;
        RECT -40.965 -33.71 -40.635 -33.38 ;
        RECT -40.965 -34.845 -40.635 -34.515 ;
        RECT -40.965 -36.205 -40.635 -35.875 ;
        RECT -40.965 -38.925 -40.635 -38.595 ;
        RECT -40.965 -39.75 -40.635 -39.42 ;
        RECT -40.965 -41.645 -40.635 -41.315 ;
        RECT -40.965 -44.365 -40.635 -44.035 ;
        RECT -40.965 -49.805 -40.635 -49.475 ;
        RECT -40.965 -51.165 -40.635 -50.835 ;
        RECT -40.965 -53.885 -40.635 -53.555 ;
        RECT -40.965 -55.245 -40.635 -54.915 ;
        RECT -40.965 -59.325 -40.635 -58.995 ;
        RECT -40.965 -60.685 -40.635 -60.355 ;
        RECT -40.965 -63.405 -40.635 -63.075 ;
        RECT -40.965 -67.485 -40.635 -67.155 ;
        RECT -40.965 -70.205 -40.635 -69.875 ;
        RECT -40.965 -71.565 -40.635 -71.235 ;
        RECT -40.965 -72.925 -40.635 -72.595 ;
        RECT -40.965 -74.285 -40.635 -73.955 ;
        RECT -40.965 -75.645 -40.635 -75.315 ;
        RECT -40.965 -77.005 -40.635 -76.675 ;
        RECT -40.965 -78.365 -40.635 -78.035 ;
        RECT -40.965 -79.725 -40.635 -79.395 ;
        RECT -40.965 -81.085 -40.635 -80.755 ;
        RECT -40.965 -82.445 -40.635 -82.115 ;
        RECT -40.965 -83.805 -40.635 -83.475 ;
        RECT -40.965 -85.165 -40.635 -84.835 ;
        RECT -40.965 -86.525 -40.635 -86.195 ;
        RECT -40.965 -87.885 -40.635 -87.555 ;
        RECT -40.965 -89.245 -40.635 -88.915 ;
        RECT -40.965 -90.605 -40.635 -90.275 ;
        RECT -40.965 -91.77 -40.635 -91.44 ;
        RECT -40.965 -93.325 -40.635 -92.995 ;
        RECT -40.965 -94.685 -40.635 -94.355 ;
        RECT -40.965 -96.045 -40.635 -95.715 ;
        RECT -40.965 -97.405 -40.635 -97.075 ;
        RECT -40.965 -98.765 -40.635 -98.435 ;
        RECT -40.965 -101.485 -40.635 -101.155 ;
        RECT -40.965 -102.31 -40.635 -101.98 ;
        RECT -40.965 -104.205 -40.635 -103.875 ;
        RECT -40.965 -105.565 -40.635 -105.235 ;
        RECT -40.965 -106.925 -40.635 -106.595 ;
        RECT -40.965 -109.645 -40.635 -109.315 ;
        RECT -40.965 -111.005 -40.635 -110.675 ;
        RECT -40.965 -113.725 -40.635 -113.395 ;
        RECT -40.965 -115.085 -40.635 -114.755 ;
        RECT -40.965 -116.445 -40.635 -116.115 ;
        RECT -40.965 -117.805 -40.635 -117.475 ;
        RECT -40.965 -119.165 -40.635 -118.835 ;
        RECT -40.965 -120.525 -40.635 -120.195 ;
        RECT -40.965 -123.245 -40.635 -122.915 ;
        RECT -40.965 -124.605 -40.635 -124.275 ;
        RECT -40.965 -125.965 -40.635 -125.635 ;
        RECT -40.965 -127.325 -40.635 -126.995 ;
        RECT -40.965 -128.685 -40.635 -128.355 ;
        RECT -40.965 -130.045 -40.635 -129.715 ;
        RECT -40.965 -131.405 -40.635 -131.075 ;
        RECT -40.965 -132.765 -40.635 -132.435 ;
        RECT -40.965 -134.125 -40.635 -133.795 ;
        RECT -40.965 -135.485 -40.635 -135.155 ;
        RECT -40.965 -136.845 -40.635 -136.515 ;
        RECT -40.965 -138.205 -40.635 -137.875 ;
        RECT -40.965 -139.565 -40.635 -139.235 ;
        RECT -40.965 -140.925 -40.635 -140.595 ;
        RECT -40.965 -142.285 -40.635 -141.955 ;
        RECT -40.965 -143.645 -40.635 -143.315 ;
        RECT -40.965 -145.005 -40.635 -144.675 ;
        RECT -40.965 -146.365 -40.635 -146.035 ;
        RECT -40.965 -147.725 -40.635 -147.395 ;
        RECT -40.965 -149.085 -40.635 -148.755 ;
        RECT -40.965 -151.805 -40.635 -151.475 ;
        RECT -40.965 -153.165 -40.635 -152.835 ;
        RECT -40.965 -154.525 -40.635 -154.195 ;
        RECT -40.965 -155.885 -40.635 -155.555 ;
        RECT -40.965 -158.605 -40.635 -158.275 ;
        RECT -40.965 -159.965 -40.635 -159.635 ;
        RECT -40.965 -161.325 -40.635 -160.995 ;
        RECT -40.965 -162.685 -40.635 -162.355 ;
        RECT -40.965 -164.045 -40.635 -163.715 ;
        RECT -40.965 -165.405 -40.635 -165.075 ;
        RECT -40.965 -166.765 -40.635 -166.435 ;
        RECT -40.965 -170.845 -40.635 -170.515 ;
        RECT -40.965 -172.205 -40.635 -171.875 ;
        RECT -40.965 -174.925 -40.635 -174.595 ;
        RECT -40.965 -177.645 -40.635 -177.315 ;
        RECT -40.965 -179.005 -40.635 -178.675 ;
        RECT -40.965 -184.65 -40.635 -183.52 ;
        RECT -40.96 -184.765 -40.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -39.605 244.04 -39.275 245.17 ;
        RECT -39.605 239.875 -39.275 240.205 ;
        RECT -39.605 238.515 -39.275 238.845 ;
        RECT -39.605 237.155 -39.275 237.485 ;
        RECT -39.605 235.795 -39.275 236.125 ;
        RECT -39.605 234.435 -39.275 234.765 ;
        RECT -39.605 233.075 -39.275 233.405 ;
        RECT -39.605 231.715 -39.275 232.045 ;
        RECT -39.605 230.355 -39.275 230.685 ;
        RECT -39.605 228.995 -39.275 229.325 ;
        RECT -39.605 227.635 -39.275 227.965 ;
        RECT -39.605 226.275 -39.275 226.605 ;
        RECT -39.605 224.915 -39.275 225.245 ;
        RECT -39.605 223.555 -39.275 223.885 ;
        RECT -39.605 222.195 -39.275 222.525 ;
        RECT -39.605 220.835 -39.275 221.165 ;
        RECT -39.605 219.475 -39.275 219.805 ;
        RECT -39.605 218.115 -39.275 218.445 ;
        RECT -39.605 216.755 -39.275 217.085 ;
        RECT -39.605 215.395 -39.275 215.725 ;
        RECT -39.605 214.035 -39.275 214.365 ;
        RECT -39.605 212.675 -39.275 213.005 ;
        RECT -39.605 211.315 -39.275 211.645 ;
        RECT -39.605 209.955 -39.275 210.285 ;
        RECT -39.605 208.595 -39.275 208.925 ;
        RECT -39.605 207.235 -39.275 207.565 ;
        RECT -39.605 205.875 -39.275 206.205 ;
        RECT -39.605 204.515 -39.275 204.845 ;
        RECT -39.605 203.155 -39.275 203.485 ;
        RECT -39.605 201.795 -39.275 202.125 ;
        RECT -39.605 200.435 -39.275 200.765 ;
        RECT -39.605 199.075 -39.275 199.405 ;
        RECT -39.605 197.715 -39.275 198.045 ;
        RECT -39.605 196.355 -39.275 196.685 ;
        RECT -39.605 194.995 -39.275 195.325 ;
        RECT -39.605 193.635 -39.275 193.965 ;
        RECT -39.605 192.275 -39.275 192.605 ;
        RECT -39.605 190.915 -39.275 191.245 ;
        RECT -39.605 189.555 -39.275 189.885 ;
        RECT -39.605 188.195 -39.275 188.525 ;
        RECT -39.605 186.835 -39.275 187.165 ;
        RECT -39.605 185.475 -39.275 185.805 ;
        RECT -39.605 184.115 -39.275 184.445 ;
        RECT -39.605 182.755 -39.275 183.085 ;
        RECT -39.605 181.395 -39.275 181.725 ;
        RECT -39.605 180.035 -39.275 180.365 ;
        RECT -39.605 178.675 -39.275 179.005 ;
        RECT -39.605 177.315 -39.275 177.645 ;
        RECT -39.605 175.955 -39.275 176.285 ;
        RECT -39.605 174.595 -39.275 174.925 ;
        RECT -39.605 173.235 -39.275 173.565 ;
        RECT -39.605 171.875 -39.275 172.205 ;
        RECT -39.605 170.515 -39.275 170.845 ;
        RECT -39.605 169.155 -39.275 169.485 ;
        RECT -39.605 167.795 -39.275 168.125 ;
        RECT -39.605 166.435 -39.275 166.765 ;
        RECT -39.605 165.075 -39.275 165.405 ;
        RECT -39.605 163.715 -39.275 164.045 ;
        RECT -39.605 162.355 -39.275 162.685 ;
        RECT -39.605 160.995 -39.275 161.325 ;
        RECT -39.605 159.635 -39.275 159.965 ;
        RECT -39.605 158.275 -39.275 158.605 ;
        RECT -39.605 156.915 -39.275 157.245 ;
        RECT -39.605 155.555 -39.275 155.885 ;
        RECT -39.605 154.195 -39.275 154.525 ;
        RECT -39.605 152.835 -39.275 153.165 ;
        RECT -39.605 151.475 -39.275 151.805 ;
        RECT -39.605 150.115 -39.275 150.445 ;
        RECT -39.605 148.755 -39.275 149.085 ;
        RECT -39.605 147.395 -39.275 147.725 ;
        RECT -39.605 146.035 -39.275 146.365 ;
        RECT -39.605 144.675 -39.275 145.005 ;
        RECT -39.605 143.315 -39.275 143.645 ;
        RECT -39.605 141.955 -39.275 142.285 ;
        RECT -39.605 140.595 -39.275 140.925 ;
        RECT -39.605 139.235 -39.275 139.565 ;
        RECT -39.605 137.875 -39.275 138.205 ;
        RECT -39.605 136.515 -39.275 136.845 ;
        RECT -39.605 135.155 -39.275 135.485 ;
        RECT -39.605 133.795 -39.275 134.125 ;
        RECT -39.605 132.435 -39.275 132.765 ;
        RECT -39.605 131.075 -39.275 131.405 ;
        RECT -39.605 129.715 -39.275 130.045 ;
        RECT -39.605 128.355 -39.275 128.685 ;
        RECT -39.605 126.995 -39.275 127.325 ;
        RECT -39.605 125.635 -39.275 125.965 ;
        RECT -39.605 124.275 -39.275 124.605 ;
        RECT -39.605 122.915 -39.275 123.245 ;
        RECT -39.605 121.555 -39.275 121.885 ;
        RECT -39.605 120.195 -39.275 120.525 ;
        RECT -39.605 118.835 -39.275 119.165 ;
        RECT -39.605 117.475 -39.275 117.805 ;
        RECT -39.605 116.115 -39.275 116.445 ;
        RECT -39.605 114.755 -39.275 115.085 ;
        RECT -39.605 113.395 -39.275 113.725 ;
        RECT -39.605 112.035 -39.275 112.365 ;
        RECT -39.605 110.675 -39.275 111.005 ;
        RECT -39.605 109.315 -39.275 109.645 ;
        RECT -39.605 107.955 -39.275 108.285 ;
        RECT -39.605 106.595 -39.275 106.925 ;
        RECT -39.605 105.235 -39.275 105.565 ;
        RECT -39.605 103.875 -39.275 104.205 ;
        RECT -39.605 102.515 -39.275 102.845 ;
        RECT -39.605 101.155 -39.275 101.485 ;
        RECT -39.605 99.795 -39.275 100.125 ;
        RECT -39.605 98.435 -39.275 98.765 ;
        RECT -39.605 97.075 -39.275 97.405 ;
        RECT -39.605 95.715 -39.275 96.045 ;
        RECT -39.605 94.355 -39.275 94.685 ;
        RECT -39.605 92.995 -39.275 93.325 ;
        RECT -39.605 91.635 -39.275 91.965 ;
        RECT -39.605 90.275 -39.275 90.605 ;
        RECT -39.605 88.915 -39.275 89.245 ;
        RECT -39.605 87.555 -39.275 87.885 ;
        RECT -39.605 86.195 -39.275 86.525 ;
        RECT -39.605 84.835 -39.275 85.165 ;
        RECT -39.605 83.475 -39.275 83.805 ;
        RECT -39.605 82.115 -39.275 82.445 ;
        RECT -39.605 80.755 -39.275 81.085 ;
        RECT -39.605 79.395 -39.275 79.725 ;
        RECT -39.605 78.035 -39.275 78.365 ;
        RECT -39.605 76.675 -39.275 77.005 ;
        RECT -39.605 75.315 -39.275 75.645 ;
        RECT -39.605 73.955 -39.275 74.285 ;
        RECT -39.605 72.595 -39.275 72.925 ;
        RECT -39.605 71.235 -39.275 71.565 ;
        RECT -39.605 69.875 -39.275 70.205 ;
        RECT -39.605 68.515 -39.275 68.845 ;
        RECT -39.605 67.155 -39.275 67.485 ;
        RECT -39.605 65.795 -39.275 66.125 ;
        RECT -39.605 64.435 -39.275 64.765 ;
        RECT -39.605 63.075 -39.275 63.405 ;
        RECT -39.605 61.715 -39.275 62.045 ;
        RECT -39.605 60.355 -39.275 60.685 ;
        RECT -39.605 58.995 -39.275 59.325 ;
        RECT -39.605 57.635 -39.275 57.965 ;
        RECT -39.605 56.275 -39.275 56.605 ;
        RECT -39.605 54.915 -39.275 55.245 ;
        RECT -39.605 53.555 -39.275 53.885 ;
        RECT -39.605 52.195 -39.275 52.525 ;
        RECT -39.605 50.835 -39.275 51.165 ;
        RECT -39.605 49.475 -39.275 49.805 ;
        RECT -39.605 48.115 -39.275 48.445 ;
        RECT -39.605 46.755 -39.275 47.085 ;
        RECT -39.605 45.395 -39.275 45.725 ;
        RECT -39.605 44.035 -39.275 44.365 ;
        RECT -39.605 42.675 -39.275 43.005 ;
        RECT -39.605 41.315 -39.275 41.645 ;
        RECT -39.605 39.955 -39.275 40.285 ;
        RECT -39.605 38.595 -39.275 38.925 ;
        RECT -39.605 37.235 -39.275 37.565 ;
        RECT -39.605 35.875 -39.275 36.205 ;
        RECT -39.605 34.515 -39.275 34.845 ;
        RECT -39.605 33.155 -39.275 33.485 ;
        RECT -39.605 31.795 -39.275 32.125 ;
        RECT -39.605 30.435 -39.275 30.765 ;
        RECT -39.605 29.075 -39.275 29.405 ;
        RECT -39.605 27.715 -39.275 28.045 ;
        RECT -39.605 26.355 -39.275 26.685 ;
        RECT -39.605 24.995 -39.275 25.325 ;
        RECT -39.605 23.635 -39.275 23.965 ;
        RECT -39.605 22.275 -39.275 22.605 ;
        RECT -39.605 20.915 -39.275 21.245 ;
        RECT -39.605 19.555 -39.275 19.885 ;
        RECT -39.605 18.195 -39.275 18.525 ;
        RECT -39.605 16.835 -39.275 17.165 ;
        RECT -39.605 15.475 -39.275 15.805 ;
        RECT -39.605 14.115 -39.275 14.445 ;
        RECT -39.605 12.755 -39.275 13.085 ;
        RECT -39.605 11.395 -39.275 11.725 ;
        RECT -39.605 10.035 -39.275 10.365 ;
        RECT -39.605 8.675 -39.275 9.005 ;
        RECT -39.605 7.315 -39.275 7.645 ;
        RECT -39.605 5.955 -39.275 6.285 ;
        RECT -39.605 4.595 -39.275 4.925 ;
        RECT -39.605 3.235 -39.275 3.565 ;
        RECT -39.605 1.875 -39.275 2.205 ;
        RECT -39.605 0.515 -39.275 0.845 ;
        RECT -39.605 -0.845 -39.275 -0.515 ;
        RECT -39.605 -2.205 -39.275 -1.875 ;
        RECT -39.605 -3.565 -39.275 -3.235 ;
        RECT -39.605 -4.925 -39.275 -4.595 ;
        RECT -39.605 -10.365 -39.275 -10.035 ;
        RECT -39.605 -14.445 -39.275 -14.115 ;
        RECT -39.605 -17.165 -39.275 -16.835 ;
        RECT -39.605 -18.525 -39.275 -18.195 ;
        RECT -39.605 -19.885 -39.275 -19.555 ;
        RECT -39.605 -21.245 -39.275 -20.915 ;
        RECT -39.605 -22.605 -39.275 -22.275 ;
        RECT -39.605 -23.965 -39.275 -23.635 ;
        RECT -39.605 -25.325 -39.275 -24.995 ;
        RECT -39.605 -32.125 -39.275 -31.795 ;
        RECT -39.605 -33.71 -39.275 -33.38 ;
        RECT -39.605 -34.845 -39.275 -34.515 ;
        RECT -39.605 -36.205 -39.275 -35.875 ;
        RECT -39.605 -38.925 -39.275 -38.595 ;
        RECT -39.605 -39.75 -39.275 -39.42 ;
        RECT -39.605 -41.645 -39.275 -41.315 ;
        RECT -39.605 -44.365 -39.275 -44.035 ;
        RECT -39.605 -49.805 -39.275 -49.475 ;
        RECT -39.605 -51.165 -39.275 -50.835 ;
        RECT -39.605 -53.885 -39.275 -53.555 ;
        RECT -39.605 -55.245 -39.275 -54.915 ;
        RECT -39.605 -59.325 -39.275 -58.995 ;
        RECT -39.605 -60.685 -39.275 -60.355 ;
        RECT -39.605 -63.405 -39.275 -63.075 ;
        RECT -39.605 -67.485 -39.275 -67.155 ;
        RECT -39.605 -70.205 -39.275 -69.875 ;
        RECT -39.605 -71.565 -39.275 -71.235 ;
        RECT -39.605 -72.925 -39.275 -72.595 ;
        RECT -39.605 -74.285 -39.275 -73.955 ;
        RECT -39.605 -75.645 -39.275 -75.315 ;
        RECT -39.605 -77.005 -39.275 -76.675 ;
        RECT -39.605 -78.365 -39.275 -78.035 ;
        RECT -39.605 -79.725 -39.275 -79.395 ;
        RECT -39.605 -81.085 -39.275 -80.755 ;
        RECT -39.605 -82.445 -39.275 -82.115 ;
        RECT -39.605 -83.805 -39.275 -83.475 ;
        RECT -39.605 -85.165 -39.275 -84.835 ;
        RECT -39.605 -86.525 -39.275 -86.195 ;
        RECT -39.605 -87.885 -39.275 -87.555 ;
        RECT -39.605 -89.245 -39.275 -88.915 ;
        RECT -39.605 -90.605 -39.275 -90.275 ;
        RECT -39.605 -91.77 -39.275 -91.44 ;
        RECT -39.605 -93.325 -39.275 -92.995 ;
        RECT -39.605 -94.685 -39.275 -94.355 ;
        RECT -39.605 -96.045 -39.275 -95.715 ;
        RECT -39.605 -97.405 -39.275 -97.075 ;
        RECT -39.605 -98.765 -39.275 -98.435 ;
        RECT -39.605 -101.485 -39.275 -101.155 ;
        RECT -39.605 -102.31 -39.275 -101.98 ;
        RECT -39.605 -104.205 -39.275 -103.875 ;
        RECT -39.605 -105.565 -39.275 -105.235 ;
        RECT -39.605 -106.925 -39.275 -106.595 ;
        RECT -39.605 -109.645 -39.275 -109.315 ;
        RECT -39.605 -111.005 -39.275 -110.675 ;
        RECT -39.605 -115.085 -39.275 -114.755 ;
        RECT -39.605 -116.445 -39.275 -116.115 ;
        RECT -39.605 -117.805 -39.275 -117.475 ;
        RECT -39.605 -119.165 -39.275 -118.835 ;
        RECT -39.605 -120.525 -39.275 -120.195 ;
        RECT -39.605 -123.245 -39.275 -122.915 ;
        RECT -39.605 -124.605 -39.275 -124.275 ;
        RECT -39.605 -125.965 -39.275 -125.635 ;
        RECT -39.605 -127.325 -39.275 -126.995 ;
        RECT -39.605 -128.685 -39.275 -128.355 ;
        RECT -39.605 -130.045 -39.275 -129.715 ;
        RECT -39.605 -131.405 -39.275 -131.075 ;
        RECT -39.605 -134.125 -39.275 -133.795 ;
        RECT -39.605 -135.485 -39.275 -135.155 ;
        RECT -39.605 -136.845 -39.275 -136.515 ;
        RECT -39.605 -138.205 -39.275 -137.875 ;
        RECT -39.605 -139.565 -39.275 -139.235 ;
        RECT -39.605 -140.925 -39.275 -140.595 ;
        RECT -39.605 -142.285 -39.275 -141.955 ;
        RECT -39.605 -143.645 -39.275 -143.315 ;
        RECT -39.605 -145.005 -39.275 -144.675 ;
        RECT -39.605 -146.365 -39.275 -146.035 ;
        RECT -39.605 -147.725 -39.275 -147.395 ;
        RECT -39.605 -149.085 -39.275 -148.755 ;
        RECT -39.605 -151.805 -39.275 -151.475 ;
        RECT -39.605 -153.165 -39.275 -152.835 ;
        RECT -39.605 -155.885 -39.275 -155.555 ;
        RECT -39.605 -158.605 -39.275 -158.275 ;
        RECT -39.605 -159.965 -39.275 -159.635 ;
        RECT -39.605 -161.325 -39.275 -160.995 ;
        RECT -39.605 -162.685 -39.275 -162.355 ;
        RECT -39.605 -164.045 -39.275 -163.715 ;
        RECT -39.605 -165.405 -39.275 -165.075 ;
        RECT -39.605 -166.765 -39.275 -166.435 ;
        RECT -39.605 -169.615 -39.275 -169.285 ;
        RECT -39.605 -170.845 -39.275 -170.515 ;
        RECT -39.605 -172.205 -39.275 -171.875 ;
        RECT -39.605 -174.925 -39.275 -174.595 ;
        RECT -39.605 -177.645 -39.275 -177.315 ;
        RECT -39.605 -179.005 -39.275 -178.675 ;
        RECT -39.605 -184.65 -39.275 -183.52 ;
        RECT -39.6 -184.765 -39.28 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.245 214.035 -37.915 214.365 ;
        RECT -38.245 212.675 -37.915 213.005 ;
        RECT -38.245 211.315 -37.915 211.645 ;
        RECT -38.245 209.955 -37.915 210.285 ;
        RECT -38.245 208.595 -37.915 208.925 ;
        RECT -38.245 207.235 -37.915 207.565 ;
        RECT -38.245 205.875 -37.915 206.205 ;
        RECT -38.245 204.515 -37.915 204.845 ;
        RECT -38.245 203.155 -37.915 203.485 ;
        RECT -38.245 201.795 -37.915 202.125 ;
        RECT -38.245 200.435 -37.915 200.765 ;
        RECT -38.245 199.075 -37.915 199.405 ;
        RECT -38.245 197.715 -37.915 198.045 ;
        RECT -38.245 196.355 -37.915 196.685 ;
        RECT -38.245 194.995 -37.915 195.325 ;
        RECT -38.245 193.635 -37.915 193.965 ;
        RECT -38.245 192.275 -37.915 192.605 ;
        RECT -38.245 190.915 -37.915 191.245 ;
        RECT -38.245 189.555 -37.915 189.885 ;
        RECT -38.245 188.195 -37.915 188.525 ;
        RECT -38.245 186.835 -37.915 187.165 ;
        RECT -38.245 185.475 -37.915 185.805 ;
        RECT -38.245 184.115 -37.915 184.445 ;
        RECT -38.245 182.755 -37.915 183.085 ;
        RECT -38.245 181.395 -37.915 181.725 ;
        RECT -38.245 180.035 -37.915 180.365 ;
        RECT -38.245 178.675 -37.915 179.005 ;
        RECT -38.245 177.315 -37.915 177.645 ;
        RECT -38.245 175.955 -37.915 176.285 ;
        RECT -38.245 174.595 -37.915 174.925 ;
        RECT -38.245 173.235 -37.915 173.565 ;
        RECT -38.245 171.875 -37.915 172.205 ;
        RECT -38.245 170.515 -37.915 170.845 ;
        RECT -38.245 169.155 -37.915 169.485 ;
        RECT -38.245 167.795 -37.915 168.125 ;
        RECT -38.245 166.435 -37.915 166.765 ;
        RECT -38.245 165.075 -37.915 165.405 ;
        RECT -38.245 163.715 -37.915 164.045 ;
        RECT -38.245 162.355 -37.915 162.685 ;
        RECT -38.245 160.995 -37.915 161.325 ;
        RECT -38.245 159.635 -37.915 159.965 ;
        RECT -38.245 158.275 -37.915 158.605 ;
        RECT -38.245 156.915 -37.915 157.245 ;
        RECT -38.245 155.555 -37.915 155.885 ;
        RECT -38.245 154.195 -37.915 154.525 ;
        RECT -38.245 152.835 -37.915 153.165 ;
        RECT -38.245 151.475 -37.915 151.805 ;
        RECT -38.245 150.115 -37.915 150.445 ;
        RECT -38.245 148.755 -37.915 149.085 ;
        RECT -38.245 147.395 -37.915 147.725 ;
        RECT -38.245 146.035 -37.915 146.365 ;
        RECT -38.245 144.675 -37.915 145.005 ;
        RECT -38.245 143.315 -37.915 143.645 ;
        RECT -38.245 141.955 -37.915 142.285 ;
        RECT -38.245 140.595 -37.915 140.925 ;
        RECT -38.245 139.235 -37.915 139.565 ;
        RECT -38.245 137.875 -37.915 138.205 ;
        RECT -38.245 136.515 -37.915 136.845 ;
        RECT -38.245 135.155 -37.915 135.485 ;
        RECT -38.245 133.795 -37.915 134.125 ;
        RECT -38.245 132.435 -37.915 132.765 ;
        RECT -38.245 131.075 -37.915 131.405 ;
        RECT -38.245 129.715 -37.915 130.045 ;
        RECT -38.245 128.355 -37.915 128.685 ;
        RECT -38.245 126.995 -37.915 127.325 ;
        RECT -38.245 125.635 -37.915 125.965 ;
        RECT -38.245 124.275 -37.915 124.605 ;
        RECT -38.245 122.915 -37.915 123.245 ;
        RECT -38.245 121.555 -37.915 121.885 ;
        RECT -38.245 120.195 -37.915 120.525 ;
        RECT -38.245 118.835 -37.915 119.165 ;
        RECT -38.245 117.475 -37.915 117.805 ;
        RECT -38.245 116.115 -37.915 116.445 ;
        RECT -38.245 114.755 -37.915 115.085 ;
        RECT -38.245 113.395 -37.915 113.725 ;
        RECT -38.245 112.035 -37.915 112.365 ;
        RECT -38.245 110.675 -37.915 111.005 ;
        RECT -38.245 109.315 -37.915 109.645 ;
        RECT -38.245 107.955 -37.915 108.285 ;
        RECT -38.245 106.595 -37.915 106.925 ;
        RECT -38.245 105.235 -37.915 105.565 ;
        RECT -38.245 103.875 -37.915 104.205 ;
        RECT -38.245 102.515 -37.915 102.845 ;
        RECT -38.245 101.155 -37.915 101.485 ;
        RECT -38.245 99.795 -37.915 100.125 ;
        RECT -38.245 98.435 -37.915 98.765 ;
        RECT -38.245 97.075 -37.915 97.405 ;
        RECT -38.245 95.715 -37.915 96.045 ;
        RECT -38.245 94.355 -37.915 94.685 ;
        RECT -38.245 92.995 -37.915 93.325 ;
        RECT -38.245 91.635 -37.915 91.965 ;
        RECT -38.245 90.275 -37.915 90.605 ;
        RECT -38.245 88.915 -37.915 89.245 ;
        RECT -38.245 87.555 -37.915 87.885 ;
        RECT -38.245 86.195 -37.915 86.525 ;
        RECT -38.245 84.835 -37.915 85.165 ;
        RECT -38.245 83.475 -37.915 83.805 ;
        RECT -38.245 82.115 -37.915 82.445 ;
        RECT -38.245 80.755 -37.915 81.085 ;
        RECT -38.245 79.395 -37.915 79.725 ;
        RECT -38.245 78.035 -37.915 78.365 ;
        RECT -38.245 76.675 -37.915 77.005 ;
        RECT -38.245 75.315 -37.915 75.645 ;
        RECT -38.245 73.955 -37.915 74.285 ;
        RECT -38.245 72.595 -37.915 72.925 ;
        RECT -38.245 71.235 -37.915 71.565 ;
        RECT -38.245 69.875 -37.915 70.205 ;
        RECT -38.245 68.515 -37.915 68.845 ;
        RECT -38.245 67.155 -37.915 67.485 ;
        RECT -38.245 65.795 -37.915 66.125 ;
        RECT -38.245 64.435 -37.915 64.765 ;
        RECT -38.245 63.075 -37.915 63.405 ;
        RECT -38.245 61.715 -37.915 62.045 ;
        RECT -38.245 60.355 -37.915 60.685 ;
        RECT -38.245 58.995 -37.915 59.325 ;
        RECT -38.245 57.635 -37.915 57.965 ;
        RECT -38.245 56.275 -37.915 56.605 ;
        RECT -38.245 54.915 -37.915 55.245 ;
        RECT -38.245 53.555 -37.915 53.885 ;
        RECT -38.245 52.195 -37.915 52.525 ;
        RECT -38.245 50.835 -37.915 51.165 ;
        RECT -38.245 49.475 -37.915 49.805 ;
        RECT -38.245 48.115 -37.915 48.445 ;
        RECT -38.245 46.755 -37.915 47.085 ;
        RECT -38.245 45.395 -37.915 45.725 ;
        RECT -38.245 44.035 -37.915 44.365 ;
        RECT -38.245 42.675 -37.915 43.005 ;
        RECT -38.245 41.315 -37.915 41.645 ;
        RECT -38.245 39.955 -37.915 40.285 ;
        RECT -38.245 38.595 -37.915 38.925 ;
        RECT -38.245 37.235 -37.915 37.565 ;
        RECT -38.245 35.875 -37.915 36.205 ;
        RECT -38.245 34.515 -37.915 34.845 ;
        RECT -38.245 33.155 -37.915 33.485 ;
        RECT -38.245 31.795 -37.915 32.125 ;
        RECT -38.245 30.435 -37.915 30.765 ;
        RECT -38.245 29.075 -37.915 29.405 ;
        RECT -38.245 27.715 -37.915 28.045 ;
        RECT -38.245 26.355 -37.915 26.685 ;
        RECT -38.245 24.995 -37.915 25.325 ;
        RECT -38.245 23.635 -37.915 23.965 ;
        RECT -38.245 22.275 -37.915 22.605 ;
        RECT -38.245 20.915 -37.915 21.245 ;
        RECT -38.245 19.555 -37.915 19.885 ;
        RECT -38.245 18.195 -37.915 18.525 ;
        RECT -38.245 16.835 -37.915 17.165 ;
        RECT -38.245 15.475 -37.915 15.805 ;
        RECT -38.245 14.115 -37.915 14.445 ;
        RECT -38.245 12.755 -37.915 13.085 ;
        RECT -38.245 11.395 -37.915 11.725 ;
        RECT -38.245 10.035 -37.915 10.365 ;
        RECT -38.245 8.675 -37.915 9.005 ;
        RECT -38.245 7.315 -37.915 7.645 ;
        RECT -38.245 5.955 -37.915 6.285 ;
        RECT -38.245 4.595 -37.915 4.925 ;
        RECT -38.245 3.235 -37.915 3.565 ;
        RECT -38.245 1.875 -37.915 2.205 ;
        RECT -38.245 0.515 -37.915 0.845 ;
        RECT -38.245 -0.845 -37.915 -0.515 ;
        RECT -38.245 -2.205 -37.915 -1.875 ;
        RECT -38.245 -3.565 -37.915 -3.235 ;
        RECT -38.245 -10.365 -37.915 -10.035 ;
        RECT -38.245 -14.445 -37.915 -14.115 ;
        RECT -38.245 -17.165 -37.915 -16.835 ;
        RECT -38.245 -18.525 -37.915 -18.195 ;
        RECT -38.245 -19.885 -37.915 -19.555 ;
        RECT -38.245 -21.245 -37.915 -20.915 ;
        RECT -38.245 -22.605 -37.915 -22.275 ;
        RECT -38.245 -23.965 -37.915 -23.635 ;
        RECT -38.245 -25.325 -37.915 -24.995 ;
        RECT -38.245 -32.125 -37.915 -31.795 ;
        RECT -38.245 -33.71 -37.915 -33.38 ;
        RECT -38.245 -34.845 -37.915 -34.515 ;
        RECT -38.245 -36.205 -37.915 -35.875 ;
        RECT -38.245 -38.925 -37.915 -38.595 ;
        RECT -38.245 -39.75 -37.915 -39.42 ;
        RECT -38.245 -41.645 -37.915 -41.315 ;
        RECT -38.245 -44.365 -37.915 -44.035 ;
        RECT -38.245 -49.805 -37.915 -49.475 ;
        RECT -38.245 -51.165 -37.915 -50.835 ;
        RECT -38.245 -52.525 -37.915 -52.195 ;
        RECT -38.245 -53.885 -37.915 -53.555 ;
        RECT -38.245 -55.245 -37.915 -54.915 ;
        RECT -38.245 -56.605 -37.915 -56.275 ;
        RECT -38.245 -57.965 -37.915 -57.635 ;
        RECT -38.245 -59.325 -37.915 -58.995 ;
        RECT -38.245 -60.685 -37.915 -60.355 ;
        RECT -38.245 -62.045 -37.915 -61.715 ;
        RECT -38.245 -63.405 -37.915 -63.075 ;
        RECT -38.245 -64.765 -37.915 -64.435 ;
        RECT -38.245 -66.125 -37.915 -65.795 ;
        RECT -38.245 -70.205 -37.915 -69.875 ;
        RECT -38.245 -71.565 -37.915 -71.235 ;
        RECT -38.245 -72.925 -37.915 -72.595 ;
        RECT -38.245 -74.285 -37.915 -73.955 ;
        RECT -38.245 -75.645 -37.915 -75.315 ;
        RECT -38.245 -77.005 -37.915 -76.675 ;
        RECT -38.245 -78.365 -37.915 -78.035 ;
        RECT -38.245 -79.725 -37.915 -79.395 ;
        RECT -38.245 -81.085 -37.915 -80.755 ;
        RECT -38.245 -82.445 -37.915 -82.115 ;
        RECT -38.245 -83.805 -37.915 -83.475 ;
        RECT -38.245 -85.165 -37.915 -84.835 ;
        RECT -38.245 -86.525 -37.915 -86.195 ;
        RECT -38.245 -87.885 -37.915 -87.555 ;
        RECT -38.245 -89.245 -37.915 -88.915 ;
        RECT -38.245 -90.605 -37.915 -90.275 ;
        RECT -38.245 -91.77 -37.915 -91.44 ;
        RECT -38.245 -93.325 -37.915 -92.995 ;
        RECT -38.245 -94.685 -37.915 -94.355 ;
        RECT -38.245 -96.045 -37.915 -95.715 ;
        RECT -38.245 -97.405 -37.915 -97.075 ;
        RECT -38.245 -98.765 -37.915 -98.435 ;
        RECT -38.245 -101.485 -37.915 -101.155 ;
        RECT -38.245 -102.31 -37.915 -101.98 ;
        RECT -38.245 -104.205 -37.915 -103.875 ;
        RECT -38.245 -105.565 -37.915 -105.235 ;
        RECT -38.245 -106.925 -37.915 -106.595 ;
        RECT -38.245 -109.645 -37.915 -109.315 ;
        RECT -38.245 -111.005 -37.915 -110.675 ;
        RECT -38.24 -113.04 -37.92 245.285 ;
        RECT -38.245 244.04 -37.915 245.17 ;
        RECT -38.245 239.875 -37.915 240.205 ;
        RECT -38.245 238.515 -37.915 238.845 ;
        RECT -38.245 237.155 -37.915 237.485 ;
        RECT -38.245 235.795 -37.915 236.125 ;
        RECT -38.245 234.435 -37.915 234.765 ;
        RECT -38.245 233.075 -37.915 233.405 ;
        RECT -38.245 231.715 -37.915 232.045 ;
        RECT -38.245 230.355 -37.915 230.685 ;
        RECT -38.245 228.995 -37.915 229.325 ;
        RECT -38.245 227.635 -37.915 227.965 ;
        RECT -38.245 226.275 -37.915 226.605 ;
        RECT -38.245 224.915 -37.915 225.245 ;
        RECT -38.245 223.555 -37.915 223.885 ;
        RECT -38.245 222.195 -37.915 222.525 ;
        RECT -38.245 220.835 -37.915 221.165 ;
        RECT -38.245 219.475 -37.915 219.805 ;
        RECT -38.245 218.115 -37.915 218.445 ;
        RECT -38.245 216.755 -37.915 217.085 ;
        RECT -38.245 215.395 -37.915 215.725 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.765 -177.645 -47.435 -177.315 ;
        RECT -47.765 -179.005 -47.435 -178.675 ;
        RECT -47.765 -184.65 -47.435 -183.52 ;
        RECT -47.76 -184.765 -47.44 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.405 244.04 -46.075 245.17 ;
        RECT -46.405 239.875 -46.075 240.205 ;
        RECT -46.405 238.515 -46.075 238.845 ;
        RECT -46.405 237.155 -46.075 237.485 ;
        RECT -46.405 235.795 -46.075 236.125 ;
        RECT -46.405 234.435 -46.075 234.765 ;
        RECT -46.405 233.075 -46.075 233.405 ;
        RECT -46.405 231.715 -46.075 232.045 ;
        RECT -46.405 230.355 -46.075 230.685 ;
        RECT -46.405 228.995 -46.075 229.325 ;
        RECT -46.405 227.635 -46.075 227.965 ;
        RECT -46.405 226.275 -46.075 226.605 ;
        RECT -46.405 224.915 -46.075 225.245 ;
        RECT -46.405 223.555 -46.075 223.885 ;
        RECT -46.405 222.195 -46.075 222.525 ;
        RECT -46.405 220.835 -46.075 221.165 ;
        RECT -46.405 219.475 -46.075 219.805 ;
        RECT -46.405 218.115 -46.075 218.445 ;
        RECT -46.405 216.755 -46.075 217.085 ;
        RECT -46.405 215.395 -46.075 215.725 ;
        RECT -46.405 214.035 -46.075 214.365 ;
        RECT -46.405 212.675 -46.075 213.005 ;
        RECT -46.405 211.315 -46.075 211.645 ;
        RECT -46.405 209.955 -46.075 210.285 ;
        RECT -46.405 208.595 -46.075 208.925 ;
        RECT -46.405 207.235 -46.075 207.565 ;
        RECT -46.405 205.875 -46.075 206.205 ;
        RECT -46.405 204.515 -46.075 204.845 ;
        RECT -46.405 203.155 -46.075 203.485 ;
        RECT -46.405 201.795 -46.075 202.125 ;
        RECT -46.405 200.435 -46.075 200.765 ;
        RECT -46.405 199.075 -46.075 199.405 ;
        RECT -46.405 197.715 -46.075 198.045 ;
        RECT -46.405 196.355 -46.075 196.685 ;
        RECT -46.405 194.995 -46.075 195.325 ;
        RECT -46.405 193.635 -46.075 193.965 ;
        RECT -46.405 192.275 -46.075 192.605 ;
        RECT -46.405 190.915 -46.075 191.245 ;
        RECT -46.405 189.555 -46.075 189.885 ;
        RECT -46.405 188.195 -46.075 188.525 ;
        RECT -46.405 186.835 -46.075 187.165 ;
        RECT -46.405 185.475 -46.075 185.805 ;
        RECT -46.405 184.115 -46.075 184.445 ;
        RECT -46.405 182.755 -46.075 183.085 ;
        RECT -46.405 181.395 -46.075 181.725 ;
        RECT -46.405 180.035 -46.075 180.365 ;
        RECT -46.405 178.675 -46.075 179.005 ;
        RECT -46.405 177.315 -46.075 177.645 ;
        RECT -46.405 175.955 -46.075 176.285 ;
        RECT -46.405 174.595 -46.075 174.925 ;
        RECT -46.405 173.235 -46.075 173.565 ;
        RECT -46.405 171.875 -46.075 172.205 ;
        RECT -46.405 170.515 -46.075 170.845 ;
        RECT -46.405 169.155 -46.075 169.485 ;
        RECT -46.405 167.795 -46.075 168.125 ;
        RECT -46.405 166.435 -46.075 166.765 ;
        RECT -46.405 165.075 -46.075 165.405 ;
        RECT -46.405 163.715 -46.075 164.045 ;
        RECT -46.405 162.355 -46.075 162.685 ;
        RECT -46.405 160.995 -46.075 161.325 ;
        RECT -46.405 159.635 -46.075 159.965 ;
        RECT -46.405 158.275 -46.075 158.605 ;
        RECT -46.405 156.915 -46.075 157.245 ;
        RECT -46.405 155.555 -46.075 155.885 ;
        RECT -46.405 154.195 -46.075 154.525 ;
        RECT -46.405 152.835 -46.075 153.165 ;
        RECT -46.405 151.475 -46.075 151.805 ;
        RECT -46.405 150.115 -46.075 150.445 ;
        RECT -46.405 148.755 -46.075 149.085 ;
        RECT -46.405 147.395 -46.075 147.725 ;
        RECT -46.405 146.035 -46.075 146.365 ;
        RECT -46.405 144.675 -46.075 145.005 ;
        RECT -46.405 143.315 -46.075 143.645 ;
        RECT -46.405 141.955 -46.075 142.285 ;
        RECT -46.405 140.595 -46.075 140.925 ;
        RECT -46.405 139.235 -46.075 139.565 ;
        RECT -46.405 137.875 -46.075 138.205 ;
        RECT -46.405 136.515 -46.075 136.845 ;
        RECT -46.405 135.155 -46.075 135.485 ;
        RECT -46.405 133.795 -46.075 134.125 ;
        RECT -46.405 132.435 -46.075 132.765 ;
        RECT -46.405 131.075 -46.075 131.405 ;
        RECT -46.405 129.715 -46.075 130.045 ;
        RECT -46.405 128.355 -46.075 128.685 ;
        RECT -46.405 126.995 -46.075 127.325 ;
        RECT -46.405 125.635 -46.075 125.965 ;
        RECT -46.405 124.275 -46.075 124.605 ;
        RECT -46.405 122.915 -46.075 123.245 ;
        RECT -46.405 121.555 -46.075 121.885 ;
        RECT -46.405 120.195 -46.075 120.525 ;
        RECT -46.405 118.835 -46.075 119.165 ;
        RECT -46.405 117.475 -46.075 117.805 ;
        RECT -46.405 116.115 -46.075 116.445 ;
        RECT -46.405 114.755 -46.075 115.085 ;
        RECT -46.405 113.395 -46.075 113.725 ;
        RECT -46.405 112.035 -46.075 112.365 ;
        RECT -46.405 110.675 -46.075 111.005 ;
        RECT -46.405 109.315 -46.075 109.645 ;
        RECT -46.405 107.955 -46.075 108.285 ;
        RECT -46.405 106.595 -46.075 106.925 ;
        RECT -46.405 105.235 -46.075 105.565 ;
        RECT -46.405 103.875 -46.075 104.205 ;
        RECT -46.405 102.515 -46.075 102.845 ;
        RECT -46.405 101.155 -46.075 101.485 ;
        RECT -46.405 99.795 -46.075 100.125 ;
        RECT -46.405 98.435 -46.075 98.765 ;
        RECT -46.405 97.075 -46.075 97.405 ;
        RECT -46.405 95.715 -46.075 96.045 ;
        RECT -46.405 94.355 -46.075 94.685 ;
        RECT -46.405 92.995 -46.075 93.325 ;
        RECT -46.405 91.635 -46.075 91.965 ;
        RECT -46.405 90.275 -46.075 90.605 ;
        RECT -46.405 88.915 -46.075 89.245 ;
        RECT -46.405 87.555 -46.075 87.885 ;
        RECT -46.405 86.195 -46.075 86.525 ;
        RECT -46.405 84.835 -46.075 85.165 ;
        RECT -46.405 83.475 -46.075 83.805 ;
        RECT -46.405 82.115 -46.075 82.445 ;
        RECT -46.405 80.755 -46.075 81.085 ;
        RECT -46.405 79.395 -46.075 79.725 ;
        RECT -46.405 78.035 -46.075 78.365 ;
        RECT -46.405 76.675 -46.075 77.005 ;
        RECT -46.405 75.315 -46.075 75.645 ;
        RECT -46.405 73.955 -46.075 74.285 ;
        RECT -46.405 72.595 -46.075 72.925 ;
        RECT -46.405 71.235 -46.075 71.565 ;
        RECT -46.405 69.875 -46.075 70.205 ;
        RECT -46.405 68.515 -46.075 68.845 ;
        RECT -46.405 67.155 -46.075 67.485 ;
        RECT -46.405 65.795 -46.075 66.125 ;
        RECT -46.405 64.435 -46.075 64.765 ;
        RECT -46.405 63.075 -46.075 63.405 ;
        RECT -46.405 61.715 -46.075 62.045 ;
        RECT -46.405 60.355 -46.075 60.685 ;
        RECT -46.405 58.995 -46.075 59.325 ;
        RECT -46.405 57.635 -46.075 57.965 ;
        RECT -46.405 56.275 -46.075 56.605 ;
        RECT -46.405 54.915 -46.075 55.245 ;
        RECT -46.405 53.555 -46.075 53.885 ;
        RECT -46.405 52.195 -46.075 52.525 ;
        RECT -46.405 50.835 -46.075 51.165 ;
        RECT -46.405 49.475 -46.075 49.805 ;
        RECT -46.405 48.115 -46.075 48.445 ;
        RECT -46.405 46.755 -46.075 47.085 ;
        RECT -46.405 45.395 -46.075 45.725 ;
        RECT -46.405 44.035 -46.075 44.365 ;
        RECT -46.405 42.675 -46.075 43.005 ;
        RECT -46.405 41.315 -46.075 41.645 ;
        RECT -46.405 39.955 -46.075 40.285 ;
        RECT -46.405 38.595 -46.075 38.925 ;
        RECT -46.405 37.235 -46.075 37.565 ;
        RECT -46.405 35.875 -46.075 36.205 ;
        RECT -46.405 34.515 -46.075 34.845 ;
        RECT -46.405 33.155 -46.075 33.485 ;
        RECT -46.405 31.795 -46.075 32.125 ;
        RECT -46.405 30.435 -46.075 30.765 ;
        RECT -46.405 29.075 -46.075 29.405 ;
        RECT -46.405 27.715 -46.075 28.045 ;
        RECT -46.405 26.355 -46.075 26.685 ;
        RECT -46.405 24.995 -46.075 25.325 ;
        RECT -46.405 23.635 -46.075 23.965 ;
        RECT -46.405 22.275 -46.075 22.605 ;
        RECT -46.405 20.915 -46.075 21.245 ;
        RECT -46.405 19.555 -46.075 19.885 ;
        RECT -46.405 18.195 -46.075 18.525 ;
        RECT -46.405 16.835 -46.075 17.165 ;
        RECT -46.405 15.475 -46.075 15.805 ;
        RECT -46.405 14.115 -46.075 14.445 ;
        RECT -46.405 12.755 -46.075 13.085 ;
        RECT -46.405 11.395 -46.075 11.725 ;
        RECT -46.405 10.035 -46.075 10.365 ;
        RECT -46.405 8.675 -46.075 9.005 ;
        RECT -46.405 7.315 -46.075 7.645 ;
        RECT -46.405 5.955 -46.075 6.285 ;
        RECT -46.405 4.595 -46.075 4.925 ;
        RECT -46.405 3.235 -46.075 3.565 ;
        RECT -46.405 1.875 -46.075 2.205 ;
        RECT -46.405 0.515 -46.075 0.845 ;
        RECT -46.405 -0.845 -46.075 -0.515 ;
        RECT -46.4 -1.52 -46.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -46.405 -32.125 -46.075 -31.795 ;
        RECT -46.405 -33.71 -46.075 -33.38 ;
        RECT -46.405 -34.845 -46.075 -34.515 ;
        RECT -46.405 -36.205 -46.075 -35.875 ;
        RECT -46.405 -38.925 -46.075 -38.595 ;
        RECT -46.405 -39.75 -46.075 -39.42 ;
        RECT -46.405 -41.645 -46.075 -41.315 ;
        RECT -46.405 -44.365 -46.075 -44.035 ;
        RECT -46.405 -49.805 -46.075 -49.475 ;
        RECT -46.405 -51.165 -46.075 -50.835 ;
        RECT -46.405 -53.885 -46.075 -53.555 ;
        RECT -46.405 -55.245 -46.075 -54.915 ;
        RECT -46.405 -59.325 -46.075 -58.995 ;
        RECT -46.405 -60.685 -46.075 -60.355 ;
        RECT -46.405 -63.405 -46.075 -63.075 ;
        RECT -46.405 -70.205 -46.075 -69.875 ;
        RECT -46.405 -71.565 -46.075 -71.235 ;
        RECT -46.405 -72.925 -46.075 -72.595 ;
        RECT -46.405 -74.285 -46.075 -73.955 ;
        RECT -46.405 -75.645 -46.075 -75.315 ;
        RECT -46.405 -77.005 -46.075 -76.675 ;
        RECT -46.405 -78.365 -46.075 -78.035 ;
        RECT -46.405 -79.725 -46.075 -79.395 ;
        RECT -46.405 -81.085 -46.075 -80.755 ;
        RECT -46.405 -82.445 -46.075 -82.115 ;
        RECT -46.405 -83.805 -46.075 -83.475 ;
        RECT -46.405 -85.165 -46.075 -84.835 ;
        RECT -46.405 -86.525 -46.075 -86.195 ;
        RECT -46.405 -87.885 -46.075 -87.555 ;
        RECT -46.405 -89.245 -46.075 -88.915 ;
        RECT -46.405 -90.605 -46.075 -90.275 ;
        RECT -46.405 -91.77 -46.075 -91.44 ;
        RECT -46.405 -93.325 -46.075 -92.995 ;
        RECT -46.405 -94.685 -46.075 -94.355 ;
        RECT -46.405 -96.045 -46.075 -95.715 ;
        RECT -46.405 -97.405 -46.075 -97.075 ;
        RECT -46.405 -98.765 -46.075 -98.435 ;
        RECT -46.405 -101.485 -46.075 -101.155 ;
        RECT -46.405 -102.31 -46.075 -101.98 ;
        RECT -46.405 -104.205 -46.075 -103.875 ;
        RECT -46.405 -105.565 -46.075 -105.235 ;
        RECT -46.405 -106.925 -46.075 -106.595 ;
        RECT -46.405 -109.645 -46.075 -109.315 ;
        RECT -46.405 -111.005 -46.075 -110.675 ;
        RECT -46.405 -113.725 -46.075 -113.395 ;
        RECT -46.405 -115.085 -46.075 -114.755 ;
        RECT -46.405 -116.445 -46.075 -116.115 ;
        RECT -46.405 -117.805 -46.075 -117.475 ;
        RECT -46.405 -119.165 -46.075 -118.835 ;
        RECT -46.405 -120.525 -46.075 -120.195 ;
        RECT -46.405 -123.245 -46.075 -122.915 ;
        RECT -46.405 -124.605 -46.075 -124.275 ;
        RECT -46.405 -125.965 -46.075 -125.635 ;
        RECT -46.405 -127.325 -46.075 -126.995 ;
        RECT -46.405 -128.685 -46.075 -128.355 ;
        RECT -46.405 -130.045 -46.075 -129.715 ;
        RECT -46.405 -131.405 -46.075 -131.075 ;
        RECT -46.405 -132.765 -46.075 -132.435 ;
        RECT -46.405 -134.125 -46.075 -133.795 ;
        RECT -46.405 -135.485 -46.075 -135.155 ;
        RECT -46.405 -136.845 -46.075 -136.515 ;
        RECT -46.405 -138.205 -46.075 -137.875 ;
        RECT -46.405 -139.565 -46.075 -139.235 ;
        RECT -46.405 -140.925 -46.075 -140.595 ;
        RECT -46.405 -142.285 -46.075 -141.955 ;
        RECT -46.405 -143.645 -46.075 -143.315 ;
        RECT -46.405 -145.005 -46.075 -144.675 ;
        RECT -46.405 -146.365 -46.075 -146.035 ;
        RECT -46.405 -147.725 -46.075 -147.395 ;
        RECT -46.405 -149.085 -46.075 -148.755 ;
        RECT -46.405 -150.445 -46.075 -150.115 ;
        RECT -46.405 -151.805 -46.075 -151.475 ;
        RECT -46.405 -153.165 -46.075 -152.835 ;
        RECT -46.405 -154.525 -46.075 -154.195 ;
        RECT -46.405 -155.885 -46.075 -155.555 ;
        RECT -46.405 -157.245 -46.075 -156.915 ;
        RECT -46.405 -158.605 -46.075 -158.275 ;
        RECT -46.405 -159.965 -46.075 -159.635 ;
        RECT -46.405 -161.325 -46.075 -160.995 ;
        RECT -46.405 -162.685 -46.075 -162.355 ;
        RECT -46.405 -164.045 -46.075 -163.715 ;
        RECT -46.405 -165.405 -46.075 -165.075 ;
        RECT -46.405 -166.765 -46.075 -166.435 ;
        RECT -46.405 -169.615 -46.075 -169.285 ;
        RECT -46.405 -170.845 -46.075 -170.515 ;
        RECT -46.405 -172.205 -46.075 -171.875 ;
        RECT -46.4 -172.88 -46.08 -30.44 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.045 244.04 -44.715 245.17 ;
        RECT -45.045 239.875 -44.715 240.205 ;
        RECT -45.045 238.515 -44.715 238.845 ;
        RECT -45.045 237.155 -44.715 237.485 ;
        RECT -45.045 235.795 -44.715 236.125 ;
        RECT -45.045 234.435 -44.715 234.765 ;
        RECT -45.045 233.075 -44.715 233.405 ;
        RECT -45.045 231.715 -44.715 232.045 ;
        RECT -45.045 230.355 -44.715 230.685 ;
        RECT -45.045 228.995 -44.715 229.325 ;
        RECT -45.045 227.635 -44.715 227.965 ;
        RECT -45.045 226.275 -44.715 226.605 ;
        RECT -45.045 224.915 -44.715 225.245 ;
        RECT -45.045 223.555 -44.715 223.885 ;
        RECT -45.045 222.195 -44.715 222.525 ;
        RECT -45.045 220.835 -44.715 221.165 ;
        RECT -45.045 219.475 -44.715 219.805 ;
        RECT -45.045 218.115 -44.715 218.445 ;
        RECT -45.045 216.755 -44.715 217.085 ;
        RECT -45.045 215.395 -44.715 215.725 ;
        RECT -45.045 214.035 -44.715 214.365 ;
        RECT -45.045 212.675 -44.715 213.005 ;
        RECT -45.045 211.315 -44.715 211.645 ;
        RECT -45.045 209.955 -44.715 210.285 ;
        RECT -45.045 208.595 -44.715 208.925 ;
        RECT -45.045 207.235 -44.715 207.565 ;
        RECT -45.045 205.875 -44.715 206.205 ;
        RECT -45.045 204.515 -44.715 204.845 ;
        RECT -45.045 203.155 -44.715 203.485 ;
        RECT -45.045 201.795 -44.715 202.125 ;
        RECT -45.045 200.435 -44.715 200.765 ;
        RECT -45.045 199.075 -44.715 199.405 ;
        RECT -45.045 197.715 -44.715 198.045 ;
        RECT -45.045 196.355 -44.715 196.685 ;
        RECT -45.045 194.995 -44.715 195.325 ;
        RECT -45.045 193.635 -44.715 193.965 ;
        RECT -45.045 192.275 -44.715 192.605 ;
        RECT -45.045 190.915 -44.715 191.245 ;
        RECT -45.045 189.555 -44.715 189.885 ;
        RECT -45.045 188.195 -44.715 188.525 ;
        RECT -45.045 186.835 -44.715 187.165 ;
        RECT -45.045 185.475 -44.715 185.805 ;
        RECT -45.045 184.115 -44.715 184.445 ;
        RECT -45.045 182.755 -44.715 183.085 ;
        RECT -45.045 181.395 -44.715 181.725 ;
        RECT -45.045 180.035 -44.715 180.365 ;
        RECT -45.045 178.675 -44.715 179.005 ;
        RECT -45.045 177.315 -44.715 177.645 ;
        RECT -45.045 175.955 -44.715 176.285 ;
        RECT -45.045 174.595 -44.715 174.925 ;
        RECT -45.045 173.235 -44.715 173.565 ;
        RECT -45.045 171.875 -44.715 172.205 ;
        RECT -45.045 170.515 -44.715 170.845 ;
        RECT -45.045 169.155 -44.715 169.485 ;
        RECT -45.045 167.795 -44.715 168.125 ;
        RECT -45.045 166.435 -44.715 166.765 ;
        RECT -45.045 165.075 -44.715 165.405 ;
        RECT -45.045 163.715 -44.715 164.045 ;
        RECT -45.045 162.355 -44.715 162.685 ;
        RECT -45.045 160.995 -44.715 161.325 ;
        RECT -45.045 159.635 -44.715 159.965 ;
        RECT -45.045 158.275 -44.715 158.605 ;
        RECT -45.045 156.915 -44.715 157.245 ;
        RECT -45.045 155.555 -44.715 155.885 ;
        RECT -45.045 154.195 -44.715 154.525 ;
        RECT -45.045 152.835 -44.715 153.165 ;
        RECT -45.045 151.475 -44.715 151.805 ;
        RECT -45.045 150.115 -44.715 150.445 ;
        RECT -45.045 148.755 -44.715 149.085 ;
        RECT -45.045 147.395 -44.715 147.725 ;
        RECT -45.045 146.035 -44.715 146.365 ;
        RECT -45.045 144.675 -44.715 145.005 ;
        RECT -45.045 143.315 -44.715 143.645 ;
        RECT -45.045 141.955 -44.715 142.285 ;
        RECT -45.045 140.595 -44.715 140.925 ;
        RECT -45.045 139.235 -44.715 139.565 ;
        RECT -45.045 137.875 -44.715 138.205 ;
        RECT -45.045 136.515 -44.715 136.845 ;
        RECT -45.045 135.155 -44.715 135.485 ;
        RECT -45.045 133.795 -44.715 134.125 ;
        RECT -45.045 132.435 -44.715 132.765 ;
        RECT -45.045 131.075 -44.715 131.405 ;
        RECT -45.045 129.715 -44.715 130.045 ;
        RECT -45.045 128.355 -44.715 128.685 ;
        RECT -45.045 126.995 -44.715 127.325 ;
        RECT -45.045 125.635 -44.715 125.965 ;
        RECT -45.045 124.275 -44.715 124.605 ;
        RECT -45.045 122.915 -44.715 123.245 ;
        RECT -45.045 121.555 -44.715 121.885 ;
        RECT -45.045 120.195 -44.715 120.525 ;
        RECT -45.045 118.835 -44.715 119.165 ;
        RECT -45.045 117.475 -44.715 117.805 ;
        RECT -45.045 116.115 -44.715 116.445 ;
        RECT -45.045 114.755 -44.715 115.085 ;
        RECT -45.045 113.395 -44.715 113.725 ;
        RECT -45.045 112.035 -44.715 112.365 ;
        RECT -45.045 110.675 -44.715 111.005 ;
        RECT -45.045 109.315 -44.715 109.645 ;
        RECT -45.045 107.955 -44.715 108.285 ;
        RECT -45.045 106.595 -44.715 106.925 ;
        RECT -45.045 105.235 -44.715 105.565 ;
        RECT -45.045 103.875 -44.715 104.205 ;
        RECT -45.045 102.515 -44.715 102.845 ;
        RECT -45.045 101.155 -44.715 101.485 ;
        RECT -45.045 99.795 -44.715 100.125 ;
        RECT -45.045 98.435 -44.715 98.765 ;
        RECT -45.045 97.075 -44.715 97.405 ;
        RECT -45.045 95.715 -44.715 96.045 ;
        RECT -45.045 94.355 -44.715 94.685 ;
        RECT -45.045 92.995 -44.715 93.325 ;
        RECT -45.045 91.635 -44.715 91.965 ;
        RECT -45.045 90.275 -44.715 90.605 ;
        RECT -45.045 88.915 -44.715 89.245 ;
        RECT -45.045 87.555 -44.715 87.885 ;
        RECT -45.045 86.195 -44.715 86.525 ;
        RECT -45.045 84.835 -44.715 85.165 ;
        RECT -45.045 83.475 -44.715 83.805 ;
        RECT -45.045 82.115 -44.715 82.445 ;
        RECT -45.045 80.755 -44.715 81.085 ;
        RECT -45.045 79.395 -44.715 79.725 ;
        RECT -45.045 78.035 -44.715 78.365 ;
        RECT -45.045 76.675 -44.715 77.005 ;
        RECT -45.045 75.315 -44.715 75.645 ;
        RECT -45.045 73.955 -44.715 74.285 ;
        RECT -45.045 72.595 -44.715 72.925 ;
        RECT -45.045 71.235 -44.715 71.565 ;
        RECT -45.045 69.875 -44.715 70.205 ;
        RECT -45.045 68.515 -44.715 68.845 ;
        RECT -45.045 67.155 -44.715 67.485 ;
        RECT -45.045 65.795 -44.715 66.125 ;
        RECT -45.045 64.435 -44.715 64.765 ;
        RECT -45.045 63.075 -44.715 63.405 ;
        RECT -45.045 61.715 -44.715 62.045 ;
        RECT -45.045 60.355 -44.715 60.685 ;
        RECT -45.045 58.995 -44.715 59.325 ;
        RECT -45.045 57.635 -44.715 57.965 ;
        RECT -45.045 56.275 -44.715 56.605 ;
        RECT -45.045 54.915 -44.715 55.245 ;
        RECT -45.045 53.555 -44.715 53.885 ;
        RECT -45.045 52.195 -44.715 52.525 ;
        RECT -45.045 50.835 -44.715 51.165 ;
        RECT -45.045 49.475 -44.715 49.805 ;
        RECT -45.045 48.115 -44.715 48.445 ;
        RECT -45.045 46.755 -44.715 47.085 ;
        RECT -45.045 45.395 -44.715 45.725 ;
        RECT -45.045 44.035 -44.715 44.365 ;
        RECT -45.045 42.675 -44.715 43.005 ;
        RECT -45.045 41.315 -44.715 41.645 ;
        RECT -45.045 39.955 -44.715 40.285 ;
        RECT -45.045 38.595 -44.715 38.925 ;
        RECT -45.045 37.235 -44.715 37.565 ;
        RECT -45.045 35.875 -44.715 36.205 ;
        RECT -45.045 34.515 -44.715 34.845 ;
        RECT -45.045 33.155 -44.715 33.485 ;
        RECT -45.045 31.795 -44.715 32.125 ;
        RECT -45.045 30.435 -44.715 30.765 ;
        RECT -45.045 29.075 -44.715 29.405 ;
        RECT -45.045 27.715 -44.715 28.045 ;
        RECT -45.045 26.355 -44.715 26.685 ;
        RECT -45.045 24.995 -44.715 25.325 ;
        RECT -45.045 23.635 -44.715 23.965 ;
        RECT -45.045 22.275 -44.715 22.605 ;
        RECT -45.045 20.915 -44.715 21.245 ;
        RECT -45.045 19.555 -44.715 19.885 ;
        RECT -45.045 18.195 -44.715 18.525 ;
        RECT -45.045 16.835 -44.715 17.165 ;
        RECT -45.045 15.475 -44.715 15.805 ;
        RECT -45.045 14.115 -44.715 14.445 ;
        RECT -45.045 12.755 -44.715 13.085 ;
        RECT -45.045 11.395 -44.715 11.725 ;
        RECT -45.045 10.035 -44.715 10.365 ;
        RECT -45.045 8.675 -44.715 9.005 ;
        RECT -45.045 7.315 -44.715 7.645 ;
        RECT -45.045 5.955 -44.715 6.285 ;
        RECT -45.045 4.595 -44.715 4.925 ;
        RECT -45.045 3.235 -44.715 3.565 ;
        RECT -45.045 1.875 -44.715 2.205 ;
        RECT -45.045 0.515 -44.715 0.845 ;
        RECT -45.045 -0.845 -44.715 -0.515 ;
        RECT -45.045 -2.205 -44.715 -1.875 ;
        RECT -45.045 -4.925 -44.715 -4.595 ;
        RECT -45.045 -6.285 -44.715 -5.955 ;
        RECT -45.045 -7.645 -44.715 -7.315 ;
        RECT -45.045 -10.365 -44.715 -10.035 ;
        RECT -45.045 -14.445 -44.715 -14.115 ;
        RECT -45.045 -17.165 -44.715 -16.835 ;
        RECT -45.045 -18.525 -44.715 -18.195 ;
        RECT -45.045 -19.885 -44.715 -19.555 ;
        RECT -45.045 -21.245 -44.715 -20.915 ;
        RECT -45.045 -22.605 -44.715 -22.275 ;
        RECT -45.045 -23.965 -44.715 -23.635 ;
        RECT -45.045 -25.325 -44.715 -24.995 ;
        RECT -45.045 -32.125 -44.715 -31.795 ;
        RECT -45.045 -33.71 -44.715 -33.38 ;
        RECT -45.045 -34.845 -44.715 -34.515 ;
        RECT -45.045 -36.205 -44.715 -35.875 ;
        RECT -45.045 -38.925 -44.715 -38.595 ;
        RECT -45.045 -39.75 -44.715 -39.42 ;
        RECT -45.045 -41.645 -44.715 -41.315 ;
        RECT -45.045 -44.365 -44.715 -44.035 ;
        RECT -45.045 -49.805 -44.715 -49.475 ;
        RECT -45.045 -51.165 -44.715 -50.835 ;
        RECT -45.045 -53.885 -44.715 -53.555 ;
        RECT -45.045 -55.245 -44.715 -54.915 ;
        RECT -45.045 -59.325 -44.715 -58.995 ;
        RECT -45.045 -60.685 -44.715 -60.355 ;
        RECT -45.045 -63.405 -44.715 -63.075 ;
        RECT -45.04 -64.76 -44.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.045 -70.205 -44.715 -69.875 ;
        RECT -45.045 -71.565 -44.715 -71.235 ;
        RECT -45.045 -72.925 -44.715 -72.595 ;
        RECT -45.045 -74.285 -44.715 -73.955 ;
        RECT -45.045 -75.645 -44.715 -75.315 ;
        RECT -45.045 -77.005 -44.715 -76.675 ;
        RECT -45.045 -78.365 -44.715 -78.035 ;
        RECT -45.045 -79.725 -44.715 -79.395 ;
        RECT -45.045 -81.085 -44.715 -80.755 ;
        RECT -45.045 -82.445 -44.715 -82.115 ;
        RECT -45.045 -83.805 -44.715 -83.475 ;
        RECT -45.045 -85.165 -44.715 -84.835 ;
        RECT -45.045 -86.525 -44.715 -86.195 ;
        RECT -45.045 -87.885 -44.715 -87.555 ;
        RECT -45.045 -89.245 -44.715 -88.915 ;
        RECT -45.045 -90.605 -44.715 -90.275 ;
        RECT -45.045 -91.77 -44.715 -91.44 ;
        RECT -45.045 -93.325 -44.715 -92.995 ;
        RECT -45.045 -94.685 -44.715 -94.355 ;
        RECT -45.045 -96.045 -44.715 -95.715 ;
        RECT -45.045 -97.405 -44.715 -97.075 ;
        RECT -45.045 -98.765 -44.715 -98.435 ;
        RECT -45.045 -101.485 -44.715 -101.155 ;
        RECT -45.045 -102.31 -44.715 -101.98 ;
        RECT -45.045 -104.205 -44.715 -103.875 ;
        RECT -45.045 -105.565 -44.715 -105.235 ;
        RECT -45.045 -106.925 -44.715 -106.595 ;
        RECT -45.045 -109.645 -44.715 -109.315 ;
        RECT -45.045 -111.005 -44.715 -110.675 ;
        RECT -45.045 -113.725 -44.715 -113.395 ;
        RECT -45.045 -115.085 -44.715 -114.755 ;
        RECT -45.045 -116.445 -44.715 -116.115 ;
        RECT -45.045 -117.805 -44.715 -117.475 ;
        RECT -45.045 -119.165 -44.715 -118.835 ;
        RECT -45.045 -120.525 -44.715 -120.195 ;
        RECT -45.045 -123.245 -44.715 -122.915 ;
        RECT -45.045 -124.605 -44.715 -124.275 ;
        RECT -45.045 -125.965 -44.715 -125.635 ;
        RECT -45.045 -127.325 -44.715 -126.995 ;
        RECT -45.045 -128.685 -44.715 -128.355 ;
        RECT -45.045 -130.045 -44.715 -129.715 ;
        RECT -45.045 -131.405 -44.715 -131.075 ;
        RECT -45.045 -132.765 -44.715 -132.435 ;
        RECT -45.045 -134.125 -44.715 -133.795 ;
        RECT -45.045 -135.485 -44.715 -135.155 ;
        RECT -45.045 -136.845 -44.715 -136.515 ;
        RECT -45.045 -138.205 -44.715 -137.875 ;
        RECT -45.045 -139.565 -44.715 -139.235 ;
        RECT -45.045 -140.925 -44.715 -140.595 ;
        RECT -45.045 -142.285 -44.715 -141.955 ;
        RECT -45.045 -143.645 -44.715 -143.315 ;
        RECT -45.045 -145.005 -44.715 -144.675 ;
        RECT -45.045 -146.365 -44.715 -146.035 ;
        RECT -45.045 -147.725 -44.715 -147.395 ;
        RECT -45.045 -149.085 -44.715 -148.755 ;
        RECT -45.045 -150.445 -44.715 -150.115 ;
        RECT -45.045 -151.805 -44.715 -151.475 ;
        RECT -45.045 -153.165 -44.715 -152.835 ;
        RECT -45.045 -154.525 -44.715 -154.195 ;
        RECT -45.045 -155.885 -44.715 -155.555 ;
        RECT -45.045 -157.245 -44.715 -156.915 ;
        RECT -45.045 -158.605 -44.715 -158.275 ;
        RECT -45.045 -159.965 -44.715 -159.635 ;
        RECT -45.045 -161.325 -44.715 -160.995 ;
        RECT -45.045 -162.685 -44.715 -162.355 ;
        RECT -45.045 -164.045 -44.715 -163.715 ;
        RECT -45.045 -165.405 -44.715 -165.075 ;
        RECT -45.045 -166.765 -44.715 -166.435 ;
        RECT -45.04 -167.44 -44.72 -69.2 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.045 -174.925 -44.715 -174.595 ;
        RECT -45.045 -177.645 -44.715 -177.315 ;
        RECT -45.045 -179.005 -44.715 -178.675 ;
        RECT -45.045 -184.65 -44.715 -183.52 ;
        RECT -45.04 -184.765 -44.72 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.685 244.04 -43.355 245.17 ;
        RECT -43.685 239.875 -43.355 240.205 ;
        RECT -43.685 238.515 -43.355 238.845 ;
        RECT -43.685 237.155 -43.355 237.485 ;
        RECT -43.685 235.795 -43.355 236.125 ;
        RECT -43.685 234.435 -43.355 234.765 ;
        RECT -43.685 233.075 -43.355 233.405 ;
        RECT -43.685 231.715 -43.355 232.045 ;
        RECT -43.685 230.355 -43.355 230.685 ;
        RECT -43.685 228.995 -43.355 229.325 ;
        RECT -43.685 227.635 -43.355 227.965 ;
        RECT -43.685 226.275 -43.355 226.605 ;
        RECT -43.685 224.915 -43.355 225.245 ;
        RECT -43.685 223.555 -43.355 223.885 ;
        RECT -43.685 222.195 -43.355 222.525 ;
        RECT -43.685 220.835 -43.355 221.165 ;
        RECT -43.685 219.475 -43.355 219.805 ;
        RECT -43.685 218.115 -43.355 218.445 ;
        RECT -43.685 216.755 -43.355 217.085 ;
        RECT -43.685 215.395 -43.355 215.725 ;
        RECT -43.685 214.035 -43.355 214.365 ;
        RECT -43.685 212.675 -43.355 213.005 ;
        RECT -43.685 211.315 -43.355 211.645 ;
        RECT -43.685 209.955 -43.355 210.285 ;
        RECT -43.685 208.595 -43.355 208.925 ;
        RECT -43.685 207.235 -43.355 207.565 ;
        RECT -43.685 205.875 -43.355 206.205 ;
        RECT -43.685 204.515 -43.355 204.845 ;
        RECT -43.685 203.155 -43.355 203.485 ;
        RECT -43.685 201.795 -43.355 202.125 ;
        RECT -43.685 200.435 -43.355 200.765 ;
        RECT -43.685 199.075 -43.355 199.405 ;
        RECT -43.685 197.715 -43.355 198.045 ;
        RECT -43.685 196.355 -43.355 196.685 ;
        RECT -43.685 194.995 -43.355 195.325 ;
        RECT -43.685 193.635 -43.355 193.965 ;
        RECT -43.685 192.275 -43.355 192.605 ;
        RECT -43.685 190.915 -43.355 191.245 ;
        RECT -43.685 189.555 -43.355 189.885 ;
        RECT -43.685 188.195 -43.355 188.525 ;
        RECT -43.685 186.835 -43.355 187.165 ;
        RECT -43.685 185.475 -43.355 185.805 ;
        RECT -43.685 184.115 -43.355 184.445 ;
        RECT -43.685 182.755 -43.355 183.085 ;
        RECT -43.685 181.395 -43.355 181.725 ;
        RECT -43.685 180.035 -43.355 180.365 ;
        RECT -43.685 178.675 -43.355 179.005 ;
        RECT -43.685 177.315 -43.355 177.645 ;
        RECT -43.685 175.955 -43.355 176.285 ;
        RECT -43.685 174.595 -43.355 174.925 ;
        RECT -43.685 173.235 -43.355 173.565 ;
        RECT -43.685 171.875 -43.355 172.205 ;
        RECT -43.685 170.515 -43.355 170.845 ;
        RECT -43.685 169.155 -43.355 169.485 ;
        RECT -43.685 167.795 -43.355 168.125 ;
        RECT -43.685 166.435 -43.355 166.765 ;
        RECT -43.685 165.075 -43.355 165.405 ;
        RECT -43.685 163.715 -43.355 164.045 ;
        RECT -43.685 162.355 -43.355 162.685 ;
        RECT -43.685 160.995 -43.355 161.325 ;
        RECT -43.685 159.635 -43.355 159.965 ;
        RECT -43.685 158.275 -43.355 158.605 ;
        RECT -43.685 156.915 -43.355 157.245 ;
        RECT -43.685 155.555 -43.355 155.885 ;
        RECT -43.685 154.195 -43.355 154.525 ;
        RECT -43.685 152.835 -43.355 153.165 ;
        RECT -43.685 151.475 -43.355 151.805 ;
        RECT -43.685 150.115 -43.355 150.445 ;
        RECT -43.685 148.755 -43.355 149.085 ;
        RECT -43.685 147.395 -43.355 147.725 ;
        RECT -43.685 146.035 -43.355 146.365 ;
        RECT -43.685 144.675 -43.355 145.005 ;
        RECT -43.685 143.315 -43.355 143.645 ;
        RECT -43.685 141.955 -43.355 142.285 ;
        RECT -43.685 140.595 -43.355 140.925 ;
        RECT -43.685 139.235 -43.355 139.565 ;
        RECT -43.685 137.875 -43.355 138.205 ;
        RECT -43.685 136.515 -43.355 136.845 ;
        RECT -43.685 135.155 -43.355 135.485 ;
        RECT -43.685 133.795 -43.355 134.125 ;
        RECT -43.685 132.435 -43.355 132.765 ;
        RECT -43.685 131.075 -43.355 131.405 ;
        RECT -43.685 129.715 -43.355 130.045 ;
        RECT -43.685 128.355 -43.355 128.685 ;
        RECT -43.685 126.995 -43.355 127.325 ;
        RECT -43.685 125.635 -43.355 125.965 ;
        RECT -43.685 124.275 -43.355 124.605 ;
        RECT -43.685 122.915 -43.355 123.245 ;
        RECT -43.685 121.555 -43.355 121.885 ;
        RECT -43.685 120.195 -43.355 120.525 ;
        RECT -43.685 118.835 -43.355 119.165 ;
        RECT -43.685 117.475 -43.355 117.805 ;
        RECT -43.685 116.115 -43.355 116.445 ;
        RECT -43.685 114.755 -43.355 115.085 ;
        RECT -43.685 113.395 -43.355 113.725 ;
        RECT -43.685 112.035 -43.355 112.365 ;
        RECT -43.685 110.675 -43.355 111.005 ;
        RECT -43.685 109.315 -43.355 109.645 ;
        RECT -43.685 107.955 -43.355 108.285 ;
        RECT -43.685 106.595 -43.355 106.925 ;
        RECT -43.685 105.235 -43.355 105.565 ;
        RECT -43.685 103.875 -43.355 104.205 ;
        RECT -43.685 102.515 -43.355 102.845 ;
        RECT -43.685 101.155 -43.355 101.485 ;
        RECT -43.685 99.795 -43.355 100.125 ;
        RECT -43.685 98.435 -43.355 98.765 ;
        RECT -43.685 97.075 -43.355 97.405 ;
        RECT -43.685 95.715 -43.355 96.045 ;
        RECT -43.685 94.355 -43.355 94.685 ;
        RECT -43.685 92.995 -43.355 93.325 ;
        RECT -43.685 91.635 -43.355 91.965 ;
        RECT -43.685 90.275 -43.355 90.605 ;
        RECT -43.685 88.915 -43.355 89.245 ;
        RECT -43.685 87.555 -43.355 87.885 ;
        RECT -43.685 86.195 -43.355 86.525 ;
        RECT -43.685 84.835 -43.355 85.165 ;
        RECT -43.685 83.475 -43.355 83.805 ;
        RECT -43.685 82.115 -43.355 82.445 ;
        RECT -43.685 80.755 -43.355 81.085 ;
        RECT -43.685 79.395 -43.355 79.725 ;
        RECT -43.685 78.035 -43.355 78.365 ;
        RECT -43.685 76.675 -43.355 77.005 ;
        RECT -43.685 75.315 -43.355 75.645 ;
        RECT -43.685 73.955 -43.355 74.285 ;
        RECT -43.685 72.595 -43.355 72.925 ;
        RECT -43.685 71.235 -43.355 71.565 ;
        RECT -43.685 69.875 -43.355 70.205 ;
        RECT -43.685 68.515 -43.355 68.845 ;
        RECT -43.685 67.155 -43.355 67.485 ;
        RECT -43.685 65.795 -43.355 66.125 ;
        RECT -43.685 64.435 -43.355 64.765 ;
        RECT -43.685 63.075 -43.355 63.405 ;
        RECT -43.685 61.715 -43.355 62.045 ;
        RECT -43.685 60.355 -43.355 60.685 ;
        RECT -43.685 58.995 -43.355 59.325 ;
        RECT -43.685 57.635 -43.355 57.965 ;
        RECT -43.685 56.275 -43.355 56.605 ;
        RECT -43.685 54.915 -43.355 55.245 ;
        RECT -43.685 53.555 -43.355 53.885 ;
        RECT -43.685 52.195 -43.355 52.525 ;
        RECT -43.685 50.835 -43.355 51.165 ;
        RECT -43.685 49.475 -43.355 49.805 ;
        RECT -43.685 48.115 -43.355 48.445 ;
        RECT -43.685 46.755 -43.355 47.085 ;
        RECT -43.685 45.395 -43.355 45.725 ;
        RECT -43.685 44.035 -43.355 44.365 ;
        RECT -43.685 42.675 -43.355 43.005 ;
        RECT -43.685 41.315 -43.355 41.645 ;
        RECT -43.685 39.955 -43.355 40.285 ;
        RECT -43.685 38.595 -43.355 38.925 ;
        RECT -43.685 37.235 -43.355 37.565 ;
        RECT -43.685 35.875 -43.355 36.205 ;
        RECT -43.685 34.515 -43.355 34.845 ;
        RECT -43.685 33.155 -43.355 33.485 ;
        RECT -43.685 31.795 -43.355 32.125 ;
        RECT -43.685 30.435 -43.355 30.765 ;
        RECT -43.685 29.075 -43.355 29.405 ;
        RECT -43.685 27.715 -43.355 28.045 ;
        RECT -43.685 26.355 -43.355 26.685 ;
        RECT -43.685 24.995 -43.355 25.325 ;
        RECT -43.685 23.635 -43.355 23.965 ;
        RECT -43.685 22.275 -43.355 22.605 ;
        RECT -43.685 20.915 -43.355 21.245 ;
        RECT -43.685 19.555 -43.355 19.885 ;
        RECT -43.685 18.195 -43.355 18.525 ;
        RECT -43.685 16.835 -43.355 17.165 ;
        RECT -43.685 15.475 -43.355 15.805 ;
        RECT -43.685 14.115 -43.355 14.445 ;
        RECT -43.685 12.755 -43.355 13.085 ;
        RECT -43.685 11.395 -43.355 11.725 ;
        RECT -43.685 10.035 -43.355 10.365 ;
        RECT -43.685 8.675 -43.355 9.005 ;
        RECT -43.685 7.315 -43.355 7.645 ;
        RECT -43.685 5.955 -43.355 6.285 ;
        RECT -43.685 4.595 -43.355 4.925 ;
        RECT -43.685 3.235 -43.355 3.565 ;
        RECT -43.685 1.875 -43.355 2.205 ;
        RECT -43.685 0.515 -43.355 0.845 ;
        RECT -43.685 -0.845 -43.355 -0.515 ;
        RECT -43.685 -2.205 -43.355 -1.875 ;
        RECT -43.685 -4.925 -43.355 -4.595 ;
        RECT -43.685 -6.285 -43.355 -5.955 ;
        RECT -43.685 -10.365 -43.355 -10.035 ;
        RECT -43.685 -14.445 -43.355 -14.115 ;
        RECT -43.685 -17.165 -43.355 -16.835 ;
        RECT -43.685 -18.525 -43.355 -18.195 ;
        RECT -43.685 -19.885 -43.355 -19.555 ;
        RECT -43.685 -21.245 -43.355 -20.915 ;
        RECT -43.685 -22.605 -43.355 -22.275 ;
        RECT -43.685 -23.965 -43.355 -23.635 ;
        RECT -43.685 -25.325 -43.355 -24.995 ;
        RECT -43.685 -32.125 -43.355 -31.795 ;
        RECT -43.685 -33.71 -43.355 -33.38 ;
        RECT -43.685 -34.845 -43.355 -34.515 ;
        RECT -43.685 -36.205 -43.355 -35.875 ;
        RECT -43.685 -38.925 -43.355 -38.595 ;
        RECT -43.685 -39.75 -43.355 -39.42 ;
        RECT -43.685 -41.645 -43.355 -41.315 ;
        RECT -43.685 -44.365 -43.355 -44.035 ;
        RECT -43.685 -49.805 -43.355 -49.475 ;
        RECT -43.685 -51.165 -43.355 -50.835 ;
        RECT -43.685 -53.885 -43.355 -53.555 ;
        RECT -43.685 -55.245 -43.355 -54.915 ;
        RECT -43.685 -59.325 -43.355 -58.995 ;
        RECT -43.685 -60.685 -43.355 -60.355 ;
        RECT -43.685 -63.405 -43.355 -63.075 ;
        RECT -43.68 -64.08 -43.36 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.685 -70.205 -43.355 -69.875 ;
        RECT -43.685 -71.565 -43.355 -71.235 ;
        RECT -43.685 -72.925 -43.355 -72.595 ;
        RECT -43.685 -74.285 -43.355 -73.955 ;
        RECT -43.685 -75.645 -43.355 -75.315 ;
        RECT -43.685 -77.005 -43.355 -76.675 ;
        RECT -43.685 -78.365 -43.355 -78.035 ;
        RECT -43.685 -79.725 -43.355 -79.395 ;
        RECT -43.685 -81.085 -43.355 -80.755 ;
        RECT -43.685 -82.445 -43.355 -82.115 ;
        RECT -43.685 -83.805 -43.355 -83.475 ;
        RECT -43.685 -85.165 -43.355 -84.835 ;
        RECT -43.685 -86.525 -43.355 -86.195 ;
        RECT -43.685 -87.885 -43.355 -87.555 ;
        RECT -43.685 -89.245 -43.355 -88.915 ;
        RECT -43.685 -90.605 -43.355 -90.275 ;
        RECT -43.685 -91.77 -43.355 -91.44 ;
        RECT -43.685 -93.325 -43.355 -92.995 ;
        RECT -43.685 -94.685 -43.355 -94.355 ;
        RECT -43.685 -96.045 -43.355 -95.715 ;
        RECT -43.685 -97.405 -43.355 -97.075 ;
        RECT -43.685 -98.765 -43.355 -98.435 ;
        RECT -43.685 -101.485 -43.355 -101.155 ;
        RECT -43.685 -102.31 -43.355 -101.98 ;
        RECT -43.685 -104.205 -43.355 -103.875 ;
        RECT -43.685 -105.565 -43.355 -105.235 ;
        RECT -43.685 -106.925 -43.355 -106.595 ;
        RECT -43.685 -109.645 -43.355 -109.315 ;
        RECT -43.685 -111.005 -43.355 -110.675 ;
        RECT -43.68 -113.04 -43.36 -67.84 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.685 -177.645 -43.355 -177.315 ;
        RECT -43.685 -179.005 -43.355 -178.675 ;
        RECT -43.685 -184.65 -43.355 -183.52 ;
        RECT -43.68 -184.765 -43.36 -175.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -42.325 -87.885 -41.995 -87.555 ;
        RECT -42.325 -89.245 -41.995 -88.915 ;
        RECT -42.325 -90.605 -41.995 -90.275 ;
        RECT -42.325 -91.77 -41.995 -91.44 ;
        RECT -42.325 -93.325 -41.995 -92.995 ;
        RECT -42.325 -94.685 -41.995 -94.355 ;
        RECT -42.325 -96.045 -41.995 -95.715 ;
        RECT -42.325 -97.405 -41.995 -97.075 ;
        RECT -42.325 -98.765 -41.995 -98.435 ;
        RECT -42.325 -101.485 -41.995 -101.155 ;
        RECT -42.325 -102.31 -41.995 -101.98 ;
        RECT -42.325 -104.205 -41.995 -103.875 ;
        RECT -42.325 -105.565 -41.995 -105.235 ;
        RECT -42.325 -106.925 -41.995 -106.595 ;
        RECT -42.325 -109.645 -41.995 -109.315 ;
        RECT -42.325 -111.005 -41.995 -110.675 ;
        RECT -42.325 -113.725 -41.995 -113.395 ;
        RECT -42.325 -115.085 -41.995 -114.755 ;
        RECT -42.325 -116.445 -41.995 -116.115 ;
        RECT -42.325 -117.805 -41.995 -117.475 ;
        RECT -42.325 -119.165 -41.995 -118.835 ;
        RECT -42.325 -120.525 -41.995 -120.195 ;
        RECT -42.325 -123.245 -41.995 -122.915 ;
        RECT -42.325 -124.605 -41.995 -124.275 ;
        RECT -42.325 -125.965 -41.995 -125.635 ;
        RECT -42.325 -127.325 -41.995 -126.995 ;
        RECT -42.325 -128.685 -41.995 -128.355 ;
        RECT -42.325 -130.045 -41.995 -129.715 ;
        RECT -42.325 -131.405 -41.995 -131.075 ;
        RECT -42.325 -132.765 -41.995 -132.435 ;
        RECT -42.325 -134.125 -41.995 -133.795 ;
        RECT -42.325 -135.485 -41.995 -135.155 ;
        RECT -42.325 -136.845 -41.995 -136.515 ;
        RECT -42.325 -138.205 -41.995 -137.875 ;
        RECT -42.325 -139.565 -41.995 -139.235 ;
        RECT -42.325 -140.925 -41.995 -140.595 ;
        RECT -42.325 -142.285 -41.995 -141.955 ;
        RECT -42.325 -143.645 -41.995 -143.315 ;
        RECT -42.325 -145.005 -41.995 -144.675 ;
        RECT -42.325 -146.365 -41.995 -146.035 ;
        RECT -42.325 -147.725 -41.995 -147.395 ;
        RECT -42.325 -149.085 -41.995 -148.755 ;
        RECT -42.325 -150.445 -41.995 -150.115 ;
        RECT -42.325 -151.805 -41.995 -151.475 ;
        RECT -42.325 -153.165 -41.995 -152.835 ;
        RECT -42.325 -154.525 -41.995 -154.195 ;
        RECT -42.325 -155.885 -41.995 -155.555 ;
        RECT -42.325 -157.245 -41.995 -156.915 ;
        RECT -42.325 -158.605 -41.995 -158.275 ;
        RECT -42.325 -159.965 -41.995 -159.635 ;
        RECT -42.325 -161.325 -41.995 -160.995 ;
        RECT -42.325 -162.685 -41.995 -162.355 ;
        RECT -42.325 -164.045 -41.995 -163.715 ;
        RECT -42.325 -165.405 -41.995 -165.075 ;
        RECT -42.325 -166.765 -41.995 -166.435 ;
        RECT -42.325 -169.615 -41.995 -169.285 ;
        RECT -42.325 -170.845 -41.995 -170.515 ;
        RECT -42.325 -172.205 -41.995 -171.875 ;
        RECT -42.325 -173.565 -41.995 -173.235 ;
        RECT -42.325 -177.645 -41.995 -177.315 ;
        RECT -42.325 -179.005 -41.995 -178.675 ;
        RECT -42.325 -184.65 -41.995 -183.52 ;
        RECT -42.32 -184.765 -42 245.285 ;
        RECT -42.325 244.04 -41.995 245.17 ;
        RECT -42.325 239.875 -41.995 240.205 ;
        RECT -42.325 238.515 -41.995 238.845 ;
        RECT -42.325 237.155 -41.995 237.485 ;
        RECT -42.325 235.795 -41.995 236.125 ;
        RECT -42.325 234.435 -41.995 234.765 ;
        RECT -42.325 233.075 -41.995 233.405 ;
        RECT -42.325 231.715 -41.995 232.045 ;
        RECT -42.325 230.355 -41.995 230.685 ;
        RECT -42.325 228.995 -41.995 229.325 ;
        RECT -42.325 227.635 -41.995 227.965 ;
        RECT -42.325 226.275 -41.995 226.605 ;
        RECT -42.325 224.915 -41.995 225.245 ;
        RECT -42.325 223.555 -41.995 223.885 ;
        RECT -42.325 222.195 -41.995 222.525 ;
        RECT -42.325 220.835 -41.995 221.165 ;
        RECT -42.325 219.475 -41.995 219.805 ;
        RECT -42.325 218.115 -41.995 218.445 ;
        RECT -42.325 216.755 -41.995 217.085 ;
        RECT -42.325 215.395 -41.995 215.725 ;
        RECT -42.325 214.035 -41.995 214.365 ;
        RECT -42.325 212.675 -41.995 213.005 ;
        RECT -42.325 211.315 -41.995 211.645 ;
        RECT -42.325 209.955 -41.995 210.285 ;
        RECT -42.325 208.595 -41.995 208.925 ;
        RECT -42.325 207.235 -41.995 207.565 ;
        RECT -42.325 205.875 -41.995 206.205 ;
        RECT -42.325 204.515 -41.995 204.845 ;
        RECT -42.325 203.155 -41.995 203.485 ;
        RECT -42.325 201.795 -41.995 202.125 ;
        RECT -42.325 200.435 -41.995 200.765 ;
        RECT -42.325 199.075 -41.995 199.405 ;
        RECT -42.325 197.715 -41.995 198.045 ;
        RECT -42.325 196.355 -41.995 196.685 ;
        RECT -42.325 194.995 -41.995 195.325 ;
        RECT -42.325 193.635 -41.995 193.965 ;
        RECT -42.325 192.275 -41.995 192.605 ;
        RECT -42.325 190.915 -41.995 191.245 ;
        RECT -42.325 189.555 -41.995 189.885 ;
        RECT -42.325 188.195 -41.995 188.525 ;
        RECT -42.325 186.835 -41.995 187.165 ;
        RECT -42.325 185.475 -41.995 185.805 ;
        RECT -42.325 184.115 -41.995 184.445 ;
        RECT -42.325 182.755 -41.995 183.085 ;
        RECT -42.325 181.395 -41.995 181.725 ;
        RECT -42.325 180.035 -41.995 180.365 ;
        RECT -42.325 178.675 -41.995 179.005 ;
        RECT -42.325 177.315 -41.995 177.645 ;
        RECT -42.325 175.955 -41.995 176.285 ;
        RECT -42.325 174.595 -41.995 174.925 ;
        RECT -42.325 173.235 -41.995 173.565 ;
        RECT -42.325 171.875 -41.995 172.205 ;
        RECT -42.325 170.515 -41.995 170.845 ;
        RECT -42.325 169.155 -41.995 169.485 ;
        RECT -42.325 167.795 -41.995 168.125 ;
        RECT -42.325 166.435 -41.995 166.765 ;
        RECT -42.325 165.075 -41.995 165.405 ;
        RECT -42.325 163.715 -41.995 164.045 ;
        RECT -42.325 162.355 -41.995 162.685 ;
        RECT -42.325 160.995 -41.995 161.325 ;
        RECT -42.325 159.635 -41.995 159.965 ;
        RECT -42.325 158.275 -41.995 158.605 ;
        RECT -42.325 156.915 -41.995 157.245 ;
        RECT -42.325 155.555 -41.995 155.885 ;
        RECT -42.325 154.195 -41.995 154.525 ;
        RECT -42.325 152.835 -41.995 153.165 ;
        RECT -42.325 151.475 -41.995 151.805 ;
        RECT -42.325 150.115 -41.995 150.445 ;
        RECT -42.325 148.755 -41.995 149.085 ;
        RECT -42.325 147.395 -41.995 147.725 ;
        RECT -42.325 146.035 -41.995 146.365 ;
        RECT -42.325 144.675 -41.995 145.005 ;
        RECT -42.325 143.315 -41.995 143.645 ;
        RECT -42.325 141.955 -41.995 142.285 ;
        RECT -42.325 140.595 -41.995 140.925 ;
        RECT -42.325 139.235 -41.995 139.565 ;
        RECT -42.325 137.875 -41.995 138.205 ;
        RECT -42.325 136.515 -41.995 136.845 ;
        RECT -42.325 135.155 -41.995 135.485 ;
        RECT -42.325 133.795 -41.995 134.125 ;
        RECT -42.325 132.435 -41.995 132.765 ;
        RECT -42.325 131.075 -41.995 131.405 ;
        RECT -42.325 129.715 -41.995 130.045 ;
        RECT -42.325 128.355 -41.995 128.685 ;
        RECT -42.325 126.995 -41.995 127.325 ;
        RECT -42.325 125.635 -41.995 125.965 ;
        RECT -42.325 124.275 -41.995 124.605 ;
        RECT -42.325 122.915 -41.995 123.245 ;
        RECT -42.325 121.555 -41.995 121.885 ;
        RECT -42.325 120.195 -41.995 120.525 ;
        RECT -42.325 118.835 -41.995 119.165 ;
        RECT -42.325 117.475 -41.995 117.805 ;
        RECT -42.325 116.115 -41.995 116.445 ;
        RECT -42.325 114.755 -41.995 115.085 ;
        RECT -42.325 113.395 -41.995 113.725 ;
        RECT -42.325 112.035 -41.995 112.365 ;
        RECT -42.325 110.675 -41.995 111.005 ;
        RECT -42.325 109.315 -41.995 109.645 ;
        RECT -42.325 107.955 -41.995 108.285 ;
        RECT -42.325 106.595 -41.995 106.925 ;
        RECT -42.325 105.235 -41.995 105.565 ;
        RECT -42.325 103.875 -41.995 104.205 ;
        RECT -42.325 102.515 -41.995 102.845 ;
        RECT -42.325 101.155 -41.995 101.485 ;
        RECT -42.325 99.795 -41.995 100.125 ;
        RECT -42.325 98.435 -41.995 98.765 ;
        RECT -42.325 97.075 -41.995 97.405 ;
        RECT -42.325 95.715 -41.995 96.045 ;
        RECT -42.325 94.355 -41.995 94.685 ;
        RECT -42.325 92.995 -41.995 93.325 ;
        RECT -42.325 91.635 -41.995 91.965 ;
        RECT -42.325 90.275 -41.995 90.605 ;
        RECT -42.325 88.915 -41.995 89.245 ;
        RECT -42.325 87.555 -41.995 87.885 ;
        RECT -42.325 86.195 -41.995 86.525 ;
        RECT -42.325 84.835 -41.995 85.165 ;
        RECT -42.325 83.475 -41.995 83.805 ;
        RECT -42.325 82.115 -41.995 82.445 ;
        RECT -42.325 80.755 -41.995 81.085 ;
        RECT -42.325 79.395 -41.995 79.725 ;
        RECT -42.325 78.035 -41.995 78.365 ;
        RECT -42.325 76.675 -41.995 77.005 ;
        RECT -42.325 75.315 -41.995 75.645 ;
        RECT -42.325 73.955 -41.995 74.285 ;
        RECT -42.325 72.595 -41.995 72.925 ;
        RECT -42.325 71.235 -41.995 71.565 ;
        RECT -42.325 69.875 -41.995 70.205 ;
        RECT -42.325 68.515 -41.995 68.845 ;
        RECT -42.325 67.155 -41.995 67.485 ;
        RECT -42.325 65.795 -41.995 66.125 ;
        RECT -42.325 64.435 -41.995 64.765 ;
        RECT -42.325 63.075 -41.995 63.405 ;
        RECT -42.325 61.715 -41.995 62.045 ;
        RECT -42.325 60.355 -41.995 60.685 ;
        RECT -42.325 58.995 -41.995 59.325 ;
        RECT -42.325 57.635 -41.995 57.965 ;
        RECT -42.325 56.275 -41.995 56.605 ;
        RECT -42.325 54.915 -41.995 55.245 ;
        RECT -42.325 53.555 -41.995 53.885 ;
        RECT -42.325 52.195 -41.995 52.525 ;
        RECT -42.325 50.835 -41.995 51.165 ;
        RECT -42.325 49.475 -41.995 49.805 ;
        RECT -42.325 48.115 -41.995 48.445 ;
        RECT -42.325 46.755 -41.995 47.085 ;
        RECT -42.325 45.395 -41.995 45.725 ;
        RECT -42.325 44.035 -41.995 44.365 ;
        RECT -42.325 42.675 -41.995 43.005 ;
        RECT -42.325 41.315 -41.995 41.645 ;
        RECT -42.325 39.955 -41.995 40.285 ;
        RECT -42.325 38.595 -41.995 38.925 ;
        RECT -42.325 37.235 -41.995 37.565 ;
        RECT -42.325 35.875 -41.995 36.205 ;
        RECT -42.325 34.515 -41.995 34.845 ;
        RECT -42.325 33.155 -41.995 33.485 ;
        RECT -42.325 31.795 -41.995 32.125 ;
        RECT -42.325 30.435 -41.995 30.765 ;
        RECT -42.325 29.075 -41.995 29.405 ;
        RECT -42.325 27.715 -41.995 28.045 ;
        RECT -42.325 26.355 -41.995 26.685 ;
        RECT -42.325 24.995 -41.995 25.325 ;
        RECT -42.325 23.635 -41.995 23.965 ;
        RECT -42.325 22.275 -41.995 22.605 ;
        RECT -42.325 20.915 -41.995 21.245 ;
        RECT -42.325 19.555 -41.995 19.885 ;
        RECT -42.325 18.195 -41.995 18.525 ;
        RECT -42.325 16.835 -41.995 17.165 ;
        RECT -42.325 15.475 -41.995 15.805 ;
        RECT -42.325 14.115 -41.995 14.445 ;
        RECT -42.325 12.755 -41.995 13.085 ;
        RECT -42.325 11.395 -41.995 11.725 ;
        RECT -42.325 10.035 -41.995 10.365 ;
        RECT -42.325 8.675 -41.995 9.005 ;
        RECT -42.325 7.315 -41.995 7.645 ;
        RECT -42.325 5.955 -41.995 6.285 ;
        RECT -42.325 4.595 -41.995 4.925 ;
        RECT -42.325 3.235 -41.995 3.565 ;
        RECT -42.325 1.875 -41.995 2.205 ;
        RECT -42.325 0.515 -41.995 0.845 ;
        RECT -42.325 -0.845 -41.995 -0.515 ;
        RECT -42.325 -2.205 -41.995 -1.875 ;
        RECT -42.325 -4.925 -41.995 -4.595 ;
        RECT -42.325 -6.285 -41.995 -5.955 ;
        RECT -42.325 -10.365 -41.995 -10.035 ;
        RECT -42.325 -14.445 -41.995 -14.115 ;
        RECT -42.325 -17.165 -41.995 -16.835 ;
        RECT -42.325 -18.525 -41.995 -18.195 ;
        RECT -42.325 -19.885 -41.995 -19.555 ;
        RECT -42.325 -21.245 -41.995 -20.915 ;
        RECT -42.325 -22.605 -41.995 -22.275 ;
        RECT -42.325 -23.965 -41.995 -23.635 ;
        RECT -42.325 -25.325 -41.995 -24.995 ;
        RECT -42.325 -32.125 -41.995 -31.795 ;
        RECT -42.325 -33.71 -41.995 -33.38 ;
        RECT -42.325 -34.845 -41.995 -34.515 ;
        RECT -42.325 -36.205 -41.995 -35.875 ;
        RECT -42.325 -38.925 -41.995 -38.595 ;
        RECT -42.325 -39.75 -41.995 -39.42 ;
        RECT -42.325 -41.645 -41.995 -41.315 ;
        RECT -42.325 -44.365 -41.995 -44.035 ;
        RECT -42.325 -49.805 -41.995 -49.475 ;
        RECT -42.325 -51.165 -41.995 -50.835 ;
        RECT -42.325 -53.885 -41.995 -53.555 ;
        RECT -42.325 -55.245 -41.995 -54.915 ;
        RECT -42.325 -59.325 -41.995 -58.995 ;
        RECT -42.325 -60.685 -41.995 -60.355 ;
        RECT -42.325 -63.405 -41.995 -63.075 ;
        RECT -42.325 -67.485 -41.995 -67.155 ;
        RECT -42.325 -70.205 -41.995 -69.875 ;
        RECT -42.325 -71.565 -41.995 -71.235 ;
        RECT -42.325 -72.925 -41.995 -72.595 ;
        RECT -42.325 -74.285 -41.995 -73.955 ;
        RECT -42.325 -75.645 -41.995 -75.315 ;
        RECT -42.325 -77.005 -41.995 -76.675 ;
        RECT -42.325 -78.365 -41.995 -78.035 ;
        RECT -42.325 -79.725 -41.995 -79.395 ;
        RECT -42.325 -81.085 -41.995 -80.755 ;
        RECT -42.325 -82.445 -41.995 -82.115 ;
        RECT -42.325 -83.805 -41.995 -83.475 ;
        RECT -42.325 -85.165 -41.995 -84.835 ;
        RECT -42.325 -86.525 -41.995 -86.195 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.845 244.04 -51.515 245.17 ;
        RECT -51.845 239.875 -51.515 240.205 ;
        RECT -51.845 238.515 -51.515 238.845 ;
        RECT -51.845 237.155 -51.515 237.485 ;
        RECT -51.845 235.795 -51.515 236.125 ;
        RECT -51.845 234.435 -51.515 234.765 ;
        RECT -51.845 233.075 -51.515 233.405 ;
        RECT -51.845 231.715 -51.515 232.045 ;
        RECT -51.845 230.355 -51.515 230.685 ;
        RECT -51.845 228.995 -51.515 229.325 ;
        RECT -51.845 227.635 -51.515 227.965 ;
        RECT -51.845 226.275 -51.515 226.605 ;
        RECT -51.845 224.915 -51.515 225.245 ;
        RECT -51.845 223.555 -51.515 223.885 ;
        RECT -51.845 222.195 -51.515 222.525 ;
        RECT -51.845 220.835 -51.515 221.165 ;
        RECT -51.845 219.475 -51.515 219.805 ;
        RECT -51.845 218.115 -51.515 218.445 ;
        RECT -51.845 216.755 -51.515 217.085 ;
        RECT -51.845 215.395 -51.515 215.725 ;
        RECT -51.845 214.035 -51.515 214.365 ;
        RECT -51.845 212.675 -51.515 213.005 ;
        RECT -51.845 211.315 -51.515 211.645 ;
        RECT -51.845 209.955 -51.515 210.285 ;
        RECT -51.845 208.595 -51.515 208.925 ;
        RECT -51.845 207.235 -51.515 207.565 ;
        RECT -51.845 205.875 -51.515 206.205 ;
        RECT -51.845 204.515 -51.515 204.845 ;
        RECT -51.845 203.155 -51.515 203.485 ;
        RECT -51.845 201.795 -51.515 202.125 ;
        RECT -51.845 200.435 -51.515 200.765 ;
        RECT -51.845 199.075 -51.515 199.405 ;
        RECT -51.845 197.715 -51.515 198.045 ;
        RECT -51.845 196.355 -51.515 196.685 ;
        RECT -51.845 194.995 -51.515 195.325 ;
        RECT -51.845 193.635 -51.515 193.965 ;
        RECT -51.845 192.275 -51.515 192.605 ;
        RECT -51.845 190.915 -51.515 191.245 ;
        RECT -51.845 189.555 -51.515 189.885 ;
        RECT -51.845 188.195 -51.515 188.525 ;
        RECT -51.845 186.835 -51.515 187.165 ;
        RECT -51.845 185.475 -51.515 185.805 ;
        RECT -51.845 184.115 -51.515 184.445 ;
        RECT -51.845 182.755 -51.515 183.085 ;
        RECT -51.845 181.395 -51.515 181.725 ;
        RECT -51.845 180.035 -51.515 180.365 ;
        RECT -51.845 178.675 -51.515 179.005 ;
        RECT -51.845 177.315 -51.515 177.645 ;
        RECT -51.845 175.955 -51.515 176.285 ;
        RECT -51.845 174.595 -51.515 174.925 ;
        RECT -51.845 173.235 -51.515 173.565 ;
        RECT -51.845 171.875 -51.515 172.205 ;
        RECT -51.845 170.515 -51.515 170.845 ;
        RECT -51.845 169.155 -51.515 169.485 ;
        RECT -51.845 167.795 -51.515 168.125 ;
        RECT -51.845 166.435 -51.515 166.765 ;
        RECT -51.845 165.075 -51.515 165.405 ;
        RECT -51.845 163.715 -51.515 164.045 ;
        RECT -51.845 162.355 -51.515 162.685 ;
        RECT -51.845 160.995 -51.515 161.325 ;
        RECT -51.845 159.635 -51.515 159.965 ;
        RECT -51.845 158.275 -51.515 158.605 ;
        RECT -51.845 156.915 -51.515 157.245 ;
        RECT -51.845 155.555 -51.515 155.885 ;
        RECT -51.845 154.195 -51.515 154.525 ;
        RECT -51.845 152.835 -51.515 153.165 ;
        RECT -51.845 151.475 -51.515 151.805 ;
        RECT -51.845 150.115 -51.515 150.445 ;
        RECT -51.845 148.755 -51.515 149.085 ;
        RECT -51.845 147.395 -51.515 147.725 ;
        RECT -51.845 146.035 -51.515 146.365 ;
        RECT -51.845 144.675 -51.515 145.005 ;
        RECT -51.845 143.315 -51.515 143.645 ;
        RECT -51.845 141.955 -51.515 142.285 ;
        RECT -51.845 140.595 -51.515 140.925 ;
        RECT -51.845 139.235 -51.515 139.565 ;
        RECT -51.845 136.42 -51.515 136.75 ;
        RECT -51.845 134.245 -51.515 134.575 ;
        RECT -51.845 133.395 -51.515 133.725 ;
        RECT -51.845 131.085 -51.515 131.415 ;
        RECT -51.845 130.235 -51.515 130.565 ;
        RECT -51.845 127.925 -51.515 128.255 ;
        RECT -51.845 127.075 -51.515 127.405 ;
        RECT -51.845 124.765 -51.515 125.095 ;
        RECT -51.845 123.915 -51.515 124.245 ;
        RECT -51.845 121.605 -51.515 121.935 ;
        RECT -51.845 120.755 -51.515 121.085 ;
        RECT -51.845 118.445 -51.515 118.775 ;
        RECT -51.845 117.595 -51.515 117.925 ;
        RECT -51.845 115.285 -51.515 115.615 ;
        RECT -51.845 114.435 -51.515 114.765 ;
        RECT -51.845 112.125 -51.515 112.455 ;
        RECT -51.845 111.275 -51.515 111.605 ;
        RECT -51.845 108.965 -51.515 109.295 ;
        RECT -51.845 108.115 -51.515 108.445 ;
        RECT -51.845 105.805 -51.515 106.135 ;
        RECT -51.845 104.955 -51.515 105.285 ;
        RECT -51.845 102.645 -51.515 102.975 ;
        RECT -51.845 101.795 -51.515 102.125 ;
        RECT -51.845 99.62 -51.515 99.95 ;
        RECT -51.845 97.075 -51.515 97.405 ;
        RECT -51.845 95.715 -51.515 96.045 ;
        RECT -51.845 94.355 -51.515 94.685 ;
        RECT -51.845 92.995 -51.515 93.325 ;
        RECT -51.845 91.635 -51.515 91.965 ;
        RECT -51.845 90.275 -51.515 90.605 ;
        RECT -51.845 88.915 -51.515 89.245 ;
        RECT -51.845 87.555 -51.515 87.885 ;
        RECT -51.845 86.195 -51.515 86.525 ;
        RECT -51.845 84.835 -51.515 85.165 ;
        RECT -51.845 83.475 -51.515 83.805 ;
        RECT -51.845 82.115 -51.515 82.445 ;
        RECT -51.845 80.755 -51.515 81.085 ;
        RECT -51.845 79.395 -51.515 79.725 ;
        RECT -51.845 78.035 -51.515 78.365 ;
        RECT -51.845 76.675 -51.515 77.005 ;
        RECT -51.845 75.315 -51.515 75.645 ;
        RECT -51.845 73.955 -51.515 74.285 ;
        RECT -51.845 72.595 -51.515 72.925 ;
        RECT -51.845 71.235 -51.515 71.565 ;
        RECT -51.845 69.875 -51.515 70.205 ;
        RECT -51.845 68.515 -51.515 68.845 ;
        RECT -51.845 67.155 -51.515 67.485 ;
        RECT -51.845 65.795 -51.515 66.125 ;
        RECT -51.845 64.435 -51.515 64.765 ;
        RECT -51.845 63.075 -51.515 63.405 ;
        RECT -51.845 61.715 -51.515 62.045 ;
        RECT -51.845 60.355 -51.515 60.685 ;
        RECT -51.845 58.995 -51.515 59.325 ;
        RECT -51.845 57.635 -51.515 57.965 ;
        RECT -51.845 56.275 -51.515 56.605 ;
        RECT -51.845 54.915 -51.515 55.245 ;
        RECT -51.845 53.555 -51.515 53.885 ;
        RECT -51.845 52.195 -51.515 52.525 ;
        RECT -51.845 50.835 -51.515 51.165 ;
        RECT -51.845 49.475 -51.515 49.805 ;
        RECT -51.845 48.115 -51.515 48.445 ;
        RECT -51.845 46.755 -51.515 47.085 ;
        RECT -51.845 45.395 -51.515 45.725 ;
        RECT -51.845 44.035 -51.515 44.365 ;
        RECT -51.845 42.675 -51.515 43.005 ;
        RECT -51.845 41.315 -51.515 41.645 ;
        RECT -51.845 39.955 -51.515 40.285 ;
        RECT -51.845 38.595 -51.515 38.925 ;
        RECT -51.845 37.235 -51.515 37.565 ;
        RECT -51.845 35.875 -51.515 36.205 ;
        RECT -51.845 34.515 -51.515 34.845 ;
        RECT -51.845 33.155 -51.515 33.485 ;
        RECT -51.845 31.795 -51.515 32.125 ;
        RECT -51.845 30.435 -51.515 30.765 ;
        RECT -51.845 29.075 -51.515 29.405 ;
        RECT -51.845 27.715 -51.515 28.045 ;
        RECT -51.845 26.355 -51.515 26.685 ;
        RECT -51.845 24.995 -51.515 25.325 ;
        RECT -51.845 23.635 -51.515 23.965 ;
        RECT -51.845 22.275 -51.515 22.605 ;
        RECT -51.845 20.915 -51.515 21.245 ;
        RECT -51.845 19.555 -51.515 19.885 ;
        RECT -51.845 18.195 -51.515 18.525 ;
        RECT -51.845 16.835 -51.515 17.165 ;
        RECT -51.845 15.475 -51.515 15.805 ;
        RECT -51.845 14.115 -51.515 14.445 ;
        RECT -51.845 12.755 -51.515 13.085 ;
        RECT -51.845 11.395 -51.515 11.725 ;
        RECT -51.845 10.035 -51.515 10.365 ;
        RECT -51.845 8.675 -51.515 9.005 ;
        RECT -51.845 7.315 -51.515 7.645 ;
        RECT -51.845 5.955 -51.515 6.285 ;
        RECT -51.845 4.595 -51.515 4.925 ;
        RECT -51.845 3.235 -51.515 3.565 ;
        RECT -51.845 1.875 -51.515 2.205 ;
        RECT -51.845 0.515 -51.515 0.845 ;
        RECT -51.845 -0.845 -51.515 -0.515 ;
        RECT -51.845 -2.205 -51.515 -1.875 ;
        RECT -51.845 -3.565 -51.515 -3.235 ;
        RECT -51.845 -4.925 -51.515 -4.595 ;
        RECT -51.845 -6.285 -51.515 -5.955 ;
        RECT -51.845 -7.645 -51.515 -7.315 ;
        RECT -51.845 -9.005 -51.515 -8.675 ;
        RECT -51.845 -10.365 -51.515 -10.035 ;
        RECT -51.845 -11.725 -51.515 -11.395 ;
        RECT -51.845 -13.085 -51.515 -12.755 ;
        RECT -51.845 -14.445 -51.515 -14.115 ;
        RECT -51.845 -15.805 -51.515 -15.475 ;
        RECT -51.845 -17.165 -51.515 -16.835 ;
        RECT -51.845 -18.525 -51.515 -18.195 ;
        RECT -51.845 -19.885 -51.515 -19.555 ;
        RECT -51.845 -21.245 -51.515 -20.915 ;
        RECT -51.845 -22.605 -51.515 -22.275 ;
        RECT -51.845 -23.965 -51.515 -23.635 ;
        RECT -51.845 -25.325 -51.515 -24.995 ;
        RECT -51.845 -30.765 -51.515 -30.435 ;
        RECT -51.845 -32.125 -51.515 -31.795 ;
        RECT -51.845 -33.485 -51.515 -33.155 ;
        RECT -51.845 -34.845 -51.515 -34.515 ;
        RECT -51.845 -36.205 -51.515 -35.875 ;
        RECT -51.845 -37.565 -51.515 -37.235 ;
        RECT -51.845 -38.925 -51.515 -38.595 ;
        RECT -51.845 -40.285 -51.515 -39.955 ;
        RECT -51.845 -41.645 -51.515 -41.315 ;
        RECT -51.845 -43.005 -51.515 -42.675 ;
        RECT -51.845 -44.365 -51.515 -44.035 ;
        RECT -51.845 -45.725 -51.515 -45.395 ;
        RECT -51.845 -47.085 -51.515 -46.755 ;
        RECT -51.845 -48.445 -51.515 -48.115 ;
        RECT -51.845 -49.805 -51.515 -49.475 ;
        RECT -51.845 -51.165 -51.515 -50.835 ;
        RECT -51.845 -52.525 -51.515 -52.195 ;
        RECT -51.845 -53.885 -51.515 -53.555 ;
        RECT -51.845 -55.245 -51.515 -54.915 ;
        RECT -51.845 -56.605 -51.515 -56.275 ;
        RECT -51.845 -57.965 -51.515 -57.635 ;
        RECT -51.845 -59.325 -51.515 -58.995 ;
        RECT -51.845 -60.685 -51.515 -60.355 ;
        RECT -51.845 -62.045 -51.515 -61.715 ;
        RECT -51.845 -63.405 -51.515 -63.075 ;
        RECT -51.845 -64.765 -51.515 -64.435 ;
        RECT -51.845 -66.125 -51.515 -65.795 ;
        RECT -51.845 -68.845 -51.515 -68.515 ;
        RECT -51.845 -70.205 -51.515 -69.875 ;
        RECT -51.845 -71.565 -51.515 -71.235 ;
        RECT -51.845 -72.925 -51.515 -72.595 ;
        RECT -51.845 -74.285 -51.515 -73.955 ;
        RECT -51.845 -75.645 -51.515 -75.315 ;
        RECT -51.845 -77.005 -51.515 -76.675 ;
        RECT -51.845 -78.365 -51.515 -78.035 ;
        RECT -51.845 -79.725 -51.515 -79.395 ;
        RECT -51.845 -81.085 -51.515 -80.755 ;
        RECT -51.845 -82.445 -51.515 -82.115 ;
        RECT -51.845 -83.805 -51.515 -83.475 ;
        RECT -51.845 -85.165 -51.515 -84.835 ;
        RECT -51.845 -86.525 -51.515 -86.195 ;
        RECT -51.845 -87.885 -51.515 -87.555 ;
        RECT -51.845 -89.245 -51.515 -88.915 ;
        RECT -51.845 -90.605 -51.515 -90.275 ;
        RECT -51.845 -91.77 -51.515 -91.44 ;
        RECT -51.845 -93.325 -51.515 -92.995 ;
        RECT -51.845 -94.685 -51.515 -94.355 ;
        RECT -51.845 -96.045 -51.515 -95.715 ;
        RECT -51.845 -97.405 -51.515 -97.075 ;
        RECT -51.845 -98.765 -51.515 -98.435 ;
        RECT -51.845 -101.485 -51.515 -101.155 ;
        RECT -51.845 -102.31 -51.515 -101.98 ;
        RECT -51.845 -104.205 -51.515 -103.875 ;
        RECT -51.845 -105.565 -51.515 -105.235 ;
        RECT -51.845 -106.925 -51.515 -106.595 ;
        RECT -51.845 -109.645 -51.515 -109.315 ;
        RECT -51.845 -111.005 -51.515 -110.675 ;
        RECT -51.845 -113.725 -51.515 -113.395 ;
        RECT -51.845 -115.085 -51.515 -114.755 ;
        RECT -51.845 -116.445 -51.515 -116.115 ;
        RECT -51.845 -117.805 -51.515 -117.475 ;
        RECT -51.845 -119.165 -51.515 -118.835 ;
        RECT -51.845 -120.525 -51.515 -120.195 ;
        RECT -51.845 -123.245 -51.515 -122.915 ;
        RECT -51.845 -124.605 -51.515 -124.275 ;
        RECT -51.845 -125.965 -51.515 -125.635 ;
        RECT -51.845 -127.325 -51.515 -126.995 ;
        RECT -51.845 -128.685 -51.515 -128.355 ;
        RECT -51.845 -130.045 -51.515 -129.715 ;
        RECT -51.845 -131.405 -51.515 -131.075 ;
        RECT -51.845 -132.765 -51.515 -132.435 ;
        RECT -51.845 -134.125 -51.515 -133.795 ;
        RECT -51.845 -135.485 -51.515 -135.155 ;
        RECT -51.845 -136.845 -51.515 -136.515 ;
        RECT -51.845 -138.205 -51.515 -137.875 ;
        RECT -51.845 -139.565 -51.515 -139.235 ;
        RECT -51.845 -140.925 -51.515 -140.595 ;
        RECT -51.845 -142.285 -51.515 -141.955 ;
        RECT -51.845 -143.645 -51.515 -143.315 ;
        RECT -51.845 -145.005 -51.515 -144.675 ;
        RECT -51.845 -146.365 -51.515 -146.035 ;
        RECT -51.845 -147.725 -51.515 -147.395 ;
        RECT -51.845 -149.085 -51.515 -148.755 ;
        RECT -51.845 -150.445 -51.515 -150.115 ;
        RECT -51.845 -151.805 -51.515 -151.475 ;
        RECT -51.845 -153.165 -51.515 -152.835 ;
        RECT -51.845 -154.525 -51.515 -154.195 ;
        RECT -51.845 -155.885 -51.515 -155.555 ;
        RECT -51.845 -157.245 -51.515 -156.915 ;
        RECT -51.845 -158.605 -51.515 -158.275 ;
        RECT -51.845 -159.965 -51.515 -159.635 ;
        RECT -51.845 -161.325 -51.515 -160.995 ;
        RECT -51.845 -162.685 -51.515 -162.355 ;
        RECT -51.845 -164.045 -51.515 -163.715 ;
        RECT -51.845 -165.405 -51.515 -165.075 ;
        RECT -51.845 -166.765 -51.515 -166.435 ;
        RECT -51.845 -169.615 -51.515 -169.285 ;
        RECT -51.845 -170.845 -51.515 -170.515 ;
        RECT -51.845 -172.205 -51.515 -171.875 ;
        RECT -51.845 -174.925 -51.515 -174.595 ;
        RECT -51.845 -177.645 -51.515 -177.315 ;
        RECT -51.845 -179.005 -51.515 -178.675 ;
        RECT -51.845 -184.65 -51.515 -183.52 ;
        RECT -51.84 -184.765 -51.52 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -50.485 244.04 -50.155 245.17 ;
        RECT -50.485 239.875 -50.155 240.205 ;
        RECT -50.485 238.515 -50.155 238.845 ;
        RECT -50.485 237.155 -50.155 237.485 ;
        RECT -50.485 235.795 -50.155 236.125 ;
        RECT -50.485 234.435 -50.155 234.765 ;
        RECT -50.485 233.075 -50.155 233.405 ;
        RECT -50.485 231.715 -50.155 232.045 ;
        RECT -50.485 230.355 -50.155 230.685 ;
        RECT -50.485 228.995 -50.155 229.325 ;
        RECT -50.485 227.635 -50.155 227.965 ;
        RECT -50.485 226.275 -50.155 226.605 ;
        RECT -50.485 224.915 -50.155 225.245 ;
        RECT -50.485 223.555 -50.155 223.885 ;
        RECT -50.485 222.195 -50.155 222.525 ;
        RECT -50.485 220.835 -50.155 221.165 ;
        RECT -50.485 219.475 -50.155 219.805 ;
        RECT -50.485 218.115 -50.155 218.445 ;
        RECT -50.485 216.755 -50.155 217.085 ;
        RECT -50.485 215.395 -50.155 215.725 ;
        RECT -50.485 214.035 -50.155 214.365 ;
        RECT -50.485 212.675 -50.155 213.005 ;
        RECT -50.485 211.315 -50.155 211.645 ;
        RECT -50.485 209.955 -50.155 210.285 ;
        RECT -50.485 208.595 -50.155 208.925 ;
        RECT -50.485 207.235 -50.155 207.565 ;
        RECT -50.485 205.875 -50.155 206.205 ;
        RECT -50.485 204.515 -50.155 204.845 ;
        RECT -50.485 203.155 -50.155 203.485 ;
        RECT -50.485 201.795 -50.155 202.125 ;
        RECT -50.485 200.435 -50.155 200.765 ;
        RECT -50.485 199.075 -50.155 199.405 ;
        RECT -50.485 197.715 -50.155 198.045 ;
        RECT -50.485 196.355 -50.155 196.685 ;
        RECT -50.485 194.995 -50.155 195.325 ;
        RECT -50.485 193.635 -50.155 193.965 ;
        RECT -50.485 192.275 -50.155 192.605 ;
        RECT -50.485 190.915 -50.155 191.245 ;
        RECT -50.485 189.555 -50.155 189.885 ;
        RECT -50.485 188.195 -50.155 188.525 ;
        RECT -50.485 186.835 -50.155 187.165 ;
        RECT -50.485 185.475 -50.155 185.805 ;
        RECT -50.485 184.115 -50.155 184.445 ;
        RECT -50.485 182.755 -50.155 183.085 ;
        RECT -50.485 181.395 -50.155 181.725 ;
        RECT -50.485 180.035 -50.155 180.365 ;
        RECT -50.485 178.675 -50.155 179.005 ;
        RECT -50.485 177.315 -50.155 177.645 ;
        RECT -50.485 175.955 -50.155 176.285 ;
        RECT -50.485 174.595 -50.155 174.925 ;
        RECT -50.485 173.235 -50.155 173.565 ;
        RECT -50.485 171.875 -50.155 172.205 ;
        RECT -50.485 170.515 -50.155 170.845 ;
        RECT -50.485 169.155 -50.155 169.485 ;
        RECT -50.485 167.795 -50.155 168.125 ;
        RECT -50.485 166.435 -50.155 166.765 ;
        RECT -50.485 165.075 -50.155 165.405 ;
        RECT -50.485 163.715 -50.155 164.045 ;
        RECT -50.485 162.355 -50.155 162.685 ;
        RECT -50.485 160.995 -50.155 161.325 ;
        RECT -50.485 159.635 -50.155 159.965 ;
        RECT -50.485 158.275 -50.155 158.605 ;
        RECT -50.485 156.915 -50.155 157.245 ;
        RECT -50.485 155.555 -50.155 155.885 ;
        RECT -50.485 154.195 -50.155 154.525 ;
        RECT -50.485 152.835 -50.155 153.165 ;
        RECT -50.485 151.475 -50.155 151.805 ;
        RECT -50.485 150.115 -50.155 150.445 ;
        RECT -50.485 148.755 -50.155 149.085 ;
        RECT -50.485 147.395 -50.155 147.725 ;
        RECT -50.485 146.035 -50.155 146.365 ;
        RECT -50.485 144.675 -50.155 145.005 ;
        RECT -50.485 143.315 -50.155 143.645 ;
        RECT -50.485 141.955 -50.155 142.285 ;
        RECT -50.485 140.595 -50.155 140.925 ;
        RECT -50.485 139.235 -50.155 139.565 ;
        RECT -50.485 136.42 -50.155 136.75 ;
        RECT -50.485 134.245 -50.155 134.575 ;
        RECT -50.485 133.395 -50.155 133.725 ;
        RECT -50.485 131.085 -50.155 131.415 ;
        RECT -50.485 130.235 -50.155 130.565 ;
        RECT -50.485 127.925 -50.155 128.255 ;
        RECT -50.485 127.075 -50.155 127.405 ;
        RECT -50.485 124.765 -50.155 125.095 ;
        RECT -50.485 123.915 -50.155 124.245 ;
        RECT -50.485 121.605 -50.155 121.935 ;
        RECT -50.485 120.755 -50.155 121.085 ;
        RECT -50.485 118.445 -50.155 118.775 ;
        RECT -50.485 117.595 -50.155 117.925 ;
        RECT -50.485 115.285 -50.155 115.615 ;
        RECT -50.485 114.435 -50.155 114.765 ;
        RECT -50.485 112.125 -50.155 112.455 ;
        RECT -50.485 111.275 -50.155 111.605 ;
        RECT -50.485 108.965 -50.155 109.295 ;
        RECT -50.485 108.115 -50.155 108.445 ;
        RECT -50.485 105.805 -50.155 106.135 ;
        RECT -50.485 104.955 -50.155 105.285 ;
        RECT -50.485 102.645 -50.155 102.975 ;
        RECT -50.485 101.795 -50.155 102.125 ;
        RECT -50.485 99.62 -50.155 99.95 ;
        RECT -50.485 97.075 -50.155 97.405 ;
        RECT -50.485 95.715 -50.155 96.045 ;
        RECT -50.485 94.355 -50.155 94.685 ;
        RECT -50.485 92.995 -50.155 93.325 ;
        RECT -50.485 91.635 -50.155 91.965 ;
        RECT -50.485 90.275 -50.155 90.605 ;
        RECT -50.485 88.915 -50.155 89.245 ;
        RECT -50.485 87.555 -50.155 87.885 ;
        RECT -50.485 86.195 -50.155 86.525 ;
        RECT -50.485 84.835 -50.155 85.165 ;
        RECT -50.485 83.475 -50.155 83.805 ;
        RECT -50.485 82.115 -50.155 82.445 ;
        RECT -50.485 80.755 -50.155 81.085 ;
        RECT -50.485 79.395 -50.155 79.725 ;
        RECT -50.485 78.035 -50.155 78.365 ;
        RECT -50.485 76.675 -50.155 77.005 ;
        RECT -50.485 75.315 -50.155 75.645 ;
        RECT -50.485 73.955 -50.155 74.285 ;
        RECT -50.485 72.595 -50.155 72.925 ;
        RECT -50.485 71.235 -50.155 71.565 ;
        RECT -50.485 69.875 -50.155 70.205 ;
        RECT -50.485 68.515 -50.155 68.845 ;
        RECT -50.485 67.155 -50.155 67.485 ;
        RECT -50.485 65.795 -50.155 66.125 ;
        RECT -50.485 64.435 -50.155 64.765 ;
        RECT -50.485 63.075 -50.155 63.405 ;
        RECT -50.485 61.715 -50.155 62.045 ;
        RECT -50.485 60.355 -50.155 60.685 ;
        RECT -50.485 58.995 -50.155 59.325 ;
        RECT -50.485 57.635 -50.155 57.965 ;
        RECT -50.485 56.275 -50.155 56.605 ;
        RECT -50.485 54.915 -50.155 55.245 ;
        RECT -50.485 53.555 -50.155 53.885 ;
        RECT -50.485 52.195 -50.155 52.525 ;
        RECT -50.485 50.835 -50.155 51.165 ;
        RECT -50.485 49.475 -50.155 49.805 ;
        RECT -50.485 48.115 -50.155 48.445 ;
        RECT -50.485 46.755 -50.155 47.085 ;
        RECT -50.485 45.395 -50.155 45.725 ;
        RECT -50.485 44.035 -50.155 44.365 ;
        RECT -50.485 42.675 -50.155 43.005 ;
        RECT -50.485 41.315 -50.155 41.645 ;
        RECT -50.485 39.955 -50.155 40.285 ;
        RECT -50.485 38.595 -50.155 38.925 ;
        RECT -50.485 37.235 -50.155 37.565 ;
        RECT -50.485 35.875 -50.155 36.205 ;
        RECT -50.485 34.515 -50.155 34.845 ;
        RECT -50.485 33.155 -50.155 33.485 ;
        RECT -50.485 31.795 -50.155 32.125 ;
        RECT -50.485 30.435 -50.155 30.765 ;
        RECT -50.485 29.075 -50.155 29.405 ;
        RECT -50.485 27.715 -50.155 28.045 ;
        RECT -50.485 26.355 -50.155 26.685 ;
        RECT -50.485 24.995 -50.155 25.325 ;
        RECT -50.485 23.635 -50.155 23.965 ;
        RECT -50.485 22.275 -50.155 22.605 ;
        RECT -50.485 20.915 -50.155 21.245 ;
        RECT -50.485 19.555 -50.155 19.885 ;
        RECT -50.485 18.195 -50.155 18.525 ;
        RECT -50.485 16.835 -50.155 17.165 ;
        RECT -50.485 15.475 -50.155 15.805 ;
        RECT -50.485 14.115 -50.155 14.445 ;
        RECT -50.485 12.755 -50.155 13.085 ;
        RECT -50.485 11.395 -50.155 11.725 ;
        RECT -50.485 10.035 -50.155 10.365 ;
        RECT -50.485 8.675 -50.155 9.005 ;
        RECT -50.485 7.315 -50.155 7.645 ;
        RECT -50.485 5.955 -50.155 6.285 ;
        RECT -50.485 4.595 -50.155 4.925 ;
        RECT -50.485 3.235 -50.155 3.565 ;
        RECT -50.485 1.875 -50.155 2.205 ;
        RECT -50.485 0.515 -50.155 0.845 ;
        RECT -50.485 -0.845 -50.155 -0.515 ;
        RECT -50.485 -2.205 -50.155 -1.875 ;
        RECT -50.485 -3.565 -50.155 -3.235 ;
        RECT -50.485 -4.925 -50.155 -4.595 ;
        RECT -50.485 -6.285 -50.155 -5.955 ;
        RECT -50.485 -7.645 -50.155 -7.315 ;
        RECT -50.485 -9.005 -50.155 -8.675 ;
        RECT -50.485 -10.365 -50.155 -10.035 ;
        RECT -50.485 -11.725 -50.155 -11.395 ;
        RECT -50.485 -13.085 -50.155 -12.755 ;
        RECT -50.485 -14.445 -50.155 -14.115 ;
        RECT -50.485 -17.165 -50.155 -16.835 ;
        RECT -50.485 -18.525 -50.155 -18.195 ;
        RECT -50.485 -19.885 -50.155 -19.555 ;
        RECT -50.485 -21.245 -50.155 -20.915 ;
        RECT -50.485 -22.605 -50.155 -22.275 ;
        RECT -50.485 -23.965 -50.155 -23.635 ;
        RECT -50.485 -25.325 -50.155 -24.995 ;
        RECT -50.485 -30.765 -50.155 -30.435 ;
        RECT -50.485 -32.125 -50.155 -31.795 ;
        RECT -50.485 -33.485 -50.155 -33.155 ;
        RECT -50.485 -34.845 -50.155 -34.515 ;
        RECT -50.485 -36.205 -50.155 -35.875 ;
        RECT -50.485 -37.565 -50.155 -37.235 ;
        RECT -50.485 -38.925 -50.155 -38.595 ;
        RECT -50.485 -40.285 -50.155 -39.955 ;
        RECT -50.485 -41.645 -50.155 -41.315 ;
        RECT -50.485 -43.005 -50.155 -42.675 ;
        RECT -50.485 -44.365 -50.155 -44.035 ;
        RECT -50.485 -45.725 -50.155 -45.395 ;
        RECT -50.485 -47.085 -50.155 -46.755 ;
        RECT -50.485 -48.445 -50.155 -48.115 ;
        RECT -50.485 -49.805 -50.155 -49.475 ;
        RECT -50.485 -51.165 -50.155 -50.835 ;
        RECT -50.485 -52.525 -50.155 -52.195 ;
        RECT -50.485 -53.885 -50.155 -53.555 ;
        RECT -50.485 -55.245 -50.155 -54.915 ;
        RECT -50.485 -56.605 -50.155 -56.275 ;
        RECT -50.485 -57.965 -50.155 -57.635 ;
        RECT -50.485 -59.325 -50.155 -58.995 ;
        RECT -50.485 -60.685 -50.155 -60.355 ;
        RECT -50.485 -62.045 -50.155 -61.715 ;
        RECT -50.485 -63.405 -50.155 -63.075 ;
        RECT -50.485 -64.765 -50.155 -64.435 ;
        RECT -50.485 -66.125 -50.155 -65.795 ;
        RECT -50.485 -68.845 -50.155 -68.515 ;
        RECT -50.485 -70.205 -50.155 -69.875 ;
        RECT -50.485 -71.565 -50.155 -71.235 ;
        RECT -50.485 -72.925 -50.155 -72.595 ;
        RECT -50.485 -74.285 -50.155 -73.955 ;
        RECT -50.485 -75.645 -50.155 -75.315 ;
        RECT -50.485 -77.005 -50.155 -76.675 ;
        RECT -50.485 -78.365 -50.155 -78.035 ;
        RECT -50.485 -79.725 -50.155 -79.395 ;
        RECT -50.485 -81.085 -50.155 -80.755 ;
        RECT -50.485 -82.445 -50.155 -82.115 ;
        RECT -50.485 -83.805 -50.155 -83.475 ;
        RECT -50.485 -85.165 -50.155 -84.835 ;
        RECT -50.485 -86.525 -50.155 -86.195 ;
        RECT -50.485 -87.885 -50.155 -87.555 ;
        RECT -50.485 -89.245 -50.155 -88.915 ;
        RECT -50.485 -90.605 -50.155 -90.275 ;
        RECT -50.485 -91.77 -50.155 -91.44 ;
        RECT -50.485 -93.325 -50.155 -92.995 ;
        RECT -50.485 -94.685 -50.155 -94.355 ;
        RECT -50.485 -96.045 -50.155 -95.715 ;
        RECT -50.485 -97.405 -50.155 -97.075 ;
        RECT -50.485 -98.765 -50.155 -98.435 ;
        RECT -50.485 -101.485 -50.155 -101.155 ;
        RECT -50.485 -102.31 -50.155 -101.98 ;
        RECT -50.485 -104.205 -50.155 -103.875 ;
        RECT -50.485 -105.565 -50.155 -105.235 ;
        RECT -50.485 -106.925 -50.155 -106.595 ;
        RECT -50.485 -109.645 -50.155 -109.315 ;
        RECT -50.485 -111.005 -50.155 -110.675 ;
        RECT -50.485 -113.725 -50.155 -113.395 ;
        RECT -50.485 -115.085 -50.155 -114.755 ;
        RECT -50.485 -116.445 -50.155 -116.115 ;
        RECT -50.485 -117.805 -50.155 -117.475 ;
        RECT -50.485 -119.165 -50.155 -118.835 ;
        RECT -50.485 -120.525 -50.155 -120.195 ;
        RECT -50.485 -123.245 -50.155 -122.915 ;
        RECT -50.485 -124.605 -50.155 -124.275 ;
        RECT -50.485 -125.965 -50.155 -125.635 ;
        RECT -50.485 -127.325 -50.155 -126.995 ;
        RECT -50.485 -128.685 -50.155 -128.355 ;
        RECT -50.485 -130.045 -50.155 -129.715 ;
        RECT -50.485 -131.405 -50.155 -131.075 ;
        RECT -50.485 -132.765 -50.155 -132.435 ;
        RECT -50.485 -134.125 -50.155 -133.795 ;
        RECT -50.485 -135.485 -50.155 -135.155 ;
        RECT -50.485 -136.845 -50.155 -136.515 ;
        RECT -50.485 -138.205 -50.155 -137.875 ;
        RECT -50.485 -139.565 -50.155 -139.235 ;
        RECT -50.485 -140.925 -50.155 -140.595 ;
        RECT -50.485 -142.285 -50.155 -141.955 ;
        RECT -50.485 -143.645 -50.155 -143.315 ;
        RECT -50.485 -145.005 -50.155 -144.675 ;
        RECT -50.485 -146.365 -50.155 -146.035 ;
        RECT -50.485 -147.725 -50.155 -147.395 ;
        RECT -50.485 -149.085 -50.155 -148.755 ;
        RECT -50.485 -150.445 -50.155 -150.115 ;
        RECT -50.485 -151.805 -50.155 -151.475 ;
        RECT -50.485 -153.165 -50.155 -152.835 ;
        RECT -50.485 -154.525 -50.155 -154.195 ;
        RECT -50.485 -155.885 -50.155 -155.555 ;
        RECT -50.485 -157.245 -50.155 -156.915 ;
        RECT -50.485 -158.605 -50.155 -158.275 ;
        RECT -50.485 -159.965 -50.155 -159.635 ;
        RECT -50.485 -161.325 -50.155 -160.995 ;
        RECT -50.485 -162.685 -50.155 -162.355 ;
        RECT -50.485 -164.045 -50.155 -163.715 ;
        RECT -50.485 -165.405 -50.155 -165.075 ;
        RECT -50.485 -166.765 -50.155 -166.435 ;
        RECT -50.485 -169.615 -50.155 -169.285 ;
        RECT -50.485 -170.845 -50.155 -170.515 ;
        RECT -50.485 -172.205 -50.155 -171.875 ;
        RECT -50.485 -173.565 -50.155 -173.235 ;
        RECT -50.485 -174.925 -50.155 -174.595 ;
        RECT -50.485 -177.645 -50.155 -177.315 ;
        RECT -50.485 -179.005 -50.155 -178.675 ;
        RECT -50.485 -184.65 -50.155 -183.52 ;
        RECT -50.48 -184.765 -50.16 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.125 244.04 -48.795 245.17 ;
        RECT -49.125 239.875 -48.795 240.205 ;
        RECT -49.125 238.515 -48.795 238.845 ;
        RECT -49.125 237.155 -48.795 237.485 ;
        RECT -49.125 235.795 -48.795 236.125 ;
        RECT -49.125 234.435 -48.795 234.765 ;
        RECT -49.125 233.075 -48.795 233.405 ;
        RECT -49.125 231.715 -48.795 232.045 ;
        RECT -49.125 230.355 -48.795 230.685 ;
        RECT -49.125 228.995 -48.795 229.325 ;
        RECT -49.125 227.635 -48.795 227.965 ;
        RECT -49.125 226.275 -48.795 226.605 ;
        RECT -49.125 224.915 -48.795 225.245 ;
        RECT -49.125 223.555 -48.795 223.885 ;
        RECT -49.125 222.195 -48.795 222.525 ;
        RECT -49.125 220.835 -48.795 221.165 ;
        RECT -49.125 219.475 -48.795 219.805 ;
        RECT -49.125 218.115 -48.795 218.445 ;
        RECT -49.125 216.755 -48.795 217.085 ;
        RECT -49.125 215.395 -48.795 215.725 ;
        RECT -49.125 214.035 -48.795 214.365 ;
        RECT -49.125 212.675 -48.795 213.005 ;
        RECT -49.125 211.315 -48.795 211.645 ;
        RECT -49.125 209.955 -48.795 210.285 ;
        RECT -49.125 208.595 -48.795 208.925 ;
        RECT -49.125 207.235 -48.795 207.565 ;
        RECT -49.125 205.875 -48.795 206.205 ;
        RECT -49.125 204.515 -48.795 204.845 ;
        RECT -49.125 203.155 -48.795 203.485 ;
        RECT -49.125 201.795 -48.795 202.125 ;
        RECT -49.125 200.435 -48.795 200.765 ;
        RECT -49.125 199.075 -48.795 199.405 ;
        RECT -49.125 197.715 -48.795 198.045 ;
        RECT -49.125 196.355 -48.795 196.685 ;
        RECT -49.125 194.995 -48.795 195.325 ;
        RECT -49.125 193.635 -48.795 193.965 ;
        RECT -49.125 192.275 -48.795 192.605 ;
        RECT -49.125 190.915 -48.795 191.245 ;
        RECT -49.125 189.555 -48.795 189.885 ;
        RECT -49.125 188.195 -48.795 188.525 ;
        RECT -49.125 186.835 -48.795 187.165 ;
        RECT -49.125 185.475 -48.795 185.805 ;
        RECT -49.125 184.115 -48.795 184.445 ;
        RECT -49.125 182.755 -48.795 183.085 ;
        RECT -49.125 181.395 -48.795 181.725 ;
        RECT -49.125 180.035 -48.795 180.365 ;
        RECT -49.125 178.675 -48.795 179.005 ;
        RECT -49.125 177.315 -48.795 177.645 ;
        RECT -49.125 175.955 -48.795 176.285 ;
        RECT -49.125 174.595 -48.795 174.925 ;
        RECT -49.125 173.235 -48.795 173.565 ;
        RECT -49.125 171.875 -48.795 172.205 ;
        RECT -49.125 170.515 -48.795 170.845 ;
        RECT -49.125 169.155 -48.795 169.485 ;
        RECT -49.125 167.795 -48.795 168.125 ;
        RECT -49.125 166.435 -48.795 166.765 ;
        RECT -49.125 165.075 -48.795 165.405 ;
        RECT -49.125 163.715 -48.795 164.045 ;
        RECT -49.125 162.355 -48.795 162.685 ;
        RECT -49.125 160.995 -48.795 161.325 ;
        RECT -49.125 159.635 -48.795 159.965 ;
        RECT -49.125 158.275 -48.795 158.605 ;
        RECT -49.125 156.915 -48.795 157.245 ;
        RECT -49.125 155.555 -48.795 155.885 ;
        RECT -49.125 154.195 -48.795 154.525 ;
        RECT -49.125 152.835 -48.795 153.165 ;
        RECT -49.125 151.475 -48.795 151.805 ;
        RECT -49.125 150.115 -48.795 150.445 ;
        RECT -49.125 148.755 -48.795 149.085 ;
        RECT -49.125 147.395 -48.795 147.725 ;
        RECT -49.125 146.035 -48.795 146.365 ;
        RECT -49.125 144.675 -48.795 145.005 ;
        RECT -49.125 143.315 -48.795 143.645 ;
        RECT -49.125 141.955 -48.795 142.285 ;
        RECT -49.125 140.595 -48.795 140.925 ;
        RECT -49.125 139.235 -48.795 139.565 ;
        RECT -49.125 136.42 -48.795 136.75 ;
        RECT -49.125 134.245 -48.795 134.575 ;
        RECT -49.125 133.395 -48.795 133.725 ;
        RECT -49.125 131.085 -48.795 131.415 ;
        RECT -49.125 130.235 -48.795 130.565 ;
        RECT -49.125 127.925 -48.795 128.255 ;
        RECT -49.125 127.075 -48.795 127.405 ;
        RECT -49.125 124.765 -48.795 125.095 ;
        RECT -49.125 123.915 -48.795 124.245 ;
        RECT -49.125 121.605 -48.795 121.935 ;
        RECT -49.125 120.755 -48.795 121.085 ;
        RECT -49.125 118.445 -48.795 118.775 ;
        RECT -49.125 117.595 -48.795 117.925 ;
        RECT -49.125 115.285 -48.795 115.615 ;
        RECT -49.125 114.435 -48.795 114.765 ;
        RECT -49.125 112.125 -48.795 112.455 ;
        RECT -49.125 111.275 -48.795 111.605 ;
        RECT -49.125 108.965 -48.795 109.295 ;
        RECT -49.125 108.115 -48.795 108.445 ;
        RECT -49.125 105.805 -48.795 106.135 ;
        RECT -49.125 104.955 -48.795 105.285 ;
        RECT -49.125 102.645 -48.795 102.975 ;
        RECT -49.125 101.795 -48.795 102.125 ;
        RECT -49.125 99.62 -48.795 99.95 ;
        RECT -49.125 97.075 -48.795 97.405 ;
        RECT -49.125 95.715 -48.795 96.045 ;
        RECT -49.125 94.355 -48.795 94.685 ;
        RECT -49.125 92.995 -48.795 93.325 ;
        RECT -49.125 91.635 -48.795 91.965 ;
        RECT -49.125 90.275 -48.795 90.605 ;
        RECT -49.125 88.915 -48.795 89.245 ;
        RECT -49.125 87.555 -48.795 87.885 ;
        RECT -49.125 86.195 -48.795 86.525 ;
        RECT -49.125 84.835 -48.795 85.165 ;
        RECT -49.125 83.475 -48.795 83.805 ;
        RECT -49.125 82.115 -48.795 82.445 ;
        RECT -49.125 80.755 -48.795 81.085 ;
        RECT -49.125 79.395 -48.795 79.725 ;
        RECT -49.125 78.035 -48.795 78.365 ;
        RECT -49.125 76.675 -48.795 77.005 ;
        RECT -49.125 75.315 -48.795 75.645 ;
        RECT -49.125 73.955 -48.795 74.285 ;
        RECT -49.125 72.595 -48.795 72.925 ;
        RECT -49.125 71.235 -48.795 71.565 ;
        RECT -49.125 69.875 -48.795 70.205 ;
        RECT -49.125 68.515 -48.795 68.845 ;
        RECT -49.125 67.155 -48.795 67.485 ;
        RECT -49.125 65.795 -48.795 66.125 ;
        RECT -49.125 64.435 -48.795 64.765 ;
        RECT -49.125 63.075 -48.795 63.405 ;
        RECT -49.125 61.715 -48.795 62.045 ;
        RECT -49.125 60.355 -48.795 60.685 ;
        RECT -49.125 58.995 -48.795 59.325 ;
        RECT -49.125 57.635 -48.795 57.965 ;
        RECT -49.125 56.275 -48.795 56.605 ;
        RECT -49.125 54.915 -48.795 55.245 ;
        RECT -49.125 53.555 -48.795 53.885 ;
        RECT -49.125 52.195 -48.795 52.525 ;
        RECT -49.125 50.835 -48.795 51.165 ;
        RECT -49.125 49.475 -48.795 49.805 ;
        RECT -49.125 48.115 -48.795 48.445 ;
        RECT -49.125 46.755 -48.795 47.085 ;
        RECT -49.125 45.395 -48.795 45.725 ;
        RECT -49.125 44.035 -48.795 44.365 ;
        RECT -49.125 42.675 -48.795 43.005 ;
        RECT -49.125 41.315 -48.795 41.645 ;
        RECT -49.125 39.955 -48.795 40.285 ;
        RECT -49.125 38.595 -48.795 38.925 ;
        RECT -49.125 37.235 -48.795 37.565 ;
        RECT -49.125 35.875 -48.795 36.205 ;
        RECT -49.125 34.515 -48.795 34.845 ;
        RECT -49.125 33.155 -48.795 33.485 ;
        RECT -49.125 31.795 -48.795 32.125 ;
        RECT -49.125 30.435 -48.795 30.765 ;
        RECT -49.125 29.075 -48.795 29.405 ;
        RECT -49.125 27.715 -48.795 28.045 ;
        RECT -49.125 26.355 -48.795 26.685 ;
        RECT -49.125 24.995 -48.795 25.325 ;
        RECT -49.125 23.635 -48.795 23.965 ;
        RECT -49.125 22.275 -48.795 22.605 ;
        RECT -49.125 20.915 -48.795 21.245 ;
        RECT -49.125 19.555 -48.795 19.885 ;
        RECT -49.125 18.195 -48.795 18.525 ;
        RECT -49.125 16.835 -48.795 17.165 ;
        RECT -49.125 15.475 -48.795 15.805 ;
        RECT -49.125 14.115 -48.795 14.445 ;
        RECT -49.125 12.755 -48.795 13.085 ;
        RECT -49.125 11.395 -48.795 11.725 ;
        RECT -49.125 10.035 -48.795 10.365 ;
        RECT -49.125 8.675 -48.795 9.005 ;
        RECT -49.125 7.315 -48.795 7.645 ;
        RECT -49.125 5.955 -48.795 6.285 ;
        RECT -49.125 4.595 -48.795 4.925 ;
        RECT -49.125 3.235 -48.795 3.565 ;
        RECT -49.125 1.875 -48.795 2.205 ;
        RECT -49.125 0.515 -48.795 0.845 ;
        RECT -49.125 -0.845 -48.795 -0.515 ;
        RECT -49.125 -2.205 -48.795 -1.875 ;
        RECT -49.125 -3.565 -48.795 -3.235 ;
        RECT -49.125 -4.925 -48.795 -4.595 ;
        RECT -49.125 -6.285 -48.795 -5.955 ;
        RECT -49.125 -7.645 -48.795 -7.315 ;
        RECT -49.125 -9.005 -48.795 -8.675 ;
        RECT -49.125 -10.365 -48.795 -10.035 ;
        RECT -49.125 -11.725 -48.795 -11.395 ;
        RECT -49.125 -14.445 -48.795 -14.115 ;
        RECT -49.125 -17.165 -48.795 -16.835 ;
        RECT -49.125 -18.525 -48.795 -18.195 ;
        RECT -49.125 -19.885 -48.795 -19.555 ;
        RECT -49.125 -21.245 -48.795 -20.915 ;
        RECT -49.125 -22.605 -48.795 -22.275 ;
        RECT -49.125 -23.965 -48.795 -23.635 ;
        RECT -49.125 -25.325 -48.795 -24.995 ;
        RECT -49.125 -30.765 -48.795 -30.435 ;
        RECT -49.125 -32.125 -48.795 -31.795 ;
        RECT -49.125 -33.71 -48.795 -33.38 ;
        RECT -49.125 -34.845 -48.795 -34.515 ;
        RECT -49.125 -36.205 -48.795 -35.875 ;
        RECT -49.125 -38.925 -48.795 -38.595 ;
        RECT -49.125 -39.75 -48.795 -39.42 ;
        RECT -49.125 -41.645 -48.795 -41.315 ;
        RECT -49.125 -44.365 -48.795 -44.035 ;
        RECT -49.125 -49.805 -48.795 -49.475 ;
        RECT -49.125 -51.165 -48.795 -50.835 ;
        RECT -49.125 -53.885 -48.795 -53.555 ;
        RECT -49.125 -55.245 -48.795 -54.915 ;
        RECT -49.125 -59.325 -48.795 -58.995 ;
        RECT -49.125 -60.685 -48.795 -60.355 ;
        RECT -49.125 -63.405 -48.795 -63.075 ;
        RECT -49.125 -68.845 -48.795 -68.515 ;
        RECT -49.125 -70.205 -48.795 -69.875 ;
        RECT -49.125 -71.565 -48.795 -71.235 ;
        RECT -49.125 -72.925 -48.795 -72.595 ;
        RECT -49.125 -74.285 -48.795 -73.955 ;
        RECT -49.125 -75.645 -48.795 -75.315 ;
        RECT -49.125 -77.005 -48.795 -76.675 ;
        RECT -49.125 -78.365 -48.795 -78.035 ;
        RECT -49.125 -79.725 -48.795 -79.395 ;
        RECT -49.125 -81.085 -48.795 -80.755 ;
        RECT -49.125 -82.445 -48.795 -82.115 ;
        RECT -49.125 -83.805 -48.795 -83.475 ;
        RECT -49.125 -85.165 -48.795 -84.835 ;
        RECT -49.125 -86.525 -48.795 -86.195 ;
        RECT -49.125 -87.885 -48.795 -87.555 ;
        RECT -49.125 -89.245 -48.795 -88.915 ;
        RECT -49.125 -90.605 -48.795 -90.275 ;
        RECT -49.125 -91.77 -48.795 -91.44 ;
        RECT -49.125 -93.325 -48.795 -92.995 ;
        RECT -49.125 -94.685 -48.795 -94.355 ;
        RECT -49.125 -96.045 -48.795 -95.715 ;
        RECT -49.125 -97.405 -48.795 -97.075 ;
        RECT -49.125 -98.765 -48.795 -98.435 ;
        RECT -49.125 -101.485 -48.795 -101.155 ;
        RECT -49.125 -102.31 -48.795 -101.98 ;
        RECT -49.125 -104.205 -48.795 -103.875 ;
        RECT -49.125 -105.565 -48.795 -105.235 ;
        RECT -49.125 -106.925 -48.795 -106.595 ;
        RECT -49.125 -109.645 -48.795 -109.315 ;
        RECT -49.125 -111.005 -48.795 -110.675 ;
        RECT -49.125 -115.085 -48.795 -114.755 ;
        RECT -49.125 -116.445 -48.795 -116.115 ;
        RECT -49.125 -117.805 -48.795 -117.475 ;
        RECT -49.125 -119.165 -48.795 -118.835 ;
        RECT -49.125 -120.525 -48.795 -120.195 ;
        RECT -49.125 -123.245 -48.795 -122.915 ;
        RECT -49.125 -124.605 -48.795 -124.275 ;
        RECT -49.125 -125.965 -48.795 -125.635 ;
        RECT -49.125 -127.325 -48.795 -126.995 ;
        RECT -49.125 -128.685 -48.795 -128.355 ;
        RECT -49.125 -130.045 -48.795 -129.715 ;
        RECT -49.125 -131.405 -48.795 -131.075 ;
        RECT -49.125 -132.765 -48.795 -132.435 ;
        RECT -49.125 -134.125 -48.795 -133.795 ;
        RECT -49.125 -135.485 -48.795 -135.155 ;
        RECT -49.125 -136.845 -48.795 -136.515 ;
        RECT -49.125 -138.205 -48.795 -137.875 ;
        RECT -49.125 -139.565 -48.795 -139.235 ;
        RECT -49.125 -140.925 -48.795 -140.595 ;
        RECT -49.125 -142.285 -48.795 -141.955 ;
        RECT -49.125 -143.645 -48.795 -143.315 ;
        RECT -49.125 -145.005 -48.795 -144.675 ;
        RECT -49.125 -146.365 -48.795 -146.035 ;
        RECT -49.125 -147.725 -48.795 -147.395 ;
        RECT -49.125 -149.085 -48.795 -148.755 ;
        RECT -49.125 -150.445 -48.795 -150.115 ;
        RECT -49.125 -151.805 -48.795 -151.475 ;
        RECT -49.125 -153.165 -48.795 -152.835 ;
        RECT -49.125 -154.525 -48.795 -154.195 ;
        RECT -49.125 -155.885 -48.795 -155.555 ;
        RECT -49.125 -157.245 -48.795 -156.915 ;
        RECT -49.125 -158.605 -48.795 -158.275 ;
        RECT -49.125 -159.965 -48.795 -159.635 ;
        RECT -49.125 -161.325 -48.795 -160.995 ;
        RECT -49.125 -162.685 -48.795 -162.355 ;
        RECT -49.125 -164.045 -48.795 -163.715 ;
        RECT -49.125 -165.405 -48.795 -165.075 ;
        RECT -49.125 -166.765 -48.795 -166.435 ;
        RECT -49.125 -169.615 -48.795 -169.285 ;
        RECT -49.125 -170.845 -48.795 -170.515 ;
        RECT -49.125 -172.205 -48.795 -171.875 ;
        RECT -49.125 -173.565 -48.795 -173.235 ;
        RECT -49.125 -174.925 -48.795 -174.595 ;
        RECT -49.125 -177.645 -48.795 -177.315 ;
        RECT -49.125 -179.005 -48.795 -178.675 ;
        RECT -49.125 -184.65 -48.795 -183.52 ;
        RECT -49.12 -184.765 -48.8 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.765 5.955 -47.435 6.285 ;
        RECT -47.765 4.595 -47.435 4.925 ;
        RECT -47.765 3.235 -47.435 3.565 ;
        RECT -47.765 1.875 -47.435 2.205 ;
        RECT -47.765 0.515 -47.435 0.845 ;
        RECT -47.765 -0.845 -47.435 -0.515 ;
        RECT -47.765 -2.205 -47.435 -1.875 ;
        RECT -47.765 -3.565 -47.435 -3.235 ;
        RECT -47.765 -4.925 -47.435 -4.595 ;
        RECT -47.765 -6.285 -47.435 -5.955 ;
        RECT -47.765 -7.645 -47.435 -7.315 ;
        RECT -47.765 -9.005 -47.435 -8.675 ;
        RECT -47.765 -10.365 -47.435 -10.035 ;
        RECT -47.765 -14.445 -47.435 -14.115 ;
        RECT -47.765 -17.165 -47.435 -16.835 ;
        RECT -47.765 -18.525 -47.435 -18.195 ;
        RECT -47.765 -19.885 -47.435 -19.555 ;
        RECT -47.765 -21.245 -47.435 -20.915 ;
        RECT -47.765 -22.605 -47.435 -22.275 ;
        RECT -47.765 -23.965 -47.435 -23.635 ;
        RECT -47.765 -25.325 -47.435 -24.995 ;
        RECT -47.765 -30.765 -47.435 -30.435 ;
        RECT -47.765 -32.125 -47.435 -31.795 ;
        RECT -47.765 -33.71 -47.435 -33.38 ;
        RECT -47.765 -34.845 -47.435 -34.515 ;
        RECT -47.765 -36.205 -47.435 -35.875 ;
        RECT -47.765 -38.925 -47.435 -38.595 ;
        RECT -47.765 -39.75 -47.435 -39.42 ;
        RECT -47.765 -41.645 -47.435 -41.315 ;
        RECT -47.765 -44.365 -47.435 -44.035 ;
        RECT -47.765 -49.805 -47.435 -49.475 ;
        RECT -47.765 -51.165 -47.435 -50.835 ;
        RECT -47.765 -53.885 -47.435 -53.555 ;
        RECT -47.765 -55.245 -47.435 -54.915 ;
        RECT -47.765 -59.325 -47.435 -58.995 ;
        RECT -47.765 -60.685 -47.435 -60.355 ;
        RECT -47.765 -63.405 -47.435 -63.075 ;
        RECT -47.765 -70.205 -47.435 -69.875 ;
        RECT -47.765 -71.565 -47.435 -71.235 ;
        RECT -47.765 -72.925 -47.435 -72.595 ;
        RECT -47.765 -74.285 -47.435 -73.955 ;
        RECT -47.765 -75.645 -47.435 -75.315 ;
        RECT -47.765 -77.005 -47.435 -76.675 ;
        RECT -47.765 -78.365 -47.435 -78.035 ;
        RECT -47.765 -79.725 -47.435 -79.395 ;
        RECT -47.765 -81.085 -47.435 -80.755 ;
        RECT -47.765 -82.445 -47.435 -82.115 ;
        RECT -47.765 -83.805 -47.435 -83.475 ;
        RECT -47.765 -85.165 -47.435 -84.835 ;
        RECT -47.765 -86.525 -47.435 -86.195 ;
        RECT -47.765 -87.885 -47.435 -87.555 ;
        RECT -47.765 -89.245 -47.435 -88.915 ;
        RECT -47.765 -90.605 -47.435 -90.275 ;
        RECT -47.765 -91.77 -47.435 -91.44 ;
        RECT -47.765 -93.325 -47.435 -92.995 ;
        RECT -47.765 -94.685 -47.435 -94.355 ;
        RECT -47.765 -96.045 -47.435 -95.715 ;
        RECT -47.765 -97.405 -47.435 -97.075 ;
        RECT -47.765 -98.765 -47.435 -98.435 ;
        RECT -47.765 -101.485 -47.435 -101.155 ;
        RECT -47.765 -102.31 -47.435 -101.98 ;
        RECT -47.765 -104.205 -47.435 -103.875 ;
        RECT -47.765 -105.565 -47.435 -105.235 ;
        RECT -47.765 -106.925 -47.435 -106.595 ;
        RECT -47.765 -109.645 -47.435 -109.315 ;
        RECT -47.765 -111.005 -47.435 -110.675 ;
        RECT -47.76 -113.04 -47.44 245.285 ;
        RECT -47.765 244.04 -47.435 245.17 ;
        RECT -47.765 239.875 -47.435 240.205 ;
        RECT -47.765 238.515 -47.435 238.845 ;
        RECT -47.765 237.155 -47.435 237.485 ;
        RECT -47.765 235.795 -47.435 236.125 ;
        RECT -47.765 234.435 -47.435 234.765 ;
        RECT -47.765 233.075 -47.435 233.405 ;
        RECT -47.765 231.715 -47.435 232.045 ;
        RECT -47.765 230.355 -47.435 230.685 ;
        RECT -47.765 228.995 -47.435 229.325 ;
        RECT -47.765 227.635 -47.435 227.965 ;
        RECT -47.765 226.275 -47.435 226.605 ;
        RECT -47.765 224.915 -47.435 225.245 ;
        RECT -47.765 223.555 -47.435 223.885 ;
        RECT -47.765 222.195 -47.435 222.525 ;
        RECT -47.765 220.835 -47.435 221.165 ;
        RECT -47.765 219.475 -47.435 219.805 ;
        RECT -47.765 218.115 -47.435 218.445 ;
        RECT -47.765 216.755 -47.435 217.085 ;
        RECT -47.765 215.395 -47.435 215.725 ;
        RECT -47.765 214.035 -47.435 214.365 ;
        RECT -47.765 212.675 -47.435 213.005 ;
        RECT -47.765 211.315 -47.435 211.645 ;
        RECT -47.765 209.955 -47.435 210.285 ;
        RECT -47.765 208.595 -47.435 208.925 ;
        RECT -47.765 207.235 -47.435 207.565 ;
        RECT -47.765 205.875 -47.435 206.205 ;
        RECT -47.765 204.515 -47.435 204.845 ;
        RECT -47.765 203.155 -47.435 203.485 ;
        RECT -47.765 201.795 -47.435 202.125 ;
        RECT -47.765 200.435 -47.435 200.765 ;
        RECT -47.765 199.075 -47.435 199.405 ;
        RECT -47.765 197.715 -47.435 198.045 ;
        RECT -47.765 196.355 -47.435 196.685 ;
        RECT -47.765 194.995 -47.435 195.325 ;
        RECT -47.765 193.635 -47.435 193.965 ;
        RECT -47.765 192.275 -47.435 192.605 ;
        RECT -47.765 190.915 -47.435 191.245 ;
        RECT -47.765 189.555 -47.435 189.885 ;
        RECT -47.765 188.195 -47.435 188.525 ;
        RECT -47.765 186.835 -47.435 187.165 ;
        RECT -47.765 185.475 -47.435 185.805 ;
        RECT -47.765 184.115 -47.435 184.445 ;
        RECT -47.765 182.755 -47.435 183.085 ;
        RECT -47.765 181.395 -47.435 181.725 ;
        RECT -47.765 180.035 -47.435 180.365 ;
        RECT -47.765 178.675 -47.435 179.005 ;
        RECT -47.765 177.315 -47.435 177.645 ;
        RECT -47.765 175.955 -47.435 176.285 ;
        RECT -47.765 174.595 -47.435 174.925 ;
        RECT -47.765 173.235 -47.435 173.565 ;
        RECT -47.765 171.875 -47.435 172.205 ;
        RECT -47.765 170.515 -47.435 170.845 ;
        RECT -47.765 169.155 -47.435 169.485 ;
        RECT -47.765 167.795 -47.435 168.125 ;
        RECT -47.765 166.435 -47.435 166.765 ;
        RECT -47.765 165.075 -47.435 165.405 ;
        RECT -47.765 163.715 -47.435 164.045 ;
        RECT -47.765 162.355 -47.435 162.685 ;
        RECT -47.765 160.995 -47.435 161.325 ;
        RECT -47.765 159.635 -47.435 159.965 ;
        RECT -47.765 158.275 -47.435 158.605 ;
        RECT -47.765 156.915 -47.435 157.245 ;
        RECT -47.765 155.555 -47.435 155.885 ;
        RECT -47.765 154.195 -47.435 154.525 ;
        RECT -47.765 152.835 -47.435 153.165 ;
        RECT -47.765 151.475 -47.435 151.805 ;
        RECT -47.765 150.115 -47.435 150.445 ;
        RECT -47.765 148.755 -47.435 149.085 ;
        RECT -47.765 147.395 -47.435 147.725 ;
        RECT -47.765 146.035 -47.435 146.365 ;
        RECT -47.765 144.675 -47.435 145.005 ;
        RECT -47.765 143.315 -47.435 143.645 ;
        RECT -47.765 141.955 -47.435 142.285 ;
        RECT -47.765 140.595 -47.435 140.925 ;
        RECT -47.765 139.235 -47.435 139.565 ;
        RECT -47.765 97.075 -47.435 97.405 ;
        RECT -47.765 95.715 -47.435 96.045 ;
        RECT -47.765 94.355 -47.435 94.685 ;
        RECT -47.765 92.995 -47.435 93.325 ;
        RECT -47.765 91.635 -47.435 91.965 ;
        RECT -47.765 90.275 -47.435 90.605 ;
        RECT -47.765 88.915 -47.435 89.245 ;
        RECT -47.765 87.555 -47.435 87.885 ;
        RECT -47.765 86.195 -47.435 86.525 ;
        RECT -47.765 84.835 -47.435 85.165 ;
        RECT -47.765 83.475 -47.435 83.805 ;
        RECT -47.765 82.115 -47.435 82.445 ;
        RECT -47.765 80.755 -47.435 81.085 ;
        RECT -47.765 79.395 -47.435 79.725 ;
        RECT -47.765 78.035 -47.435 78.365 ;
        RECT -47.765 76.675 -47.435 77.005 ;
        RECT -47.765 75.315 -47.435 75.645 ;
        RECT -47.765 73.955 -47.435 74.285 ;
        RECT -47.765 72.595 -47.435 72.925 ;
        RECT -47.765 71.235 -47.435 71.565 ;
        RECT -47.765 69.875 -47.435 70.205 ;
        RECT -47.765 68.515 -47.435 68.845 ;
        RECT -47.765 67.155 -47.435 67.485 ;
        RECT -47.765 65.795 -47.435 66.125 ;
        RECT -47.765 64.435 -47.435 64.765 ;
        RECT -47.765 63.075 -47.435 63.405 ;
        RECT -47.765 61.715 -47.435 62.045 ;
        RECT -47.765 60.355 -47.435 60.685 ;
        RECT -47.765 58.995 -47.435 59.325 ;
        RECT -47.765 57.635 -47.435 57.965 ;
        RECT -47.765 56.275 -47.435 56.605 ;
        RECT -47.765 54.915 -47.435 55.245 ;
        RECT -47.765 53.555 -47.435 53.885 ;
        RECT -47.765 52.195 -47.435 52.525 ;
        RECT -47.765 50.835 -47.435 51.165 ;
        RECT -47.765 49.475 -47.435 49.805 ;
        RECT -47.765 48.115 -47.435 48.445 ;
        RECT -47.765 46.755 -47.435 47.085 ;
        RECT -47.765 45.395 -47.435 45.725 ;
        RECT -47.765 44.035 -47.435 44.365 ;
        RECT -47.765 42.675 -47.435 43.005 ;
        RECT -47.765 41.315 -47.435 41.645 ;
        RECT -47.765 39.955 -47.435 40.285 ;
        RECT -47.765 38.595 -47.435 38.925 ;
        RECT -47.765 37.235 -47.435 37.565 ;
        RECT -47.765 35.875 -47.435 36.205 ;
        RECT -47.765 34.515 -47.435 34.845 ;
        RECT -47.765 33.155 -47.435 33.485 ;
        RECT -47.765 31.795 -47.435 32.125 ;
        RECT -47.765 30.435 -47.435 30.765 ;
        RECT -47.765 29.075 -47.435 29.405 ;
        RECT -47.765 27.715 -47.435 28.045 ;
        RECT -47.765 26.355 -47.435 26.685 ;
        RECT -47.765 24.995 -47.435 25.325 ;
        RECT -47.765 23.635 -47.435 23.965 ;
        RECT -47.765 22.275 -47.435 22.605 ;
        RECT -47.765 20.915 -47.435 21.245 ;
        RECT -47.765 19.555 -47.435 19.885 ;
        RECT -47.765 18.195 -47.435 18.525 ;
        RECT -47.765 16.835 -47.435 17.165 ;
        RECT -47.765 15.475 -47.435 15.805 ;
        RECT -47.765 14.115 -47.435 14.445 ;
        RECT -47.765 12.755 -47.435 13.085 ;
        RECT -47.765 11.395 -47.435 11.725 ;
        RECT -47.765 10.035 -47.435 10.365 ;
        RECT -47.765 8.675 -47.435 9.005 ;
        RECT -47.765 7.315 -47.435 7.645 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.285 244.04 -56.955 245.17 ;
        RECT -57.285 239.875 -56.955 240.205 ;
        RECT -57.285 238.515 -56.955 238.845 ;
        RECT -57.285 237.155 -56.955 237.485 ;
        RECT -57.285 235.795 -56.955 236.125 ;
        RECT -57.285 234.435 -56.955 234.765 ;
        RECT -57.285 233.075 -56.955 233.405 ;
        RECT -57.285 231.715 -56.955 232.045 ;
        RECT -57.285 230.355 -56.955 230.685 ;
        RECT -57.285 228.995 -56.955 229.325 ;
        RECT -57.285 227.635 -56.955 227.965 ;
        RECT -57.285 226.275 -56.955 226.605 ;
        RECT -57.285 224.915 -56.955 225.245 ;
        RECT -57.285 223.555 -56.955 223.885 ;
        RECT -57.285 222.195 -56.955 222.525 ;
        RECT -57.285 220.835 -56.955 221.165 ;
        RECT -57.285 219.475 -56.955 219.805 ;
        RECT -57.285 218.115 -56.955 218.445 ;
        RECT -57.285 216.755 -56.955 217.085 ;
        RECT -57.285 215.395 -56.955 215.725 ;
        RECT -57.285 214.035 -56.955 214.365 ;
        RECT -57.285 212.675 -56.955 213.005 ;
        RECT -57.285 211.315 -56.955 211.645 ;
        RECT -57.285 209.955 -56.955 210.285 ;
        RECT -57.285 208.595 -56.955 208.925 ;
        RECT -57.285 207.235 -56.955 207.565 ;
        RECT -57.285 205.875 -56.955 206.205 ;
        RECT -57.285 204.515 -56.955 204.845 ;
        RECT -57.285 203.155 -56.955 203.485 ;
        RECT -57.285 201.795 -56.955 202.125 ;
        RECT -57.285 200.435 -56.955 200.765 ;
        RECT -57.285 199.075 -56.955 199.405 ;
        RECT -57.285 197.715 -56.955 198.045 ;
        RECT -57.285 196.355 -56.955 196.685 ;
        RECT -57.285 194.995 -56.955 195.325 ;
        RECT -57.285 193.635 -56.955 193.965 ;
        RECT -57.285 192.275 -56.955 192.605 ;
        RECT -57.285 190.915 -56.955 191.245 ;
        RECT -57.285 189.555 -56.955 189.885 ;
        RECT -57.285 188.195 -56.955 188.525 ;
        RECT -57.285 186.835 -56.955 187.165 ;
        RECT -57.285 185.475 -56.955 185.805 ;
        RECT -57.285 184.115 -56.955 184.445 ;
        RECT -57.285 182.755 -56.955 183.085 ;
        RECT -57.285 181.395 -56.955 181.725 ;
        RECT -57.285 180.035 -56.955 180.365 ;
        RECT -57.285 178.675 -56.955 179.005 ;
        RECT -57.285 177.315 -56.955 177.645 ;
        RECT -57.285 175.955 -56.955 176.285 ;
        RECT -57.285 174.595 -56.955 174.925 ;
        RECT -57.285 173.235 -56.955 173.565 ;
        RECT -57.285 171.875 -56.955 172.205 ;
        RECT -57.285 170.515 -56.955 170.845 ;
        RECT -57.285 169.155 -56.955 169.485 ;
        RECT -57.285 167.795 -56.955 168.125 ;
        RECT -57.285 166.435 -56.955 166.765 ;
        RECT -57.285 165.075 -56.955 165.405 ;
        RECT -57.285 163.715 -56.955 164.045 ;
        RECT -57.285 162.355 -56.955 162.685 ;
        RECT -57.285 160.995 -56.955 161.325 ;
        RECT -57.285 159.635 -56.955 159.965 ;
        RECT -57.285 158.275 -56.955 158.605 ;
        RECT -57.285 156.915 -56.955 157.245 ;
        RECT -57.285 155.555 -56.955 155.885 ;
        RECT -57.285 154.195 -56.955 154.525 ;
        RECT -57.285 152.835 -56.955 153.165 ;
        RECT -57.285 151.475 -56.955 151.805 ;
        RECT -57.285 150.115 -56.955 150.445 ;
        RECT -57.285 148.755 -56.955 149.085 ;
        RECT -57.285 147.395 -56.955 147.725 ;
        RECT -57.285 146.035 -56.955 146.365 ;
        RECT -57.285 144.675 -56.955 145.005 ;
        RECT -57.285 143.315 -56.955 143.645 ;
        RECT -57.285 141.955 -56.955 142.285 ;
        RECT -57.285 140.595 -56.955 140.925 ;
        RECT -57.285 139.235 -56.955 139.565 ;
        RECT -57.28 138.56 -56.96 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.285 97.075 -56.955 97.405 ;
        RECT -57.285 95.715 -56.955 96.045 ;
        RECT -57.285 94.355 -56.955 94.685 ;
        RECT -57.285 92.995 -56.955 93.325 ;
        RECT -57.285 88.915 -56.955 89.245 ;
        RECT -57.285 84.835 -56.955 85.165 ;
        RECT -57.285 83.475 -56.955 83.805 ;
        RECT -57.285 82.115 -56.955 82.445 ;
        RECT -57.285 80.755 -56.955 81.085 ;
        RECT -57.285 79.395 -56.955 79.725 ;
        RECT -57.285 78.035 -56.955 78.365 ;
        RECT -57.285 76.675 -56.955 77.005 ;
        RECT -57.285 75.315 -56.955 75.645 ;
        RECT -57.285 73.955 -56.955 74.285 ;
        RECT -57.285 72.595 -56.955 72.925 ;
        RECT -57.285 71.235 -56.955 71.565 ;
        RECT -57.285 69.875 -56.955 70.205 ;
        RECT -57.285 68.515 -56.955 68.845 ;
        RECT -57.285 67.155 -56.955 67.485 ;
        RECT -57.285 65.795 -56.955 66.125 ;
        RECT -57.285 64.435 -56.955 64.765 ;
        RECT -57.285 63.075 -56.955 63.405 ;
        RECT -57.285 61.715 -56.955 62.045 ;
        RECT -57.285 60.355 -56.955 60.685 ;
        RECT -57.285 58.995 -56.955 59.325 ;
        RECT -57.285 57.635 -56.955 57.965 ;
        RECT -57.285 56.275 -56.955 56.605 ;
        RECT -57.285 54.915 -56.955 55.245 ;
        RECT -57.285 53.555 -56.955 53.885 ;
        RECT -57.285 52.195 -56.955 52.525 ;
        RECT -57.285 50.835 -56.955 51.165 ;
        RECT -57.285 49.475 -56.955 49.805 ;
        RECT -57.285 48.115 -56.955 48.445 ;
        RECT -57.285 46.755 -56.955 47.085 ;
        RECT -57.285 45.395 -56.955 45.725 ;
        RECT -57.285 44.035 -56.955 44.365 ;
        RECT -57.285 42.675 -56.955 43.005 ;
        RECT -57.285 41.315 -56.955 41.645 ;
        RECT -57.285 39.955 -56.955 40.285 ;
        RECT -57.285 38.595 -56.955 38.925 ;
        RECT -57.285 37.235 -56.955 37.565 ;
        RECT -57.285 35.875 -56.955 36.205 ;
        RECT -57.285 34.515 -56.955 34.845 ;
        RECT -57.285 33.155 -56.955 33.485 ;
        RECT -57.285 31.795 -56.955 32.125 ;
        RECT -57.285 30.435 -56.955 30.765 ;
        RECT -57.285 29.075 -56.955 29.405 ;
        RECT -57.285 27.715 -56.955 28.045 ;
        RECT -57.285 26.355 -56.955 26.685 ;
        RECT -57.285 24.995 -56.955 25.325 ;
        RECT -57.285 23.635 -56.955 23.965 ;
        RECT -57.285 22.275 -56.955 22.605 ;
        RECT -57.285 20.915 -56.955 21.245 ;
        RECT -57.285 19.555 -56.955 19.885 ;
        RECT -57.285 18.195 -56.955 18.525 ;
        RECT -57.285 16.835 -56.955 17.165 ;
        RECT -57.285 15.475 -56.955 15.805 ;
        RECT -57.285 14.115 -56.955 14.445 ;
        RECT -57.285 12.755 -56.955 13.085 ;
        RECT -57.285 11.395 -56.955 11.725 ;
        RECT -57.285 10.035 -56.955 10.365 ;
        RECT -57.285 8.675 -56.955 9.005 ;
        RECT -57.285 7.315 -56.955 7.645 ;
        RECT -57.285 5.955 -56.955 6.285 ;
        RECT -57.285 4.595 -56.955 4.925 ;
        RECT -57.285 3.235 -56.955 3.565 ;
        RECT -57.285 1.875 -56.955 2.205 ;
        RECT -57.285 0.515 -56.955 0.845 ;
        RECT -57.285 -0.845 -56.955 -0.515 ;
        RECT -57.285 -2.205 -56.955 -1.875 ;
        RECT -57.285 -3.565 -56.955 -3.235 ;
        RECT -57.285 -4.925 -56.955 -4.595 ;
        RECT -57.285 -6.285 -56.955 -5.955 ;
        RECT -57.285 -7.645 -56.955 -7.315 ;
        RECT -57.285 -9.005 -56.955 -8.675 ;
        RECT -57.285 -10.365 -56.955 -10.035 ;
        RECT -57.285 -11.725 -56.955 -11.395 ;
        RECT -57.285 -13.085 -56.955 -12.755 ;
        RECT -57.285 -14.445 -56.955 -14.115 ;
        RECT -57.285 -15.805 -56.955 -15.475 ;
        RECT -57.285 -17.165 -56.955 -16.835 ;
        RECT -57.285 -18.525 -56.955 -18.195 ;
        RECT -57.285 -19.885 -56.955 -19.555 ;
        RECT -57.285 -21.245 -56.955 -20.915 ;
        RECT -57.285 -22.605 -56.955 -22.275 ;
        RECT -57.285 -23.965 -56.955 -23.635 ;
        RECT -57.285 -25.325 -56.955 -24.995 ;
        RECT -57.285 -30.765 -56.955 -30.435 ;
        RECT -57.285 -32.125 -56.955 -31.795 ;
        RECT -57.285 -33.485 -56.955 -33.155 ;
        RECT -57.285 -34.845 -56.955 -34.515 ;
        RECT -57.285 -36.205 -56.955 -35.875 ;
        RECT -57.285 -37.565 -56.955 -37.235 ;
        RECT -57.285 -38.925 -56.955 -38.595 ;
        RECT -57.285 -40.285 -56.955 -39.955 ;
        RECT -57.285 -41.645 -56.955 -41.315 ;
        RECT -57.285 -43.005 -56.955 -42.675 ;
        RECT -57.285 -44.365 -56.955 -44.035 ;
        RECT -57.285 -45.725 -56.955 -45.395 ;
        RECT -57.285 -47.085 -56.955 -46.755 ;
        RECT -57.285 -48.445 -56.955 -48.115 ;
        RECT -57.285 -49.805 -56.955 -49.475 ;
        RECT -57.285 -51.165 -56.955 -50.835 ;
        RECT -57.285 -52.525 -56.955 -52.195 ;
        RECT -57.285 -53.885 -56.955 -53.555 ;
        RECT -57.285 -55.245 -56.955 -54.915 ;
        RECT -57.285 -56.605 -56.955 -56.275 ;
        RECT -57.285 -57.965 -56.955 -57.635 ;
        RECT -57.285 -59.325 -56.955 -58.995 ;
        RECT -57.285 -60.685 -56.955 -60.355 ;
        RECT -57.285 -62.045 -56.955 -61.715 ;
        RECT -57.285 -63.405 -56.955 -63.075 ;
        RECT -57.285 -64.765 -56.955 -64.435 ;
        RECT -57.285 -66.125 -56.955 -65.795 ;
        RECT -57.285 -67.485 -56.955 -67.155 ;
        RECT -57.285 -68.845 -56.955 -68.515 ;
        RECT -57.285 -70.205 -56.955 -69.875 ;
        RECT -57.285 -71.565 -56.955 -71.235 ;
        RECT -57.285 -72.925 -56.955 -72.595 ;
        RECT -57.285 -74.285 -56.955 -73.955 ;
        RECT -57.285 -75.645 -56.955 -75.315 ;
        RECT -57.285 -77.005 -56.955 -76.675 ;
        RECT -57.285 -78.365 -56.955 -78.035 ;
        RECT -57.285 -79.725 -56.955 -79.395 ;
        RECT -57.285 -81.085 -56.955 -80.755 ;
        RECT -57.285 -82.445 -56.955 -82.115 ;
        RECT -57.285 -83.805 -56.955 -83.475 ;
        RECT -57.285 -85.165 -56.955 -84.835 ;
        RECT -57.285 -86.525 -56.955 -86.195 ;
        RECT -57.285 -87.885 -56.955 -87.555 ;
        RECT -57.285 -89.245 -56.955 -88.915 ;
        RECT -57.285 -90.605 -56.955 -90.275 ;
        RECT -57.285 -91.77 -56.955 -91.44 ;
        RECT -57.285 -93.325 -56.955 -92.995 ;
        RECT -57.285 -94.685 -56.955 -94.355 ;
        RECT -57.285 -96.045 -56.955 -95.715 ;
        RECT -57.285 -97.405 -56.955 -97.075 ;
        RECT -57.285 -98.765 -56.955 -98.435 ;
        RECT -57.285 -101.485 -56.955 -101.155 ;
        RECT -57.285 -102.31 -56.955 -101.98 ;
        RECT -57.285 -104.205 -56.955 -103.875 ;
        RECT -57.285 -105.565 -56.955 -105.235 ;
        RECT -57.285 -106.925 -56.955 -106.595 ;
        RECT -57.285 -109.645 -56.955 -109.315 ;
        RECT -57.285 -111.005 -56.955 -110.675 ;
        RECT -57.285 -113.725 -56.955 -113.395 ;
        RECT -57.285 -115.085 -56.955 -114.755 ;
        RECT -57.285 -116.445 -56.955 -116.115 ;
        RECT -57.285 -117.805 -56.955 -117.475 ;
        RECT -57.285 -119.165 -56.955 -118.835 ;
        RECT -57.285 -120.525 -56.955 -120.195 ;
        RECT -57.285 -123.245 -56.955 -122.915 ;
        RECT -57.285 -124.605 -56.955 -124.275 ;
        RECT -57.285 -125.965 -56.955 -125.635 ;
        RECT -57.285 -127.325 -56.955 -126.995 ;
        RECT -57.285 -128.685 -56.955 -128.355 ;
        RECT -57.285 -130.045 -56.955 -129.715 ;
        RECT -57.285 -131.405 -56.955 -131.075 ;
        RECT -57.285 -132.765 -56.955 -132.435 ;
        RECT -57.285 -134.125 -56.955 -133.795 ;
        RECT -57.285 -135.485 -56.955 -135.155 ;
        RECT -57.285 -136.845 -56.955 -136.515 ;
        RECT -57.285 -138.205 -56.955 -137.875 ;
        RECT -57.285 -139.565 -56.955 -139.235 ;
        RECT -57.285 -140.925 -56.955 -140.595 ;
        RECT -57.285 -142.285 -56.955 -141.955 ;
        RECT -57.285 -143.645 -56.955 -143.315 ;
        RECT -57.285 -145.005 -56.955 -144.675 ;
        RECT -57.285 -146.365 -56.955 -146.035 ;
        RECT -57.285 -147.725 -56.955 -147.395 ;
        RECT -57.285 -149.085 -56.955 -148.755 ;
        RECT -57.285 -150.445 -56.955 -150.115 ;
        RECT -57.285 -151.805 -56.955 -151.475 ;
        RECT -57.285 -153.165 -56.955 -152.835 ;
        RECT -57.285 -154.525 -56.955 -154.195 ;
        RECT -57.285 -155.885 -56.955 -155.555 ;
        RECT -57.285 -157.245 -56.955 -156.915 ;
        RECT -57.285 -158.605 -56.955 -158.275 ;
        RECT -57.285 -159.965 -56.955 -159.635 ;
        RECT -57.285 -161.325 -56.955 -160.995 ;
        RECT -57.285 -162.685 -56.955 -162.355 ;
        RECT -57.285 -164.045 -56.955 -163.715 ;
        RECT -57.285 -165.405 -56.955 -165.075 ;
        RECT -57.285 -166.765 -56.955 -166.435 ;
        RECT -57.28 -167.44 -56.96 98.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.285 -174.925 -56.955 -174.595 ;
        RECT -57.285 -177.645 -56.955 -177.315 ;
        RECT -57.285 -179.005 -56.955 -178.675 ;
        RECT -57.285 -184.65 -56.955 -183.52 ;
        RECT -57.28 -184.765 -56.96 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.925 244.04 -55.595 245.17 ;
        RECT -55.925 239.875 -55.595 240.205 ;
        RECT -55.925 238.515 -55.595 238.845 ;
        RECT -55.925 237.155 -55.595 237.485 ;
        RECT -55.925 235.795 -55.595 236.125 ;
        RECT -55.925 234.435 -55.595 234.765 ;
        RECT -55.925 233.075 -55.595 233.405 ;
        RECT -55.925 231.715 -55.595 232.045 ;
        RECT -55.925 230.355 -55.595 230.685 ;
        RECT -55.925 228.995 -55.595 229.325 ;
        RECT -55.925 227.635 -55.595 227.965 ;
        RECT -55.925 226.275 -55.595 226.605 ;
        RECT -55.925 224.915 -55.595 225.245 ;
        RECT -55.925 223.555 -55.595 223.885 ;
        RECT -55.925 222.195 -55.595 222.525 ;
        RECT -55.925 220.835 -55.595 221.165 ;
        RECT -55.925 219.475 -55.595 219.805 ;
        RECT -55.925 218.115 -55.595 218.445 ;
        RECT -55.925 216.755 -55.595 217.085 ;
        RECT -55.925 215.395 -55.595 215.725 ;
        RECT -55.925 214.035 -55.595 214.365 ;
        RECT -55.925 212.675 -55.595 213.005 ;
        RECT -55.925 211.315 -55.595 211.645 ;
        RECT -55.925 209.955 -55.595 210.285 ;
        RECT -55.925 208.595 -55.595 208.925 ;
        RECT -55.925 207.235 -55.595 207.565 ;
        RECT -55.925 205.875 -55.595 206.205 ;
        RECT -55.925 204.515 -55.595 204.845 ;
        RECT -55.925 203.155 -55.595 203.485 ;
        RECT -55.925 201.795 -55.595 202.125 ;
        RECT -55.925 200.435 -55.595 200.765 ;
        RECT -55.925 199.075 -55.595 199.405 ;
        RECT -55.925 197.715 -55.595 198.045 ;
        RECT -55.925 196.355 -55.595 196.685 ;
        RECT -55.925 194.995 -55.595 195.325 ;
        RECT -55.925 193.635 -55.595 193.965 ;
        RECT -55.925 192.275 -55.595 192.605 ;
        RECT -55.925 190.915 -55.595 191.245 ;
        RECT -55.925 189.555 -55.595 189.885 ;
        RECT -55.925 188.195 -55.595 188.525 ;
        RECT -55.925 186.835 -55.595 187.165 ;
        RECT -55.925 185.475 -55.595 185.805 ;
        RECT -55.925 184.115 -55.595 184.445 ;
        RECT -55.925 182.755 -55.595 183.085 ;
        RECT -55.925 181.395 -55.595 181.725 ;
        RECT -55.925 180.035 -55.595 180.365 ;
        RECT -55.925 178.675 -55.595 179.005 ;
        RECT -55.925 177.315 -55.595 177.645 ;
        RECT -55.925 175.955 -55.595 176.285 ;
        RECT -55.925 174.595 -55.595 174.925 ;
        RECT -55.925 173.235 -55.595 173.565 ;
        RECT -55.925 171.875 -55.595 172.205 ;
        RECT -55.925 170.515 -55.595 170.845 ;
        RECT -55.925 169.155 -55.595 169.485 ;
        RECT -55.925 167.795 -55.595 168.125 ;
        RECT -55.925 166.435 -55.595 166.765 ;
        RECT -55.925 165.075 -55.595 165.405 ;
        RECT -55.925 163.715 -55.595 164.045 ;
        RECT -55.925 162.355 -55.595 162.685 ;
        RECT -55.925 160.995 -55.595 161.325 ;
        RECT -55.925 159.635 -55.595 159.965 ;
        RECT -55.925 158.275 -55.595 158.605 ;
        RECT -55.925 156.915 -55.595 157.245 ;
        RECT -55.925 155.555 -55.595 155.885 ;
        RECT -55.925 154.195 -55.595 154.525 ;
        RECT -55.925 152.835 -55.595 153.165 ;
        RECT -55.925 151.475 -55.595 151.805 ;
        RECT -55.925 150.115 -55.595 150.445 ;
        RECT -55.925 148.755 -55.595 149.085 ;
        RECT -55.925 147.395 -55.595 147.725 ;
        RECT -55.925 146.035 -55.595 146.365 ;
        RECT -55.925 144.675 -55.595 145.005 ;
        RECT -55.925 143.315 -55.595 143.645 ;
        RECT -55.925 141.955 -55.595 142.285 ;
        RECT -55.925 140.595 -55.595 140.925 ;
        RECT -55.925 139.235 -55.595 139.565 ;
        RECT -55.92 138.56 -55.6 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.925 97.075 -55.595 97.405 ;
        RECT -55.925 95.715 -55.595 96.045 ;
        RECT -55.925 94.355 -55.595 94.685 ;
        RECT -55.925 92.995 -55.595 93.325 ;
        RECT -55.925 88.915 -55.595 89.245 ;
        RECT -55.925 84.835 -55.595 85.165 ;
        RECT -55.925 83.475 -55.595 83.805 ;
        RECT -55.925 82.115 -55.595 82.445 ;
        RECT -55.925 80.755 -55.595 81.085 ;
        RECT -55.925 79.395 -55.595 79.725 ;
        RECT -55.925 78.035 -55.595 78.365 ;
        RECT -55.925 76.675 -55.595 77.005 ;
        RECT -55.925 75.315 -55.595 75.645 ;
        RECT -55.925 73.955 -55.595 74.285 ;
        RECT -55.925 72.595 -55.595 72.925 ;
        RECT -55.925 71.235 -55.595 71.565 ;
        RECT -55.925 69.875 -55.595 70.205 ;
        RECT -55.925 68.515 -55.595 68.845 ;
        RECT -55.925 67.155 -55.595 67.485 ;
        RECT -55.925 65.795 -55.595 66.125 ;
        RECT -55.925 64.435 -55.595 64.765 ;
        RECT -55.925 63.075 -55.595 63.405 ;
        RECT -55.925 61.715 -55.595 62.045 ;
        RECT -55.925 60.355 -55.595 60.685 ;
        RECT -55.925 58.995 -55.595 59.325 ;
        RECT -55.925 57.635 -55.595 57.965 ;
        RECT -55.925 56.275 -55.595 56.605 ;
        RECT -55.925 54.915 -55.595 55.245 ;
        RECT -55.925 53.555 -55.595 53.885 ;
        RECT -55.925 52.195 -55.595 52.525 ;
        RECT -55.925 50.835 -55.595 51.165 ;
        RECT -55.925 49.475 -55.595 49.805 ;
        RECT -55.925 48.115 -55.595 48.445 ;
        RECT -55.925 46.755 -55.595 47.085 ;
        RECT -55.925 45.395 -55.595 45.725 ;
        RECT -55.925 44.035 -55.595 44.365 ;
        RECT -55.925 42.675 -55.595 43.005 ;
        RECT -55.925 41.315 -55.595 41.645 ;
        RECT -55.925 39.955 -55.595 40.285 ;
        RECT -55.925 38.595 -55.595 38.925 ;
        RECT -55.925 37.235 -55.595 37.565 ;
        RECT -55.925 35.875 -55.595 36.205 ;
        RECT -55.925 34.515 -55.595 34.845 ;
        RECT -55.925 33.155 -55.595 33.485 ;
        RECT -55.925 31.795 -55.595 32.125 ;
        RECT -55.925 30.435 -55.595 30.765 ;
        RECT -55.925 29.075 -55.595 29.405 ;
        RECT -55.925 27.715 -55.595 28.045 ;
        RECT -55.925 26.355 -55.595 26.685 ;
        RECT -55.925 24.995 -55.595 25.325 ;
        RECT -55.925 23.635 -55.595 23.965 ;
        RECT -55.925 22.275 -55.595 22.605 ;
        RECT -55.925 20.915 -55.595 21.245 ;
        RECT -55.925 19.555 -55.595 19.885 ;
        RECT -55.925 18.195 -55.595 18.525 ;
        RECT -55.925 16.835 -55.595 17.165 ;
        RECT -55.925 15.475 -55.595 15.805 ;
        RECT -55.925 14.115 -55.595 14.445 ;
        RECT -55.925 12.755 -55.595 13.085 ;
        RECT -55.925 11.395 -55.595 11.725 ;
        RECT -55.925 10.035 -55.595 10.365 ;
        RECT -55.925 8.675 -55.595 9.005 ;
        RECT -55.925 7.315 -55.595 7.645 ;
        RECT -55.925 5.955 -55.595 6.285 ;
        RECT -55.925 4.595 -55.595 4.925 ;
        RECT -55.925 3.235 -55.595 3.565 ;
        RECT -55.925 1.875 -55.595 2.205 ;
        RECT -55.925 0.515 -55.595 0.845 ;
        RECT -55.925 -0.845 -55.595 -0.515 ;
        RECT -55.925 -2.205 -55.595 -1.875 ;
        RECT -55.925 -3.565 -55.595 -3.235 ;
        RECT -55.925 -4.925 -55.595 -4.595 ;
        RECT -55.925 -6.285 -55.595 -5.955 ;
        RECT -55.925 -7.645 -55.595 -7.315 ;
        RECT -55.925 -9.005 -55.595 -8.675 ;
        RECT -55.925 -10.365 -55.595 -10.035 ;
        RECT -55.925 -11.725 -55.595 -11.395 ;
        RECT -55.925 -13.085 -55.595 -12.755 ;
        RECT -55.925 -14.445 -55.595 -14.115 ;
        RECT -55.925 -15.805 -55.595 -15.475 ;
        RECT -55.925 -17.165 -55.595 -16.835 ;
        RECT -55.925 -18.525 -55.595 -18.195 ;
        RECT -55.925 -19.885 -55.595 -19.555 ;
        RECT -55.925 -21.245 -55.595 -20.915 ;
        RECT -55.925 -22.605 -55.595 -22.275 ;
        RECT -55.925 -23.965 -55.595 -23.635 ;
        RECT -55.925 -25.325 -55.595 -24.995 ;
        RECT -55.925 -30.765 -55.595 -30.435 ;
        RECT -55.925 -32.125 -55.595 -31.795 ;
        RECT -55.925 -33.485 -55.595 -33.155 ;
        RECT -55.925 -34.845 -55.595 -34.515 ;
        RECT -55.925 -36.205 -55.595 -35.875 ;
        RECT -55.925 -37.565 -55.595 -37.235 ;
        RECT -55.925 -38.925 -55.595 -38.595 ;
        RECT -55.925 -40.285 -55.595 -39.955 ;
        RECT -55.925 -41.645 -55.595 -41.315 ;
        RECT -55.925 -43.005 -55.595 -42.675 ;
        RECT -55.925 -44.365 -55.595 -44.035 ;
        RECT -55.925 -45.725 -55.595 -45.395 ;
        RECT -55.925 -47.085 -55.595 -46.755 ;
        RECT -55.925 -48.445 -55.595 -48.115 ;
        RECT -55.925 -49.805 -55.595 -49.475 ;
        RECT -55.925 -51.165 -55.595 -50.835 ;
        RECT -55.925 -52.525 -55.595 -52.195 ;
        RECT -55.925 -53.885 -55.595 -53.555 ;
        RECT -55.925 -55.245 -55.595 -54.915 ;
        RECT -55.925 -56.605 -55.595 -56.275 ;
        RECT -55.925 -57.965 -55.595 -57.635 ;
        RECT -55.925 -59.325 -55.595 -58.995 ;
        RECT -55.925 -60.685 -55.595 -60.355 ;
        RECT -55.925 -62.045 -55.595 -61.715 ;
        RECT -55.925 -63.405 -55.595 -63.075 ;
        RECT -55.925 -64.765 -55.595 -64.435 ;
        RECT -55.925 -66.125 -55.595 -65.795 ;
        RECT -55.925 -67.485 -55.595 -67.155 ;
        RECT -55.925 -68.845 -55.595 -68.515 ;
        RECT -55.925 -70.205 -55.595 -69.875 ;
        RECT -55.925 -71.565 -55.595 -71.235 ;
        RECT -55.925 -72.925 -55.595 -72.595 ;
        RECT -55.925 -74.285 -55.595 -73.955 ;
        RECT -55.925 -75.645 -55.595 -75.315 ;
        RECT -55.925 -77.005 -55.595 -76.675 ;
        RECT -55.925 -78.365 -55.595 -78.035 ;
        RECT -55.925 -79.725 -55.595 -79.395 ;
        RECT -55.925 -81.085 -55.595 -80.755 ;
        RECT -55.925 -82.445 -55.595 -82.115 ;
        RECT -55.925 -83.805 -55.595 -83.475 ;
        RECT -55.925 -85.165 -55.595 -84.835 ;
        RECT -55.925 -86.525 -55.595 -86.195 ;
        RECT -55.925 -87.885 -55.595 -87.555 ;
        RECT -55.925 -89.245 -55.595 -88.915 ;
        RECT -55.925 -90.605 -55.595 -90.275 ;
        RECT -55.925 -91.77 -55.595 -91.44 ;
        RECT -55.925 -93.325 -55.595 -92.995 ;
        RECT -55.925 -94.685 -55.595 -94.355 ;
        RECT -55.925 -96.045 -55.595 -95.715 ;
        RECT -55.925 -97.405 -55.595 -97.075 ;
        RECT -55.925 -98.765 -55.595 -98.435 ;
        RECT -55.925 -101.485 -55.595 -101.155 ;
        RECT -55.925 -102.31 -55.595 -101.98 ;
        RECT -55.925 -104.205 -55.595 -103.875 ;
        RECT -55.925 -105.565 -55.595 -105.235 ;
        RECT -55.925 -106.925 -55.595 -106.595 ;
        RECT -55.925 -109.645 -55.595 -109.315 ;
        RECT -55.925 -111.005 -55.595 -110.675 ;
        RECT -55.925 -113.725 -55.595 -113.395 ;
        RECT -55.925 -115.085 -55.595 -114.755 ;
        RECT -55.925 -116.445 -55.595 -116.115 ;
        RECT -55.925 -117.805 -55.595 -117.475 ;
        RECT -55.925 -119.165 -55.595 -118.835 ;
        RECT -55.925 -120.525 -55.595 -120.195 ;
        RECT -55.925 -123.245 -55.595 -122.915 ;
        RECT -55.925 -124.605 -55.595 -124.275 ;
        RECT -55.925 -125.965 -55.595 -125.635 ;
        RECT -55.925 -127.325 -55.595 -126.995 ;
        RECT -55.925 -128.685 -55.595 -128.355 ;
        RECT -55.925 -130.045 -55.595 -129.715 ;
        RECT -55.925 -131.405 -55.595 -131.075 ;
        RECT -55.925 -132.765 -55.595 -132.435 ;
        RECT -55.925 -134.125 -55.595 -133.795 ;
        RECT -55.925 -135.485 -55.595 -135.155 ;
        RECT -55.925 -136.845 -55.595 -136.515 ;
        RECT -55.925 -138.205 -55.595 -137.875 ;
        RECT -55.925 -139.565 -55.595 -139.235 ;
        RECT -55.925 -140.925 -55.595 -140.595 ;
        RECT -55.925 -142.285 -55.595 -141.955 ;
        RECT -55.925 -143.645 -55.595 -143.315 ;
        RECT -55.925 -145.005 -55.595 -144.675 ;
        RECT -55.925 -146.365 -55.595 -146.035 ;
        RECT -55.925 -147.725 -55.595 -147.395 ;
        RECT -55.925 -149.085 -55.595 -148.755 ;
        RECT -55.925 -150.445 -55.595 -150.115 ;
        RECT -55.925 -151.805 -55.595 -151.475 ;
        RECT -55.925 -153.165 -55.595 -152.835 ;
        RECT -55.925 -154.525 -55.595 -154.195 ;
        RECT -55.925 -155.885 -55.595 -155.555 ;
        RECT -55.925 -157.245 -55.595 -156.915 ;
        RECT -55.925 -158.605 -55.595 -158.275 ;
        RECT -55.925 -159.965 -55.595 -159.635 ;
        RECT -55.925 -161.325 -55.595 -160.995 ;
        RECT -55.925 -162.685 -55.595 -162.355 ;
        RECT -55.925 -164.045 -55.595 -163.715 ;
        RECT -55.925 -165.405 -55.595 -165.075 ;
        RECT -55.925 -166.765 -55.595 -166.435 ;
        RECT -55.925 -169.615 -55.595 -169.285 ;
        RECT -55.925 -170.845 -55.595 -170.515 ;
        RECT -55.925 -172.205 -55.595 -171.875 ;
        RECT -55.925 -173.565 -55.595 -173.235 ;
        RECT -55.925 -174.925 -55.595 -174.595 ;
        RECT -55.925 -177.645 -55.595 -177.315 ;
        RECT -55.925 -179.005 -55.595 -178.675 ;
        RECT -55.925 -184.65 -55.595 -183.52 ;
        RECT -55.92 -184.765 -55.6 98.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 244.04 -54.235 245.17 ;
        RECT -54.565 239.875 -54.235 240.205 ;
        RECT -54.565 238.515 -54.235 238.845 ;
        RECT -54.565 237.155 -54.235 237.485 ;
        RECT -54.565 235.795 -54.235 236.125 ;
        RECT -54.565 234.435 -54.235 234.765 ;
        RECT -54.565 233.075 -54.235 233.405 ;
        RECT -54.565 231.715 -54.235 232.045 ;
        RECT -54.565 230.355 -54.235 230.685 ;
        RECT -54.565 228.995 -54.235 229.325 ;
        RECT -54.565 227.635 -54.235 227.965 ;
        RECT -54.565 226.275 -54.235 226.605 ;
        RECT -54.565 224.915 -54.235 225.245 ;
        RECT -54.565 223.555 -54.235 223.885 ;
        RECT -54.565 222.195 -54.235 222.525 ;
        RECT -54.565 220.835 -54.235 221.165 ;
        RECT -54.565 219.475 -54.235 219.805 ;
        RECT -54.565 218.115 -54.235 218.445 ;
        RECT -54.565 216.755 -54.235 217.085 ;
        RECT -54.565 215.395 -54.235 215.725 ;
        RECT -54.565 214.035 -54.235 214.365 ;
        RECT -54.565 212.675 -54.235 213.005 ;
        RECT -54.565 211.315 -54.235 211.645 ;
        RECT -54.565 209.955 -54.235 210.285 ;
        RECT -54.565 208.595 -54.235 208.925 ;
        RECT -54.565 207.235 -54.235 207.565 ;
        RECT -54.565 205.875 -54.235 206.205 ;
        RECT -54.565 204.515 -54.235 204.845 ;
        RECT -54.565 203.155 -54.235 203.485 ;
        RECT -54.565 201.795 -54.235 202.125 ;
        RECT -54.565 200.435 -54.235 200.765 ;
        RECT -54.565 199.075 -54.235 199.405 ;
        RECT -54.565 197.715 -54.235 198.045 ;
        RECT -54.565 196.355 -54.235 196.685 ;
        RECT -54.565 194.995 -54.235 195.325 ;
        RECT -54.565 193.635 -54.235 193.965 ;
        RECT -54.565 192.275 -54.235 192.605 ;
        RECT -54.565 190.915 -54.235 191.245 ;
        RECT -54.565 189.555 -54.235 189.885 ;
        RECT -54.565 188.195 -54.235 188.525 ;
        RECT -54.565 186.835 -54.235 187.165 ;
        RECT -54.565 185.475 -54.235 185.805 ;
        RECT -54.565 184.115 -54.235 184.445 ;
        RECT -54.565 182.755 -54.235 183.085 ;
        RECT -54.565 181.395 -54.235 181.725 ;
        RECT -54.565 180.035 -54.235 180.365 ;
        RECT -54.565 178.675 -54.235 179.005 ;
        RECT -54.565 177.315 -54.235 177.645 ;
        RECT -54.565 175.955 -54.235 176.285 ;
        RECT -54.565 174.595 -54.235 174.925 ;
        RECT -54.565 173.235 -54.235 173.565 ;
        RECT -54.565 171.875 -54.235 172.205 ;
        RECT -54.565 170.515 -54.235 170.845 ;
        RECT -54.565 169.155 -54.235 169.485 ;
        RECT -54.565 167.795 -54.235 168.125 ;
        RECT -54.565 166.435 -54.235 166.765 ;
        RECT -54.565 165.075 -54.235 165.405 ;
        RECT -54.565 163.715 -54.235 164.045 ;
        RECT -54.565 162.355 -54.235 162.685 ;
        RECT -54.565 160.995 -54.235 161.325 ;
        RECT -54.565 159.635 -54.235 159.965 ;
        RECT -54.565 158.275 -54.235 158.605 ;
        RECT -54.565 156.915 -54.235 157.245 ;
        RECT -54.565 155.555 -54.235 155.885 ;
        RECT -54.565 154.195 -54.235 154.525 ;
        RECT -54.565 152.835 -54.235 153.165 ;
        RECT -54.565 151.475 -54.235 151.805 ;
        RECT -54.565 150.115 -54.235 150.445 ;
        RECT -54.565 148.755 -54.235 149.085 ;
        RECT -54.565 147.395 -54.235 147.725 ;
        RECT -54.565 146.035 -54.235 146.365 ;
        RECT -54.565 144.675 -54.235 145.005 ;
        RECT -54.565 143.315 -54.235 143.645 ;
        RECT -54.565 141.955 -54.235 142.285 ;
        RECT -54.565 140.595 -54.235 140.925 ;
        RECT -54.565 139.235 -54.235 139.565 ;
        RECT -54.56 138.56 -54.24 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 97.075 -54.235 97.405 ;
        RECT -54.565 95.715 -54.235 96.045 ;
        RECT -54.565 94.355 -54.235 94.685 ;
        RECT -54.565 92.995 -54.235 93.325 ;
        RECT -54.565 88.915 -54.235 89.245 ;
        RECT -54.565 84.835 -54.235 85.165 ;
        RECT -54.565 83.475 -54.235 83.805 ;
        RECT -54.565 82.115 -54.235 82.445 ;
        RECT -54.565 80.755 -54.235 81.085 ;
        RECT -54.565 79.395 -54.235 79.725 ;
        RECT -54.565 78.035 -54.235 78.365 ;
        RECT -54.565 76.675 -54.235 77.005 ;
        RECT -54.565 75.315 -54.235 75.645 ;
        RECT -54.565 73.955 -54.235 74.285 ;
        RECT -54.565 72.595 -54.235 72.925 ;
        RECT -54.565 71.235 -54.235 71.565 ;
        RECT -54.565 69.875 -54.235 70.205 ;
        RECT -54.565 68.515 -54.235 68.845 ;
        RECT -54.565 67.155 -54.235 67.485 ;
        RECT -54.565 65.795 -54.235 66.125 ;
        RECT -54.565 64.435 -54.235 64.765 ;
        RECT -54.565 63.075 -54.235 63.405 ;
        RECT -54.565 61.715 -54.235 62.045 ;
        RECT -54.565 60.355 -54.235 60.685 ;
        RECT -54.565 58.995 -54.235 59.325 ;
        RECT -54.565 57.635 -54.235 57.965 ;
        RECT -54.565 56.275 -54.235 56.605 ;
        RECT -54.565 54.915 -54.235 55.245 ;
        RECT -54.565 53.555 -54.235 53.885 ;
        RECT -54.565 52.195 -54.235 52.525 ;
        RECT -54.565 50.835 -54.235 51.165 ;
        RECT -54.565 49.475 -54.235 49.805 ;
        RECT -54.565 48.115 -54.235 48.445 ;
        RECT -54.565 46.755 -54.235 47.085 ;
        RECT -54.565 45.395 -54.235 45.725 ;
        RECT -54.565 44.035 -54.235 44.365 ;
        RECT -54.565 42.675 -54.235 43.005 ;
        RECT -54.565 41.315 -54.235 41.645 ;
        RECT -54.565 39.955 -54.235 40.285 ;
        RECT -54.565 38.595 -54.235 38.925 ;
        RECT -54.565 37.235 -54.235 37.565 ;
        RECT -54.565 35.875 -54.235 36.205 ;
        RECT -54.565 34.515 -54.235 34.845 ;
        RECT -54.565 33.155 -54.235 33.485 ;
        RECT -54.565 31.795 -54.235 32.125 ;
        RECT -54.565 30.435 -54.235 30.765 ;
        RECT -54.565 29.075 -54.235 29.405 ;
        RECT -54.565 27.715 -54.235 28.045 ;
        RECT -54.565 26.355 -54.235 26.685 ;
        RECT -54.565 24.995 -54.235 25.325 ;
        RECT -54.565 23.635 -54.235 23.965 ;
        RECT -54.565 22.275 -54.235 22.605 ;
        RECT -54.565 20.915 -54.235 21.245 ;
        RECT -54.565 19.555 -54.235 19.885 ;
        RECT -54.565 18.195 -54.235 18.525 ;
        RECT -54.565 16.835 -54.235 17.165 ;
        RECT -54.565 15.475 -54.235 15.805 ;
        RECT -54.565 14.115 -54.235 14.445 ;
        RECT -54.565 12.755 -54.235 13.085 ;
        RECT -54.565 11.395 -54.235 11.725 ;
        RECT -54.565 10.035 -54.235 10.365 ;
        RECT -54.565 8.675 -54.235 9.005 ;
        RECT -54.565 7.315 -54.235 7.645 ;
        RECT -54.565 5.955 -54.235 6.285 ;
        RECT -54.565 4.595 -54.235 4.925 ;
        RECT -54.565 3.235 -54.235 3.565 ;
        RECT -54.565 1.875 -54.235 2.205 ;
        RECT -54.565 0.515 -54.235 0.845 ;
        RECT -54.565 -0.845 -54.235 -0.515 ;
        RECT -54.565 -2.205 -54.235 -1.875 ;
        RECT -54.565 -3.565 -54.235 -3.235 ;
        RECT -54.565 -4.925 -54.235 -4.595 ;
        RECT -54.565 -6.285 -54.235 -5.955 ;
        RECT -54.565 -7.645 -54.235 -7.315 ;
        RECT -54.565 -9.005 -54.235 -8.675 ;
        RECT -54.565 -10.365 -54.235 -10.035 ;
        RECT -54.565 -11.725 -54.235 -11.395 ;
        RECT -54.565 -13.085 -54.235 -12.755 ;
        RECT -54.565 -14.445 -54.235 -14.115 ;
        RECT -54.565 -15.805 -54.235 -15.475 ;
        RECT -54.565 -17.165 -54.235 -16.835 ;
        RECT -54.565 -18.525 -54.235 -18.195 ;
        RECT -54.565 -19.885 -54.235 -19.555 ;
        RECT -54.565 -21.245 -54.235 -20.915 ;
        RECT -54.565 -22.605 -54.235 -22.275 ;
        RECT -54.565 -23.965 -54.235 -23.635 ;
        RECT -54.565 -25.325 -54.235 -24.995 ;
        RECT -54.565 -30.765 -54.235 -30.435 ;
        RECT -54.565 -32.125 -54.235 -31.795 ;
        RECT -54.565 -33.485 -54.235 -33.155 ;
        RECT -54.565 -34.845 -54.235 -34.515 ;
        RECT -54.565 -36.205 -54.235 -35.875 ;
        RECT -54.565 -37.565 -54.235 -37.235 ;
        RECT -54.565 -38.925 -54.235 -38.595 ;
        RECT -54.565 -40.285 -54.235 -39.955 ;
        RECT -54.565 -41.645 -54.235 -41.315 ;
        RECT -54.565 -43.005 -54.235 -42.675 ;
        RECT -54.565 -44.365 -54.235 -44.035 ;
        RECT -54.565 -45.725 -54.235 -45.395 ;
        RECT -54.565 -47.085 -54.235 -46.755 ;
        RECT -54.565 -48.445 -54.235 -48.115 ;
        RECT -54.565 -49.805 -54.235 -49.475 ;
        RECT -54.565 -51.165 -54.235 -50.835 ;
        RECT -54.565 -52.525 -54.235 -52.195 ;
        RECT -54.565 -53.885 -54.235 -53.555 ;
        RECT -54.565 -55.245 -54.235 -54.915 ;
        RECT -54.565 -56.605 -54.235 -56.275 ;
        RECT -54.565 -57.965 -54.235 -57.635 ;
        RECT -54.565 -59.325 -54.235 -58.995 ;
        RECT -54.565 -60.685 -54.235 -60.355 ;
        RECT -54.565 -62.045 -54.235 -61.715 ;
        RECT -54.565 -63.405 -54.235 -63.075 ;
        RECT -54.565 -64.765 -54.235 -64.435 ;
        RECT -54.565 -66.125 -54.235 -65.795 ;
        RECT -54.565 -67.485 -54.235 -67.155 ;
        RECT -54.565 -68.845 -54.235 -68.515 ;
        RECT -54.565 -70.205 -54.235 -69.875 ;
        RECT -54.565 -71.565 -54.235 -71.235 ;
        RECT -54.565 -72.925 -54.235 -72.595 ;
        RECT -54.565 -74.285 -54.235 -73.955 ;
        RECT -54.565 -75.645 -54.235 -75.315 ;
        RECT -54.565 -77.005 -54.235 -76.675 ;
        RECT -54.565 -78.365 -54.235 -78.035 ;
        RECT -54.565 -79.725 -54.235 -79.395 ;
        RECT -54.565 -81.085 -54.235 -80.755 ;
        RECT -54.565 -82.445 -54.235 -82.115 ;
        RECT -54.565 -83.805 -54.235 -83.475 ;
        RECT -54.565 -85.165 -54.235 -84.835 ;
        RECT -54.565 -86.525 -54.235 -86.195 ;
        RECT -54.565 -87.885 -54.235 -87.555 ;
        RECT -54.565 -89.245 -54.235 -88.915 ;
        RECT -54.565 -90.605 -54.235 -90.275 ;
        RECT -54.565 -91.77 -54.235 -91.44 ;
        RECT -54.565 -93.325 -54.235 -92.995 ;
        RECT -54.565 -94.685 -54.235 -94.355 ;
        RECT -54.565 -96.045 -54.235 -95.715 ;
        RECT -54.565 -97.405 -54.235 -97.075 ;
        RECT -54.565 -98.765 -54.235 -98.435 ;
        RECT -54.565 -101.485 -54.235 -101.155 ;
        RECT -54.565 -102.31 -54.235 -101.98 ;
        RECT -54.565 -104.205 -54.235 -103.875 ;
        RECT -54.565 -105.565 -54.235 -105.235 ;
        RECT -54.565 -106.925 -54.235 -106.595 ;
        RECT -54.565 -109.645 -54.235 -109.315 ;
        RECT -54.565 -111.005 -54.235 -110.675 ;
        RECT -54.565 -113.725 -54.235 -113.395 ;
        RECT -54.56 -113.725 -54.24 98.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -54.565 -177.645 -54.235 -177.315 ;
        RECT -54.565 -179.005 -54.235 -178.675 ;
        RECT -54.565 -184.65 -54.235 -183.52 ;
        RECT -54.56 -184.765 -54.24 -175.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.205 244.04 -52.875 245.17 ;
        RECT -53.205 239.875 -52.875 240.205 ;
        RECT -53.205 238.515 -52.875 238.845 ;
        RECT -53.205 237.155 -52.875 237.485 ;
        RECT -53.205 235.795 -52.875 236.125 ;
        RECT -53.205 234.435 -52.875 234.765 ;
        RECT -53.205 233.075 -52.875 233.405 ;
        RECT -53.205 231.715 -52.875 232.045 ;
        RECT -53.205 230.355 -52.875 230.685 ;
        RECT -53.205 228.995 -52.875 229.325 ;
        RECT -53.205 227.635 -52.875 227.965 ;
        RECT -53.205 226.275 -52.875 226.605 ;
        RECT -53.205 224.915 -52.875 225.245 ;
        RECT -53.205 223.555 -52.875 223.885 ;
        RECT -53.205 222.195 -52.875 222.525 ;
        RECT -53.205 220.835 -52.875 221.165 ;
        RECT -53.205 219.475 -52.875 219.805 ;
        RECT -53.205 218.115 -52.875 218.445 ;
        RECT -53.205 216.755 -52.875 217.085 ;
        RECT -53.205 215.395 -52.875 215.725 ;
        RECT -53.205 214.035 -52.875 214.365 ;
        RECT -53.205 212.675 -52.875 213.005 ;
        RECT -53.205 211.315 -52.875 211.645 ;
        RECT -53.205 209.955 -52.875 210.285 ;
        RECT -53.205 208.595 -52.875 208.925 ;
        RECT -53.205 207.235 -52.875 207.565 ;
        RECT -53.205 205.875 -52.875 206.205 ;
        RECT -53.205 204.515 -52.875 204.845 ;
        RECT -53.205 203.155 -52.875 203.485 ;
        RECT -53.205 201.795 -52.875 202.125 ;
        RECT -53.205 200.435 -52.875 200.765 ;
        RECT -53.205 199.075 -52.875 199.405 ;
        RECT -53.205 197.715 -52.875 198.045 ;
        RECT -53.205 196.355 -52.875 196.685 ;
        RECT -53.205 194.995 -52.875 195.325 ;
        RECT -53.205 193.635 -52.875 193.965 ;
        RECT -53.205 192.275 -52.875 192.605 ;
        RECT -53.205 190.915 -52.875 191.245 ;
        RECT -53.205 189.555 -52.875 189.885 ;
        RECT -53.205 188.195 -52.875 188.525 ;
        RECT -53.205 186.835 -52.875 187.165 ;
        RECT -53.205 185.475 -52.875 185.805 ;
        RECT -53.205 184.115 -52.875 184.445 ;
        RECT -53.205 182.755 -52.875 183.085 ;
        RECT -53.205 181.395 -52.875 181.725 ;
        RECT -53.205 180.035 -52.875 180.365 ;
        RECT -53.205 178.675 -52.875 179.005 ;
        RECT -53.205 177.315 -52.875 177.645 ;
        RECT -53.205 175.955 -52.875 176.285 ;
        RECT -53.205 174.595 -52.875 174.925 ;
        RECT -53.205 173.235 -52.875 173.565 ;
        RECT -53.205 171.875 -52.875 172.205 ;
        RECT -53.205 170.515 -52.875 170.845 ;
        RECT -53.205 169.155 -52.875 169.485 ;
        RECT -53.205 167.795 -52.875 168.125 ;
        RECT -53.205 166.435 -52.875 166.765 ;
        RECT -53.205 165.075 -52.875 165.405 ;
        RECT -53.205 163.715 -52.875 164.045 ;
        RECT -53.205 162.355 -52.875 162.685 ;
        RECT -53.205 160.995 -52.875 161.325 ;
        RECT -53.205 159.635 -52.875 159.965 ;
        RECT -53.205 158.275 -52.875 158.605 ;
        RECT -53.205 156.915 -52.875 157.245 ;
        RECT -53.205 155.555 -52.875 155.885 ;
        RECT -53.205 154.195 -52.875 154.525 ;
        RECT -53.205 152.835 -52.875 153.165 ;
        RECT -53.205 151.475 -52.875 151.805 ;
        RECT -53.205 150.115 -52.875 150.445 ;
        RECT -53.205 148.755 -52.875 149.085 ;
        RECT -53.205 147.395 -52.875 147.725 ;
        RECT -53.205 146.035 -52.875 146.365 ;
        RECT -53.205 144.675 -52.875 145.005 ;
        RECT -53.205 143.315 -52.875 143.645 ;
        RECT -53.205 141.955 -52.875 142.285 ;
        RECT -53.205 140.595 -52.875 140.925 ;
        RECT -53.205 139.235 -52.875 139.565 ;
        RECT -53.2 138.56 -52.88 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.205 8.675 -52.875 9.005 ;
        RECT -53.205 7.315 -52.875 7.645 ;
        RECT -53.205 5.955 -52.875 6.285 ;
        RECT -53.205 4.595 -52.875 4.925 ;
        RECT -53.205 3.235 -52.875 3.565 ;
        RECT -53.205 1.875 -52.875 2.205 ;
        RECT -53.205 0.515 -52.875 0.845 ;
        RECT -53.205 -0.845 -52.875 -0.515 ;
        RECT -53.205 -2.205 -52.875 -1.875 ;
        RECT -53.205 -3.565 -52.875 -3.235 ;
        RECT -53.205 -4.925 -52.875 -4.595 ;
        RECT -53.205 -6.285 -52.875 -5.955 ;
        RECT -53.205 -7.645 -52.875 -7.315 ;
        RECT -53.205 -9.005 -52.875 -8.675 ;
        RECT -53.205 -10.365 -52.875 -10.035 ;
        RECT -53.205 -11.725 -52.875 -11.395 ;
        RECT -53.205 -13.085 -52.875 -12.755 ;
        RECT -53.205 -14.445 -52.875 -14.115 ;
        RECT -53.205 -15.805 -52.875 -15.475 ;
        RECT -53.205 -17.165 -52.875 -16.835 ;
        RECT -53.205 -18.525 -52.875 -18.195 ;
        RECT -53.205 -19.885 -52.875 -19.555 ;
        RECT -53.205 -21.245 -52.875 -20.915 ;
        RECT -53.205 -22.605 -52.875 -22.275 ;
        RECT -53.205 -23.965 -52.875 -23.635 ;
        RECT -53.205 -25.325 -52.875 -24.995 ;
        RECT -53.205 -30.765 -52.875 -30.435 ;
        RECT -53.205 -32.125 -52.875 -31.795 ;
        RECT -53.205 -33.485 -52.875 -33.155 ;
        RECT -53.205 -34.845 -52.875 -34.515 ;
        RECT -53.205 -36.205 -52.875 -35.875 ;
        RECT -53.205 -37.565 -52.875 -37.235 ;
        RECT -53.205 -38.925 -52.875 -38.595 ;
        RECT -53.205 -40.285 -52.875 -39.955 ;
        RECT -53.205 -41.645 -52.875 -41.315 ;
        RECT -53.205 -43.005 -52.875 -42.675 ;
        RECT -53.205 -44.365 -52.875 -44.035 ;
        RECT -53.205 -45.725 -52.875 -45.395 ;
        RECT -53.205 -47.085 -52.875 -46.755 ;
        RECT -53.205 -48.445 -52.875 -48.115 ;
        RECT -53.205 -49.805 -52.875 -49.475 ;
        RECT -53.205 -51.165 -52.875 -50.835 ;
        RECT -53.205 -52.525 -52.875 -52.195 ;
        RECT -53.205 -53.885 -52.875 -53.555 ;
        RECT -53.205 -55.245 -52.875 -54.915 ;
        RECT -53.205 -56.605 -52.875 -56.275 ;
        RECT -53.205 -57.965 -52.875 -57.635 ;
        RECT -53.205 -59.325 -52.875 -58.995 ;
        RECT -53.205 -60.685 -52.875 -60.355 ;
        RECT -53.205 -62.045 -52.875 -61.715 ;
        RECT -53.205 -63.405 -52.875 -63.075 ;
        RECT -53.205 -64.765 -52.875 -64.435 ;
        RECT -53.205 -66.125 -52.875 -65.795 ;
        RECT -53.205 -68.845 -52.875 -68.515 ;
        RECT -53.205 -70.205 -52.875 -69.875 ;
        RECT -53.205 -71.565 -52.875 -71.235 ;
        RECT -53.205 -72.925 -52.875 -72.595 ;
        RECT -53.205 -74.285 -52.875 -73.955 ;
        RECT -53.205 -75.645 -52.875 -75.315 ;
        RECT -53.205 -77.005 -52.875 -76.675 ;
        RECT -53.205 -78.365 -52.875 -78.035 ;
        RECT -53.205 -79.725 -52.875 -79.395 ;
        RECT -53.205 -81.085 -52.875 -80.755 ;
        RECT -53.205 -82.445 -52.875 -82.115 ;
        RECT -53.205 -83.805 -52.875 -83.475 ;
        RECT -53.205 -85.165 -52.875 -84.835 ;
        RECT -53.205 -86.525 -52.875 -86.195 ;
        RECT -53.205 -87.885 -52.875 -87.555 ;
        RECT -53.205 -89.245 -52.875 -88.915 ;
        RECT -53.205 -90.605 -52.875 -90.275 ;
        RECT -53.205 -91.77 -52.875 -91.44 ;
        RECT -53.205 -93.325 -52.875 -92.995 ;
        RECT -53.205 -94.685 -52.875 -94.355 ;
        RECT -53.205 -96.045 -52.875 -95.715 ;
        RECT -53.205 -97.405 -52.875 -97.075 ;
        RECT -53.205 -98.765 -52.875 -98.435 ;
        RECT -53.205 -101.485 -52.875 -101.155 ;
        RECT -53.205 -102.31 -52.875 -101.98 ;
        RECT -53.205 -104.205 -52.875 -103.875 ;
        RECT -53.205 -105.565 -52.875 -105.235 ;
        RECT -53.205 -106.925 -52.875 -106.595 ;
        RECT -53.205 -109.645 -52.875 -109.315 ;
        RECT -53.205 -111.005 -52.875 -110.675 ;
        RECT -53.205 -113.725 -52.875 -113.395 ;
        RECT -53.205 -115.085 -52.875 -114.755 ;
        RECT -53.205 -116.445 -52.875 -116.115 ;
        RECT -53.205 -117.805 -52.875 -117.475 ;
        RECT -53.205 -119.165 -52.875 -118.835 ;
        RECT -53.205 -120.525 -52.875 -120.195 ;
        RECT -53.205 -123.245 -52.875 -122.915 ;
        RECT -53.205 -124.605 -52.875 -124.275 ;
        RECT -53.205 -125.965 -52.875 -125.635 ;
        RECT -53.205 -127.325 -52.875 -126.995 ;
        RECT -53.205 -128.685 -52.875 -128.355 ;
        RECT -53.205 -130.045 -52.875 -129.715 ;
        RECT -53.205 -131.405 -52.875 -131.075 ;
        RECT -53.205 -132.765 -52.875 -132.435 ;
        RECT -53.205 -134.125 -52.875 -133.795 ;
        RECT -53.205 -135.485 -52.875 -135.155 ;
        RECT -53.205 -136.845 -52.875 -136.515 ;
        RECT -53.205 -138.205 -52.875 -137.875 ;
        RECT -53.205 -139.565 -52.875 -139.235 ;
        RECT -53.205 -140.925 -52.875 -140.595 ;
        RECT -53.205 -142.285 -52.875 -141.955 ;
        RECT -53.205 -143.645 -52.875 -143.315 ;
        RECT -53.205 -145.005 -52.875 -144.675 ;
        RECT -53.205 -146.365 -52.875 -146.035 ;
        RECT -53.205 -147.725 -52.875 -147.395 ;
        RECT -53.205 -149.085 -52.875 -148.755 ;
        RECT -53.205 -150.445 -52.875 -150.115 ;
        RECT -53.205 -151.805 -52.875 -151.475 ;
        RECT -53.205 -153.165 -52.875 -152.835 ;
        RECT -53.205 -154.525 -52.875 -154.195 ;
        RECT -53.205 -155.885 -52.875 -155.555 ;
        RECT -53.205 -157.245 -52.875 -156.915 ;
        RECT -53.205 -158.605 -52.875 -158.275 ;
        RECT -53.205 -159.965 -52.875 -159.635 ;
        RECT -53.205 -161.325 -52.875 -160.995 ;
        RECT -53.205 -162.685 -52.875 -162.355 ;
        RECT -53.205 -164.045 -52.875 -163.715 ;
        RECT -53.205 -165.405 -52.875 -165.075 ;
        RECT -53.205 -166.765 -52.875 -166.435 ;
        RECT -53.205 -169.615 -52.875 -169.285 ;
        RECT -53.205 -170.845 -52.875 -170.515 ;
        RECT -53.205 -172.205 -52.875 -171.875 ;
        RECT -53.205 -174.925 -52.875 -174.595 ;
        RECT -53.205 -177.645 -52.875 -177.315 ;
        RECT -53.205 -179.005 -52.875 -178.675 ;
        RECT -53.205 -184.65 -52.875 -183.52 ;
        RECT -53.2 -184.765 -52.88 98.08 ;
        RECT -53.205 97.075 -52.875 97.405 ;
        RECT -53.205 95.715 -52.875 96.045 ;
        RECT -53.205 94.355 -52.875 94.685 ;
        RECT -53.205 92.995 -52.875 93.325 ;
        RECT -53.205 88.915 -52.875 89.245 ;
        RECT -53.205 84.835 -52.875 85.165 ;
        RECT -53.205 83.475 -52.875 83.805 ;
        RECT -53.205 82.115 -52.875 82.445 ;
        RECT -53.205 80.755 -52.875 81.085 ;
        RECT -53.205 79.395 -52.875 79.725 ;
        RECT -53.205 78.035 -52.875 78.365 ;
        RECT -53.205 76.675 -52.875 77.005 ;
        RECT -53.205 75.315 -52.875 75.645 ;
        RECT -53.205 73.955 -52.875 74.285 ;
        RECT -53.205 72.595 -52.875 72.925 ;
        RECT -53.205 71.235 -52.875 71.565 ;
        RECT -53.205 69.875 -52.875 70.205 ;
        RECT -53.205 68.515 -52.875 68.845 ;
        RECT -53.205 67.155 -52.875 67.485 ;
        RECT -53.205 65.795 -52.875 66.125 ;
        RECT -53.205 64.435 -52.875 64.765 ;
        RECT -53.205 63.075 -52.875 63.405 ;
        RECT -53.205 61.715 -52.875 62.045 ;
        RECT -53.205 60.355 -52.875 60.685 ;
        RECT -53.205 58.995 -52.875 59.325 ;
        RECT -53.205 57.635 -52.875 57.965 ;
        RECT -53.205 56.275 -52.875 56.605 ;
        RECT -53.205 54.915 -52.875 55.245 ;
        RECT -53.205 53.555 -52.875 53.885 ;
        RECT -53.205 52.195 -52.875 52.525 ;
        RECT -53.205 50.835 -52.875 51.165 ;
        RECT -53.205 49.475 -52.875 49.805 ;
        RECT -53.205 48.115 -52.875 48.445 ;
        RECT -53.205 46.755 -52.875 47.085 ;
        RECT -53.205 45.395 -52.875 45.725 ;
        RECT -53.205 44.035 -52.875 44.365 ;
        RECT -53.205 42.675 -52.875 43.005 ;
        RECT -53.205 41.315 -52.875 41.645 ;
        RECT -53.205 39.955 -52.875 40.285 ;
        RECT -53.205 38.595 -52.875 38.925 ;
        RECT -53.205 37.235 -52.875 37.565 ;
        RECT -53.205 35.875 -52.875 36.205 ;
        RECT -53.205 34.515 -52.875 34.845 ;
        RECT -53.205 33.155 -52.875 33.485 ;
        RECT -53.205 31.795 -52.875 32.125 ;
        RECT -53.205 30.435 -52.875 30.765 ;
        RECT -53.205 29.075 -52.875 29.405 ;
        RECT -53.205 27.715 -52.875 28.045 ;
        RECT -53.205 26.355 -52.875 26.685 ;
        RECT -53.205 24.995 -52.875 25.325 ;
        RECT -53.205 23.635 -52.875 23.965 ;
        RECT -53.205 22.275 -52.875 22.605 ;
        RECT -53.205 20.915 -52.875 21.245 ;
        RECT -53.205 19.555 -52.875 19.885 ;
        RECT -53.205 18.195 -52.875 18.525 ;
        RECT -53.205 16.835 -52.875 17.165 ;
        RECT -53.205 15.475 -52.875 15.805 ;
        RECT -53.205 14.115 -52.875 14.445 ;
        RECT -53.205 12.755 -52.875 13.085 ;
        RECT -53.205 11.395 -52.875 11.725 ;
        RECT -53.205 10.035 -52.875 10.365 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.085 -177.645 -63.755 -177.315 ;
        RECT -64.085 -179.005 -63.755 -178.675 ;
        RECT -64.085 -184.65 -63.755 -183.52 ;
        RECT -64.08 -184.765 -63.76 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.725 244.04 -62.395 245.17 ;
        RECT -62.725 239.875 -62.395 240.205 ;
        RECT -62.725 238.515 -62.395 238.845 ;
        RECT -62.725 237.155 -62.395 237.485 ;
        RECT -62.725 235.795 -62.395 236.125 ;
        RECT -62.725 234.435 -62.395 234.765 ;
        RECT -62.725 233.075 -62.395 233.405 ;
        RECT -62.725 231.715 -62.395 232.045 ;
        RECT -62.725 230.355 -62.395 230.685 ;
        RECT -62.725 228.995 -62.395 229.325 ;
        RECT -62.725 227.635 -62.395 227.965 ;
        RECT -62.725 226.275 -62.395 226.605 ;
        RECT -62.725 224.915 -62.395 225.245 ;
        RECT -62.725 223.555 -62.395 223.885 ;
        RECT -62.725 222.195 -62.395 222.525 ;
        RECT -62.725 220.835 -62.395 221.165 ;
        RECT -62.725 219.475 -62.395 219.805 ;
        RECT -62.725 218.115 -62.395 218.445 ;
        RECT -62.725 216.755 -62.395 217.085 ;
        RECT -62.725 215.395 -62.395 215.725 ;
        RECT -62.725 214.035 -62.395 214.365 ;
        RECT -62.725 212.675 -62.395 213.005 ;
        RECT -62.725 211.315 -62.395 211.645 ;
        RECT -62.725 209.955 -62.395 210.285 ;
        RECT -62.725 208.595 -62.395 208.925 ;
        RECT -62.725 207.235 -62.395 207.565 ;
        RECT -62.725 205.875 -62.395 206.205 ;
        RECT -62.725 204.515 -62.395 204.845 ;
        RECT -62.725 203.155 -62.395 203.485 ;
        RECT -62.725 201.795 -62.395 202.125 ;
        RECT -62.725 200.435 -62.395 200.765 ;
        RECT -62.725 199.075 -62.395 199.405 ;
        RECT -62.725 197.715 -62.395 198.045 ;
        RECT -62.725 196.355 -62.395 196.685 ;
        RECT -62.725 194.995 -62.395 195.325 ;
        RECT -62.725 193.635 -62.395 193.965 ;
        RECT -62.725 192.275 -62.395 192.605 ;
        RECT -62.725 190.915 -62.395 191.245 ;
        RECT -62.725 189.555 -62.395 189.885 ;
        RECT -62.725 188.195 -62.395 188.525 ;
        RECT -62.725 186.835 -62.395 187.165 ;
        RECT -62.725 185.475 -62.395 185.805 ;
        RECT -62.725 184.115 -62.395 184.445 ;
        RECT -62.725 182.755 -62.395 183.085 ;
        RECT -62.725 181.395 -62.395 181.725 ;
        RECT -62.725 180.035 -62.395 180.365 ;
        RECT -62.725 178.675 -62.395 179.005 ;
        RECT -62.725 177.315 -62.395 177.645 ;
        RECT -62.725 175.955 -62.395 176.285 ;
        RECT -62.725 174.595 -62.395 174.925 ;
        RECT -62.725 173.235 -62.395 173.565 ;
        RECT -62.725 171.875 -62.395 172.205 ;
        RECT -62.725 170.515 -62.395 170.845 ;
        RECT -62.725 169.155 -62.395 169.485 ;
        RECT -62.725 167.795 -62.395 168.125 ;
        RECT -62.725 166.435 -62.395 166.765 ;
        RECT -62.725 165.075 -62.395 165.405 ;
        RECT -62.725 163.715 -62.395 164.045 ;
        RECT -62.725 162.355 -62.395 162.685 ;
        RECT -62.725 160.995 -62.395 161.325 ;
        RECT -62.725 159.635 -62.395 159.965 ;
        RECT -62.725 158.275 -62.395 158.605 ;
        RECT -62.725 156.915 -62.395 157.245 ;
        RECT -62.725 155.555 -62.395 155.885 ;
        RECT -62.725 154.195 -62.395 154.525 ;
        RECT -62.725 152.835 -62.395 153.165 ;
        RECT -62.725 151.475 -62.395 151.805 ;
        RECT -62.725 150.115 -62.395 150.445 ;
        RECT -62.725 148.755 -62.395 149.085 ;
        RECT -62.725 147.395 -62.395 147.725 ;
        RECT -62.725 146.035 -62.395 146.365 ;
        RECT -62.725 144.675 -62.395 145.005 ;
        RECT -62.725 143.315 -62.395 143.645 ;
        RECT -62.725 141.955 -62.395 142.285 ;
        RECT -62.725 140.595 -62.395 140.925 ;
        RECT -62.725 139.235 -62.395 139.565 ;
        RECT -62.725 136.42 -62.395 136.75 ;
        RECT -62.725 134.245 -62.395 134.575 ;
        RECT -62.725 133.395 -62.395 133.725 ;
        RECT -62.725 131.085 -62.395 131.415 ;
        RECT -62.725 130.235 -62.395 130.565 ;
        RECT -62.725 127.925 -62.395 128.255 ;
        RECT -62.725 127.075 -62.395 127.405 ;
        RECT -62.725 124.765 -62.395 125.095 ;
        RECT -62.725 123.915 -62.395 124.245 ;
        RECT -62.725 121.605 -62.395 121.935 ;
        RECT -62.725 120.755 -62.395 121.085 ;
        RECT -62.725 118.445 -62.395 118.775 ;
        RECT -62.725 117.595 -62.395 117.925 ;
        RECT -62.725 115.285 -62.395 115.615 ;
        RECT -62.725 114.435 -62.395 114.765 ;
        RECT -62.725 112.125 -62.395 112.455 ;
        RECT -62.725 111.275 -62.395 111.605 ;
        RECT -62.725 108.965 -62.395 109.295 ;
        RECT -62.725 108.115 -62.395 108.445 ;
        RECT -62.725 105.805 -62.395 106.135 ;
        RECT -62.725 104.955 -62.395 105.285 ;
        RECT -62.725 102.645 -62.395 102.975 ;
        RECT -62.725 101.795 -62.395 102.125 ;
        RECT -62.725 99.62 -62.395 99.95 ;
        RECT -62.725 97.075 -62.395 97.405 ;
        RECT -62.725 95.715 -62.395 96.045 ;
        RECT -62.725 94.355 -62.395 94.685 ;
        RECT -62.725 92.995 -62.395 93.325 ;
        RECT -62.725 91.635 -62.395 91.965 ;
        RECT -62.725 90.275 -62.395 90.605 ;
        RECT -62.725 88.915 -62.395 89.245 ;
        RECT -62.725 87.555 -62.395 87.885 ;
        RECT -62.725 86.195 -62.395 86.525 ;
        RECT -62.725 84.835 -62.395 85.165 ;
        RECT -62.725 83.475 -62.395 83.805 ;
        RECT -62.725 82.115 -62.395 82.445 ;
        RECT -62.725 80.755 -62.395 81.085 ;
        RECT -62.725 79.395 -62.395 79.725 ;
        RECT -62.725 78.035 -62.395 78.365 ;
        RECT -62.725 76.675 -62.395 77.005 ;
        RECT -62.725 75.315 -62.395 75.645 ;
        RECT -62.725 73.955 -62.395 74.285 ;
        RECT -62.725 72.595 -62.395 72.925 ;
        RECT -62.725 71.235 -62.395 71.565 ;
        RECT -62.725 69.875 -62.395 70.205 ;
        RECT -62.725 68.515 -62.395 68.845 ;
        RECT -62.725 67.155 -62.395 67.485 ;
        RECT -62.725 65.795 -62.395 66.125 ;
        RECT -62.725 64.435 -62.395 64.765 ;
        RECT -62.725 63.075 -62.395 63.405 ;
        RECT -62.725 61.715 -62.395 62.045 ;
        RECT -62.725 60.355 -62.395 60.685 ;
        RECT -62.725 58.995 -62.395 59.325 ;
        RECT -62.725 57.635 -62.395 57.965 ;
        RECT -62.725 56.275 -62.395 56.605 ;
        RECT -62.725 54.915 -62.395 55.245 ;
        RECT -62.725 53.555 -62.395 53.885 ;
        RECT -62.725 52.195 -62.395 52.525 ;
        RECT -62.725 50.835 -62.395 51.165 ;
        RECT -62.725 49.475 -62.395 49.805 ;
        RECT -62.725 48.115 -62.395 48.445 ;
        RECT -62.725 46.755 -62.395 47.085 ;
        RECT -62.725 45.395 -62.395 45.725 ;
        RECT -62.725 44.035 -62.395 44.365 ;
        RECT -62.725 42.675 -62.395 43.005 ;
        RECT -62.725 41.315 -62.395 41.645 ;
        RECT -62.725 39.955 -62.395 40.285 ;
        RECT -62.725 38.595 -62.395 38.925 ;
        RECT -62.725 37.235 -62.395 37.565 ;
        RECT -62.725 35.875 -62.395 36.205 ;
        RECT -62.725 34.515 -62.395 34.845 ;
        RECT -62.725 33.155 -62.395 33.485 ;
        RECT -62.725 31.795 -62.395 32.125 ;
        RECT -62.725 30.435 -62.395 30.765 ;
        RECT -62.725 29.075 -62.395 29.405 ;
        RECT -62.725 27.715 -62.395 28.045 ;
        RECT -62.725 26.355 -62.395 26.685 ;
        RECT -62.725 24.995 -62.395 25.325 ;
        RECT -62.725 23.635 -62.395 23.965 ;
        RECT -62.725 22.275 -62.395 22.605 ;
        RECT -62.725 20.915 -62.395 21.245 ;
        RECT -62.725 19.555 -62.395 19.885 ;
        RECT -62.725 18.195 -62.395 18.525 ;
        RECT -62.725 16.835 -62.395 17.165 ;
        RECT -62.725 15.475 -62.395 15.805 ;
        RECT -62.725 14.115 -62.395 14.445 ;
        RECT -62.725 12.755 -62.395 13.085 ;
        RECT -62.725 11.395 -62.395 11.725 ;
        RECT -62.725 10.035 -62.395 10.365 ;
        RECT -62.725 8.675 -62.395 9.005 ;
        RECT -62.725 7.315 -62.395 7.645 ;
        RECT -62.725 5.955 -62.395 6.285 ;
        RECT -62.725 4.595 -62.395 4.925 ;
        RECT -62.725 3.235 -62.395 3.565 ;
        RECT -62.725 1.875 -62.395 2.205 ;
        RECT -62.725 0.515 -62.395 0.845 ;
        RECT -62.725 -0.845 -62.395 -0.515 ;
        RECT -62.725 -2.205 -62.395 -1.875 ;
        RECT -62.725 -3.565 -62.395 -3.235 ;
        RECT -62.725 -4.925 -62.395 -4.595 ;
        RECT -62.725 -6.285 -62.395 -5.955 ;
        RECT -62.725 -7.645 -62.395 -7.315 ;
        RECT -62.725 -9.005 -62.395 -8.675 ;
        RECT -62.725 -10.365 -62.395 -10.035 ;
        RECT -62.725 -11.725 -62.395 -11.395 ;
        RECT -62.725 -13.085 -62.395 -12.755 ;
        RECT -62.725 -14.445 -62.395 -14.115 ;
        RECT -62.725 -15.805 -62.395 -15.475 ;
        RECT -62.725 -17.165 -62.395 -16.835 ;
        RECT -62.725 -18.525 -62.395 -18.195 ;
        RECT -62.725 -19.885 -62.395 -19.555 ;
        RECT -62.725 -21.245 -62.395 -20.915 ;
        RECT -62.725 -22.605 -62.395 -22.275 ;
        RECT -62.725 -23.965 -62.395 -23.635 ;
        RECT -62.725 -25.325 -62.395 -24.995 ;
        RECT -62.725 -29.405 -62.395 -29.075 ;
        RECT -62.725 -30.765 -62.395 -30.435 ;
        RECT -62.725 -32.125 -62.395 -31.795 ;
        RECT -62.725 -33.485 -62.395 -33.155 ;
        RECT -62.725 -34.845 -62.395 -34.515 ;
        RECT -62.725 -36.205 -62.395 -35.875 ;
        RECT -62.725 -37.565 -62.395 -37.235 ;
        RECT -62.725 -38.925 -62.395 -38.595 ;
        RECT -62.725 -40.285 -62.395 -39.955 ;
        RECT -62.725 -41.645 -62.395 -41.315 ;
        RECT -62.725 -43.005 -62.395 -42.675 ;
        RECT -62.725 -44.365 -62.395 -44.035 ;
        RECT -62.725 -45.725 -62.395 -45.395 ;
        RECT -62.725 -47.085 -62.395 -46.755 ;
        RECT -62.725 -48.445 -62.395 -48.115 ;
        RECT -62.725 -49.805 -62.395 -49.475 ;
        RECT -62.725 -51.165 -62.395 -50.835 ;
        RECT -62.725 -52.525 -62.395 -52.195 ;
        RECT -62.725 -53.885 -62.395 -53.555 ;
        RECT -62.725 -55.245 -62.395 -54.915 ;
        RECT -62.725 -56.605 -62.395 -56.275 ;
        RECT -62.725 -57.965 -62.395 -57.635 ;
        RECT -62.725 -59.325 -62.395 -58.995 ;
        RECT -62.725 -60.685 -62.395 -60.355 ;
        RECT -62.725 -62.045 -62.395 -61.715 ;
        RECT -62.725 -63.405 -62.395 -63.075 ;
        RECT -62.725 -64.765 -62.395 -64.435 ;
        RECT -62.725 -66.125 -62.395 -65.795 ;
        RECT -62.725 -67.485 -62.395 -67.155 ;
        RECT -62.725 -68.845 -62.395 -68.515 ;
        RECT -62.725 -70.205 -62.395 -69.875 ;
        RECT -62.725 -71.565 -62.395 -71.235 ;
        RECT -62.725 -72.925 -62.395 -72.595 ;
        RECT -62.725 -74.285 -62.395 -73.955 ;
        RECT -62.725 -75.645 -62.395 -75.315 ;
        RECT -62.725 -77.005 -62.395 -76.675 ;
        RECT -62.725 -78.365 -62.395 -78.035 ;
        RECT -62.725 -79.725 -62.395 -79.395 ;
        RECT -62.725 -81.085 -62.395 -80.755 ;
        RECT -62.725 -82.445 -62.395 -82.115 ;
        RECT -62.725 -83.805 -62.395 -83.475 ;
        RECT -62.725 -85.165 -62.395 -84.835 ;
        RECT -62.725 -86.525 -62.395 -86.195 ;
        RECT -62.725 -87.885 -62.395 -87.555 ;
        RECT -62.725 -89.245 -62.395 -88.915 ;
        RECT -62.725 -90.605 -62.395 -90.275 ;
        RECT -62.725 -91.77 -62.395 -91.44 ;
        RECT -62.725 -93.325 -62.395 -92.995 ;
        RECT -62.725 -94.685 -62.395 -94.355 ;
        RECT -62.725 -96.045 -62.395 -95.715 ;
        RECT -62.725 -97.405 -62.395 -97.075 ;
        RECT -62.725 -98.765 -62.395 -98.435 ;
        RECT -62.725 -101.485 -62.395 -101.155 ;
        RECT -62.725 -102.31 -62.395 -101.98 ;
        RECT -62.725 -104.205 -62.395 -103.875 ;
        RECT -62.725 -105.565 -62.395 -105.235 ;
        RECT -62.725 -106.925 -62.395 -106.595 ;
        RECT -62.725 -109.645 -62.395 -109.315 ;
        RECT -62.725 -111.005 -62.395 -110.675 ;
        RECT -62.72 -113.04 -62.4 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.725 -177.645 -62.395 -177.315 ;
        RECT -62.725 -179.005 -62.395 -178.675 ;
        RECT -62.725 -184.65 -62.395 -183.52 ;
        RECT -62.72 -184.765 -62.4 -175.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -61.365 244.04 -61.035 245.17 ;
        RECT -61.365 239.875 -61.035 240.205 ;
        RECT -61.365 238.515 -61.035 238.845 ;
        RECT -61.365 237.155 -61.035 237.485 ;
        RECT -61.365 235.795 -61.035 236.125 ;
        RECT -61.365 234.435 -61.035 234.765 ;
        RECT -61.365 233.075 -61.035 233.405 ;
        RECT -61.365 231.715 -61.035 232.045 ;
        RECT -61.365 230.355 -61.035 230.685 ;
        RECT -61.365 228.995 -61.035 229.325 ;
        RECT -61.365 227.635 -61.035 227.965 ;
        RECT -61.365 226.275 -61.035 226.605 ;
        RECT -61.365 224.915 -61.035 225.245 ;
        RECT -61.365 223.555 -61.035 223.885 ;
        RECT -61.365 222.195 -61.035 222.525 ;
        RECT -61.365 220.835 -61.035 221.165 ;
        RECT -61.365 219.475 -61.035 219.805 ;
        RECT -61.365 218.115 -61.035 218.445 ;
        RECT -61.365 216.755 -61.035 217.085 ;
        RECT -61.365 215.395 -61.035 215.725 ;
        RECT -61.365 214.035 -61.035 214.365 ;
        RECT -61.365 212.675 -61.035 213.005 ;
        RECT -61.365 211.315 -61.035 211.645 ;
        RECT -61.365 209.955 -61.035 210.285 ;
        RECT -61.365 208.595 -61.035 208.925 ;
        RECT -61.365 207.235 -61.035 207.565 ;
        RECT -61.365 205.875 -61.035 206.205 ;
        RECT -61.365 204.515 -61.035 204.845 ;
        RECT -61.365 203.155 -61.035 203.485 ;
        RECT -61.365 201.795 -61.035 202.125 ;
        RECT -61.365 200.435 -61.035 200.765 ;
        RECT -61.365 199.075 -61.035 199.405 ;
        RECT -61.365 197.715 -61.035 198.045 ;
        RECT -61.365 196.355 -61.035 196.685 ;
        RECT -61.365 194.995 -61.035 195.325 ;
        RECT -61.365 193.635 -61.035 193.965 ;
        RECT -61.365 192.275 -61.035 192.605 ;
        RECT -61.365 190.915 -61.035 191.245 ;
        RECT -61.365 189.555 -61.035 189.885 ;
        RECT -61.365 188.195 -61.035 188.525 ;
        RECT -61.365 186.835 -61.035 187.165 ;
        RECT -61.365 185.475 -61.035 185.805 ;
        RECT -61.365 184.115 -61.035 184.445 ;
        RECT -61.365 182.755 -61.035 183.085 ;
        RECT -61.365 181.395 -61.035 181.725 ;
        RECT -61.365 180.035 -61.035 180.365 ;
        RECT -61.365 178.675 -61.035 179.005 ;
        RECT -61.365 177.315 -61.035 177.645 ;
        RECT -61.365 175.955 -61.035 176.285 ;
        RECT -61.365 174.595 -61.035 174.925 ;
        RECT -61.365 173.235 -61.035 173.565 ;
        RECT -61.365 171.875 -61.035 172.205 ;
        RECT -61.365 170.515 -61.035 170.845 ;
        RECT -61.365 169.155 -61.035 169.485 ;
        RECT -61.365 167.795 -61.035 168.125 ;
        RECT -61.365 166.435 -61.035 166.765 ;
        RECT -61.365 165.075 -61.035 165.405 ;
        RECT -61.365 163.715 -61.035 164.045 ;
        RECT -61.365 162.355 -61.035 162.685 ;
        RECT -61.365 160.995 -61.035 161.325 ;
        RECT -61.365 159.635 -61.035 159.965 ;
        RECT -61.365 158.275 -61.035 158.605 ;
        RECT -61.365 156.915 -61.035 157.245 ;
        RECT -61.365 155.555 -61.035 155.885 ;
        RECT -61.365 154.195 -61.035 154.525 ;
        RECT -61.365 152.835 -61.035 153.165 ;
        RECT -61.365 151.475 -61.035 151.805 ;
        RECT -61.365 150.115 -61.035 150.445 ;
        RECT -61.365 148.755 -61.035 149.085 ;
        RECT -61.365 147.395 -61.035 147.725 ;
        RECT -61.365 146.035 -61.035 146.365 ;
        RECT -61.365 144.675 -61.035 145.005 ;
        RECT -61.365 143.315 -61.035 143.645 ;
        RECT -61.365 141.955 -61.035 142.285 ;
        RECT -61.365 140.595 -61.035 140.925 ;
        RECT -61.365 139.235 -61.035 139.565 ;
        RECT -61.365 136.42 -61.035 136.75 ;
        RECT -61.365 134.245 -61.035 134.575 ;
        RECT -61.365 133.395 -61.035 133.725 ;
        RECT -61.365 131.085 -61.035 131.415 ;
        RECT -61.365 130.235 -61.035 130.565 ;
        RECT -61.365 127.925 -61.035 128.255 ;
        RECT -61.365 127.075 -61.035 127.405 ;
        RECT -61.365 124.765 -61.035 125.095 ;
        RECT -61.365 123.915 -61.035 124.245 ;
        RECT -61.365 121.605 -61.035 121.935 ;
        RECT -61.365 120.755 -61.035 121.085 ;
        RECT -61.365 118.445 -61.035 118.775 ;
        RECT -61.365 117.595 -61.035 117.925 ;
        RECT -61.365 115.285 -61.035 115.615 ;
        RECT -61.365 114.435 -61.035 114.765 ;
        RECT -61.365 112.125 -61.035 112.455 ;
        RECT -61.365 111.275 -61.035 111.605 ;
        RECT -61.365 108.965 -61.035 109.295 ;
        RECT -61.365 108.115 -61.035 108.445 ;
        RECT -61.365 105.805 -61.035 106.135 ;
        RECT -61.365 104.955 -61.035 105.285 ;
        RECT -61.365 102.645 -61.035 102.975 ;
        RECT -61.365 101.795 -61.035 102.125 ;
        RECT -61.365 99.62 -61.035 99.95 ;
        RECT -61.365 97.075 -61.035 97.405 ;
        RECT -61.365 95.715 -61.035 96.045 ;
        RECT -61.365 94.355 -61.035 94.685 ;
        RECT -61.365 92.995 -61.035 93.325 ;
        RECT -61.365 91.635 -61.035 91.965 ;
        RECT -61.365 90.275 -61.035 90.605 ;
        RECT -61.365 88.915 -61.035 89.245 ;
        RECT -61.365 87.555 -61.035 87.885 ;
        RECT -61.365 86.195 -61.035 86.525 ;
        RECT -61.365 84.835 -61.035 85.165 ;
        RECT -61.365 83.475 -61.035 83.805 ;
        RECT -61.365 82.115 -61.035 82.445 ;
        RECT -61.365 80.755 -61.035 81.085 ;
        RECT -61.365 79.395 -61.035 79.725 ;
        RECT -61.365 78.035 -61.035 78.365 ;
        RECT -61.365 76.675 -61.035 77.005 ;
        RECT -61.365 75.315 -61.035 75.645 ;
        RECT -61.365 73.955 -61.035 74.285 ;
        RECT -61.365 72.595 -61.035 72.925 ;
        RECT -61.365 71.235 -61.035 71.565 ;
        RECT -61.365 69.875 -61.035 70.205 ;
        RECT -61.365 68.515 -61.035 68.845 ;
        RECT -61.365 67.155 -61.035 67.485 ;
        RECT -61.365 65.795 -61.035 66.125 ;
        RECT -61.365 64.435 -61.035 64.765 ;
        RECT -61.365 63.075 -61.035 63.405 ;
        RECT -61.365 61.715 -61.035 62.045 ;
        RECT -61.365 60.355 -61.035 60.685 ;
        RECT -61.365 58.995 -61.035 59.325 ;
        RECT -61.365 57.635 -61.035 57.965 ;
        RECT -61.365 56.275 -61.035 56.605 ;
        RECT -61.365 54.915 -61.035 55.245 ;
        RECT -61.365 53.555 -61.035 53.885 ;
        RECT -61.365 52.195 -61.035 52.525 ;
        RECT -61.365 50.835 -61.035 51.165 ;
        RECT -61.365 49.475 -61.035 49.805 ;
        RECT -61.365 48.115 -61.035 48.445 ;
        RECT -61.365 46.755 -61.035 47.085 ;
        RECT -61.365 45.395 -61.035 45.725 ;
        RECT -61.365 44.035 -61.035 44.365 ;
        RECT -61.365 42.675 -61.035 43.005 ;
        RECT -61.365 41.315 -61.035 41.645 ;
        RECT -61.365 39.955 -61.035 40.285 ;
        RECT -61.365 38.595 -61.035 38.925 ;
        RECT -61.365 37.235 -61.035 37.565 ;
        RECT -61.365 35.875 -61.035 36.205 ;
        RECT -61.365 34.515 -61.035 34.845 ;
        RECT -61.365 33.155 -61.035 33.485 ;
        RECT -61.365 31.795 -61.035 32.125 ;
        RECT -61.365 30.435 -61.035 30.765 ;
        RECT -61.365 29.075 -61.035 29.405 ;
        RECT -61.365 27.715 -61.035 28.045 ;
        RECT -61.365 26.355 -61.035 26.685 ;
        RECT -61.365 24.995 -61.035 25.325 ;
        RECT -61.365 23.635 -61.035 23.965 ;
        RECT -61.365 22.275 -61.035 22.605 ;
        RECT -61.365 20.915 -61.035 21.245 ;
        RECT -61.365 19.555 -61.035 19.885 ;
        RECT -61.365 18.195 -61.035 18.525 ;
        RECT -61.365 16.835 -61.035 17.165 ;
        RECT -61.365 15.475 -61.035 15.805 ;
        RECT -61.365 14.115 -61.035 14.445 ;
        RECT -61.365 12.755 -61.035 13.085 ;
        RECT -61.365 11.395 -61.035 11.725 ;
        RECT -61.365 10.035 -61.035 10.365 ;
        RECT -61.365 8.675 -61.035 9.005 ;
        RECT -61.365 7.315 -61.035 7.645 ;
        RECT -61.365 5.955 -61.035 6.285 ;
        RECT -61.365 4.595 -61.035 4.925 ;
        RECT -61.365 3.235 -61.035 3.565 ;
        RECT -61.365 1.875 -61.035 2.205 ;
        RECT -61.365 0.515 -61.035 0.845 ;
        RECT -61.365 -0.845 -61.035 -0.515 ;
        RECT -61.365 -2.205 -61.035 -1.875 ;
        RECT -61.365 -3.565 -61.035 -3.235 ;
        RECT -61.365 -4.925 -61.035 -4.595 ;
        RECT -61.365 -6.285 -61.035 -5.955 ;
        RECT -61.365 -7.645 -61.035 -7.315 ;
        RECT -61.365 -9.005 -61.035 -8.675 ;
        RECT -61.365 -10.365 -61.035 -10.035 ;
        RECT -61.365 -11.725 -61.035 -11.395 ;
        RECT -61.365 -13.085 -61.035 -12.755 ;
        RECT -61.365 -14.445 -61.035 -14.115 ;
        RECT -61.365 -15.805 -61.035 -15.475 ;
        RECT -61.365 -17.165 -61.035 -16.835 ;
        RECT -61.365 -18.525 -61.035 -18.195 ;
        RECT -61.365 -19.885 -61.035 -19.555 ;
        RECT -61.365 -21.245 -61.035 -20.915 ;
        RECT -61.365 -22.605 -61.035 -22.275 ;
        RECT -61.365 -23.965 -61.035 -23.635 ;
        RECT -61.365 -25.325 -61.035 -24.995 ;
        RECT -61.365 -29.405 -61.035 -29.075 ;
        RECT -61.365 -30.765 -61.035 -30.435 ;
        RECT -61.365 -32.125 -61.035 -31.795 ;
        RECT -61.365 -33.485 -61.035 -33.155 ;
        RECT -61.365 -34.845 -61.035 -34.515 ;
        RECT -61.365 -36.205 -61.035 -35.875 ;
        RECT -61.365 -37.565 -61.035 -37.235 ;
        RECT -61.365 -38.925 -61.035 -38.595 ;
        RECT -61.365 -40.285 -61.035 -39.955 ;
        RECT -61.365 -41.645 -61.035 -41.315 ;
        RECT -61.365 -43.005 -61.035 -42.675 ;
        RECT -61.365 -44.365 -61.035 -44.035 ;
        RECT -61.365 -45.725 -61.035 -45.395 ;
        RECT -61.365 -47.085 -61.035 -46.755 ;
        RECT -61.365 -48.445 -61.035 -48.115 ;
        RECT -61.365 -49.805 -61.035 -49.475 ;
        RECT -61.365 -51.165 -61.035 -50.835 ;
        RECT -61.365 -52.525 -61.035 -52.195 ;
        RECT -61.365 -53.885 -61.035 -53.555 ;
        RECT -61.365 -55.245 -61.035 -54.915 ;
        RECT -61.365 -56.605 -61.035 -56.275 ;
        RECT -61.365 -57.965 -61.035 -57.635 ;
        RECT -61.365 -59.325 -61.035 -58.995 ;
        RECT -61.365 -60.685 -61.035 -60.355 ;
        RECT -61.365 -62.045 -61.035 -61.715 ;
        RECT -61.365 -63.405 -61.035 -63.075 ;
        RECT -61.365 -64.765 -61.035 -64.435 ;
        RECT -61.365 -66.125 -61.035 -65.795 ;
        RECT -61.365 -67.485 -61.035 -67.155 ;
        RECT -61.365 -68.845 -61.035 -68.515 ;
        RECT -61.365 -70.205 -61.035 -69.875 ;
        RECT -61.365 -71.565 -61.035 -71.235 ;
        RECT -61.365 -72.925 -61.035 -72.595 ;
        RECT -61.365 -74.285 -61.035 -73.955 ;
        RECT -61.365 -75.645 -61.035 -75.315 ;
        RECT -61.365 -77.005 -61.035 -76.675 ;
        RECT -61.365 -78.365 -61.035 -78.035 ;
        RECT -61.365 -79.725 -61.035 -79.395 ;
        RECT -61.365 -81.085 -61.035 -80.755 ;
        RECT -61.365 -82.445 -61.035 -82.115 ;
        RECT -61.365 -83.805 -61.035 -83.475 ;
        RECT -61.365 -85.165 -61.035 -84.835 ;
        RECT -61.365 -86.525 -61.035 -86.195 ;
        RECT -61.365 -87.885 -61.035 -87.555 ;
        RECT -61.365 -89.245 -61.035 -88.915 ;
        RECT -61.365 -90.605 -61.035 -90.275 ;
        RECT -61.365 -91.77 -61.035 -91.44 ;
        RECT -61.365 -93.325 -61.035 -92.995 ;
        RECT -61.365 -94.685 -61.035 -94.355 ;
        RECT -61.365 -96.045 -61.035 -95.715 ;
        RECT -61.365 -97.405 -61.035 -97.075 ;
        RECT -61.365 -98.765 -61.035 -98.435 ;
        RECT -61.365 -101.485 -61.035 -101.155 ;
        RECT -61.365 -102.31 -61.035 -101.98 ;
        RECT -61.365 -104.205 -61.035 -103.875 ;
        RECT -61.365 -105.565 -61.035 -105.235 ;
        RECT -61.365 -106.925 -61.035 -106.595 ;
        RECT -61.365 -109.645 -61.035 -109.315 ;
        RECT -61.365 -111.005 -61.035 -110.675 ;
        RECT -61.365 -113.725 -61.035 -113.395 ;
        RECT -61.365 -115.085 -61.035 -114.755 ;
        RECT -61.365 -116.445 -61.035 -116.115 ;
        RECT -61.365 -117.805 -61.035 -117.475 ;
        RECT -61.365 -119.165 -61.035 -118.835 ;
        RECT -61.365 -120.525 -61.035 -120.195 ;
        RECT -61.365 -123.245 -61.035 -122.915 ;
        RECT -61.365 -124.605 -61.035 -124.275 ;
        RECT -61.365 -125.965 -61.035 -125.635 ;
        RECT -61.365 -127.325 -61.035 -126.995 ;
        RECT -61.365 -128.685 -61.035 -128.355 ;
        RECT -61.365 -130.045 -61.035 -129.715 ;
        RECT -61.365 -131.405 -61.035 -131.075 ;
        RECT -61.365 -132.765 -61.035 -132.435 ;
        RECT -61.365 -134.125 -61.035 -133.795 ;
        RECT -61.365 -135.485 -61.035 -135.155 ;
        RECT -61.365 -136.845 -61.035 -136.515 ;
        RECT -61.365 -138.205 -61.035 -137.875 ;
        RECT -61.365 -139.565 -61.035 -139.235 ;
        RECT -61.365 -140.925 -61.035 -140.595 ;
        RECT -61.365 -142.285 -61.035 -141.955 ;
        RECT -61.365 -143.645 -61.035 -143.315 ;
        RECT -61.365 -145.005 -61.035 -144.675 ;
        RECT -61.365 -146.365 -61.035 -146.035 ;
        RECT -61.365 -147.725 -61.035 -147.395 ;
        RECT -61.365 -149.085 -61.035 -148.755 ;
        RECT -61.365 -150.445 -61.035 -150.115 ;
        RECT -61.365 -151.805 -61.035 -151.475 ;
        RECT -61.365 -153.165 -61.035 -152.835 ;
        RECT -61.365 -154.525 -61.035 -154.195 ;
        RECT -61.365 -155.885 -61.035 -155.555 ;
        RECT -61.365 -157.245 -61.035 -156.915 ;
        RECT -61.365 -158.605 -61.035 -158.275 ;
        RECT -61.365 -159.965 -61.035 -159.635 ;
        RECT -61.365 -161.325 -61.035 -160.995 ;
        RECT -61.365 -162.685 -61.035 -162.355 ;
        RECT -61.365 -164.045 -61.035 -163.715 ;
        RECT -61.365 -165.405 -61.035 -165.075 ;
        RECT -61.365 -166.765 -61.035 -166.435 ;
        RECT -61.365 -169.615 -61.035 -169.285 ;
        RECT -61.365 -170.845 -61.035 -170.515 ;
        RECT -61.365 -172.205 -61.035 -171.875 ;
        RECT -61.365 -173.565 -61.035 -173.235 ;
        RECT -61.365 -174.925 -61.035 -174.595 ;
        RECT -61.365 -177.645 -61.035 -177.315 ;
        RECT -61.365 -179.005 -61.035 -178.675 ;
        RECT -61.365 -184.65 -61.035 -183.52 ;
        RECT -61.36 -184.765 -61.04 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.005 244.04 -59.675 245.17 ;
        RECT -60.005 239.875 -59.675 240.205 ;
        RECT -60.005 238.515 -59.675 238.845 ;
        RECT -60.005 237.155 -59.675 237.485 ;
        RECT -60.005 235.795 -59.675 236.125 ;
        RECT -60.005 234.435 -59.675 234.765 ;
        RECT -60.005 233.075 -59.675 233.405 ;
        RECT -60.005 231.715 -59.675 232.045 ;
        RECT -60.005 230.355 -59.675 230.685 ;
        RECT -60.005 228.995 -59.675 229.325 ;
        RECT -60.005 227.635 -59.675 227.965 ;
        RECT -60.005 226.275 -59.675 226.605 ;
        RECT -60.005 224.915 -59.675 225.245 ;
        RECT -60.005 223.555 -59.675 223.885 ;
        RECT -60.005 222.195 -59.675 222.525 ;
        RECT -60.005 220.835 -59.675 221.165 ;
        RECT -60.005 219.475 -59.675 219.805 ;
        RECT -60.005 218.115 -59.675 218.445 ;
        RECT -60.005 216.755 -59.675 217.085 ;
        RECT -60.005 215.395 -59.675 215.725 ;
        RECT -60.005 214.035 -59.675 214.365 ;
        RECT -60.005 212.675 -59.675 213.005 ;
        RECT -60.005 211.315 -59.675 211.645 ;
        RECT -60.005 209.955 -59.675 210.285 ;
        RECT -60.005 208.595 -59.675 208.925 ;
        RECT -60.005 207.235 -59.675 207.565 ;
        RECT -60.005 205.875 -59.675 206.205 ;
        RECT -60.005 204.515 -59.675 204.845 ;
        RECT -60.005 203.155 -59.675 203.485 ;
        RECT -60.005 201.795 -59.675 202.125 ;
        RECT -60.005 200.435 -59.675 200.765 ;
        RECT -60.005 199.075 -59.675 199.405 ;
        RECT -60.005 197.715 -59.675 198.045 ;
        RECT -60.005 196.355 -59.675 196.685 ;
        RECT -60.005 194.995 -59.675 195.325 ;
        RECT -60.005 193.635 -59.675 193.965 ;
        RECT -60.005 192.275 -59.675 192.605 ;
        RECT -60.005 190.915 -59.675 191.245 ;
        RECT -60.005 189.555 -59.675 189.885 ;
        RECT -60.005 188.195 -59.675 188.525 ;
        RECT -60.005 186.835 -59.675 187.165 ;
        RECT -60.005 185.475 -59.675 185.805 ;
        RECT -60.005 184.115 -59.675 184.445 ;
        RECT -60.005 182.755 -59.675 183.085 ;
        RECT -60.005 181.395 -59.675 181.725 ;
        RECT -60.005 180.035 -59.675 180.365 ;
        RECT -60.005 178.675 -59.675 179.005 ;
        RECT -60.005 177.315 -59.675 177.645 ;
        RECT -60.005 175.955 -59.675 176.285 ;
        RECT -60.005 174.595 -59.675 174.925 ;
        RECT -60.005 173.235 -59.675 173.565 ;
        RECT -60.005 171.875 -59.675 172.205 ;
        RECT -60.005 170.515 -59.675 170.845 ;
        RECT -60.005 169.155 -59.675 169.485 ;
        RECT -60.005 167.795 -59.675 168.125 ;
        RECT -60.005 166.435 -59.675 166.765 ;
        RECT -60.005 165.075 -59.675 165.405 ;
        RECT -60.005 163.715 -59.675 164.045 ;
        RECT -60.005 162.355 -59.675 162.685 ;
        RECT -60.005 160.995 -59.675 161.325 ;
        RECT -60.005 159.635 -59.675 159.965 ;
        RECT -60.005 158.275 -59.675 158.605 ;
        RECT -60.005 156.915 -59.675 157.245 ;
        RECT -60.005 155.555 -59.675 155.885 ;
        RECT -60.005 154.195 -59.675 154.525 ;
        RECT -60.005 152.835 -59.675 153.165 ;
        RECT -60.005 151.475 -59.675 151.805 ;
        RECT -60.005 150.115 -59.675 150.445 ;
        RECT -60.005 148.755 -59.675 149.085 ;
        RECT -60.005 147.395 -59.675 147.725 ;
        RECT -60.005 146.035 -59.675 146.365 ;
        RECT -60.005 144.675 -59.675 145.005 ;
        RECT -60.005 143.315 -59.675 143.645 ;
        RECT -60.005 141.955 -59.675 142.285 ;
        RECT -60.005 140.595 -59.675 140.925 ;
        RECT -60.005 139.235 -59.675 139.565 ;
        RECT -60.005 136.42 -59.675 136.75 ;
        RECT -60.005 134.245 -59.675 134.575 ;
        RECT -60.005 133.395 -59.675 133.725 ;
        RECT -60.005 131.085 -59.675 131.415 ;
        RECT -60.005 130.235 -59.675 130.565 ;
        RECT -60.005 127.925 -59.675 128.255 ;
        RECT -60.005 127.075 -59.675 127.405 ;
        RECT -60.005 124.765 -59.675 125.095 ;
        RECT -60.005 123.915 -59.675 124.245 ;
        RECT -60.005 121.605 -59.675 121.935 ;
        RECT -60.005 120.755 -59.675 121.085 ;
        RECT -60.005 118.445 -59.675 118.775 ;
        RECT -60.005 117.595 -59.675 117.925 ;
        RECT -60.005 115.285 -59.675 115.615 ;
        RECT -60.005 114.435 -59.675 114.765 ;
        RECT -60.005 112.125 -59.675 112.455 ;
        RECT -60.005 111.275 -59.675 111.605 ;
        RECT -60.005 108.965 -59.675 109.295 ;
        RECT -60.005 108.115 -59.675 108.445 ;
        RECT -60.005 105.805 -59.675 106.135 ;
        RECT -60.005 104.955 -59.675 105.285 ;
        RECT -60.005 102.645 -59.675 102.975 ;
        RECT -60.005 101.795 -59.675 102.125 ;
        RECT -60.005 99.62 -59.675 99.95 ;
        RECT -60.005 97.075 -59.675 97.405 ;
        RECT -60.005 95.715 -59.675 96.045 ;
        RECT -60.005 94.355 -59.675 94.685 ;
        RECT -60.005 92.995 -59.675 93.325 ;
        RECT -60.005 91.635 -59.675 91.965 ;
        RECT -60.005 90.275 -59.675 90.605 ;
        RECT -60.005 88.915 -59.675 89.245 ;
        RECT -60 86.88 -59.68 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.005 -123.245 -59.675 -122.915 ;
        RECT -60.005 -124.605 -59.675 -124.275 ;
        RECT -60.005 -125.965 -59.675 -125.635 ;
        RECT -60.005 -127.325 -59.675 -126.995 ;
        RECT -60.005 -128.685 -59.675 -128.355 ;
        RECT -60.005 -130.045 -59.675 -129.715 ;
        RECT -60.005 -131.405 -59.675 -131.075 ;
        RECT -60.005 -132.765 -59.675 -132.435 ;
        RECT -60.005 -134.125 -59.675 -133.795 ;
        RECT -60.005 -135.485 -59.675 -135.155 ;
        RECT -60.005 -136.845 -59.675 -136.515 ;
        RECT -60.005 -138.205 -59.675 -137.875 ;
        RECT -60.005 -139.565 -59.675 -139.235 ;
        RECT -60.005 -140.925 -59.675 -140.595 ;
        RECT -60.005 -142.285 -59.675 -141.955 ;
        RECT -60.005 -143.645 -59.675 -143.315 ;
        RECT -60.005 -145.005 -59.675 -144.675 ;
        RECT -60.005 -146.365 -59.675 -146.035 ;
        RECT -60.005 -147.725 -59.675 -147.395 ;
        RECT -60.005 -149.085 -59.675 -148.755 ;
        RECT -60.005 -150.445 -59.675 -150.115 ;
        RECT -60.005 -151.805 -59.675 -151.475 ;
        RECT -60.005 -153.165 -59.675 -152.835 ;
        RECT -60.005 -154.525 -59.675 -154.195 ;
        RECT -60.005 -155.885 -59.675 -155.555 ;
        RECT -60.005 -157.245 -59.675 -156.915 ;
        RECT -60.005 -158.605 -59.675 -158.275 ;
        RECT -60.005 -159.965 -59.675 -159.635 ;
        RECT -60.005 -161.325 -59.675 -160.995 ;
        RECT -60.005 -162.685 -59.675 -162.355 ;
        RECT -60.005 -164.045 -59.675 -163.715 ;
        RECT -60.005 -165.405 -59.675 -165.075 ;
        RECT -60.005 -166.765 -59.675 -166.435 ;
        RECT -60.005 -170.845 -59.675 -170.515 ;
        RECT -60.005 -172.205 -59.675 -171.875 ;
        RECT -60.005 -177.645 -59.675 -177.315 ;
        RECT -60.005 -179.005 -59.675 -178.675 ;
        RECT -60.005 -184.65 -59.675 -183.52 ;
        RECT -60 -184.765 -59.68 -122.915 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.645 244.04 -58.315 245.17 ;
        RECT -58.645 239.875 -58.315 240.205 ;
        RECT -58.645 238.515 -58.315 238.845 ;
        RECT -58.645 237.155 -58.315 237.485 ;
        RECT -58.645 235.795 -58.315 236.125 ;
        RECT -58.645 234.435 -58.315 234.765 ;
        RECT -58.645 233.075 -58.315 233.405 ;
        RECT -58.645 231.715 -58.315 232.045 ;
        RECT -58.645 230.355 -58.315 230.685 ;
        RECT -58.645 228.995 -58.315 229.325 ;
        RECT -58.645 227.635 -58.315 227.965 ;
        RECT -58.645 226.275 -58.315 226.605 ;
        RECT -58.645 224.915 -58.315 225.245 ;
        RECT -58.645 223.555 -58.315 223.885 ;
        RECT -58.645 222.195 -58.315 222.525 ;
        RECT -58.645 220.835 -58.315 221.165 ;
        RECT -58.645 219.475 -58.315 219.805 ;
        RECT -58.645 218.115 -58.315 218.445 ;
        RECT -58.645 216.755 -58.315 217.085 ;
        RECT -58.645 215.395 -58.315 215.725 ;
        RECT -58.645 214.035 -58.315 214.365 ;
        RECT -58.645 212.675 -58.315 213.005 ;
        RECT -58.645 211.315 -58.315 211.645 ;
        RECT -58.645 209.955 -58.315 210.285 ;
        RECT -58.645 208.595 -58.315 208.925 ;
        RECT -58.645 207.235 -58.315 207.565 ;
        RECT -58.645 205.875 -58.315 206.205 ;
        RECT -58.645 204.515 -58.315 204.845 ;
        RECT -58.645 203.155 -58.315 203.485 ;
        RECT -58.645 201.795 -58.315 202.125 ;
        RECT -58.645 200.435 -58.315 200.765 ;
        RECT -58.645 199.075 -58.315 199.405 ;
        RECT -58.645 197.715 -58.315 198.045 ;
        RECT -58.645 196.355 -58.315 196.685 ;
        RECT -58.645 194.995 -58.315 195.325 ;
        RECT -58.645 193.635 -58.315 193.965 ;
        RECT -58.645 192.275 -58.315 192.605 ;
        RECT -58.645 190.915 -58.315 191.245 ;
        RECT -58.645 189.555 -58.315 189.885 ;
        RECT -58.645 188.195 -58.315 188.525 ;
        RECT -58.645 186.835 -58.315 187.165 ;
        RECT -58.645 185.475 -58.315 185.805 ;
        RECT -58.645 184.115 -58.315 184.445 ;
        RECT -58.645 182.755 -58.315 183.085 ;
        RECT -58.645 181.395 -58.315 181.725 ;
        RECT -58.645 180.035 -58.315 180.365 ;
        RECT -58.645 178.675 -58.315 179.005 ;
        RECT -58.645 177.315 -58.315 177.645 ;
        RECT -58.645 175.955 -58.315 176.285 ;
        RECT -58.645 174.595 -58.315 174.925 ;
        RECT -58.645 173.235 -58.315 173.565 ;
        RECT -58.645 171.875 -58.315 172.205 ;
        RECT -58.645 170.515 -58.315 170.845 ;
        RECT -58.645 169.155 -58.315 169.485 ;
        RECT -58.645 167.795 -58.315 168.125 ;
        RECT -58.645 166.435 -58.315 166.765 ;
        RECT -58.645 165.075 -58.315 165.405 ;
        RECT -58.645 163.715 -58.315 164.045 ;
        RECT -58.645 162.355 -58.315 162.685 ;
        RECT -58.645 160.995 -58.315 161.325 ;
        RECT -58.645 159.635 -58.315 159.965 ;
        RECT -58.645 158.275 -58.315 158.605 ;
        RECT -58.645 156.915 -58.315 157.245 ;
        RECT -58.645 155.555 -58.315 155.885 ;
        RECT -58.645 154.195 -58.315 154.525 ;
        RECT -58.645 152.835 -58.315 153.165 ;
        RECT -58.645 151.475 -58.315 151.805 ;
        RECT -58.645 150.115 -58.315 150.445 ;
        RECT -58.645 148.755 -58.315 149.085 ;
        RECT -58.645 147.395 -58.315 147.725 ;
        RECT -58.645 146.035 -58.315 146.365 ;
        RECT -58.645 144.675 -58.315 145.005 ;
        RECT -58.645 143.315 -58.315 143.645 ;
        RECT -58.645 141.955 -58.315 142.285 ;
        RECT -58.645 140.595 -58.315 140.925 ;
        RECT -58.645 139.235 -58.315 139.565 ;
        RECT -58.64 138.56 -58.32 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -58.645 53.555 -58.315 53.885 ;
        RECT -58.645 52.195 -58.315 52.525 ;
        RECT -58.645 50.835 -58.315 51.165 ;
        RECT -58.645 49.475 -58.315 49.805 ;
        RECT -58.645 48.115 -58.315 48.445 ;
        RECT -58.645 46.755 -58.315 47.085 ;
        RECT -58.645 45.395 -58.315 45.725 ;
        RECT -58.645 44.035 -58.315 44.365 ;
        RECT -58.645 42.675 -58.315 43.005 ;
        RECT -58.645 41.315 -58.315 41.645 ;
        RECT -58.645 39.955 -58.315 40.285 ;
        RECT -58.645 38.595 -58.315 38.925 ;
        RECT -58.645 37.235 -58.315 37.565 ;
        RECT -58.645 35.875 -58.315 36.205 ;
        RECT -58.645 34.515 -58.315 34.845 ;
        RECT -58.645 33.155 -58.315 33.485 ;
        RECT -58.645 31.795 -58.315 32.125 ;
        RECT -58.645 30.435 -58.315 30.765 ;
        RECT -58.645 29.075 -58.315 29.405 ;
        RECT -58.645 27.715 -58.315 28.045 ;
        RECT -58.645 26.355 -58.315 26.685 ;
        RECT -58.645 24.995 -58.315 25.325 ;
        RECT -58.645 23.635 -58.315 23.965 ;
        RECT -58.645 22.275 -58.315 22.605 ;
        RECT -58.645 20.915 -58.315 21.245 ;
        RECT -58.645 19.555 -58.315 19.885 ;
        RECT -58.645 18.195 -58.315 18.525 ;
        RECT -58.645 16.835 -58.315 17.165 ;
        RECT -58.645 15.475 -58.315 15.805 ;
        RECT -58.645 14.115 -58.315 14.445 ;
        RECT -58.645 12.755 -58.315 13.085 ;
        RECT -58.645 11.395 -58.315 11.725 ;
        RECT -58.645 10.035 -58.315 10.365 ;
        RECT -58.645 8.675 -58.315 9.005 ;
        RECT -58.645 7.315 -58.315 7.645 ;
        RECT -58.645 5.955 -58.315 6.285 ;
        RECT -58.645 4.595 -58.315 4.925 ;
        RECT -58.645 3.235 -58.315 3.565 ;
        RECT -58.645 1.875 -58.315 2.205 ;
        RECT -58.645 0.515 -58.315 0.845 ;
        RECT -58.645 -0.845 -58.315 -0.515 ;
        RECT -58.645 -2.205 -58.315 -1.875 ;
        RECT -58.645 -3.565 -58.315 -3.235 ;
        RECT -58.645 -4.925 -58.315 -4.595 ;
        RECT -58.645 -6.285 -58.315 -5.955 ;
        RECT -58.645 -7.645 -58.315 -7.315 ;
        RECT -58.645 -9.005 -58.315 -8.675 ;
        RECT -58.645 -10.365 -58.315 -10.035 ;
        RECT -58.645 -11.725 -58.315 -11.395 ;
        RECT -58.645 -13.085 -58.315 -12.755 ;
        RECT -58.645 -14.445 -58.315 -14.115 ;
        RECT -58.645 -15.805 -58.315 -15.475 ;
        RECT -58.645 -17.165 -58.315 -16.835 ;
        RECT -58.645 -18.525 -58.315 -18.195 ;
        RECT -58.645 -19.885 -58.315 -19.555 ;
        RECT -58.645 -21.245 -58.315 -20.915 ;
        RECT -58.645 -22.605 -58.315 -22.275 ;
        RECT -58.645 -23.965 -58.315 -23.635 ;
        RECT -58.645 -25.325 -58.315 -24.995 ;
        RECT -58.645 -29.405 -58.315 -29.075 ;
        RECT -58.645 -30.765 -58.315 -30.435 ;
        RECT -58.645 -32.125 -58.315 -31.795 ;
        RECT -58.645 -33.485 -58.315 -33.155 ;
        RECT -58.645 -34.845 -58.315 -34.515 ;
        RECT -58.645 -36.205 -58.315 -35.875 ;
        RECT -58.645 -37.565 -58.315 -37.235 ;
        RECT -58.645 -38.925 -58.315 -38.595 ;
        RECT -58.645 -40.285 -58.315 -39.955 ;
        RECT -58.645 -41.645 -58.315 -41.315 ;
        RECT -58.645 -43.005 -58.315 -42.675 ;
        RECT -58.645 -44.365 -58.315 -44.035 ;
        RECT -58.645 -45.725 -58.315 -45.395 ;
        RECT -58.645 -47.085 -58.315 -46.755 ;
        RECT -58.645 -48.445 -58.315 -48.115 ;
        RECT -58.645 -49.805 -58.315 -49.475 ;
        RECT -58.645 -51.165 -58.315 -50.835 ;
        RECT -58.645 -52.525 -58.315 -52.195 ;
        RECT -58.645 -53.885 -58.315 -53.555 ;
        RECT -58.645 -55.245 -58.315 -54.915 ;
        RECT -58.645 -56.605 -58.315 -56.275 ;
        RECT -58.645 -57.965 -58.315 -57.635 ;
        RECT -58.645 -59.325 -58.315 -58.995 ;
        RECT -58.645 -60.685 -58.315 -60.355 ;
        RECT -58.645 -62.045 -58.315 -61.715 ;
        RECT -58.645 -63.405 -58.315 -63.075 ;
        RECT -58.645 -64.765 -58.315 -64.435 ;
        RECT -58.645 -66.125 -58.315 -65.795 ;
        RECT -58.645 -67.485 -58.315 -67.155 ;
        RECT -58.645 -68.845 -58.315 -68.515 ;
        RECT -58.645 -70.205 -58.315 -69.875 ;
        RECT -58.645 -71.565 -58.315 -71.235 ;
        RECT -58.645 -72.925 -58.315 -72.595 ;
        RECT -58.645 -74.285 -58.315 -73.955 ;
        RECT -58.645 -75.645 -58.315 -75.315 ;
        RECT -58.645 -77.005 -58.315 -76.675 ;
        RECT -58.645 -78.365 -58.315 -78.035 ;
        RECT -58.645 -79.725 -58.315 -79.395 ;
        RECT -58.645 -81.085 -58.315 -80.755 ;
        RECT -58.645 -82.445 -58.315 -82.115 ;
        RECT -58.645 -83.805 -58.315 -83.475 ;
        RECT -58.645 -85.165 -58.315 -84.835 ;
        RECT -58.645 -86.525 -58.315 -86.195 ;
        RECT -58.645 -87.885 -58.315 -87.555 ;
        RECT -58.645 -89.245 -58.315 -88.915 ;
        RECT -58.645 -90.605 -58.315 -90.275 ;
        RECT -58.645 -91.77 -58.315 -91.44 ;
        RECT -58.645 -93.325 -58.315 -92.995 ;
        RECT -58.645 -94.685 -58.315 -94.355 ;
        RECT -58.645 -96.045 -58.315 -95.715 ;
        RECT -58.645 -97.405 -58.315 -97.075 ;
        RECT -58.645 -98.765 -58.315 -98.435 ;
        RECT -58.645 -101.485 -58.315 -101.155 ;
        RECT -58.645 -102.31 -58.315 -101.98 ;
        RECT -58.645 -104.205 -58.315 -103.875 ;
        RECT -58.645 -105.565 -58.315 -105.235 ;
        RECT -58.645 -106.925 -58.315 -106.595 ;
        RECT -58.645 -109.645 -58.315 -109.315 ;
        RECT -58.645 -111.005 -58.315 -110.675 ;
        RECT -58.64 -113.04 -58.32 98.08 ;
        RECT -58.645 97.075 -58.315 97.405 ;
        RECT -58.645 95.715 -58.315 96.045 ;
        RECT -58.645 94.355 -58.315 94.685 ;
        RECT -58.645 92.995 -58.315 93.325 ;
        RECT -58.645 88.915 -58.315 89.245 ;
        RECT -58.645 84.835 -58.315 85.165 ;
        RECT -58.645 83.475 -58.315 83.805 ;
        RECT -58.645 82.115 -58.315 82.445 ;
        RECT -58.645 80.755 -58.315 81.085 ;
        RECT -58.645 79.395 -58.315 79.725 ;
        RECT -58.645 78.035 -58.315 78.365 ;
        RECT -58.645 76.675 -58.315 77.005 ;
        RECT -58.645 75.315 -58.315 75.645 ;
        RECT -58.645 73.955 -58.315 74.285 ;
        RECT -58.645 72.595 -58.315 72.925 ;
        RECT -58.645 71.235 -58.315 71.565 ;
        RECT -58.645 69.875 -58.315 70.205 ;
        RECT -58.645 68.515 -58.315 68.845 ;
        RECT -58.645 67.155 -58.315 67.485 ;
        RECT -58.645 65.795 -58.315 66.125 ;
        RECT -58.645 64.435 -58.315 64.765 ;
        RECT -58.645 63.075 -58.315 63.405 ;
        RECT -58.645 61.715 -58.315 62.045 ;
        RECT -58.645 60.355 -58.315 60.685 ;
        RECT -58.645 58.995 -58.315 59.325 ;
        RECT -58.645 57.635 -58.315 57.965 ;
        RECT -58.645 56.275 -58.315 56.605 ;
        RECT -58.645 54.915 -58.315 55.245 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.165 -177.645 -67.835 -177.315 ;
        RECT -68.165 -179.005 -67.835 -178.675 ;
        RECT -68.165 -184.65 -67.835 -183.52 ;
        RECT -68.16 -184.765 -67.84 -175.28 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.805 244.04 -66.475 245.17 ;
        RECT -66.805 239.875 -66.475 240.205 ;
        RECT -66.805 238.515 -66.475 238.845 ;
        RECT -66.805 237.155 -66.475 237.485 ;
        RECT -66.805 235.795 -66.475 236.125 ;
        RECT -66.805 234.435 -66.475 234.765 ;
        RECT -66.805 233.075 -66.475 233.405 ;
        RECT -66.805 231.715 -66.475 232.045 ;
        RECT -66.805 230.355 -66.475 230.685 ;
        RECT -66.805 228.995 -66.475 229.325 ;
        RECT -66.805 227.635 -66.475 227.965 ;
        RECT -66.805 226.275 -66.475 226.605 ;
        RECT -66.805 224.915 -66.475 225.245 ;
        RECT -66.805 223.555 -66.475 223.885 ;
        RECT -66.805 222.195 -66.475 222.525 ;
        RECT -66.805 220.835 -66.475 221.165 ;
        RECT -66.805 219.475 -66.475 219.805 ;
        RECT -66.805 218.115 -66.475 218.445 ;
        RECT -66.805 216.755 -66.475 217.085 ;
        RECT -66.805 215.395 -66.475 215.725 ;
        RECT -66.805 214.035 -66.475 214.365 ;
        RECT -66.805 212.675 -66.475 213.005 ;
        RECT -66.805 211.315 -66.475 211.645 ;
        RECT -66.805 209.955 -66.475 210.285 ;
        RECT -66.805 208.595 -66.475 208.925 ;
        RECT -66.805 207.235 -66.475 207.565 ;
        RECT -66.805 205.875 -66.475 206.205 ;
        RECT -66.805 204.515 -66.475 204.845 ;
        RECT -66.805 203.155 -66.475 203.485 ;
        RECT -66.805 201.795 -66.475 202.125 ;
        RECT -66.805 200.435 -66.475 200.765 ;
        RECT -66.805 199.075 -66.475 199.405 ;
        RECT -66.805 197.715 -66.475 198.045 ;
        RECT -66.805 196.355 -66.475 196.685 ;
        RECT -66.805 194.995 -66.475 195.325 ;
        RECT -66.805 193.635 -66.475 193.965 ;
        RECT -66.805 192.275 -66.475 192.605 ;
        RECT -66.805 190.915 -66.475 191.245 ;
        RECT -66.805 189.555 -66.475 189.885 ;
        RECT -66.805 188.195 -66.475 188.525 ;
        RECT -66.805 186.835 -66.475 187.165 ;
        RECT -66.805 185.475 -66.475 185.805 ;
        RECT -66.805 184.115 -66.475 184.445 ;
        RECT -66.805 182.755 -66.475 183.085 ;
        RECT -66.805 181.395 -66.475 181.725 ;
        RECT -66.805 180.035 -66.475 180.365 ;
        RECT -66.805 178.675 -66.475 179.005 ;
        RECT -66.805 177.315 -66.475 177.645 ;
        RECT -66.805 175.955 -66.475 176.285 ;
        RECT -66.805 174.595 -66.475 174.925 ;
        RECT -66.805 173.235 -66.475 173.565 ;
        RECT -66.805 171.875 -66.475 172.205 ;
        RECT -66.805 170.515 -66.475 170.845 ;
        RECT -66.805 169.155 -66.475 169.485 ;
        RECT -66.805 167.795 -66.475 168.125 ;
        RECT -66.805 166.435 -66.475 166.765 ;
        RECT -66.805 165.075 -66.475 165.405 ;
        RECT -66.805 163.715 -66.475 164.045 ;
        RECT -66.805 162.355 -66.475 162.685 ;
        RECT -66.805 160.995 -66.475 161.325 ;
        RECT -66.805 159.635 -66.475 159.965 ;
        RECT -66.805 158.275 -66.475 158.605 ;
        RECT -66.805 156.915 -66.475 157.245 ;
        RECT -66.805 155.555 -66.475 155.885 ;
        RECT -66.805 154.195 -66.475 154.525 ;
        RECT -66.805 152.835 -66.475 153.165 ;
        RECT -66.805 151.475 -66.475 151.805 ;
        RECT -66.805 150.115 -66.475 150.445 ;
        RECT -66.805 148.755 -66.475 149.085 ;
        RECT -66.805 147.395 -66.475 147.725 ;
        RECT -66.805 146.035 -66.475 146.365 ;
        RECT -66.805 144.675 -66.475 145.005 ;
        RECT -66.805 143.315 -66.475 143.645 ;
        RECT -66.805 141.955 -66.475 142.285 ;
        RECT -66.805 140.595 -66.475 140.925 ;
        RECT -66.805 139.235 -66.475 139.565 ;
        RECT -66.805 137.875 -66.475 138.205 ;
        RECT -66.805 136.515 -66.475 136.845 ;
        RECT -66.805 135.155 -66.475 135.485 ;
        RECT -66.805 133.795 -66.475 134.125 ;
        RECT -66.805 132.435 -66.475 132.765 ;
        RECT -66.805 131.075 -66.475 131.405 ;
        RECT -66.805 129.715 -66.475 130.045 ;
        RECT -66.805 128.355 -66.475 128.685 ;
        RECT -66.805 126.995 -66.475 127.325 ;
        RECT -66.805 125.635 -66.475 125.965 ;
        RECT -66.805 124.275 -66.475 124.605 ;
        RECT -66.805 122.915 -66.475 123.245 ;
        RECT -66.805 121.555 -66.475 121.885 ;
        RECT -66.805 120.195 -66.475 120.525 ;
        RECT -66.805 118.835 -66.475 119.165 ;
        RECT -66.805 117.475 -66.475 117.805 ;
        RECT -66.805 116.115 -66.475 116.445 ;
        RECT -66.805 114.755 -66.475 115.085 ;
        RECT -66.805 113.395 -66.475 113.725 ;
        RECT -66.805 112.035 -66.475 112.365 ;
        RECT -66.805 110.675 -66.475 111.005 ;
        RECT -66.805 109.315 -66.475 109.645 ;
        RECT -66.805 107.955 -66.475 108.285 ;
        RECT -66.805 106.595 -66.475 106.925 ;
        RECT -66.805 105.235 -66.475 105.565 ;
        RECT -66.805 103.875 -66.475 104.205 ;
        RECT -66.805 102.515 -66.475 102.845 ;
        RECT -66.805 101.155 -66.475 101.485 ;
        RECT -66.805 99.795 -66.475 100.125 ;
        RECT -66.805 98.435 -66.475 98.765 ;
        RECT -66.805 97.075 -66.475 97.405 ;
        RECT -66.805 95.715 -66.475 96.045 ;
        RECT -66.805 94.355 -66.475 94.685 ;
        RECT -66.805 92.995 -66.475 93.325 ;
        RECT -66.805 91.635 -66.475 91.965 ;
        RECT -66.805 90.275 -66.475 90.605 ;
        RECT -66.805 88.915 -66.475 89.245 ;
        RECT -66.805 87.555 -66.475 87.885 ;
        RECT -66.805 86.195 -66.475 86.525 ;
        RECT -66.805 84.835 -66.475 85.165 ;
        RECT -66.805 83.475 -66.475 83.805 ;
        RECT -66.805 82.115 -66.475 82.445 ;
        RECT -66.805 80.755 -66.475 81.085 ;
        RECT -66.805 79.395 -66.475 79.725 ;
        RECT -66.805 78.035 -66.475 78.365 ;
        RECT -66.805 76.675 -66.475 77.005 ;
        RECT -66.805 75.315 -66.475 75.645 ;
        RECT -66.805 73.955 -66.475 74.285 ;
        RECT -66.805 72.595 -66.475 72.925 ;
        RECT -66.805 71.235 -66.475 71.565 ;
        RECT -66.805 69.875 -66.475 70.205 ;
        RECT -66.805 68.515 -66.475 68.845 ;
        RECT -66.805 67.155 -66.475 67.485 ;
        RECT -66.805 65.795 -66.475 66.125 ;
        RECT -66.805 64.435 -66.475 64.765 ;
        RECT -66.805 63.075 -66.475 63.405 ;
        RECT -66.805 61.715 -66.475 62.045 ;
        RECT -66.805 60.355 -66.475 60.685 ;
        RECT -66.805 58.995 -66.475 59.325 ;
        RECT -66.805 57.635 -66.475 57.965 ;
        RECT -66.805 56.275 -66.475 56.605 ;
        RECT -66.805 54.915 -66.475 55.245 ;
        RECT -66.805 53.555 -66.475 53.885 ;
        RECT -66.805 52.195 -66.475 52.525 ;
        RECT -66.805 50.835 -66.475 51.165 ;
        RECT -66.805 49.475 -66.475 49.805 ;
        RECT -66.805 48.115 -66.475 48.445 ;
        RECT -66.805 46.755 -66.475 47.085 ;
        RECT -66.805 45.395 -66.475 45.725 ;
        RECT -66.805 44.035 -66.475 44.365 ;
        RECT -66.805 42.675 -66.475 43.005 ;
        RECT -66.805 41.315 -66.475 41.645 ;
        RECT -66.805 39.955 -66.475 40.285 ;
        RECT -66.805 38.595 -66.475 38.925 ;
        RECT -66.805 37.235 -66.475 37.565 ;
        RECT -66.805 35.875 -66.475 36.205 ;
        RECT -66.805 34.515 -66.475 34.845 ;
        RECT -66.805 33.155 -66.475 33.485 ;
        RECT -66.805 31.795 -66.475 32.125 ;
        RECT -66.805 30.435 -66.475 30.765 ;
        RECT -66.805 29.075 -66.475 29.405 ;
        RECT -66.805 27.715 -66.475 28.045 ;
        RECT -66.805 26.355 -66.475 26.685 ;
        RECT -66.805 24.995 -66.475 25.325 ;
        RECT -66.805 23.635 -66.475 23.965 ;
        RECT -66.805 22.275 -66.475 22.605 ;
        RECT -66.805 20.915 -66.475 21.245 ;
        RECT -66.805 19.555 -66.475 19.885 ;
        RECT -66.805 18.195 -66.475 18.525 ;
        RECT -66.805 16.835 -66.475 17.165 ;
        RECT -66.805 15.475 -66.475 15.805 ;
        RECT -66.805 14.115 -66.475 14.445 ;
        RECT -66.805 12.755 -66.475 13.085 ;
        RECT -66.805 11.395 -66.475 11.725 ;
        RECT -66.805 10.035 -66.475 10.365 ;
        RECT -66.805 8.675 -66.475 9.005 ;
        RECT -66.805 7.315 -66.475 7.645 ;
        RECT -66.805 5.955 -66.475 6.285 ;
        RECT -66.805 4.595 -66.475 4.925 ;
        RECT -66.805 3.235 -66.475 3.565 ;
        RECT -66.805 1.875 -66.475 2.205 ;
        RECT -66.805 0.515 -66.475 0.845 ;
        RECT -66.805 -0.845 -66.475 -0.515 ;
        RECT -66.805 -2.205 -66.475 -1.875 ;
        RECT -66.805 -3.565 -66.475 -3.235 ;
        RECT -66.805 -4.925 -66.475 -4.595 ;
        RECT -66.805 -6.285 -66.475 -5.955 ;
        RECT -66.805 -7.645 -66.475 -7.315 ;
        RECT -66.805 -9.005 -66.475 -8.675 ;
        RECT -66.805 -10.365 -66.475 -10.035 ;
        RECT -66.805 -11.725 -66.475 -11.395 ;
        RECT -66.805 -13.085 -66.475 -12.755 ;
        RECT -66.805 -14.445 -66.475 -14.115 ;
        RECT -66.805 -15.805 -66.475 -15.475 ;
        RECT -66.805 -17.165 -66.475 -16.835 ;
        RECT -66.805 -18.525 -66.475 -18.195 ;
        RECT -66.805 -19.885 -66.475 -19.555 ;
        RECT -66.805 -21.245 -66.475 -20.915 ;
        RECT -66.805 -22.605 -66.475 -22.275 ;
        RECT -66.805 -23.965 -66.475 -23.635 ;
        RECT -66.805 -25.325 -66.475 -24.995 ;
        RECT -66.805 -28.045 -66.475 -27.715 ;
        RECT -66.805 -29.405 -66.475 -29.075 ;
        RECT -66.805 -30.765 -66.475 -30.435 ;
        RECT -66.805 -32.125 -66.475 -31.795 ;
        RECT -66.805 -33.485 -66.475 -33.155 ;
        RECT -66.805 -34.845 -66.475 -34.515 ;
        RECT -66.805 -36.205 -66.475 -35.875 ;
        RECT -66.805 -37.565 -66.475 -37.235 ;
        RECT -66.805 -38.925 -66.475 -38.595 ;
        RECT -66.805 -40.285 -66.475 -39.955 ;
        RECT -66.805 -41.645 -66.475 -41.315 ;
        RECT -66.805 -43.005 -66.475 -42.675 ;
        RECT -66.805 -44.365 -66.475 -44.035 ;
        RECT -66.805 -45.725 -66.475 -45.395 ;
        RECT -66.805 -47.085 -66.475 -46.755 ;
        RECT -66.805 -48.445 -66.475 -48.115 ;
        RECT -66.805 -49.805 -66.475 -49.475 ;
        RECT -66.805 -51.165 -66.475 -50.835 ;
        RECT -66.805 -52.525 -66.475 -52.195 ;
        RECT -66.805 -53.885 -66.475 -53.555 ;
        RECT -66.805 -55.245 -66.475 -54.915 ;
        RECT -66.805 -56.605 -66.475 -56.275 ;
        RECT -66.805 -57.965 -66.475 -57.635 ;
        RECT -66.805 -59.325 -66.475 -58.995 ;
        RECT -66.805 -60.685 -66.475 -60.355 ;
        RECT -66.805 -62.045 -66.475 -61.715 ;
        RECT -66.805 -63.405 -66.475 -63.075 ;
        RECT -66.805 -64.765 -66.475 -64.435 ;
        RECT -66.805 -66.125 -66.475 -65.795 ;
        RECT -66.805 -67.485 -66.475 -67.155 ;
        RECT -66.805 -68.845 -66.475 -68.515 ;
        RECT -66.805 -70.205 -66.475 -69.875 ;
        RECT -66.805 -71.565 -66.475 -71.235 ;
        RECT -66.805 -72.925 -66.475 -72.595 ;
        RECT -66.805 -74.285 -66.475 -73.955 ;
        RECT -66.805 -75.645 -66.475 -75.315 ;
        RECT -66.805 -77.005 -66.475 -76.675 ;
        RECT -66.805 -78.365 -66.475 -78.035 ;
        RECT -66.805 -79.725 -66.475 -79.395 ;
        RECT -66.805 -81.085 -66.475 -80.755 ;
        RECT -66.805 -82.445 -66.475 -82.115 ;
        RECT -66.805 -83.805 -66.475 -83.475 ;
        RECT -66.805 -85.165 -66.475 -84.835 ;
        RECT -66.805 -86.525 -66.475 -86.195 ;
        RECT -66.805 -87.885 -66.475 -87.555 ;
        RECT -66.805 -89.245 -66.475 -88.915 ;
        RECT -66.805 -90.605 -66.475 -90.275 ;
        RECT -66.805 -91.77 -66.475 -91.44 ;
        RECT -66.805 -93.325 -66.475 -92.995 ;
        RECT -66.805 -94.685 -66.475 -94.355 ;
        RECT -66.805 -96.045 -66.475 -95.715 ;
        RECT -66.805 -97.405 -66.475 -97.075 ;
        RECT -66.805 -98.765 -66.475 -98.435 ;
        RECT -66.805 -101.485 -66.475 -101.155 ;
        RECT -66.805 -102.31 -66.475 -101.98 ;
        RECT -66.805 -104.205 -66.475 -103.875 ;
        RECT -66.805 -105.565 -66.475 -105.235 ;
        RECT -66.805 -106.925 -66.475 -106.595 ;
        RECT -66.805 -109.645 -66.475 -109.315 ;
        RECT -66.805 -111.005 -66.475 -110.675 ;
        RECT -66.805 -113.725 -66.475 -113.395 ;
        RECT -66.805 -115.085 -66.475 -114.755 ;
        RECT -66.805 -116.445 -66.475 -116.115 ;
        RECT -66.805 -117.805 -66.475 -117.475 ;
        RECT -66.805 -119.165 -66.475 -118.835 ;
        RECT -66.805 -120.525 -66.475 -120.195 ;
        RECT -66.805 -123.245 -66.475 -122.915 ;
        RECT -66.805 -124.605 -66.475 -124.275 ;
        RECT -66.805 -125.965 -66.475 -125.635 ;
        RECT -66.805 -127.325 -66.475 -126.995 ;
        RECT -66.805 -128.685 -66.475 -128.355 ;
        RECT -66.805 -130.045 -66.475 -129.715 ;
        RECT -66.805 -131.405 -66.475 -131.075 ;
        RECT -66.805 -132.765 -66.475 -132.435 ;
        RECT -66.805 -134.125 -66.475 -133.795 ;
        RECT -66.805 -135.485 -66.475 -135.155 ;
        RECT -66.805 -136.845 -66.475 -136.515 ;
        RECT -66.805 -138.205 -66.475 -137.875 ;
        RECT -66.805 -139.565 -66.475 -139.235 ;
        RECT -66.805 -140.925 -66.475 -140.595 ;
        RECT -66.805 -142.285 -66.475 -141.955 ;
        RECT -66.805 -143.645 -66.475 -143.315 ;
        RECT -66.805 -145.005 -66.475 -144.675 ;
        RECT -66.805 -146.365 -66.475 -146.035 ;
        RECT -66.805 -147.725 -66.475 -147.395 ;
        RECT -66.805 -149.085 -66.475 -148.755 ;
        RECT -66.805 -150.445 -66.475 -150.115 ;
        RECT -66.805 -151.805 -66.475 -151.475 ;
        RECT -66.805 -153.165 -66.475 -152.835 ;
        RECT -66.805 -154.525 -66.475 -154.195 ;
        RECT -66.805 -155.885 -66.475 -155.555 ;
        RECT -66.805 -157.245 -66.475 -156.915 ;
        RECT -66.805 -158.605 -66.475 -158.275 ;
        RECT -66.805 -159.965 -66.475 -159.635 ;
        RECT -66.805 -161.325 -66.475 -160.995 ;
        RECT -66.805 -162.685 -66.475 -162.355 ;
        RECT -66.805 -164.045 -66.475 -163.715 ;
        RECT -66.805 -165.405 -66.475 -165.075 ;
        RECT -66.805 -166.765 -66.475 -166.435 ;
        RECT -66.805 -169.615 -66.475 -169.285 ;
        RECT -66.805 -170.845 -66.475 -170.515 ;
        RECT -66.805 -172.205 -66.475 -171.875 ;
        RECT -66.805 -177.645 -66.475 -177.315 ;
        RECT -66.805 -179.005 -66.475 -178.675 ;
        RECT -66.805 -184.65 -66.475 -183.52 ;
        RECT -66.8 -184.765 -66.48 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -65.445 244.04 -65.115 245.17 ;
        RECT -65.445 239.875 -65.115 240.205 ;
        RECT -65.445 238.515 -65.115 238.845 ;
        RECT -65.445 237.155 -65.115 237.485 ;
        RECT -65.445 235.795 -65.115 236.125 ;
        RECT -65.445 234.435 -65.115 234.765 ;
        RECT -65.445 233.075 -65.115 233.405 ;
        RECT -65.445 231.715 -65.115 232.045 ;
        RECT -65.445 230.355 -65.115 230.685 ;
        RECT -65.445 228.995 -65.115 229.325 ;
        RECT -65.445 227.635 -65.115 227.965 ;
        RECT -65.445 226.275 -65.115 226.605 ;
        RECT -65.445 224.915 -65.115 225.245 ;
        RECT -65.445 223.555 -65.115 223.885 ;
        RECT -65.445 222.195 -65.115 222.525 ;
        RECT -65.445 220.835 -65.115 221.165 ;
        RECT -65.445 219.475 -65.115 219.805 ;
        RECT -65.445 218.115 -65.115 218.445 ;
        RECT -65.445 216.755 -65.115 217.085 ;
        RECT -65.445 215.395 -65.115 215.725 ;
        RECT -65.445 214.035 -65.115 214.365 ;
        RECT -65.445 212.675 -65.115 213.005 ;
        RECT -65.445 211.315 -65.115 211.645 ;
        RECT -65.445 209.955 -65.115 210.285 ;
        RECT -65.445 208.595 -65.115 208.925 ;
        RECT -65.445 207.235 -65.115 207.565 ;
        RECT -65.445 205.875 -65.115 206.205 ;
        RECT -65.445 204.515 -65.115 204.845 ;
        RECT -65.445 203.155 -65.115 203.485 ;
        RECT -65.445 201.795 -65.115 202.125 ;
        RECT -65.445 200.435 -65.115 200.765 ;
        RECT -65.445 199.075 -65.115 199.405 ;
        RECT -65.445 197.715 -65.115 198.045 ;
        RECT -65.445 196.355 -65.115 196.685 ;
        RECT -65.445 194.995 -65.115 195.325 ;
        RECT -65.445 193.635 -65.115 193.965 ;
        RECT -65.445 192.275 -65.115 192.605 ;
        RECT -65.445 190.915 -65.115 191.245 ;
        RECT -65.445 189.555 -65.115 189.885 ;
        RECT -65.445 188.195 -65.115 188.525 ;
        RECT -65.445 186.835 -65.115 187.165 ;
        RECT -65.445 185.475 -65.115 185.805 ;
        RECT -65.445 184.115 -65.115 184.445 ;
        RECT -65.445 182.755 -65.115 183.085 ;
        RECT -65.445 181.395 -65.115 181.725 ;
        RECT -65.445 180.035 -65.115 180.365 ;
        RECT -65.445 178.675 -65.115 179.005 ;
        RECT -65.445 177.315 -65.115 177.645 ;
        RECT -65.445 175.955 -65.115 176.285 ;
        RECT -65.445 174.595 -65.115 174.925 ;
        RECT -65.445 173.235 -65.115 173.565 ;
        RECT -65.445 171.875 -65.115 172.205 ;
        RECT -65.445 170.515 -65.115 170.845 ;
        RECT -65.445 169.155 -65.115 169.485 ;
        RECT -65.445 167.795 -65.115 168.125 ;
        RECT -65.445 166.435 -65.115 166.765 ;
        RECT -65.445 165.075 -65.115 165.405 ;
        RECT -65.445 163.715 -65.115 164.045 ;
        RECT -65.445 162.355 -65.115 162.685 ;
        RECT -65.445 160.995 -65.115 161.325 ;
        RECT -65.445 159.635 -65.115 159.965 ;
        RECT -65.445 158.275 -65.115 158.605 ;
        RECT -65.445 156.915 -65.115 157.245 ;
        RECT -65.445 155.555 -65.115 155.885 ;
        RECT -65.445 154.195 -65.115 154.525 ;
        RECT -65.445 152.835 -65.115 153.165 ;
        RECT -65.445 151.475 -65.115 151.805 ;
        RECT -65.445 150.115 -65.115 150.445 ;
        RECT -65.445 148.755 -65.115 149.085 ;
        RECT -65.445 147.395 -65.115 147.725 ;
        RECT -65.445 146.035 -65.115 146.365 ;
        RECT -65.445 144.675 -65.115 145.005 ;
        RECT -65.445 143.315 -65.115 143.645 ;
        RECT -65.445 141.955 -65.115 142.285 ;
        RECT -65.445 140.595 -65.115 140.925 ;
        RECT -65.445 139.235 -65.115 139.565 ;
        RECT -65.445 137.875 -65.115 138.205 ;
        RECT -65.445 136.515 -65.115 136.845 ;
        RECT -65.445 135.155 -65.115 135.485 ;
        RECT -65.445 133.795 -65.115 134.125 ;
        RECT -65.445 132.435 -65.115 132.765 ;
        RECT -65.445 131.075 -65.115 131.405 ;
        RECT -65.445 129.715 -65.115 130.045 ;
        RECT -65.445 128.355 -65.115 128.685 ;
        RECT -65.445 126.995 -65.115 127.325 ;
        RECT -65.445 125.635 -65.115 125.965 ;
        RECT -65.445 124.275 -65.115 124.605 ;
        RECT -65.445 122.915 -65.115 123.245 ;
        RECT -65.445 121.555 -65.115 121.885 ;
        RECT -65.445 120.195 -65.115 120.525 ;
        RECT -65.445 118.835 -65.115 119.165 ;
        RECT -65.445 117.475 -65.115 117.805 ;
        RECT -65.445 116.115 -65.115 116.445 ;
        RECT -65.445 114.755 -65.115 115.085 ;
        RECT -65.445 113.395 -65.115 113.725 ;
        RECT -65.445 112.035 -65.115 112.365 ;
        RECT -65.445 110.675 -65.115 111.005 ;
        RECT -65.445 109.315 -65.115 109.645 ;
        RECT -65.445 107.955 -65.115 108.285 ;
        RECT -65.445 106.595 -65.115 106.925 ;
        RECT -65.445 105.235 -65.115 105.565 ;
        RECT -65.445 103.875 -65.115 104.205 ;
        RECT -65.445 102.515 -65.115 102.845 ;
        RECT -65.445 101.155 -65.115 101.485 ;
        RECT -65.445 99.795 -65.115 100.125 ;
        RECT -65.445 98.435 -65.115 98.765 ;
        RECT -65.445 97.075 -65.115 97.405 ;
        RECT -65.445 95.715 -65.115 96.045 ;
        RECT -65.445 94.355 -65.115 94.685 ;
        RECT -65.445 92.995 -65.115 93.325 ;
        RECT -65.445 91.635 -65.115 91.965 ;
        RECT -65.445 90.275 -65.115 90.605 ;
        RECT -65.445 88.915 -65.115 89.245 ;
        RECT -65.445 87.555 -65.115 87.885 ;
        RECT -65.445 86.195 -65.115 86.525 ;
        RECT -65.445 84.835 -65.115 85.165 ;
        RECT -65.445 83.475 -65.115 83.805 ;
        RECT -65.445 82.115 -65.115 82.445 ;
        RECT -65.445 80.755 -65.115 81.085 ;
        RECT -65.445 79.395 -65.115 79.725 ;
        RECT -65.445 78.035 -65.115 78.365 ;
        RECT -65.445 76.675 -65.115 77.005 ;
        RECT -65.445 75.315 -65.115 75.645 ;
        RECT -65.445 73.955 -65.115 74.285 ;
        RECT -65.445 72.595 -65.115 72.925 ;
        RECT -65.445 71.235 -65.115 71.565 ;
        RECT -65.445 69.875 -65.115 70.205 ;
        RECT -65.445 68.515 -65.115 68.845 ;
        RECT -65.445 67.155 -65.115 67.485 ;
        RECT -65.445 65.795 -65.115 66.125 ;
        RECT -65.445 64.435 -65.115 64.765 ;
        RECT -65.445 63.075 -65.115 63.405 ;
        RECT -65.445 61.715 -65.115 62.045 ;
        RECT -65.445 60.355 -65.115 60.685 ;
        RECT -65.445 58.995 -65.115 59.325 ;
        RECT -65.445 57.635 -65.115 57.965 ;
        RECT -65.445 56.275 -65.115 56.605 ;
        RECT -65.445 54.915 -65.115 55.245 ;
        RECT -65.445 53.555 -65.115 53.885 ;
        RECT -65.445 52.195 -65.115 52.525 ;
        RECT -65.445 50.835 -65.115 51.165 ;
        RECT -65.445 49.475 -65.115 49.805 ;
        RECT -65.445 48.115 -65.115 48.445 ;
        RECT -65.445 46.755 -65.115 47.085 ;
        RECT -65.445 45.395 -65.115 45.725 ;
        RECT -65.445 44.035 -65.115 44.365 ;
        RECT -65.445 42.675 -65.115 43.005 ;
        RECT -65.445 41.315 -65.115 41.645 ;
        RECT -65.445 39.955 -65.115 40.285 ;
        RECT -65.445 38.595 -65.115 38.925 ;
        RECT -65.445 37.235 -65.115 37.565 ;
        RECT -65.445 35.875 -65.115 36.205 ;
        RECT -65.445 34.515 -65.115 34.845 ;
        RECT -65.445 33.155 -65.115 33.485 ;
        RECT -65.445 31.795 -65.115 32.125 ;
        RECT -65.445 30.435 -65.115 30.765 ;
        RECT -65.445 29.075 -65.115 29.405 ;
        RECT -65.445 27.715 -65.115 28.045 ;
        RECT -65.445 26.355 -65.115 26.685 ;
        RECT -65.445 24.995 -65.115 25.325 ;
        RECT -65.445 23.635 -65.115 23.965 ;
        RECT -65.445 22.275 -65.115 22.605 ;
        RECT -65.445 20.915 -65.115 21.245 ;
        RECT -65.445 19.555 -65.115 19.885 ;
        RECT -65.445 18.195 -65.115 18.525 ;
        RECT -65.445 16.835 -65.115 17.165 ;
        RECT -65.445 15.475 -65.115 15.805 ;
        RECT -65.445 14.115 -65.115 14.445 ;
        RECT -65.445 12.755 -65.115 13.085 ;
        RECT -65.445 11.395 -65.115 11.725 ;
        RECT -65.445 10.035 -65.115 10.365 ;
        RECT -65.445 8.675 -65.115 9.005 ;
        RECT -65.445 7.315 -65.115 7.645 ;
        RECT -65.445 5.955 -65.115 6.285 ;
        RECT -65.445 4.595 -65.115 4.925 ;
        RECT -65.445 3.235 -65.115 3.565 ;
        RECT -65.445 1.875 -65.115 2.205 ;
        RECT -65.445 0.515 -65.115 0.845 ;
        RECT -65.445 -0.845 -65.115 -0.515 ;
        RECT -65.445 -2.205 -65.115 -1.875 ;
        RECT -65.445 -3.565 -65.115 -3.235 ;
        RECT -65.445 -4.925 -65.115 -4.595 ;
        RECT -65.445 -6.285 -65.115 -5.955 ;
        RECT -65.445 -7.645 -65.115 -7.315 ;
        RECT -65.445 -9.005 -65.115 -8.675 ;
        RECT -65.445 -10.365 -65.115 -10.035 ;
        RECT -65.445 -11.725 -65.115 -11.395 ;
        RECT -65.445 -13.085 -65.115 -12.755 ;
        RECT -65.445 -14.445 -65.115 -14.115 ;
        RECT -65.445 -15.805 -65.115 -15.475 ;
        RECT -65.445 -17.165 -65.115 -16.835 ;
        RECT -65.445 -18.525 -65.115 -18.195 ;
        RECT -65.445 -19.885 -65.115 -19.555 ;
        RECT -65.445 -21.245 -65.115 -20.915 ;
        RECT -65.445 -22.605 -65.115 -22.275 ;
        RECT -65.445 -23.965 -65.115 -23.635 ;
        RECT -65.445 -25.325 -65.115 -24.995 ;
        RECT -65.445 -28.045 -65.115 -27.715 ;
        RECT -65.445 -29.405 -65.115 -29.075 ;
        RECT -65.445 -30.765 -65.115 -30.435 ;
        RECT -65.445 -32.125 -65.115 -31.795 ;
        RECT -65.445 -33.485 -65.115 -33.155 ;
        RECT -65.445 -34.845 -65.115 -34.515 ;
        RECT -65.445 -36.205 -65.115 -35.875 ;
        RECT -65.445 -37.565 -65.115 -37.235 ;
        RECT -65.445 -38.925 -65.115 -38.595 ;
        RECT -65.445 -40.285 -65.115 -39.955 ;
        RECT -65.445 -41.645 -65.115 -41.315 ;
        RECT -65.445 -43.005 -65.115 -42.675 ;
        RECT -65.445 -44.365 -65.115 -44.035 ;
        RECT -65.445 -45.725 -65.115 -45.395 ;
        RECT -65.445 -47.085 -65.115 -46.755 ;
        RECT -65.445 -48.445 -65.115 -48.115 ;
        RECT -65.445 -49.805 -65.115 -49.475 ;
        RECT -65.445 -51.165 -65.115 -50.835 ;
        RECT -65.445 -52.525 -65.115 -52.195 ;
        RECT -65.445 -53.885 -65.115 -53.555 ;
        RECT -65.445 -55.245 -65.115 -54.915 ;
        RECT -65.445 -56.605 -65.115 -56.275 ;
        RECT -65.445 -57.965 -65.115 -57.635 ;
        RECT -65.445 -59.325 -65.115 -58.995 ;
        RECT -65.445 -60.685 -65.115 -60.355 ;
        RECT -65.445 -62.045 -65.115 -61.715 ;
        RECT -65.445 -63.405 -65.115 -63.075 ;
        RECT -65.445 -64.765 -65.115 -64.435 ;
        RECT -65.445 -66.125 -65.115 -65.795 ;
        RECT -65.445 -67.485 -65.115 -67.155 ;
        RECT -65.445 -68.845 -65.115 -68.515 ;
        RECT -65.445 -70.205 -65.115 -69.875 ;
        RECT -65.445 -71.565 -65.115 -71.235 ;
        RECT -65.445 -72.925 -65.115 -72.595 ;
        RECT -65.445 -74.285 -65.115 -73.955 ;
        RECT -65.445 -75.645 -65.115 -75.315 ;
        RECT -65.445 -77.005 -65.115 -76.675 ;
        RECT -65.445 -78.365 -65.115 -78.035 ;
        RECT -65.445 -79.725 -65.115 -79.395 ;
        RECT -65.445 -81.085 -65.115 -80.755 ;
        RECT -65.445 -82.445 -65.115 -82.115 ;
        RECT -65.445 -83.805 -65.115 -83.475 ;
        RECT -65.445 -85.165 -65.115 -84.835 ;
        RECT -65.445 -86.525 -65.115 -86.195 ;
        RECT -65.445 -87.885 -65.115 -87.555 ;
        RECT -65.445 -89.245 -65.115 -88.915 ;
        RECT -65.445 -90.605 -65.115 -90.275 ;
        RECT -65.445 -91.77 -65.115 -91.44 ;
        RECT -65.445 -93.325 -65.115 -92.995 ;
        RECT -65.445 -94.685 -65.115 -94.355 ;
        RECT -65.445 -96.045 -65.115 -95.715 ;
        RECT -65.445 -97.405 -65.115 -97.075 ;
        RECT -65.445 -98.765 -65.115 -98.435 ;
        RECT -65.445 -101.485 -65.115 -101.155 ;
        RECT -65.445 -102.31 -65.115 -101.98 ;
        RECT -65.445 -104.205 -65.115 -103.875 ;
        RECT -65.445 -105.565 -65.115 -105.235 ;
        RECT -65.445 -106.925 -65.115 -106.595 ;
        RECT -65.445 -109.645 -65.115 -109.315 ;
        RECT -65.445 -111.005 -65.115 -110.675 ;
        RECT -65.445 -113.725 -65.115 -113.395 ;
        RECT -65.445 -115.085 -65.115 -114.755 ;
        RECT -65.445 -116.445 -65.115 -116.115 ;
        RECT -65.445 -117.805 -65.115 -117.475 ;
        RECT -65.445 -119.165 -65.115 -118.835 ;
        RECT -65.445 -120.525 -65.115 -120.195 ;
        RECT -65.445 -123.245 -65.115 -122.915 ;
        RECT -65.445 -124.605 -65.115 -124.275 ;
        RECT -65.445 -125.965 -65.115 -125.635 ;
        RECT -65.445 -127.325 -65.115 -126.995 ;
        RECT -65.445 -128.685 -65.115 -128.355 ;
        RECT -65.445 -130.045 -65.115 -129.715 ;
        RECT -65.445 -131.405 -65.115 -131.075 ;
        RECT -65.445 -132.765 -65.115 -132.435 ;
        RECT -65.445 -134.125 -65.115 -133.795 ;
        RECT -65.445 -135.485 -65.115 -135.155 ;
        RECT -65.445 -136.845 -65.115 -136.515 ;
        RECT -65.445 -138.205 -65.115 -137.875 ;
        RECT -65.445 -139.565 -65.115 -139.235 ;
        RECT -65.445 -140.925 -65.115 -140.595 ;
        RECT -65.445 -142.285 -65.115 -141.955 ;
        RECT -65.445 -143.645 -65.115 -143.315 ;
        RECT -65.445 -145.005 -65.115 -144.675 ;
        RECT -65.445 -146.365 -65.115 -146.035 ;
        RECT -65.445 -147.725 -65.115 -147.395 ;
        RECT -65.445 -149.085 -65.115 -148.755 ;
        RECT -65.445 -150.445 -65.115 -150.115 ;
        RECT -65.445 -151.805 -65.115 -151.475 ;
        RECT -65.445 -153.165 -65.115 -152.835 ;
        RECT -65.445 -154.525 -65.115 -154.195 ;
        RECT -65.445 -155.885 -65.115 -155.555 ;
        RECT -65.445 -157.245 -65.115 -156.915 ;
        RECT -65.445 -158.605 -65.115 -158.275 ;
        RECT -65.445 -159.965 -65.115 -159.635 ;
        RECT -65.445 -161.325 -65.115 -160.995 ;
        RECT -65.445 -162.685 -65.115 -162.355 ;
        RECT -65.445 -164.045 -65.115 -163.715 ;
        RECT -65.445 -165.405 -65.115 -165.075 ;
        RECT -65.445 -166.765 -65.115 -166.435 ;
        RECT -65.445 -169.615 -65.115 -169.285 ;
        RECT -65.445 -170.845 -65.115 -170.515 ;
        RECT -65.445 -172.205 -65.115 -171.875 ;
        RECT -65.445 -177.645 -65.115 -177.315 ;
        RECT -65.445 -179.005 -65.115 -178.675 ;
        RECT -65.445 -184.65 -65.115 -183.52 ;
        RECT -65.44 -184.765 -65.12 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.085 97.075 -63.755 97.405 ;
        RECT -64.085 95.715 -63.755 96.045 ;
        RECT -64.085 94.355 -63.755 94.685 ;
        RECT -64.085 92.995 -63.755 93.325 ;
        RECT -64.085 91.635 -63.755 91.965 ;
        RECT -64.085 90.275 -63.755 90.605 ;
        RECT -64.085 88.915 -63.755 89.245 ;
        RECT -64.085 87.555 -63.755 87.885 ;
        RECT -64.085 86.195 -63.755 86.525 ;
        RECT -64.085 84.835 -63.755 85.165 ;
        RECT -64.085 83.475 -63.755 83.805 ;
        RECT -64.085 82.115 -63.755 82.445 ;
        RECT -64.085 80.755 -63.755 81.085 ;
        RECT -64.085 79.395 -63.755 79.725 ;
        RECT -64.085 78.035 -63.755 78.365 ;
        RECT -64.085 76.675 -63.755 77.005 ;
        RECT -64.085 75.315 -63.755 75.645 ;
        RECT -64.085 73.955 -63.755 74.285 ;
        RECT -64.085 72.595 -63.755 72.925 ;
        RECT -64.085 71.235 -63.755 71.565 ;
        RECT -64.085 69.875 -63.755 70.205 ;
        RECT -64.085 68.515 -63.755 68.845 ;
        RECT -64.085 67.155 -63.755 67.485 ;
        RECT -64.085 65.795 -63.755 66.125 ;
        RECT -64.085 64.435 -63.755 64.765 ;
        RECT -64.085 63.075 -63.755 63.405 ;
        RECT -64.085 61.715 -63.755 62.045 ;
        RECT -64.085 60.355 -63.755 60.685 ;
        RECT -64.085 58.995 -63.755 59.325 ;
        RECT -64.085 57.635 -63.755 57.965 ;
        RECT -64.085 56.275 -63.755 56.605 ;
        RECT -64.085 54.915 -63.755 55.245 ;
        RECT -64.085 53.555 -63.755 53.885 ;
        RECT -64.085 52.195 -63.755 52.525 ;
        RECT -64.085 50.835 -63.755 51.165 ;
        RECT -64.085 49.475 -63.755 49.805 ;
        RECT -64.085 48.115 -63.755 48.445 ;
        RECT -64.085 46.755 -63.755 47.085 ;
        RECT -64.085 45.395 -63.755 45.725 ;
        RECT -64.085 44.035 -63.755 44.365 ;
        RECT -64.085 42.675 -63.755 43.005 ;
        RECT -64.085 41.315 -63.755 41.645 ;
        RECT -64.085 39.955 -63.755 40.285 ;
        RECT -64.085 38.595 -63.755 38.925 ;
        RECT -64.085 37.235 -63.755 37.565 ;
        RECT -64.085 35.875 -63.755 36.205 ;
        RECT -64.085 34.515 -63.755 34.845 ;
        RECT -64.085 33.155 -63.755 33.485 ;
        RECT -64.085 31.795 -63.755 32.125 ;
        RECT -64.085 30.435 -63.755 30.765 ;
        RECT -64.085 29.075 -63.755 29.405 ;
        RECT -64.085 27.715 -63.755 28.045 ;
        RECT -64.085 26.355 -63.755 26.685 ;
        RECT -64.085 24.995 -63.755 25.325 ;
        RECT -64.085 23.635 -63.755 23.965 ;
        RECT -64.085 22.275 -63.755 22.605 ;
        RECT -64.085 20.915 -63.755 21.245 ;
        RECT -64.085 19.555 -63.755 19.885 ;
        RECT -64.085 18.195 -63.755 18.525 ;
        RECT -64.085 16.835 -63.755 17.165 ;
        RECT -64.085 15.475 -63.755 15.805 ;
        RECT -64.085 14.115 -63.755 14.445 ;
        RECT -64.085 12.755 -63.755 13.085 ;
        RECT -64.085 11.395 -63.755 11.725 ;
        RECT -64.085 10.035 -63.755 10.365 ;
        RECT -64.085 8.675 -63.755 9.005 ;
        RECT -64.085 7.315 -63.755 7.645 ;
        RECT -64.085 5.955 -63.755 6.285 ;
        RECT -64.085 4.595 -63.755 4.925 ;
        RECT -64.085 3.235 -63.755 3.565 ;
        RECT -64.085 1.875 -63.755 2.205 ;
        RECT -64.085 0.515 -63.755 0.845 ;
        RECT -64.085 -0.845 -63.755 -0.515 ;
        RECT -64.085 -2.205 -63.755 -1.875 ;
        RECT -64.085 -3.565 -63.755 -3.235 ;
        RECT -64.085 -4.925 -63.755 -4.595 ;
        RECT -64.085 -6.285 -63.755 -5.955 ;
        RECT -64.085 -7.645 -63.755 -7.315 ;
        RECT -64.085 -9.005 -63.755 -8.675 ;
        RECT -64.085 -10.365 -63.755 -10.035 ;
        RECT -64.085 -11.725 -63.755 -11.395 ;
        RECT -64.085 -13.085 -63.755 -12.755 ;
        RECT -64.085 -14.445 -63.755 -14.115 ;
        RECT -64.085 -15.805 -63.755 -15.475 ;
        RECT -64.085 -17.165 -63.755 -16.835 ;
        RECT -64.085 -18.525 -63.755 -18.195 ;
        RECT -64.085 -19.885 -63.755 -19.555 ;
        RECT -64.085 -21.245 -63.755 -20.915 ;
        RECT -64.085 -22.605 -63.755 -22.275 ;
        RECT -64.085 -23.965 -63.755 -23.635 ;
        RECT -64.085 -25.325 -63.755 -24.995 ;
        RECT -64.085 -28.045 -63.755 -27.715 ;
        RECT -64.085 -29.405 -63.755 -29.075 ;
        RECT -64.085 -30.765 -63.755 -30.435 ;
        RECT -64.085 -32.125 -63.755 -31.795 ;
        RECT -64.085 -33.485 -63.755 -33.155 ;
        RECT -64.085 -34.845 -63.755 -34.515 ;
        RECT -64.085 -36.205 -63.755 -35.875 ;
        RECT -64.085 -37.565 -63.755 -37.235 ;
        RECT -64.085 -38.925 -63.755 -38.595 ;
        RECT -64.085 -40.285 -63.755 -39.955 ;
        RECT -64.085 -41.645 -63.755 -41.315 ;
        RECT -64.085 -43.005 -63.755 -42.675 ;
        RECT -64.085 -44.365 -63.755 -44.035 ;
        RECT -64.085 -45.725 -63.755 -45.395 ;
        RECT -64.085 -47.085 -63.755 -46.755 ;
        RECT -64.085 -48.445 -63.755 -48.115 ;
        RECT -64.085 -49.805 -63.755 -49.475 ;
        RECT -64.085 -51.165 -63.755 -50.835 ;
        RECT -64.085 -52.525 -63.755 -52.195 ;
        RECT -64.085 -53.885 -63.755 -53.555 ;
        RECT -64.085 -55.245 -63.755 -54.915 ;
        RECT -64.085 -56.605 -63.755 -56.275 ;
        RECT -64.085 -57.965 -63.755 -57.635 ;
        RECT -64.085 -59.325 -63.755 -58.995 ;
        RECT -64.085 -60.685 -63.755 -60.355 ;
        RECT -64.085 -62.045 -63.755 -61.715 ;
        RECT -64.085 -63.405 -63.755 -63.075 ;
        RECT -64.085 -64.765 -63.755 -64.435 ;
        RECT -64.085 -66.125 -63.755 -65.795 ;
        RECT -64.085 -67.485 -63.755 -67.155 ;
        RECT -64.085 -68.845 -63.755 -68.515 ;
        RECT -64.085 -70.205 -63.755 -69.875 ;
        RECT -64.085 -71.565 -63.755 -71.235 ;
        RECT -64.085 -72.925 -63.755 -72.595 ;
        RECT -64.085 -74.285 -63.755 -73.955 ;
        RECT -64.085 -75.645 -63.755 -75.315 ;
        RECT -64.085 -77.005 -63.755 -76.675 ;
        RECT -64.085 -78.365 -63.755 -78.035 ;
        RECT -64.085 -79.725 -63.755 -79.395 ;
        RECT -64.085 -81.085 -63.755 -80.755 ;
        RECT -64.085 -82.445 -63.755 -82.115 ;
        RECT -64.085 -83.805 -63.755 -83.475 ;
        RECT -64.085 -85.165 -63.755 -84.835 ;
        RECT -64.085 -86.525 -63.755 -86.195 ;
        RECT -64.085 -87.885 -63.755 -87.555 ;
        RECT -64.085 -89.245 -63.755 -88.915 ;
        RECT -64.085 -90.605 -63.755 -90.275 ;
        RECT -64.085 -91.77 -63.755 -91.44 ;
        RECT -64.085 -93.325 -63.755 -92.995 ;
        RECT -64.085 -94.685 -63.755 -94.355 ;
        RECT -64.085 -96.045 -63.755 -95.715 ;
        RECT -64.085 -97.405 -63.755 -97.075 ;
        RECT -64.085 -98.765 -63.755 -98.435 ;
        RECT -64.085 -101.485 -63.755 -101.155 ;
        RECT -64.085 -102.31 -63.755 -101.98 ;
        RECT -64.085 -104.205 -63.755 -103.875 ;
        RECT -64.085 -105.565 -63.755 -105.235 ;
        RECT -64.085 -106.925 -63.755 -106.595 ;
        RECT -64.085 -109.645 -63.755 -109.315 ;
        RECT -64.085 -111.005 -63.755 -110.675 ;
        RECT -64.085 -115.085 -63.755 -114.755 ;
        RECT -64.085 -116.445 -63.755 -116.115 ;
        RECT -64.085 -117.805 -63.755 -117.475 ;
        RECT -64.085 -119.165 -63.755 -118.835 ;
        RECT -64.085 -120.525 -63.755 -120.195 ;
        RECT -64.085 -123.245 -63.755 -122.915 ;
        RECT -64.085 -124.605 -63.755 -124.275 ;
        RECT -64.085 -125.965 -63.755 -125.635 ;
        RECT -64.085 -127.325 -63.755 -126.995 ;
        RECT -64.085 -128.685 -63.755 -128.355 ;
        RECT -64.085 -130.045 -63.755 -129.715 ;
        RECT -64.085 -131.405 -63.755 -131.075 ;
        RECT -64.085 -132.765 -63.755 -132.435 ;
        RECT -64.085 -134.125 -63.755 -133.795 ;
        RECT -64.085 -135.485 -63.755 -135.155 ;
        RECT -64.085 -136.845 -63.755 -136.515 ;
        RECT -64.085 -138.205 -63.755 -137.875 ;
        RECT -64.085 -139.565 -63.755 -139.235 ;
        RECT -64.085 -140.925 -63.755 -140.595 ;
        RECT -64.085 -142.285 -63.755 -141.955 ;
        RECT -64.085 -143.645 -63.755 -143.315 ;
        RECT -64.085 -145.005 -63.755 -144.675 ;
        RECT -64.085 -146.365 -63.755 -146.035 ;
        RECT -64.085 -147.725 -63.755 -147.395 ;
        RECT -64.085 -149.085 -63.755 -148.755 ;
        RECT -64.085 -150.445 -63.755 -150.115 ;
        RECT -64.085 -151.805 -63.755 -151.475 ;
        RECT -64.085 -153.165 -63.755 -152.835 ;
        RECT -64.085 -154.525 -63.755 -154.195 ;
        RECT -64.085 -155.885 -63.755 -155.555 ;
        RECT -64.085 -157.245 -63.755 -156.915 ;
        RECT -64.085 -158.605 -63.755 -158.275 ;
        RECT -64.085 -159.965 -63.755 -159.635 ;
        RECT -64.085 -161.325 -63.755 -160.995 ;
        RECT -64.085 -162.685 -63.755 -162.355 ;
        RECT -64.085 -164.045 -63.755 -163.715 ;
        RECT -64.085 -165.405 -63.755 -165.075 ;
        RECT -64.085 -166.765 -63.755 -166.435 ;
        RECT -64.08 -167.44 -63.76 245.285 ;
        RECT -64.085 244.04 -63.755 245.17 ;
        RECT -64.085 239.875 -63.755 240.205 ;
        RECT -64.085 238.515 -63.755 238.845 ;
        RECT -64.085 237.155 -63.755 237.485 ;
        RECT -64.085 235.795 -63.755 236.125 ;
        RECT -64.085 234.435 -63.755 234.765 ;
        RECT -64.085 233.075 -63.755 233.405 ;
        RECT -64.085 231.715 -63.755 232.045 ;
        RECT -64.085 230.355 -63.755 230.685 ;
        RECT -64.085 228.995 -63.755 229.325 ;
        RECT -64.085 227.635 -63.755 227.965 ;
        RECT -64.085 226.275 -63.755 226.605 ;
        RECT -64.085 224.915 -63.755 225.245 ;
        RECT -64.085 223.555 -63.755 223.885 ;
        RECT -64.085 222.195 -63.755 222.525 ;
        RECT -64.085 220.835 -63.755 221.165 ;
        RECT -64.085 219.475 -63.755 219.805 ;
        RECT -64.085 218.115 -63.755 218.445 ;
        RECT -64.085 216.755 -63.755 217.085 ;
        RECT -64.085 215.395 -63.755 215.725 ;
        RECT -64.085 214.035 -63.755 214.365 ;
        RECT -64.085 212.675 -63.755 213.005 ;
        RECT -64.085 211.315 -63.755 211.645 ;
        RECT -64.085 209.955 -63.755 210.285 ;
        RECT -64.085 208.595 -63.755 208.925 ;
        RECT -64.085 207.235 -63.755 207.565 ;
        RECT -64.085 205.875 -63.755 206.205 ;
        RECT -64.085 204.515 -63.755 204.845 ;
        RECT -64.085 203.155 -63.755 203.485 ;
        RECT -64.085 201.795 -63.755 202.125 ;
        RECT -64.085 200.435 -63.755 200.765 ;
        RECT -64.085 199.075 -63.755 199.405 ;
        RECT -64.085 197.715 -63.755 198.045 ;
        RECT -64.085 196.355 -63.755 196.685 ;
        RECT -64.085 194.995 -63.755 195.325 ;
        RECT -64.085 193.635 -63.755 193.965 ;
        RECT -64.085 192.275 -63.755 192.605 ;
        RECT -64.085 190.915 -63.755 191.245 ;
        RECT -64.085 189.555 -63.755 189.885 ;
        RECT -64.085 188.195 -63.755 188.525 ;
        RECT -64.085 186.835 -63.755 187.165 ;
        RECT -64.085 185.475 -63.755 185.805 ;
        RECT -64.085 184.115 -63.755 184.445 ;
        RECT -64.085 182.755 -63.755 183.085 ;
        RECT -64.085 181.395 -63.755 181.725 ;
        RECT -64.085 180.035 -63.755 180.365 ;
        RECT -64.085 178.675 -63.755 179.005 ;
        RECT -64.085 177.315 -63.755 177.645 ;
        RECT -64.085 175.955 -63.755 176.285 ;
        RECT -64.085 174.595 -63.755 174.925 ;
        RECT -64.085 173.235 -63.755 173.565 ;
        RECT -64.085 171.875 -63.755 172.205 ;
        RECT -64.085 170.515 -63.755 170.845 ;
        RECT -64.085 169.155 -63.755 169.485 ;
        RECT -64.085 167.795 -63.755 168.125 ;
        RECT -64.085 166.435 -63.755 166.765 ;
        RECT -64.085 165.075 -63.755 165.405 ;
        RECT -64.085 163.715 -63.755 164.045 ;
        RECT -64.085 162.355 -63.755 162.685 ;
        RECT -64.085 160.995 -63.755 161.325 ;
        RECT -64.085 159.635 -63.755 159.965 ;
        RECT -64.085 158.275 -63.755 158.605 ;
        RECT -64.085 156.915 -63.755 157.245 ;
        RECT -64.085 155.555 -63.755 155.885 ;
        RECT -64.085 154.195 -63.755 154.525 ;
        RECT -64.085 152.835 -63.755 153.165 ;
        RECT -64.085 151.475 -63.755 151.805 ;
        RECT -64.085 150.115 -63.755 150.445 ;
        RECT -64.085 148.755 -63.755 149.085 ;
        RECT -64.085 147.395 -63.755 147.725 ;
        RECT -64.085 146.035 -63.755 146.365 ;
        RECT -64.085 144.675 -63.755 145.005 ;
        RECT -64.085 143.315 -63.755 143.645 ;
        RECT -64.085 141.955 -63.755 142.285 ;
        RECT -64.085 140.595 -63.755 140.925 ;
        RECT -64.085 139.235 -63.755 139.565 ;
        RECT -64.085 136.42 -63.755 136.75 ;
        RECT -64.085 134.245 -63.755 134.575 ;
        RECT -64.085 133.395 -63.755 133.725 ;
        RECT -64.085 131.085 -63.755 131.415 ;
        RECT -64.085 130.235 -63.755 130.565 ;
        RECT -64.085 127.925 -63.755 128.255 ;
        RECT -64.085 127.075 -63.755 127.405 ;
        RECT -64.085 124.765 -63.755 125.095 ;
        RECT -64.085 123.915 -63.755 124.245 ;
        RECT -64.085 121.605 -63.755 121.935 ;
        RECT -64.085 120.755 -63.755 121.085 ;
        RECT -64.085 118.445 -63.755 118.775 ;
        RECT -64.085 117.595 -63.755 117.925 ;
        RECT -64.085 115.285 -63.755 115.615 ;
        RECT -64.085 114.435 -63.755 114.765 ;
        RECT -64.085 112.125 -63.755 112.455 ;
        RECT -64.085 111.275 -63.755 111.605 ;
        RECT -64.085 108.965 -63.755 109.295 ;
        RECT -64.085 108.115 -63.755 108.445 ;
        RECT -64.085 105.805 -63.755 106.135 ;
        RECT -64.085 104.955 -63.755 105.285 ;
        RECT -64.085 102.645 -63.755 102.975 ;
        RECT -64.085 101.795 -63.755 102.125 ;
        RECT -64.085 99.62 -63.755 99.95 ;
    END
    PORT
      LAYER met3 ;
        RECT -73.605 -173.565 -73.275 -173.235 ;
        RECT -73.605 -177.645 -73.275 -177.315 ;
        RECT -73.605 -179.005 -73.275 -178.675 ;
        RECT -73.605 -184.65 -73.275 -183.52 ;
        RECT -73.6 -184.765 -73.28 -173.235 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.245 244.04 -71.915 245.17 ;
        RECT -72.245 239.875 -71.915 240.205 ;
        RECT -72.245 238.515 -71.915 238.845 ;
        RECT -72.245 237.155 -71.915 237.485 ;
        RECT -72.245 235.795 -71.915 236.125 ;
        RECT -72.245 234.435 -71.915 234.765 ;
        RECT -72.245 233.075 -71.915 233.405 ;
        RECT -72.245 231.715 -71.915 232.045 ;
        RECT -72.245 230.355 -71.915 230.685 ;
        RECT -72.245 228.995 -71.915 229.325 ;
        RECT -72.245 227.635 -71.915 227.965 ;
        RECT -72.245 226.275 -71.915 226.605 ;
        RECT -72.245 224.915 -71.915 225.245 ;
        RECT -72.245 223.555 -71.915 223.885 ;
        RECT -72.245 222.195 -71.915 222.525 ;
        RECT -72.245 220.835 -71.915 221.165 ;
        RECT -72.245 219.475 -71.915 219.805 ;
        RECT -72.245 218.115 -71.915 218.445 ;
        RECT -72.245 216.755 -71.915 217.085 ;
        RECT -72.245 215.395 -71.915 215.725 ;
        RECT -72.245 214.035 -71.915 214.365 ;
        RECT -72.245 212.675 -71.915 213.005 ;
        RECT -72.245 211.315 -71.915 211.645 ;
        RECT -72.245 209.955 -71.915 210.285 ;
        RECT -72.245 208.595 -71.915 208.925 ;
        RECT -72.245 207.235 -71.915 207.565 ;
        RECT -72.245 205.875 -71.915 206.205 ;
        RECT -72.245 204.515 -71.915 204.845 ;
        RECT -72.245 203.155 -71.915 203.485 ;
        RECT -72.245 201.795 -71.915 202.125 ;
        RECT -72.245 200.435 -71.915 200.765 ;
        RECT -72.245 199.075 -71.915 199.405 ;
        RECT -72.245 197.715 -71.915 198.045 ;
        RECT -72.245 196.355 -71.915 196.685 ;
        RECT -72.245 194.995 -71.915 195.325 ;
        RECT -72.245 193.635 -71.915 193.965 ;
        RECT -72.245 192.275 -71.915 192.605 ;
        RECT -72.245 190.915 -71.915 191.245 ;
        RECT -72.245 189.555 -71.915 189.885 ;
        RECT -72.245 188.195 -71.915 188.525 ;
        RECT -72.245 186.835 -71.915 187.165 ;
        RECT -72.245 185.475 -71.915 185.805 ;
        RECT -72.245 184.115 -71.915 184.445 ;
        RECT -72.245 182.755 -71.915 183.085 ;
        RECT -72.245 181.395 -71.915 181.725 ;
        RECT -72.245 180.035 -71.915 180.365 ;
        RECT -72.245 178.675 -71.915 179.005 ;
        RECT -72.245 177.315 -71.915 177.645 ;
        RECT -72.245 175.955 -71.915 176.285 ;
        RECT -72.245 174.595 -71.915 174.925 ;
        RECT -72.245 173.235 -71.915 173.565 ;
        RECT -72.245 171.875 -71.915 172.205 ;
        RECT -72.245 170.515 -71.915 170.845 ;
        RECT -72.245 169.155 -71.915 169.485 ;
        RECT -72.245 167.795 -71.915 168.125 ;
        RECT -72.245 166.435 -71.915 166.765 ;
        RECT -72.245 165.075 -71.915 165.405 ;
        RECT -72.245 163.715 -71.915 164.045 ;
        RECT -72.245 162.355 -71.915 162.685 ;
        RECT -72.245 160.995 -71.915 161.325 ;
        RECT -72.245 159.635 -71.915 159.965 ;
        RECT -72.245 158.275 -71.915 158.605 ;
        RECT -72.245 156.915 -71.915 157.245 ;
        RECT -72.245 155.555 -71.915 155.885 ;
        RECT -72.245 154.195 -71.915 154.525 ;
        RECT -72.245 152.835 -71.915 153.165 ;
        RECT -72.245 151.475 -71.915 151.805 ;
        RECT -72.245 150.115 -71.915 150.445 ;
        RECT -72.245 148.755 -71.915 149.085 ;
        RECT -72.245 147.395 -71.915 147.725 ;
        RECT -72.245 146.035 -71.915 146.365 ;
        RECT -72.245 144.675 -71.915 145.005 ;
        RECT -72.245 143.315 -71.915 143.645 ;
        RECT -72.245 141.955 -71.915 142.285 ;
        RECT -72.245 140.595 -71.915 140.925 ;
        RECT -72.245 139.235 -71.915 139.565 ;
        RECT -72.245 137.875 -71.915 138.205 ;
        RECT -72.245 136.515 -71.915 136.845 ;
        RECT -72.245 135.155 -71.915 135.485 ;
        RECT -72.245 133.795 -71.915 134.125 ;
        RECT -72.245 132.435 -71.915 132.765 ;
        RECT -72.245 131.075 -71.915 131.405 ;
        RECT -72.245 129.715 -71.915 130.045 ;
        RECT -72.245 128.355 -71.915 128.685 ;
        RECT -72.245 126.995 -71.915 127.325 ;
        RECT -72.245 125.635 -71.915 125.965 ;
        RECT -72.245 124.275 -71.915 124.605 ;
        RECT -72.245 122.915 -71.915 123.245 ;
        RECT -72.245 121.555 -71.915 121.885 ;
        RECT -72.245 120.195 -71.915 120.525 ;
        RECT -72.245 118.835 -71.915 119.165 ;
        RECT -72.245 117.475 -71.915 117.805 ;
        RECT -72.245 116.115 -71.915 116.445 ;
        RECT -72.245 114.755 -71.915 115.085 ;
        RECT -72.245 113.395 -71.915 113.725 ;
        RECT -72.245 112.035 -71.915 112.365 ;
        RECT -72.245 110.675 -71.915 111.005 ;
        RECT -72.245 109.315 -71.915 109.645 ;
        RECT -72.245 107.955 -71.915 108.285 ;
        RECT -72.245 106.595 -71.915 106.925 ;
        RECT -72.245 105.235 -71.915 105.565 ;
        RECT -72.245 103.875 -71.915 104.205 ;
        RECT -72.245 102.515 -71.915 102.845 ;
        RECT -72.245 101.155 -71.915 101.485 ;
        RECT -72.245 99.795 -71.915 100.125 ;
        RECT -72.245 98.435 -71.915 98.765 ;
        RECT -72.245 97.075 -71.915 97.405 ;
        RECT -72.245 95.715 -71.915 96.045 ;
        RECT -72.245 94.355 -71.915 94.685 ;
        RECT -72.245 92.995 -71.915 93.325 ;
        RECT -72.245 91.635 -71.915 91.965 ;
        RECT -72.245 90.275 -71.915 90.605 ;
        RECT -72.245 88.915 -71.915 89.245 ;
        RECT -72.245 87.555 -71.915 87.885 ;
        RECT -72.245 86.195 -71.915 86.525 ;
        RECT -72.245 84.835 -71.915 85.165 ;
        RECT -72.245 83.475 -71.915 83.805 ;
        RECT -72.245 82.115 -71.915 82.445 ;
        RECT -72.245 80.755 -71.915 81.085 ;
        RECT -72.245 79.395 -71.915 79.725 ;
        RECT -72.245 78.035 -71.915 78.365 ;
        RECT -72.245 76.675 -71.915 77.005 ;
        RECT -72.245 75.315 -71.915 75.645 ;
        RECT -72.245 73.955 -71.915 74.285 ;
        RECT -72.245 72.595 -71.915 72.925 ;
        RECT -72.245 71.235 -71.915 71.565 ;
        RECT -72.245 69.875 -71.915 70.205 ;
        RECT -72.245 68.515 -71.915 68.845 ;
        RECT -72.245 67.155 -71.915 67.485 ;
        RECT -72.245 65.795 -71.915 66.125 ;
        RECT -72.245 64.435 -71.915 64.765 ;
        RECT -72.245 63.075 -71.915 63.405 ;
        RECT -72.245 61.715 -71.915 62.045 ;
        RECT -72.245 60.355 -71.915 60.685 ;
        RECT -72.245 58.995 -71.915 59.325 ;
        RECT -72.245 57.635 -71.915 57.965 ;
        RECT -72.245 56.275 -71.915 56.605 ;
        RECT -72.245 54.915 -71.915 55.245 ;
        RECT -72.245 53.555 -71.915 53.885 ;
        RECT -72.245 52.195 -71.915 52.525 ;
        RECT -72.245 50.835 -71.915 51.165 ;
        RECT -72.245 49.475 -71.915 49.805 ;
        RECT -72.245 48.115 -71.915 48.445 ;
        RECT -72.245 46.755 -71.915 47.085 ;
        RECT -72.245 45.395 -71.915 45.725 ;
        RECT -72.245 44.035 -71.915 44.365 ;
        RECT -72.245 42.675 -71.915 43.005 ;
        RECT -72.245 41.315 -71.915 41.645 ;
        RECT -72.245 39.955 -71.915 40.285 ;
        RECT -72.245 38.595 -71.915 38.925 ;
        RECT -72.245 37.235 -71.915 37.565 ;
        RECT -72.245 35.875 -71.915 36.205 ;
        RECT -72.245 34.515 -71.915 34.845 ;
        RECT -72.245 33.155 -71.915 33.485 ;
        RECT -72.245 31.795 -71.915 32.125 ;
        RECT -72.245 30.435 -71.915 30.765 ;
        RECT -72.245 29.075 -71.915 29.405 ;
        RECT -72.245 27.715 -71.915 28.045 ;
        RECT -72.245 26.355 -71.915 26.685 ;
        RECT -72.245 24.995 -71.915 25.325 ;
        RECT -72.245 23.635 -71.915 23.965 ;
        RECT -72.245 22.275 -71.915 22.605 ;
        RECT -72.245 20.915 -71.915 21.245 ;
        RECT -72.245 19.555 -71.915 19.885 ;
        RECT -72.245 18.195 -71.915 18.525 ;
        RECT -72.245 16.835 -71.915 17.165 ;
        RECT -72.245 15.475 -71.915 15.805 ;
        RECT -72.245 14.115 -71.915 14.445 ;
        RECT -72.245 12.755 -71.915 13.085 ;
        RECT -72.245 11.395 -71.915 11.725 ;
        RECT -72.245 10.035 -71.915 10.365 ;
        RECT -72.245 8.675 -71.915 9.005 ;
        RECT -72.245 7.315 -71.915 7.645 ;
        RECT -72.245 5.955 -71.915 6.285 ;
        RECT -72.245 4.595 -71.915 4.925 ;
        RECT -72.245 3.235 -71.915 3.565 ;
        RECT -72.245 1.875 -71.915 2.205 ;
        RECT -72.245 0.515 -71.915 0.845 ;
        RECT -72.245 -0.845 -71.915 -0.515 ;
        RECT -72.245 -2.205 -71.915 -1.875 ;
        RECT -72.245 -3.565 -71.915 -3.235 ;
        RECT -72.245 -4.925 -71.915 -4.595 ;
        RECT -72.245 -6.285 -71.915 -5.955 ;
        RECT -72.245 -7.645 -71.915 -7.315 ;
        RECT -72.245 -9.005 -71.915 -8.675 ;
        RECT -72.245 -10.365 -71.915 -10.035 ;
        RECT -72.245 -11.725 -71.915 -11.395 ;
        RECT -72.245 -13.085 -71.915 -12.755 ;
        RECT -72.245 -14.445 -71.915 -14.115 ;
        RECT -72.245 -15.805 -71.915 -15.475 ;
        RECT -72.245 -17.165 -71.915 -16.835 ;
        RECT -72.245 -18.525 -71.915 -18.195 ;
        RECT -72.245 -19.885 -71.915 -19.555 ;
        RECT -72.245 -21.245 -71.915 -20.915 ;
        RECT -72.245 -22.605 -71.915 -22.275 ;
        RECT -72.245 -23.965 -71.915 -23.635 ;
        RECT -72.245 -25.325 -71.915 -24.995 ;
        RECT -72.245 -26.685 -71.915 -26.355 ;
        RECT -72.245 -28.045 -71.915 -27.715 ;
        RECT -72.245 -29.405 -71.915 -29.075 ;
        RECT -72.245 -30.765 -71.915 -30.435 ;
        RECT -72.245 -32.125 -71.915 -31.795 ;
        RECT -72.245 -33.485 -71.915 -33.155 ;
        RECT -72.245 -34.845 -71.915 -34.515 ;
        RECT -72.245 -36.205 -71.915 -35.875 ;
        RECT -72.245 -37.565 -71.915 -37.235 ;
        RECT -72.245 -38.925 -71.915 -38.595 ;
        RECT -72.245 -40.285 -71.915 -39.955 ;
        RECT -72.245 -41.645 -71.915 -41.315 ;
        RECT -72.245 -43.005 -71.915 -42.675 ;
        RECT -72.245 -44.365 -71.915 -44.035 ;
        RECT -72.245 -45.725 -71.915 -45.395 ;
        RECT -72.245 -47.085 -71.915 -46.755 ;
        RECT -72.245 -48.445 -71.915 -48.115 ;
        RECT -72.245 -49.805 -71.915 -49.475 ;
        RECT -72.245 -51.165 -71.915 -50.835 ;
        RECT -72.245 -52.525 -71.915 -52.195 ;
        RECT -72.245 -53.885 -71.915 -53.555 ;
        RECT -72.245 -55.245 -71.915 -54.915 ;
        RECT -72.245 -56.605 -71.915 -56.275 ;
        RECT -72.245 -57.965 -71.915 -57.635 ;
        RECT -72.245 -59.325 -71.915 -58.995 ;
        RECT -72.245 -60.685 -71.915 -60.355 ;
        RECT -72.245 -62.045 -71.915 -61.715 ;
        RECT -72.245 -63.405 -71.915 -63.075 ;
        RECT -72.245 -64.765 -71.915 -64.435 ;
        RECT -72.245 -66.125 -71.915 -65.795 ;
        RECT -72.245 -67.485 -71.915 -67.155 ;
        RECT -72.245 -68.845 -71.915 -68.515 ;
        RECT -72.245 -70.205 -71.915 -69.875 ;
        RECT -72.245 -71.565 -71.915 -71.235 ;
        RECT -72.245 -72.925 -71.915 -72.595 ;
        RECT -72.245 -74.285 -71.915 -73.955 ;
        RECT -72.245 -75.645 -71.915 -75.315 ;
        RECT -72.245 -77.005 -71.915 -76.675 ;
        RECT -72.245 -78.365 -71.915 -78.035 ;
        RECT -72.245 -79.725 -71.915 -79.395 ;
        RECT -72.245 -81.085 -71.915 -80.755 ;
        RECT -72.245 -82.445 -71.915 -82.115 ;
        RECT -72.245 -83.805 -71.915 -83.475 ;
        RECT -72.245 -85.165 -71.915 -84.835 ;
        RECT -72.245 -86.525 -71.915 -86.195 ;
        RECT -72.245 -87.885 -71.915 -87.555 ;
        RECT -72.245 -89.245 -71.915 -88.915 ;
        RECT -72.245 -90.605 -71.915 -90.275 ;
        RECT -72.245 -91.965 -71.915 -91.635 ;
        RECT -72.245 -93.325 -71.915 -92.995 ;
        RECT -72.245 -94.685 -71.915 -94.355 ;
        RECT -72.245 -96.045 -71.915 -95.715 ;
        RECT -72.245 -97.405 -71.915 -97.075 ;
        RECT -72.245 -98.765 -71.915 -98.435 ;
        RECT -72.245 -100.125 -71.915 -99.795 ;
        RECT -72.245 -101.485 -71.915 -101.155 ;
        RECT -72.245 -102.845 -71.915 -102.515 ;
        RECT -72.245 -104.205 -71.915 -103.875 ;
        RECT -72.245 -105.565 -71.915 -105.235 ;
        RECT -72.245 -106.925 -71.915 -106.595 ;
        RECT -72.245 -108.285 -71.915 -107.955 ;
        RECT -72.245 -109.645 -71.915 -109.315 ;
        RECT -72.245 -111.005 -71.915 -110.675 ;
        RECT -72.245 -112.365 -71.915 -112.035 ;
        RECT -72.245 -115.085 -71.915 -114.755 ;
        RECT -72.245 -116.445 -71.915 -116.115 ;
        RECT -72.245 -117.805 -71.915 -117.475 ;
        RECT -72.245 -119.165 -71.915 -118.835 ;
        RECT -72.245 -120.525 -71.915 -120.195 ;
        RECT -72.245 -121.885 -71.915 -121.555 ;
        RECT -72.245 -123.245 -71.915 -122.915 ;
        RECT -72.245 -124.605 -71.915 -124.275 ;
        RECT -72.245 -125.965 -71.915 -125.635 ;
        RECT -72.245 -127.325 -71.915 -126.995 ;
        RECT -72.245 -128.685 -71.915 -128.355 ;
        RECT -72.245 -130.045 -71.915 -129.715 ;
        RECT -72.245 -131.405 -71.915 -131.075 ;
        RECT -72.245 -132.765 -71.915 -132.435 ;
        RECT -72.245 -134.125 -71.915 -133.795 ;
        RECT -72.245 -135.485 -71.915 -135.155 ;
        RECT -72.245 -136.845 -71.915 -136.515 ;
        RECT -72.245 -138.205 -71.915 -137.875 ;
        RECT -72.245 -139.565 -71.915 -139.235 ;
        RECT -72.245 -140.925 -71.915 -140.595 ;
        RECT -72.245 -142.285 -71.915 -141.955 ;
        RECT -72.245 -143.645 -71.915 -143.315 ;
        RECT -72.245 -145.005 -71.915 -144.675 ;
        RECT -72.245 -146.365 -71.915 -146.035 ;
        RECT -72.245 -147.725 -71.915 -147.395 ;
        RECT -72.245 -149.085 -71.915 -148.755 ;
        RECT -72.245 -150.445 -71.915 -150.115 ;
        RECT -72.245 -151.805 -71.915 -151.475 ;
        RECT -72.245 -153.165 -71.915 -152.835 ;
        RECT -72.245 -154.525 -71.915 -154.195 ;
        RECT -72.245 -155.885 -71.915 -155.555 ;
        RECT -72.245 -157.245 -71.915 -156.915 ;
        RECT -72.245 -158.605 -71.915 -158.275 ;
        RECT -72.245 -159.965 -71.915 -159.635 ;
        RECT -72.245 -161.325 -71.915 -160.995 ;
        RECT -72.245 -162.685 -71.915 -162.355 ;
        RECT -72.245 -164.045 -71.915 -163.715 ;
        RECT -72.245 -165.405 -71.915 -165.075 ;
        RECT -72.245 -166.765 -71.915 -166.435 ;
        RECT -72.245 -170.845 -71.915 -170.515 ;
        RECT -72.245 -177.645 -71.915 -177.315 ;
        RECT -72.245 -179.005 -71.915 -178.675 ;
        RECT -72.245 -184.65 -71.915 -183.52 ;
        RECT -72.24 -184.765 -71.92 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.885 244.04 -70.555 245.17 ;
        RECT -70.885 239.875 -70.555 240.205 ;
        RECT -70.885 238.515 -70.555 238.845 ;
        RECT -70.885 237.155 -70.555 237.485 ;
        RECT -70.885 235.795 -70.555 236.125 ;
        RECT -70.885 234.435 -70.555 234.765 ;
        RECT -70.885 233.075 -70.555 233.405 ;
        RECT -70.885 231.715 -70.555 232.045 ;
        RECT -70.885 230.355 -70.555 230.685 ;
        RECT -70.885 228.995 -70.555 229.325 ;
        RECT -70.885 227.635 -70.555 227.965 ;
        RECT -70.885 226.275 -70.555 226.605 ;
        RECT -70.885 224.915 -70.555 225.245 ;
        RECT -70.885 223.555 -70.555 223.885 ;
        RECT -70.885 222.195 -70.555 222.525 ;
        RECT -70.885 220.835 -70.555 221.165 ;
        RECT -70.885 219.475 -70.555 219.805 ;
        RECT -70.885 218.115 -70.555 218.445 ;
        RECT -70.885 216.755 -70.555 217.085 ;
        RECT -70.885 215.395 -70.555 215.725 ;
        RECT -70.885 214.035 -70.555 214.365 ;
        RECT -70.885 212.675 -70.555 213.005 ;
        RECT -70.885 211.315 -70.555 211.645 ;
        RECT -70.885 209.955 -70.555 210.285 ;
        RECT -70.885 208.595 -70.555 208.925 ;
        RECT -70.885 207.235 -70.555 207.565 ;
        RECT -70.885 205.875 -70.555 206.205 ;
        RECT -70.885 204.515 -70.555 204.845 ;
        RECT -70.885 203.155 -70.555 203.485 ;
        RECT -70.885 201.795 -70.555 202.125 ;
        RECT -70.885 200.435 -70.555 200.765 ;
        RECT -70.885 199.075 -70.555 199.405 ;
        RECT -70.885 197.715 -70.555 198.045 ;
        RECT -70.885 196.355 -70.555 196.685 ;
        RECT -70.885 194.995 -70.555 195.325 ;
        RECT -70.885 193.635 -70.555 193.965 ;
        RECT -70.885 192.275 -70.555 192.605 ;
        RECT -70.885 190.915 -70.555 191.245 ;
        RECT -70.885 189.555 -70.555 189.885 ;
        RECT -70.885 188.195 -70.555 188.525 ;
        RECT -70.885 186.835 -70.555 187.165 ;
        RECT -70.885 185.475 -70.555 185.805 ;
        RECT -70.885 184.115 -70.555 184.445 ;
        RECT -70.885 182.755 -70.555 183.085 ;
        RECT -70.885 181.395 -70.555 181.725 ;
        RECT -70.885 180.035 -70.555 180.365 ;
        RECT -70.885 178.675 -70.555 179.005 ;
        RECT -70.885 177.315 -70.555 177.645 ;
        RECT -70.885 175.955 -70.555 176.285 ;
        RECT -70.885 174.595 -70.555 174.925 ;
        RECT -70.885 173.235 -70.555 173.565 ;
        RECT -70.885 171.875 -70.555 172.205 ;
        RECT -70.885 170.515 -70.555 170.845 ;
        RECT -70.885 169.155 -70.555 169.485 ;
        RECT -70.885 167.795 -70.555 168.125 ;
        RECT -70.885 166.435 -70.555 166.765 ;
        RECT -70.885 165.075 -70.555 165.405 ;
        RECT -70.885 163.715 -70.555 164.045 ;
        RECT -70.885 162.355 -70.555 162.685 ;
        RECT -70.885 160.995 -70.555 161.325 ;
        RECT -70.885 159.635 -70.555 159.965 ;
        RECT -70.885 158.275 -70.555 158.605 ;
        RECT -70.885 156.915 -70.555 157.245 ;
        RECT -70.885 155.555 -70.555 155.885 ;
        RECT -70.885 154.195 -70.555 154.525 ;
        RECT -70.885 152.835 -70.555 153.165 ;
        RECT -70.885 151.475 -70.555 151.805 ;
        RECT -70.885 150.115 -70.555 150.445 ;
        RECT -70.885 148.755 -70.555 149.085 ;
        RECT -70.885 147.395 -70.555 147.725 ;
        RECT -70.885 146.035 -70.555 146.365 ;
        RECT -70.885 144.675 -70.555 145.005 ;
        RECT -70.885 143.315 -70.555 143.645 ;
        RECT -70.885 141.955 -70.555 142.285 ;
        RECT -70.885 140.595 -70.555 140.925 ;
        RECT -70.885 139.235 -70.555 139.565 ;
        RECT -70.885 137.875 -70.555 138.205 ;
        RECT -70.885 136.515 -70.555 136.845 ;
        RECT -70.885 135.155 -70.555 135.485 ;
        RECT -70.885 133.795 -70.555 134.125 ;
        RECT -70.885 132.435 -70.555 132.765 ;
        RECT -70.885 131.075 -70.555 131.405 ;
        RECT -70.885 129.715 -70.555 130.045 ;
        RECT -70.885 128.355 -70.555 128.685 ;
        RECT -70.885 126.995 -70.555 127.325 ;
        RECT -70.885 125.635 -70.555 125.965 ;
        RECT -70.885 124.275 -70.555 124.605 ;
        RECT -70.885 122.915 -70.555 123.245 ;
        RECT -70.885 121.555 -70.555 121.885 ;
        RECT -70.885 120.195 -70.555 120.525 ;
        RECT -70.885 118.835 -70.555 119.165 ;
        RECT -70.885 117.475 -70.555 117.805 ;
        RECT -70.885 116.115 -70.555 116.445 ;
        RECT -70.885 114.755 -70.555 115.085 ;
        RECT -70.885 113.395 -70.555 113.725 ;
        RECT -70.885 112.035 -70.555 112.365 ;
        RECT -70.885 110.675 -70.555 111.005 ;
        RECT -70.885 109.315 -70.555 109.645 ;
        RECT -70.885 107.955 -70.555 108.285 ;
        RECT -70.885 106.595 -70.555 106.925 ;
        RECT -70.885 105.235 -70.555 105.565 ;
        RECT -70.885 103.875 -70.555 104.205 ;
        RECT -70.885 102.515 -70.555 102.845 ;
        RECT -70.885 101.155 -70.555 101.485 ;
        RECT -70.885 99.795 -70.555 100.125 ;
        RECT -70.885 98.435 -70.555 98.765 ;
        RECT -70.885 97.075 -70.555 97.405 ;
        RECT -70.885 95.715 -70.555 96.045 ;
        RECT -70.885 94.355 -70.555 94.685 ;
        RECT -70.885 92.995 -70.555 93.325 ;
        RECT -70.885 91.635 -70.555 91.965 ;
        RECT -70.885 90.275 -70.555 90.605 ;
        RECT -70.885 88.915 -70.555 89.245 ;
        RECT -70.885 87.555 -70.555 87.885 ;
        RECT -70.885 86.195 -70.555 86.525 ;
        RECT -70.885 84.835 -70.555 85.165 ;
        RECT -70.885 83.475 -70.555 83.805 ;
        RECT -70.885 82.115 -70.555 82.445 ;
        RECT -70.885 80.755 -70.555 81.085 ;
        RECT -70.885 79.395 -70.555 79.725 ;
        RECT -70.885 78.035 -70.555 78.365 ;
        RECT -70.885 76.675 -70.555 77.005 ;
        RECT -70.885 75.315 -70.555 75.645 ;
        RECT -70.885 73.955 -70.555 74.285 ;
        RECT -70.885 72.595 -70.555 72.925 ;
        RECT -70.885 71.235 -70.555 71.565 ;
        RECT -70.885 69.875 -70.555 70.205 ;
        RECT -70.885 68.515 -70.555 68.845 ;
        RECT -70.885 67.155 -70.555 67.485 ;
        RECT -70.885 65.795 -70.555 66.125 ;
        RECT -70.885 64.435 -70.555 64.765 ;
        RECT -70.885 63.075 -70.555 63.405 ;
        RECT -70.885 61.715 -70.555 62.045 ;
        RECT -70.885 60.355 -70.555 60.685 ;
        RECT -70.885 58.995 -70.555 59.325 ;
        RECT -70.885 57.635 -70.555 57.965 ;
        RECT -70.885 56.275 -70.555 56.605 ;
        RECT -70.885 54.915 -70.555 55.245 ;
        RECT -70.885 53.555 -70.555 53.885 ;
        RECT -70.885 52.195 -70.555 52.525 ;
        RECT -70.885 50.835 -70.555 51.165 ;
        RECT -70.885 49.475 -70.555 49.805 ;
        RECT -70.885 48.115 -70.555 48.445 ;
        RECT -70.885 46.755 -70.555 47.085 ;
        RECT -70.885 45.395 -70.555 45.725 ;
        RECT -70.885 44.035 -70.555 44.365 ;
        RECT -70.885 42.675 -70.555 43.005 ;
        RECT -70.885 41.315 -70.555 41.645 ;
        RECT -70.885 39.955 -70.555 40.285 ;
        RECT -70.885 38.595 -70.555 38.925 ;
        RECT -70.885 37.235 -70.555 37.565 ;
        RECT -70.885 35.875 -70.555 36.205 ;
        RECT -70.885 34.515 -70.555 34.845 ;
        RECT -70.885 33.155 -70.555 33.485 ;
        RECT -70.885 31.795 -70.555 32.125 ;
        RECT -70.885 30.435 -70.555 30.765 ;
        RECT -70.885 29.075 -70.555 29.405 ;
        RECT -70.885 27.715 -70.555 28.045 ;
        RECT -70.885 26.355 -70.555 26.685 ;
        RECT -70.885 24.995 -70.555 25.325 ;
        RECT -70.885 23.635 -70.555 23.965 ;
        RECT -70.885 22.275 -70.555 22.605 ;
        RECT -70.885 20.915 -70.555 21.245 ;
        RECT -70.885 19.555 -70.555 19.885 ;
        RECT -70.885 18.195 -70.555 18.525 ;
        RECT -70.885 16.835 -70.555 17.165 ;
        RECT -70.885 15.475 -70.555 15.805 ;
        RECT -70.885 14.115 -70.555 14.445 ;
        RECT -70.885 12.755 -70.555 13.085 ;
        RECT -70.885 11.395 -70.555 11.725 ;
        RECT -70.885 10.035 -70.555 10.365 ;
        RECT -70.885 8.675 -70.555 9.005 ;
        RECT -70.885 7.315 -70.555 7.645 ;
        RECT -70.885 5.955 -70.555 6.285 ;
        RECT -70.885 4.595 -70.555 4.925 ;
        RECT -70.885 3.235 -70.555 3.565 ;
        RECT -70.885 1.875 -70.555 2.205 ;
        RECT -70.885 0.515 -70.555 0.845 ;
        RECT -70.885 -0.845 -70.555 -0.515 ;
        RECT -70.885 -2.205 -70.555 -1.875 ;
        RECT -70.885 -3.565 -70.555 -3.235 ;
        RECT -70.885 -4.925 -70.555 -4.595 ;
        RECT -70.885 -6.285 -70.555 -5.955 ;
        RECT -70.885 -7.645 -70.555 -7.315 ;
        RECT -70.885 -9.005 -70.555 -8.675 ;
        RECT -70.885 -10.365 -70.555 -10.035 ;
        RECT -70.885 -11.725 -70.555 -11.395 ;
        RECT -70.885 -13.085 -70.555 -12.755 ;
        RECT -70.885 -14.445 -70.555 -14.115 ;
        RECT -70.885 -15.805 -70.555 -15.475 ;
        RECT -70.885 -17.165 -70.555 -16.835 ;
        RECT -70.885 -18.525 -70.555 -18.195 ;
        RECT -70.885 -19.885 -70.555 -19.555 ;
        RECT -70.885 -21.245 -70.555 -20.915 ;
        RECT -70.885 -22.605 -70.555 -22.275 ;
        RECT -70.885 -23.965 -70.555 -23.635 ;
        RECT -70.885 -25.325 -70.555 -24.995 ;
        RECT -70.885 -26.685 -70.555 -26.355 ;
        RECT -70.885 -28.045 -70.555 -27.715 ;
        RECT -70.885 -29.405 -70.555 -29.075 ;
        RECT -70.885 -30.765 -70.555 -30.435 ;
        RECT -70.885 -32.125 -70.555 -31.795 ;
        RECT -70.885 -33.485 -70.555 -33.155 ;
        RECT -70.885 -34.845 -70.555 -34.515 ;
        RECT -70.885 -36.205 -70.555 -35.875 ;
        RECT -70.885 -37.565 -70.555 -37.235 ;
        RECT -70.885 -38.925 -70.555 -38.595 ;
        RECT -70.885 -40.285 -70.555 -39.955 ;
        RECT -70.885 -41.645 -70.555 -41.315 ;
        RECT -70.885 -43.005 -70.555 -42.675 ;
        RECT -70.885 -44.365 -70.555 -44.035 ;
        RECT -70.885 -45.725 -70.555 -45.395 ;
        RECT -70.885 -47.085 -70.555 -46.755 ;
        RECT -70.885 -48.445 -70.555 -48.115 ;
        RECT -70.885 -49.805 -70.555 -49.475 ;
        RECT -70.885 -51.165 -70.555 -50.835 ;
        RECT -70.885 -52.525 -70.555 -52.195 ;
        RECT -70.885 -53.885 -70.555 -53.555 ;
        RECT -70.885 -55.245 -70.555 -54.915 ;
        RECT -70.885 -56.605 -70.555 -56.275 ;
        RECT -70.885 -57.965 -70.555 -57.635 ;
        RECT -70.885 -59.325 -70.555 -58.995 ;
        RECT -70.885 -60.685 -70.555 -60.355 ;
        RECT -70.885 -62.045 -70.555 -61.715 ;
        RECT -70.885 -63.405 -70.555 -63.075 ;
        RECT -70.885 -64.765 -70.555 -64.435 ;
        RECT -70.885 -66.125 -70.555 -65.795 ;
        RECT -70.885 -67.485 -70.555 -67.155 ;
        RECT -70.885 -68.845 -70.555 -68.515 ;
        RECT -70.885 -70.205 -70.555 -69.875 ;
        RECT -70.885 -71.565 -70.555 -71.235 ;
        RECT -70.885 -72.925 -70.555 -72.595 ;
        RECT -70.885 -74.285 -70.555 -73.955 ;
        RECT -70.885 -75.645 -70.555 -75.315 ;
        RECT -70.885 -77.005 -70.555 -76.675 ;
        RECT -70.885 -78.365 -70.555 -78.035 ;
        RECT -70.885 -79.725 -70.555 -79.395 ;
        RECT -70.885 -81.085 -70.555 -80.755 ;
        RECT -70.885 -82.445 -70.555 -82.115 ;
        RECT -70.885 -83.805 -70.555 -83.475 ;
        RECT -70.885 -85.165 -70.555 -84.835 ;
        RECT -70.885 -86.525 -70.555 -86.195 ;
        RECT -70.885 -87.885 -70.555 -87.555 ;
        RECT -70.885 -89.245 -70.555 -88.915 ;
        RECT -70.885 -90.605 -70.555 -90.275 ;
        RECT -70.885 -93.325 -70.555 -92.995 ;
        RECT -70.885 -94.685 -70.555 -94.355 ;
        RECT -70.885 -96.045 -70.555 -95.715 ;
        RECT -70.885 -97.405 -70.555 -97.075 ;
        RECT -70.885 -98.765 -70.555 -98.435 ;
        RECT -70.885 -101.485 -70.555 -101.155 ;
        RECT -70.885 -104.205 -70.555 -103.875 ;
        RECT -70.885 -105.565 -70.555 -105.235 ;
        RECT -70.885 -106.925 -70.555 -106.595 ;
        RECT -70.885 -109.645 -70.555 -109.315 ;
        RECT -70.885 -111.005 -70.555 -110.675 ;
        RECT -70.885 -115.085 -70.555 -114.755 ;
        RECT -70.885 -116.445 -70.555 -116.115 ;
        RECT -70.885 -117.805 -70.555 -117.475 ;
        RECT -70.885 -119.165 -70.555 -118.835 ;
        RECT -70.885 -120.525 -70.555 -120.195 ;
        RECT -70.885 -123.245 -70.555 -122.915 ;
        RECT -70.885 -124.605 -70.555 -124.275 ;
        RECT -70.885 -125.965 -70.555 -125.635 ;
        RECT -70.885 -127.325 -70.555 -126.995 ;
        RECT -70.885 -128.685 -70.555 -128.355 ;
        RECT -70.885 -130.045 -70.555 -129.715 ;
        RECT -70.885 -131.405 -70.555 -131.075 ;
        RECT -70.885 -132.765 -70.555 -132.435 ;
        RECT -70.885 -134.125 -70.555 -133.795 ;
        RECT -70.885 -135.485 -70.555 -135.155 ;
        RECT -70.885 -136.845 -70.555 -136.515 ;
        RECT -70.885 -138.205 -70.555 -137.875 ;
        RECT -70.885 -139.565 -70.555 -139.235 ;
        RECT -70.885 -140.925 -70.555 -140.595 ;
        RECT -70.885 -142.285 -70.555 -141.955 ;
        RECT -70.885 -143.645 -70.555 -143.315 ;
        RECT -70.885 -145.005 -70.555 -144.675 ;
        RECT -70.885 -146.365 -70.555 -146.035 ;
        RECT -70.885 -147.725 -70.555 -147.395 ;
        RECT -70.885 -149.085 -70.555 -148.755 ;
        RECT -70.885 -150.445 -70.555 -150.115 ;
        RECT -70.885 -151.805 -70.555 -151.475 ;
        RECT -70.885 -153.165 -70.555 -152.835 ;
        RECT -70.885 -154.525 -70.555 -154.195 ;
        RECT -70.885 -155.885 -70.555 -155.555 ;
        RECT -70.885 -157.245 -70.555 -156.915 ;
        RECT -70.885 -158.605 -70.555 -158.275 ;
        RECT -70.885 -159.965 -70.555 -159.635 ;
        RECT -70.885 -161.325 -70.555 -160.995 ;
        RECT -70.885 -162.685 -70.555 -162.355 ;
        RECT -70.885 -164.045 -70.555 -163.715 ;
        RECT -70.885 -165.405 -70.555 -165.075 ;
        RECT -70.885 -166.765 -70.555 -166.435 ;
        RECT -70.885 -169.615 -70.555 -169.285 ;
        RECT -70.885 -170.845 -70.555 -170.515 ;
        RECT -70.885 -172.205 -70.555 -171.875 ;
        RECT -70.88 -172.88 -70.56 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -69.525 244.04 -69.195 245.17 ;
        RECT -69.525 239.875 -69.195 240.205 ;
        RECT -69.525 238.515 -69.195 238.845 ;
        RECT -69.525 237.155 -69.195 237.485 ;
        RECT -69.525 235.795 -69.195 236.125 ;
        RECT -69.525 234.435 -69.195 234.765 ;
        RECT -69.525 233.075 -69.195 233.405 ;
        RECT -69.525 231.715 -69.195 232.045 ;
        RECT -69.525 230.355 -69.195 230.685 ;
        RECT -69.525 228.995 -69.195 229.325 ;
        RECT -69.525 227.635 -69.195 227.965 ;
        RECT -69.525 226.275 -69.195 226.605 ;
        RECT -69.525 224.915 -69.195 225.245 ;
        RECT -69.525 223.555 -69.195 223.885 ;
        RECT -69.525 222.195 -69.195 222.525 ;
        RECT -69.525 220.835 -69.195 221.165 ;
        RECT -69.525 219.475 -69.195 219.805 ;
        RECT -69.525 218.115 -69.195 218.445 ;
        RECT -69.525 216.755 -69.195 217.085 ;
        RECT -69.525 215.395 -69.195 215.725 ;
        RECT -69.525 214.035 -69.195 214.365 ;
        RECT -69.525 212.675 -69.195 213.005 ;
        RECT -69.525 211.315 -69.195 211.645 ;
        RECT -69.525 209.955 -69.195 210.285 ;
        RECT -69.525 208.595 -69.195 208.925 ;
        RECT -69.525 207.235 -69.195 207.565 ;
        RECT -69.525 205.875 -69.195 206.205 ;
        RECT -69.525 204.515 -69.195 204.845 ;
        RECT -69.525 203.155 -69.195 203.485 ;
        RECT -69.525 201.795 -69.195 202.125 ;
        RECT -69.525 200.435 -69.195 200.765 ;
        RECT -69.525 199.075 -69.195 199.405 ;
        RECT -69.525 197.715 -69.195 198.045 ;
        RECT -69.525 196.355 -69.195 196.685 ;
        RECT -69.525 194.995 -69.195 195.325 ;
        RECT -69.525 193.635 -69.195 193.965 ;
        RECT -69.525 192.275 -69.195 192.605 ;
        RECT -69.525 190.915 -69.195 191.245 ;
        RECT -69.525 189.555 -69.195 189.885 ;
        RECT -69.525 188.195 -69.195 188.525 ;
        RECT -69.525 186.835 -69.195 187.165 ;
        RECT -69.525 185.475 -69.195 185.805 ;
        RECT -69.525 184.115 -69.195 184.445 ;
        RECT -69.525 182.755 -69.195 183.085 ;
        RECT -69.525 181.395 -69.195 181.725 ;
        RECT -69.525 180.035 -69.195 180.365 ;
        RECT -69.525 178.675 -69.195 179.005 ;
        RECT -69.525 177.315 -69.195 177.645 ;
        RECT -69.525 175.955 -69.195 176.285 ;
        RECT -69.525 174.595 -69.195 174.925 ;
        RECT -69.525 173.235 -69.195 173.565 ;
        RECT -69.525 171.875 -69.195 172.205 ;
        RECT -69.525 170.515 -69.195 170.845 ;
        RECT -69.525 169.155 -69.195 169.485 ;
        RECT -69.525 167.795 -69.195 168.125 ;
        RECT -69.525 166.435 -69.195 166.765 ;
        RECT -69.525 165.075 -69.195 165.405 ;
        RECT -69.525 163.715 -69.195 164.045 ;
        RECT -69.525 162.355 -69.195 162.685 ;
        RECT -69.525 160.995 -69.195 161.325 ;
        RECT -69.525 159.635 -69.195 159.965 ;
        RECT -69.525 158.275 -69.195 158.605 ;
        RECT -69.525 156.915 -69.195 157.245 ;
        RECT -69.525 155.555 -69.195 155.885 ;
        RECT -69.525 154.195 -69.195 154.525 ;
        RECT -69.525 152.835 -69.195 153.165 ;
        RECT -69.525 151.475 -69.195 151.805 ;
        RECT -69.525 150.115 -69.195 150.445 ;
        RECT -69.525 148.755 -69.195 149.085 ;
        RECT -69.525 147.395 -69.195 147.725 ;
        RECT -69.525 146.035 -69.195 146.365 ;
        RECT -69.525 144.675 -69.195 145.005 ;
        RECT -69.525 143.315 -69.195 143.645 ;
        RECT -69.525 141.955 -69.195 142.285 ;
        RECT -69.525 140.595 -69.195 140.925 ;
        RECT -69.525 139.235 -69.195 139.565 ;
        RECT -69.525 137.875 -69.195 138.205 ;
        RECT -69.525 136.515 -69.195 136.845 ;
        RECT -69.525 135.155 -69.195 135.485 ;
        RECT -69.525 133.795 -69.195 134.125 ;
        RECT -69.525 132.435 -69.195 132.765 ;
        RECT -69.525 131.075 -69.195 131.405 ;
        RECT -69.525 129.715 -69.195 130.045 ;
        RECT -69.525 128.355 -69.195 128.685 ;
        RECT -69.525 126.995 -69.195 127.325 ;
        RECT -69.525 125.635 -69.195 125.965 ;
        RECT -69.525 124.275 -69.195 124.605 ;
        RECT -69.525 122.915 -69.195 123.245 ;
        RECT -69.525 121.555 -69.195 121.885 ;
        RECT -69.525 120.195 -69.195 120.525 ;
        RECT -69.525 118.835 -69.195 119.165 ;
        RECT -69.525 117.475 -69.195 117.805 ;
        RECT -69.525 116.115 -69.195 116.445 ;
        RECT -69.525 114.755 -69.195 115.085 ;
        RECT -69.525 113.395 -69.195 113.725 ;
        RECT -69.525 112.035 -69.195 112.365 ;
        RECT -69.525 110.675 -69.195 111.005 ;
        RECT -69.525 109.315 -69.195 109.645 ;
        RECT -69.525 107.955 -69.195 108.285 ;
        RECT -69.525 106.595 -69.195 106.925 ;
        RECT -69.525 105.235 -69.195 105.565 ;
        RECT -69.525 103.875 -69.195 104.205 ;
        RECT -69.525 102.515 -69.195 102.845 ;
        RECT -69.525 101.155 -69.195 101.485 ;
        RECT -69.525 99.795 -69.195 100.125 ;
        RECT -69.525 98.435 -69.195 98.765 ;
        RECT -69.525 97.075 -69.195 97.405 ;
        RECT -69.525 95.715 -69.195 96.045 ;
        RECT -69.525 94.355 -69.195 94.685 ;
        RECT -69.525 92.995 -69.195 93.325 ;
        RECT -69.525 91.635 -69.195 91.965 ;
        RECT -69.525 90.275 -69.195 90.605 ;
        RECT -69.525 88.915 -69.195 89.245 ;
        RECT -69.525 87.555 -69.195 87.885 ;
        RECT -69.525 86.195 -69.195 86.525 ;
        RECT -69.525 84.835 -69.195 85.165 ;
        RECT -69.525 83.475 -69.195 83.805 ;
        RECT -69.525 82.115 -69.195 82.445 ;
        RECT -69.525 80.755 -69.195 81.085 ;
        RECT -69.525 79.395 -69.195 79.725 ;
        RECT -69.525 78.035 -69.195 78.365 ;
        RECT -69.525 76.675 -69.195 77.005 ;
        RECT -69.525 75.315 -69.195 75.645 ;
        RECT -69.525 73.955 -69.195 74.285 ;
        RECT -69.525 72.595 -69.195 72.925 ;
        RECT -69.525 71.235 -69.195 71.565 ;
        RECT -69.525 69.875 -69.195 70.205 ;
        RECT -69.525 68.515 -69.195 68.845 ;
        RECT -69.525 67.155 -69.195 67.485 ;
        RECT -69.525 65.795 -69.195 66.125 ;
        RECT -69.525 64.435 -69.195 64.765 ;
        RECT -69.525 63.075 -69.195 63.405 ;
        RECT -69.525 61.715 -69.195 62.045 ;
        RECT -69.525 60.355 -69.195 60.685 ;
        RECT -69.525 58.995 -69.195 59.325 ;
        RECT -69.525 57.635 -69.195 57.965 ;
        RECT -69.525 56.275 -69.195 56.605 ;
        RECT -69.525 54.915 -69.195 55.245 ;
        RECT -69.525 53.555 -69.195 53.885 ;
        RECT -69.525 52.195 -69.195 52.525 ;
        RECT -69.525 50.835 -69.195 51.165 ;
        RECT -69.525 49.475 -69.195 49.805 ;
        RECT -69.525 48.115 -69.195 48.445 ;
        RECT -69.525 46.755 -69.195 47.085 ;
        RECT -69.525 45.395 -69.195 45.725 ;
        RECT -69.525 44.035 -69.195 44.365 ;
        RECT -69.525 42.675 -69.195 43.005 ;
        RECT -69.525 41.315 -69.195 41.645 ;
        RECT -69.525 39.955 -69.195 40.285 ;
        RECT -69.525 38.595 -69.195 38.925 ;
        RECT -69.525 37.235 -69.195 37.565 ;
        RECT -69.525 35.875 -69.195 36.205 ;
        RECT -69.525 34.515 -69.195 34.845 ;
        RECT -69.525 33.155 -69.195 33.485 ;
        RECT -69.525 31.795 -69.195 32.125 ;
        RECT -69.525 30.435 -69.195 30.765 ;
        RECT -69.525 29.075 -69.195 29.405 ;
        RECT -69.525 27.715 -69.195 28.045 ;
        RECT -69.525 26.355 -69.195 26.685 ;
        RECT -69.525 24.995 -69.195 25.325 ;
        RECT -69.525 23.635 -69.195 23.965 ;
        RECT -69.525 22.275 -69.195 22.605 ;
        RECT -69.525 20.915 -69.195 21.245 ;
        RECT -69.525 19.555 -69.195 19.885 ;
        RECT -69.525 18.195 -69.195 18.525 ;
        RECT -69.525 16.835 -69.195 17.165 ;
        RECT -69.525 15.475 -69.195 15.805 ;
        RECT -69.525 14.115 -69.195 14.445 ;
        RECT -69.525 12.755 -69.195 13.085 ;
        RECT -69.525 11.395 -69.195 11.725 ;
        RECT -69.525 10.035 -69.195 10.365 ;
        RECT -69.525 8.675 -69.195 9.005 ;
        RECT -69.525 7.315 -69.195 7.645 ;
        RECT -69.525 5.955 -69.195 6.285 ;
        RECT -69.525 4.595 -69.195 4.925 ;
        RECT -69.525 3.235 -69.195 3.565 ;
        RECT -69.525 1.875 -69.195 2.205 ;
        RECT -69.525 0.515 -69.195 0.845 ;
        RECT -69.525 -0.845 -69.195 -0.515 ;
        RECT -69.525 -2.205 -69.195 -1.875 ;
        RECT -69.525 -3.565 -69.195 -3.235 ;
        RECT -69.525 -4.925 -69.195 -4.595 ;
        RECT -69.525 -6.285 -69.195 -5.955 ;
        RECT -69.525 -7.645 -69.195 -7.315 ;
        RECT -69.525 -9.005 -69.195 -8.675 ;
        RECT -69.525 -10.365 -69.195 -10.035 ;
        RECT -69.525 -11.725 -69.195 -11.395 ;
        RECT -69.525 -13.085 -69.195 -12.755 ;
        RECT -69.525 -14.445 -69.195 -14.115 ;
        RECT -69.525 -15.805 -69.195 -15.475 ;
        RECT -69.525 -17.165 -69.195 -16.835 ;
        RECT -69.525 -18.525 -69.195 -18.195 ;
        RECT -69.525 -19.885 -69.195 -19.555 ;
        RECT -69.525 -21.245 -69.195 -20.915 ;
        RECT -69.525 -22.605 -69.195 -22.275 ;
        RECT -69.525 -23.965 -69.195 -23.635 ;
        RECT -69.525 -25.325 -69.195 -24.995 ;
        RECT -69.525 -26.685 -69.195 -26.355 ;
        RECT -69.525 -28.045 -69.195 -27.715 ;
        RECT -69.525 -29.405 -69.195 -29.075 ;
        RECT -69.525 -30.765 -69.195 -30.435 ;
        RECT -69.525 -32.125 -69.195 -31.795 ;
        RECT -69.525 -33.485 -69.195 -33.155 ;
        RECT -69.525 -34.845 -69.195 -34.515 ;
        RECT -69.525 -36.205 -69.195 -35.875 ;
        RECT -69.525 -37.565 -69.195 -37.235 ;
        RECT -69.525 -38.925 -69.195 -38.595 ;
        RECT -69.525 -40.285 -69.195 -39.955 ;
        RECT -69.525 -41.645 -69.195 -41.315 ;
        RECT -69.525 -43.005 -69.195 -42.675 ;
        RECT -69.525 -44.365 -69.195 -44.035 ;
        RECT -69.525 -45.725 -69.195 -45.395 ;
        RECT -69.525 -47.085 -69.195 -46.755 ;
        RECT -69.525 -48.445 -69.195 -48.115 ;
        RECT -69.525 -49.805 -69.195 -49.475 ;
        RECT -69.525 -51.165 -69.195 -50.835 ;
        RECT -69.525 -52.525 -69.195 -52.195 ;
        RECT -69.525 -53.885 -69.195 -53.555 ;
        RECT -69.525 -55.245 -69.195 -54.915 ;
        RECT -69.525 -56.605 -69.195 -56.275 ;
        RECT -69.525 -57.965 -69.195 -57.635 ;
        RECT -69.525 -59.325 -69.195 -58.995 ;
        RECT -69.525 -60.685 -69.195 -60.355 ;
        RECT -69.525 -62.045 -69.195 -61.715 ;
        RECT -69.525 -63.405 -69.195 -63.075 ;
        RECT -69.525 -64.765 -69.195 -64.435 ;
        RECT -69.525 -66.125 -69.195 -65.795 ;
        RECT -69.525 -67.485 -69.195 -67.155 ;
        RECT -69.525 -68.845 -69.195 -68.515 ;
        RECT -69.525 -70.205 -69.195 -69.875 ;
        RECT -69.525 -71.565 -69.195 -71.235 ;
        RECT -69.525 -72.925 -69.195 -72.595 ;
        RECT -69.525 -74.285 -69.195 -73.955 ;
        RECT -69.525 -75.645 -69.195 -75.315 ;
        RECT -69.525 -77.005 -69.195 -76.675 ;
        RECT -69.525 -78.365 -69.195 -78.035 ;
        RECT -69.525 -79.725 -69.195 -79.395 ;
        RECT -69.525 -81.085 -69.195 -80.755 ;
        RECT -69.525 -82.445 -69.195 -82.115 ;
        RECT -69.525 -83.805 -69.195 -83.475 ;
        RECT -69.525 -85.165 -69.195 -84.835 ;
        RECT -69.525 -86.525 -69.195 -86.195 ;
        RECT -69.525 -87.885 -69.195 -87.555 ;
        RECT -69.525 -89.245 -69.195 -88.915 ;
        RECT -69.525 -90.605 -69.195 -90.275 ;
        RECT -69.525 -91.77 -69.195 -91.44 ;
        RECT -69.525 -93.325 -69.195 -92.995 ;
        RECT -69.525 -94.685 -69.195 -94.355 ;
        RECT -69.525 -96.045 -69.195 -95.715 ;
        RECT -69.525 -97.405 -69.195 -97.075 ;
        RECT -69.525 -98.765 -69.195 -98.435 ;
        RECT -69.525 -101.485 -69.195 -101.155 ;
        RECT -69.525 -102.31 -69.195 -101.98 ;
        RECT -69.525 -104.205 -69.195 -103.875 ;
        RECT -69.525 -105.565 -69.195 -105.235 ;
        RECT -69.525 -106.925 -69.195 -106.595 ;
        RECT -69.525 -109.645 -69.195 -109.315 ;
        RECT -69.525 -111.005 -69.195 -110.675 ;
        RECT -69.525 -115.085 -69.195 -114.755 ;
        RECT -69.525 -116.445 -69.195 -116.115 ;
        RECT -69.525 -117.805 -69.195 -117.475 ;
        RECT -69.525 -119.165 -69.195 -118.835 ;
        RECT -69.525 -120.525 -69.195 -120.195 ;
        RECT -69.525 -123.245 -69.195 -122.915 ;
        RECT -69.525 -124.605 -69.195 -124.275 ;
        RECT -69.525 -125.965 -69.195 -125.635 ;
        RECT -69.525 -127.325 -69.195 -126.995 ;
        RECT -69.525 -128.685 -69.195 -128.355 ;
        RECT -69.525 -130.045 -69.195 -129.715 ;
        RECT -69.525 -131.405 -69.195 -131.075 ;
        RECT -69.525 -132.765 -69.195 -132.435 ;
        RECT -69.525 -134.125 -69.195 -133.795 ;
        RECT -69.525 -135.485 -69.195 -135.155 ;
        RECT -69.525 -136.845 -69.195 -136.515 ;
        RECT -69.525 -138.205 -69.195 -137.875 ;
        RECT -69.525 -139.565 -69.195 -139.235 ;
        RECT -69.525 -140.925 -69.195 -140.595 ;
        RECT -69.525 -142.285 -69.195 -141.955 ;
        RECT -69.525 -143.645 -69.195 -143.315 ;
        RECT -69.525 -145.005 -69.195 -144.675 ;
        RECT -69.525 -146.365 -69.195 -146.035 ;
        RECT -69.525 -147.725 -69.195 -147.395 ;
        RECT -69.525 -149.085 -69.195 -148.755 ;
        RECT -69.525 -150.445 -69.195 -150.115 ;
        RECT -69.525 -151.805 -69.195 -151.475 ;
        RECT -69.525 -153.165 -69.195 -152.835 ;
        RECT -69.525 -154.525 -69.195 -154.195 ;
        RECT -69.525 -155.885 -69.195 -155.555 ;
        RECT -69.525 -157.245 -69.195 -156.915 ;
        RECT -69.525 -158.605 -69.195 -158.275 ;
        RECT -69.525 -159.965 -69.195 -159.635 ;
        RECT -69.525 -161.325 -69.195 -160.995 ;
        RECT -69.525 -162.685 -69.195 -162.355 ;
        RECT -69.525 -164.045 -69.195 -163.715 ;
        RECT -69.525 -165.405 -69.195 -165.075 ;
        RECT -69.525 -166.765 -69.195 -166.435 ;
        RECT -69.525 -169.615 -69.195 -169.285 ;
        RECT -69.525 -170.845 -69.195 -170.515 ;
        RECT -69.525 -172.205 -69.195 -171.875 ;
        RECT -69.525 -177.645 -69.195 -177.315 ;
        RECT -69.525 -179.005 -69.195 -178.675 ;
        RECT -69.525 -184.65 -69.195 -183.52 ;
        RECT -69.52 -184.765 -69.2 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.165 -30.765 -67.835 -30.435 ;
        RECT -68.165 -32.125 -67.835 -31.795 ;
        RECT -68.165 -33.485 -67.835 -33.155 ;
        RECT -68.165 -34.845 -67.835 -34.515 ;
        RECT -68.165 -36.205 -67.835 -35.875 ;
        RECT -68.165 -37.565 -67.835 -37.235 ;
        RECT -68.165 -38.925 -67.835 -38.595 ;
        RECT -68.165 -40.285 -67.835 -39.955 ;
        RECT -68.165 -41.645 -67.835 -41.315 ;
        RECT -68.165 -43.005 -67.835 -42.675 ;
        RECT -68.165 -44.365 -67.835 -44.035 ;
        RECT -68.165 -45.725 -67.835 -45.395 ;
        RECT -68.165 -47.085 -67.835 -46.755 ;
        RECT -68.165 -48.445 -67.835 -48.115 ;
        RECT -68.165 -49.805 -67.835 -49.475 ;
        RECT -68.165 -51.165 -67.835 -50.835 ;
        RECT -68.165 -52.525 -67.835 -52.195 ;
        RECT -68.165 -53.885 -67.835 -53.555 ;
        RECT -68.165 -55.245 -67.835 -54.915 ;
        RECT -68.165 -56.605 -67.835 -56.275 ;
        RECT -68.165 -57.965 -67.835 -57.635 ;
        RECT -68.165 -59.325 -67.835 -58.995 ;
        RECT -68.165 -60.685 -67.835 -60.355 ;
        RECT -68.165 -62.045 -67.835 -61.715 ;
        RECT -68.165 -63.405 -67.835 -63.075 ;
        RECT -68.165 -64.765 -67.835 -64.435 ;
        RECT -68.165 -66.125 -67.835 -65.795 ;
        RECT -68.165 -67.485 -67.835 -67.155 ;
        RECT -68.165 -68.845 -67.835 -68.515 ;
        RECT -68.165 -70.205 -67.835 -69.875 ;
        RECT -68.165 -71.565 -67.835 -71.235 ;
        RECT -68.165 -72.925 -67.835 -72.595 ;
        RECT -68.165 -74.285 -67.835 -73.955 ;
        RECT -68.165 -75.645 -67.835 -75.315 ;
        RECT -68.165 -77.005 -67.835 -76.675 ;
        RECT -68.165 -78.365 -67.835 -78.035 ;
        RECT -68.165 -79.725 -67.835 -79.395 ;
        RECT -68.165 -81.085 -67.835 -80.755 ;
        RECT -68.165 -82.445 -67.835 -82.115 ;
        RECT -68.165 -83.805 -67.835 -83.475 ;
        RECT -68.165 -85.165 -67.835 -84.835 ;
        RECT -68.165 -86.525 -67.835 -86.195 ;
        RECT -68.165 -87.885 -67.835 -87.555 ;
        RECT -68.165 -89.245 -67.835 -88.915 ;
        RECT -68.165 -90.605 -67.835 -90.275 ;
        RECT -68.165 -91.77 -67.835 -91.44 ;
        RECT -68.165 -93.325 -67.835 -92.995 ;
        RECT -68.165 -94.685 -67.835 -94.355 ;
        RECT -68.165 -96.045 -67.835 -95.715 ;
        RECT -68.165 -97.405 -67.835 -97.075 ;
        RECT -68.165 -98.765 -67.835 -98.435 ;
        RECT -68.165 -101.485 -67.835 -101.155 ;
        RECT -68.165 -102.31 -67.835 -101.98 ;
        RECT -68.165 -104.205 -67.835 -103.875 ;
        RECT -68.165 -105.565 -67.835 -105.235 ;
        RECT -68.165 -106.925 -67.835 -106.595 ;
        RECT -68.165 -109.645 -67.835 -109.315 ;
        RECT -68.165 -111.005 -67.835 -110.675 ;
        RECT -68.16 -113.72 -67.84 245.285 ;
        RECT -68.165 244.04 -67.835 245.17 ;
        RECT -68.165 239.875 -67.835 240.205 ;
        RECT -68.165 238.515 -67.835 238.845 ;
        RECT -68.165 237.155 -67.835 237.485 ;
        RECT -68.165 235.795 -67.835 236.125 ;
        RECT -68.165 234.435 -67.835 234.765 ;
        RECT -68.165 233.075 -67.835 233.405 ;
        RECT -68.165 231.715 -67.835 232.045 ;
        RECT -68.165 230.355 -67.835 230.685 ;
        RECT -68.165 228.995 -67.835 229.325 ;
        RECT -68.165 227.635 -67.835 227.965 ;
        RECT -68.165 226.275 -67.835 226.605 ;
        RECT -68.165 224.915 -67.835 225.245 ;
        RECT -68.165 223.555 -67.835 223.885 ;
        RECT -68.165 222.195 -67.835 222.525 ;
        RECT -68.165 220.835 -67.835 221.165 ;
        RECT -68.165 219.475 -67.835 219.805 ;
        RECT -68.165 218.115 -67.835 218.445 ;
        RECT -68.165 216.755 -67.835 217.085 ;
        RECT -68.165 215.395 -67.835 215.725 ;
        RECT -68.165 214.035 -67.835 214.365 ;
        RECT -68.165 212.675 -67.835 213.005 ;
        RECT -68.165 211.315 -67.835 211.645 ;
        RECT -68.165 209.955 -67.835 210.285 ;
        RECT -68.165 208.595 -67.835 208.925 ;
        RECT -68.165 207.235 -67.835 207.565 ;
        RECT -68.165 205.875 -67.835 206.205 ;
        RECT -68.165 204.515 -67.835 204.845 ;
        RECT -68.165 203.155 -67.835 203.485 ;
        RECT -68.165 201.795 -67.835 202.125 ;
        RECT -68.165 200.435 -67.835 200.765 ;
        RECT -68.165 199.075 -67.835 199.405 ;
        RECT -68.165 197.715 -67.835 198.045 ;
        RECT -68.165 196.355 -67.835 196.685 ;
        RECT -68.165 194.995 -67.835 195.325 ;
        RECT -68.165 193.635 -67.835 193.965 ;
        RECT -68.165 192.275 -67.835 192.605 ;
        RECT -68.165 190.915 -67.835 191.245 ;
        RECT -68.165 189.555 -67.835 189.885 ;
        RECT -68.165 188.195 -67.835 188.525 ;
        RECT -68.165 186.835 -67.835 187.165 ;
        RECT -68.165 185.475 -67.835 185.805 ;
        RECT -68.165 184.115 -67.835 184.445 ;
        RECT -68.165 182.755 -67.835 183.085 ;
        RECT -68.165 181.395 -67.835 181.725 ;
        RECT -68.165 180.035 -67.835 180.365 ;
        RECT -68.165 178.675 -67.835 179.005 ;
        RECT -68.165 177.315 -67.835 177.645 ;
        RECT -68.165 175.955 -67.835 176.285 ;
        RECT -68.165 174.595 -67.835 174.925 ;
        RECT -68.165 173.235 -67.835 173.565 ;
        RECT -68.165 171.875 -67.835 172.205 ;
        RECT -68.165 170.515 -67.835 170.845 ;
        RECT -68.165 169.155 -67.835 169.485 ;
        RECT -68.165 167.795 -67.835 168.125 ;
        RECT -68.165 166.435 -67.835 166.765 ;
        RECT -68.165 165.075 -67.835 165.405 ;
        RECT -68.165 163.715 -67.835 164.045 ;
        RECT -68.165 162.355 -67.835 162.685 ;
        RECT -68.165 160.995 -67.835 161.325 ;
        RECT -68.165 159.635 -67.835 159.965 ;
        RECT -68.165 158.275 -67.835 158.605 ;
        RECT -68.165 156.915 -67.835 157.245 ;
        RECT -68.165 155.555 -67.835 155.885 ;
        RECT -68.165 154.195 -67.835 154.525 ;
        RECT -68.165 152.835 -67.835 153.165 ;
        RECT -68.165 151.475 -67.835 151.805 ;
        RECT -68.165 150.115 -67.835 150.445 ;
        RECT -68.165 148.755 -67.835 149.085 ;
        RECT -68.165 147.395 -67.835 147.725 ;
        RECT -68.165 146.035 -67.835 146.365 ;
        RECT -68.165 144.675 -67.835 145.005 ;
        RECT -68.165 143.315 -67.835 143.645 ;
        RECT -68.165 141.955 -67.835 142.285 ;
        RECT -68.165 140.595 -67.835 140.925 ;
        RECT -68.165 139.235 -67.835 139.565 ;
        RECT -68.165 137.875 -67.835 138.205 ;
        RECT -68.165 136.515 -67.835 136.845 ;
        RECT -68.165 135.155 -67.835 135.485 ;
        RECT -68.165 133.795 -67.835 134.125 ;
        RECT -68.165 132.435 -67.835 132.765 ;
        RECT -68.165 131.075 -67.835 131.405 ;
        RECT -68.165 129.715 -67.835 130.045 ;
        RECT -68.165 128.355 -67.835 128.685 ;
        RECT -68.165 126.995 -67.835 127.325 ;
        RECT -68.165 125.635 -67.835 125.965 ;
        RECT -68.165 124.275 -67.835 124.605 ;
        RECT -68.165 122.915 -67.835 123.245 ;
        RECT -68.165 121.555 -67.835 121.885 ;
        RECT -68.165 120.195 -67.835 120.525 ;
        RECT -68.165 118.835 -67.835 119.165 ;
        RECT -68.165 117.475 -67.835 117.805 ;
        RECT -68.165 116.115 -67.835 116.445 ;
        RECT -68.165 114.755 -67.835 115.085 ;
        RECT -68.165 113.395 -67.835 113.725 ;
        RECT -68.165 112.035 -67.835 112.365 ;
        RECT -68.165 110.675 -67.835 111.005 ;
        RECT -68.165 109.315 -67.835 109.645 ;
        RECT -68.165 107.955 -67.835 108.285 ;
        RECT -68.165 106.595 -67.835 106.925 ;
        RECT -68.165 105.235 -67.835 105.565 ;
        RECT -68.165 103.875 -67.835 104.205 ;
        RECT -68.165 102.515 -67.835 102.845 ;
        RECT -68.165 101.155 -67.835 101.485 ;
        RECT -68.165 99.795 -67.835 100.125 ;
        RECT -68.165 98.435 -67.835 98.765 ;
        RECT -68.165 97.075 -67.835 97.405 ;
        RECT -68.165 95.715 -67.835 96.045 ;
        RECT -68.165 94.355 -67.835 94.685 ;
        RECT -68.165 92.995 -67.835 93.325 ;
        RECT -68.165 91.635 -67.835 91.965 ;
        RECT -68.165 90.275 -67.835 90.605 ;
        RECT -68.165 88.915 -67.835 89.245 ;
        RECT -68.165 87.555 -67.835 87.885 ;
        RECT -68.165 86.195 -67.835 86.525 ;
        RECT -68.165 84.835 -67.835 85.165 ;
        RECT -68.165 83.475 -67.835 83.805 ;
        RECT -68.165 82.115 -67.835 82.445 ;
        RECT -68.165 80.755 -67.835 81.085 ;
        RECT -68.165 79.395 -67.835 79.725 ;
        RECT -68.165 78.035 -67.835 78.365 ;
        RECT -68.165 76.675 -67.835 77.005 ;
        RECT -68.165 75.315 -67.835 75.645 ;
        RECT -68.165 73.955 -67.835 74.285 ;
        RECT -68.165 72.595 -67.835 72.925 ;
        RECT -68.165 71.235 -67.835 71.565 ;
        RECT -68.165 69.875 -67.835 70.205 ;
        RECT -68.165 68.515 -67.835 68.845 ;
        RECT -68.165 67.155 -67.835 67.485 ;
        RECT -68.165 65.795 -67.835 66.125 ;
        RECT -68.165 64.435 -67.835 64.765 ;
        RECT -68.165 63.075 -67.835 63.405 ;
        RECT -68.165 61.715 -67.835 62.045 ;
        RECT -68.165 60.355 -67.835 60.685 ;
        RECT -68.165 58.995 -67.835 59.325 ;
        RECT -68.165 57.635 -67.835 57.965 ;
        RECT -68.165 56.275 -67.835 56.605 ;
        RECT -68.165 54.915 -67.835 55.245 ;
        RECT -68.165 53.555 -67.835 53.885 ;
        RECT -68.165 52.195 -67.835 52.525 ;
        RECT -68.165 50.835 -67.835 51.165 ;
        RECT -68.165 49.475 -67.835 49.805 ;
        RECT -68.165 48.115 -67.835 48.445 ;
        RECT -68.165 46.755 -67.835 47.085 ;
        RECT -68.165 45.395 -67.835 45.725 ;
        RECT -68.165 44.035 -67.835 44.365 ;
        RECT -68.165 42.675 -67.835 43.005 ;
        RECT -68.165 41.315 -67.835 41.645 ;
        RECT -68.165 39.955 -67.835 40.285 ;
        RECT -68.165 38.595 -67.835 38.925 ;
        RECT -68.165 37.235 -67.835 37.565 ;
        RECT -68.165 35.875 -67.835 36.205 ;
        RECT -68.165 34.515 -67.835 34.845 ;
        RECT -68.165 33.155 -67.835 33.485 ;
        RECT -68.165 31.795 -67.835 32.125 ;
        RECT -68.165 30.435 -67.835 30.765 ;
        RECT -68.165 29.075 -67.835 29.405 ;
        RECT -68.165 27.715 -67.835 28.045 ;
        RECT -68.165 26.355 -67.835 26.685 ;
        RECT -68.165 24.995 -67.835 25.325 ;
        RECT -68.165 23.635 -67.835 23.965 ;
        RECT -68.165 22.275 -67.835 22.605 ;
        RECT -68.165 20.915 -67.835 21.245 ;
        RECT -68.165 19.555 -67.835 19.885 ;
        RECT -68.165 18.195 -67.835 18.525 ;
        RECT -68.165 16.835 -67.835 17.165 ;
        RECT -68.165 15.475 -67.835 15.805 ;
        RECT -68.165 14.115 -67.835 14.445 ;
        RECT -68.165 12.755 -67.835 13.085 ;
        RECT -68.165 11.395 -67.835 11.725 ;
        RECT -68.165 10.035 -67.835 10.365 ;
        RECT -68.165 8.675 -67.835 9.005 ;
        RECT -68.165 7.315 -67.835 7.645 ;
        RECT -68.165 5.955 -67.835 6.285 ;
        RECT -68.165 4.595 -67.835 4.925 ;
        RECT -68.165 3.235 -67.835 3.565 ;
        RECT -68.165 1.875 -67.835 2.205 ;
        RECT -68.165 0.515 -67.835 0.845 ;
        RECT -68.165 -0.845 -67.835 -0.515 ;
        RECT -68.165 -2.205 -67.835 -1.875 ;
        RECT -68.165 -3.565 -67.835 -3.235 ;
        RECT -68.165 -4.925 -67.835 -4.595 ;
        RECT -68.165 -6.285 -67.835 -5.955 ;
        RECT -68.165 -7.645 -67.835 -7.315 ;
        RECT -68.165 -9.005 -67.835 -8.675 ;
        RECT -68.165 -10.365 -67.835 -10.035 ;
        RECT -68.165 -11.725 -67.835 -11.395 ;
        RECT -68.165 -13.085 -67.835 -12.755 ;
        RECT -68.165 -14.445 -67.835 -14.115 ;
        RECT -68.165 -15.805 -67.835 -15.475 ;
        RECT -68.165 -17.165 -67.835 -16.835 ;
        RECT -68.165 -18.525 -67.835 -18.195 ;
        RECT -68.165 -19.885 -67.835 -19.555 ;
        RECT -68.165 -21.245 -67.835 -20.915 ;
        RECT -68.165 -22.605 -67.835 -22.275 ;
        RECT -68.165 -23.965 -67.835 -23.635 ;
        RECT -68.165 -25.325 -67.835 -24.995 ;
        RECT -68.165 -26.685 -67.835 -26.355 ;
        RECT -68.165 -28.045 -67.835 -27.715 ;
        RECT -68.165 -29.405 -67.835 -29.075 ;
    END
    PORT
      LAYER met3 ;
        RECT -76.325 244.04 -75.995 245.17 ;
        RECT -76.325 239.875 -75.995 240.205 ;
        RECT -76.325 238.515 -75.995 238.845 ;
        RECT -76.325 237.155 -75.995 237.485 ;
        RECT -76.325 235.795 -75.995 236.125 ;
        RECT -76.325 234.435 -75.995 234.765 ;
        RECT -76.325 233.075 -75.995 233.405 ;
        RECT -76.325 231.715 -75.995 232.045 ;
        RECT -76.325 230.355 -75.995 230.685 ;
        RECT -76.325 228.995 -75.995 229.325 ;
        RECT -76.325 227.635 -75.995 227.965 ;
        RECT -76.325 226.275 -75.995 226.605 ;
        RECT -76.325 224.915 -75.995 225.245 ;
        RECT -76.325 223.555 -75.995 223.885 ;
        RECT -76.325 222.195 -75.995 222.525 ;
        RECT -76.325 220.835 -75.995 221.165 ;
        RECT -76.325 219.475 -75.995 219.805 ;
        RECT -76.325 218.115 -75.995 218.445 ;
        RECT -76.325 216.755 -75.995 217.085 ;
        RECT -76.325 215.395 -75.995 215.725 ;
        RECT -76.325 214.035 -75.995 214.365 ;
        RECT -76.325 212.675 -75.995 213.005 ;
        RECT -76.325 211.315 -75.995 211.645 ;
        RECT -76.325 209.955 -75.995 210.285 ;
        RECT -76.325 208.595 -75.995 208.925 ;
        RECT -76.325 207.235 -75.995 207.565 ;
        RECT -76.325 205.875 -75.995 206.205 ;
        RECT -76.325 204.515 -75.995 204.845 ;
        RECT -76.325 203.155 -75.995 203.485 ;
        RECT -76.325 201.795 -75.995 202.125 ;
        RECT -76.325 200.435 -75.995 200.765 ;
        RECT -76.325 199.075 -75.995 199.405 ;
        RECT -76.325 197.715 -75.995 198.045 ;
        RECT -76.325 196.355 -75.995 196.685 ;
        RECT -76.325 194.995 -75.995 195.325 ;
        RECT -76.325 193.635 -75.995 193.965 ;
        RECT -76.325 192.275 -75.995 192.605 ;
        RECT -76.325 190.915 -75.995 191.245 ;
        RECT -76.325 189.555 -75.995 189.885 ;
        RECT -76.325 188.195 -75.995 188.525 ;
        RECT -76.325 186.835 -75.995 187.165 ;
        RECT -76.325 185.475 -75.995 185.805 ;
        RECT -76.325 184.115 -75.995 184.445 ;
        RECT -76.325 182.755 -75.995 183.085 ;
        RECT -76.325 181.395 -75.995 181.725 ;
        RECT -76.325 180.035 -75.995 180.365 ;
        RECT -76.325 178.675 -75.995 179.005 ;
        RECT -76.325 177.315 -75.995 177.645 ;
        RECT -76.325 175.955 -75.995 176.285 ;
        RECT -76.325 174.595 -75.995 174.925 ;
        RECT -76.325 173.235 -75.995 173.565 ;
        RECT -76.325 171.875 -75.995 172.205 ;
        RECT -76.325 170.515 -75.995 170.845 ;
        RECT -76.325 169.155 -75.995 169.485 ;
        RECT -76.325 167.795 -75.995 168.125 ;
        RECT -76.325 166.435 -75.995 166.765 ;
        RECT -76.325 165.075 -75.995 165.405 ;
        RECT -76.325 163.715 -75.995 164.045 ;
        RECT -76.325 162.355 -75.995 162.685 ;
        RECT -76.325 160.995 -75.995 161.325 ;
        RECT -76.325 159.635 -75.995 159.965 ;
        RECT -76.325 158.275 -75.995 158.605 ;
        RECT -76.325 156.915 -75.995 157.245 ;
        RECT -76.325 155.555 -75.995 155.885 ;
        RECT -76.325 154.195 -75.995 154.525 ;
        RECT -76.325 152.835 -75.995 153.165 ;
        RECT -76.325 151.475 -75.995 151.805 ;
        RECT -76.325 150.115 -75.995 150.445 ;
        RECT -76.325 148.755 -75.995 149.085 ;
        RECT -76.325 147.395 -75.995 147.725 ;
        RECT -76.325 146.035 -75.995 146.365 ;
        RECT -76.325 144.675 -75.995 145.005 ;
        RECT -76.325 143.315 -75.995 143.645 ;
        RECT -76.325 141.955 -75.995 142.285 ;
        RECT -76.325 140.595 -75.995 140.925 ;
        RECT -76.325 139.235 -75.995 139.565 ;
        RECT -76.325 137.875 -75.995 138.205 ;
        RECT -76.325 136.515 -75.995 136.845 ;
        RECT -76.325 135.155 -75.995 135.485 ;
        RECT -76.325 133.795 -75.995 134.125 ;
        RECT -76.325 132.435 -75.995 132.765 ;
        RECT -76.325 131.075 -75.995 131.405 ;
        RECT -76.325 129.715 -75.995 130.045 ;
        RECT -76.325 128.355 -75.995 128.685 ;
        RECT -76.325 126.995 -75.995 127.325 ;
        RECT -76.325 125.635 -75.995 125.965 ;
        RECT -76.325 124.275 -75.995 124.605 ;
        RECT -76.325 122.915 -75.995 123.245 ;
        RECT -76.325 121.555 -75.995 121.885 ;
        RECT -76.325 120.195 -75.995 120.525 ;
        RECT -76.325 118.835 -75.995 119.165 ;
        RECT -76.325 117.475 -75.995 117.805 ;
        RECT -76.325 116.115 -75.995 116.445 ;
        RECT -76.325 114.755 -75.995 115.085 ;
        RECT -76.325 113.395 -75.995 113.725 ;
        RECT -76.325 112.035 -75.995 112.365 ;
        RECT -76.325 110.675 -75.995 111.005 ;
        RECT -76.325 109.315 -75.995 109.645 ;
        RECT -76.325 107.955 -75.995 108.285 ;
        RECT -76.325 106.595 -75.995 106.925 ;
        RECT -76.325 105.235 -75.995 105.565 ;
        RECT -76.325 103.875 -75.995 104.205 ;
        RECT -76.325 102.515 -75.995 102.845 ;
        RECT -76.325 101.155 -75.995 101.485 ;
        RECT -76.325 99.795 -75.995 100.125 ;
        RECT -76.325 98.435 -75.995 98.765 ;
        RECT -76.325 97.075 -75.995 97.405 ;
        RECT -76.325 95.715 -75.995 96.045 ;
        RECT -76.325 94.355 -75.995 94.685 ;
        RECT -76.325 92.995 -75.995 93.325 ;
        RECT -76.325 91.635 -75.995 91.965 ;
        RECT -76.325 90.275 -75.995 90.605 ;
        RECT -76.325 88.915 -75.995 89.245 ;
        RECT -76.325 87.555 -75.995 87.885 ;
        RECT -76.325 86.195 -75.995 86.525 ;
        RECT -76.325 84.835 -75.995 85.165 ;
        RECT -76.325 83.475 -75.995 83.805 ;
        RECT -76.325 82.115 -75.995 82.445 ;
        RECT -76.325 80.755 -75.995 81.085 ;
        RECT -76.325 79.395 -75.995 79.725 ;
        RECT -76.325 78.035 -75.995 78.365 ;
        RECT -76.325 76.675 -75.995 77.005 ;
        RECT -76.325 75.315 -75.995 75.645 ;
        RECT -76.325 73.955 -75.995 74.285 ;
        RECT -76.325 72.595 -75.995 72.925 ;
        RECT -76.325 71.235 -75.995 71.565 ;
        RECT -76.325 69.875 -75.995 70.205 ;
        RECT -76.325 68.515 -75.995 68.845 ;
        RECT -76.325 67.155 -75.995 67.485 ;
        RECT -76.325 65.795 -75.995 66.125 ;
        RECT -76.325 64.435 -75.995 64.765 ;
        RECT -76.325 63.075 -75.995 63.405 ;
        RECT -76.325 61.715 -75.995 62.045 ;
        RECT -76.325 60.355 -75.995 60.685 ;
        RECT -76.325 58.995 -75.995 59.325 ;
        RECT -76.325 57.635 -75.995 57.965 ;
        RECT -76.325 56.275 -75.995 56.605 ;
        RECT -76.325 54.915 -75.995 55.245 ;
        RECT -76.325 53.555 -75.995 53.885 ;
        RECT -76.325 52.195 -75.995 52.525 ;
        RECT -76.325 50.835 -75.995 51.165 ;
        RECT -76.325 49.475 -75.995 49.805 ;
        RECT -76.325 48.115 -75.995 48.445 ;
        RECT -76.325 46.755 -75.995 47.085 ;
        RECT -76.325 45.395 -75.995 45.725 ;
        RECT -76.325 44.035 -75.995 44.365 ;
        RECT -76.325 42.675 -75.995 43.005 ;
        RECT -76.325 41.315 -75.995 41.645 ;
        RECT -76.325 39.955 -75.995 40.285 ;
        RECT -76.325 38.595 -75.995 38.925 ;
        RECT -76.325 37.235 -75.995 37.565 ;
        RECT -76.325 35.875 -75.995 36.205 ;
        RECT -76.325 34.515 -75.995 34.845 ;
        RECT -76.325 33.155 -75.995 33.485 ;
        RECT -76.325 31.795 -75.995 32.125 ;
        RECT -76.325 30.435 -75.995 30.765 ;
        RECT -76.325 29.075 -75.995 29.405 ;
        RECT -76.325 27.715 -75.995 28.045 ;
        RECT -76.325 26.355 -75.995 26.685 ;
        RECT -76.325 24.995 -75.995 25.325 ;
        RECT -76.325 23.635 -75.995 23.965 ;
        RECT -76.325 22.275 -75.995 22.605 ;
        RECT -76.325 20.915 -75.995 21.245 ;
        RECT -76.325 19.555 -75.995 19.885 ;
        RECT -76.325 18.195 -75.995 18.525 ;
        RECT -76.325 16.835 -75.995 17.165 ;
        RECT -76.325 15.475 -75.995 15.805 ;
        RECT -76.325 14.115 -75.995 14.445 ;
        RECT -76.325 12.755 -75.995 13.085 ;
        RECT -76.325 11.395 -75.995 11.725 ;
        RECT -76.325 10.035 -75.995 10.365 ;
        RECT -76.325 8.675 -75.995 9.005 ;
        RECT -76.325 7.315 -75.995 7.645 ;
        RECT -76.325 5.955 -75.995 6.285 ;
        RECT -76.325 4.595 -75.995 4.925 ;
        RECT -76.325 3.235 -75.995 3.565 ;
        RECT -76.325 1.875 -75.995 2.205 ;
        RECT -76.325 0.515 -75.995 0.845 ;
        RECT -76.325 -0.845 -75.995 -0.515 ;
        RECT -76.325 -2.205 -75.995 -1.875 ;
        RECT -76.325 -3.565 -75.995 -3.235 ;
        RECT -76.325 -4.925 -75.995 -4.595 ;
        RECT -76.325 -6.285 -75.995 -5.955 ;
        RECT -76.325 -7.645 -75.995 -7.315 ;
        RECT -76.325 -9.005 -75.995 -8.675 ;
        RECT -76.325 -10.365 -75.995 -10.035 ;
        RECT -76.325 -11.725 -75.995 -11.395 ;
        RECT -76.325 -13.085 -75.995 -12.755 ;
        RECT -76.325 -14.445 -75.995 -14.115 ;
        RECT -76.325 -15.805 -75.995 -15.475 ;
        RECT -76.325 -17.165 -75.995 -16.835 ;
        RECT -76.325 -18.525 -75.995 -18.195 ;
        RECT -76.325 -19.885 -75.995 -19.555 ;
        RECT -76.325 -21.245 -75.995 -20.915 ;
        RECT -76.325 -22.605 -75.995 -22.275 ;
        RECT -76.325 -23.965 -75.995 -23.635 ;
        RECT -76.325 -25.325 -75.995 -24.995 ;
        RECT -76.325 -26.685 -75.995 -26.355 ;
        RECT -76.325 -28.045 -75.995 -27.715 ;
        RECT -76.325 -29.405 -75.995 -29.075 ;
        RECT -76.325 -30.765 -75.995 -30.435 ;
        RECT -76.325 -32.125 -75.995 -31.795 ;
        RECT -76.325 -33.485 -75.995 -33.155 ;
        RECT -76.325 -34.845 -75.995 -34.515 ;
        RECT -76.325 -36.205 -75.995 -35.875 ;
        RECT -76.325 -37.565 -75.995 -37.235 ;
        RECT -76.325 -38.925 -75.995 -38.595 ;
        RECT -76.325 -40.285 -75.995 -39.955 ;
        RECT -76.325 -41.645 -75.995 -41.315 ;
        RECT -76.325 -43.005 -75.995 -42.675 ;
        RECT -76.325 -44.365 -75.995 -44.035 ;
        RECT -76.325 -45.725 -75.995 -45.395 ;
        RECT -76.325 -47.085 -75.995 -46.755 ;
        RECT -76.325 -48.445 -75.995 -48.115 ;
        RECT -76.325 -49.805 -75.995 -49.475 ;
        RECT -76.325 -51.165 -75.995 -50.835 ;
        RECT -76.325 -52.525 -75.995 -52.195 ;
        RECT -76.325 -53.885 -75.995 -53.555 ;
        RECT -76.325 -55.245 -75.995 -54.915 ;
        RECT -76.325 -56.605 -75.995 -56.275 ;
        RECT -76.325 -57.965 -75.995 -57.635 ;
        RECT -76.325 -59.325 -75.995 -58.995 ;
        RECT -76.325 -60.685 -75.995 -60.355 ;
        RECT -76.325 -62.045 -75.995 -61.715 ;
        RECT -76.325 -63.405 -75.995 -63.075 ;
        RECT -76.325 -64.765 -75.995 -64.435 ;
        RECT -76.325 -66.125 -75.995 -65.795 ;
        RECT -76.325 -67.485 -75.995 -67.155 ;
        RECT -76.325 -68.845 -75.995 -68.515 ;
        RECT -76.325 -70.205 -75.995 -69.875 ;
        RECT -76.325 -71.565 -75.995 -71.235 ;
        RECT -76.325 -72.925 -75.995 -72.595 ;
        RECT -76.325 -74.285 -75.995 -73.955 ;
        RECT -76.325 -75.645 -75.995 -75.315 ;
        RECT -76.325 -77.005 -75.995 -76.675 ;
        RECT -76.325 -78.365 -75.995 -78.035 ;
        RECT -76.325 -79.725 -75.995 -79.395 ;
        RECT -76.325 -81.085 -75.995 -80.755 ;
        RECT -76.325 -82.445 -75.995 -82.115 ;
        RECT -76.325 -83.805 -75.995 -83.475 ;
        RECT -76.325 -85.165 -75.995 -84.835 ;
        RECT -76.325 -86.525 -75.995 -86.195 ;
        RECT -76.325 -87.885 -75.995 -87.555 ;
        RECT -76.325 -89.245 -75.995 -88.915 ;
        RECT -76.325 -90.605 -75.995 -90.275 ;
        RECT -76.325 -91.965 -75.995 -91.635 ;
        RECT -76.325 -93.325 -75.995 -92.995 ;
        RECT -76.325 -94.685 -75.995 -94.355 ;
        RECT -76.325 -96.045 -75.995 -95.715 ;
        RECT -76.325 -97.405 -75.995 -97.075 ;
        RECT -76.325 -98.765 -75.995 -98.435 ;
        RECT -76.325 -100.125 -75.995 -99.795 ;
        RECT -76.325 -101.485 -75.995 -101.155 ;
        RECT -76.325 -102.845 -75.995 -102.515 ;
        RECT -76.325 -104.205 -75.995 -103.875 ;
        RECT -76.325 -105.565 -75.995 -105.235 ;
        RECT -76.325 -106.925 -75.995 -106.595 ;
        RECT -76.325 -108.285 -75.995 -107.955 ;
        RECT -76.325 -109.645 -75.995 -109.315 ;
        RECT -76.325 -111.005 -75.995 -110.675 ;
        RECT -76.325 -112.365 -75.995 -112.035 ;
        RECT -76.325 -113.725 -75.995 -113.395 ;
        RECT -76.325 -115.085 -75.995 -114.755 ;
        RECT -76.325 -116.445 -75.995 -116.115 ;
        RECT -76.325 -117.805 -75.995 -117.475 ;
        RECT -76.325 -119.165 -75.995 -118.835 ;
        RECT -76.325 -120.525 -75.995 -120.195 ;
        RECT -76.325 -121.885 -75.995 -121.555 ;
        RECT -76.325 -123.245 -75.995 -122.915 ;
        RECT -76.325 -124.605 -75.995 -124.275 ;
        RECT -76.325 -125.965 -75.995 -125.635 ;
        RECT -76.325 -127.325 -75.995 -126.995 ;
        RECT -76.325 -128.685 -75.995 -128.355 ;
        RECT -76.325 -130.045 -75.995 -129.715 ;
        RECT -76.325 -131.405 -75.995 -131.075 ;
        RECT -76.325 -132.765 -75.995 -132.435 ;
        RECT -76.325 -134.125 -75.995 -133.795 ;
        RECT -76.325 -135.485 -75.995 -135.155 ;
        RECT -76.325 -136.845 -75.995 -136.515 ;
        RECT -76.325 -138.205 -75.995 -137.875 ;
        RECT -76.325 -139.565 -75.995 -139.235 ;
        RECT -76.325 -140.925 -75.995 -140.595 ;
        RECT -76.325 -142.285 -75.995 -141.955 ;
        RECT -76.325 -143.645 -75.995 -143.315 ;
        RECT -76.325 -145.005 -75.995 -144.675 ;
        RECT -76.325 -146.365 -75.995 -146.035 ;
        RECT -76.325 -147.725 -75.995 -147.395 ;
        RECT -76.325 -149.085 -75.995 -148.755 ;
        RECT -76.325 -150.445 -75.995 -150.115 ;
        RECT -76.325 -151.805 -75.995 -151.475 ;
        RECT -76.325 -153.165 -75.995 -152.835 ;
        RECT -76.325 -154.525 -75.995 -154.195 ;
        RECT -76.325 -155.885 -75.995 -155.555 ;
        RECT -76.325 -157.245 -75.995 -156.915 ;
        RECT -76.325 -158.605 -75.995 -158.275 ;
        RECT -76.325 -159.965 -75.995 -159.635 ;
        RECT -76.325 -161.325 -75.995 -160.995 ;
        RECT -76.325 -162.685 -75.995 -162.355 ;
        RECT -76.325 -164.045 -75.995 -163.715 ;
        RECT -76.325 -165.405 -75.995 -165.075 ;
        RECT -76.325 -166.765 -75.995 -166.435 ;
        RECT -76.325 -168.125 -75.995 -167.795 ;
        RECT -76.325 -169.615 -75.995 -169.285 ;
        RECT -76.325 -170.845 -75.995 -170.515 ;
        RECT -76.325 -172.205 -75.995 -171.875 ;
        RECT -76.325 -174.925 -75.995 -174.595 ;
        RECT -76.325 -177.645 -75.995 -177.315 ;
        RECT -76.325 -179.005 -75.995 -178.675 ;
        RECT -76.325 -184.65 -75.995 -183.52 ;
        RECT -76.32 -184.765 -76 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -74.965 244.04 -74.635 245.17 ;
        RECT -74.965 239.875 -74.635 240.205 ;
        RECT -74.965 238.515 -74.635 238.845 ;
        RECT -74.965 237.155 -74.635 237.485 ;
        RECT -74.965 235.795 -74.635 236.125 ;
        RECT -74.965 234.435 -74.635 234.765 ;
        RECT -74.965 233.075 -74.635 233.405 ;
        RECT -74.965 231.715 -74.635 232.045 ;
        RECT -74.965 230.355 -74.635 230.685 ;
        RECT -74.965 228.995 -74.635 229.325 ;
        RECT -74.965 227.635 -74.635 227.965 ;
        RECT -74.965 226.275 -74.635 226.605 ;
        RECT -74.965 224.915 -74.635 225.245 ;
        RECT -74.965 223.555 -74.635 223.885 ;
        RECT -74.965 222.195 -74.635 222.525 ;
        RECT -74.965 220.835 -74.635 221.165 ;
        RECT -74.965 219.475 -74.635 219.805 ;
        RECT -74.965 218.115 -74.635 218.445 ;
        RECT -74.965 216.755 -74.635 217.085 ;
        RECT -74.965 215.395 -74.635 215.725 ;
        RECT -74.965 214.035 -74.635 214.365 ;
        RECT -74.965 212.675 -74.635 213.005 ;
        RECT -74.965 211.315 -74.635 211.645 ;
        RECT -74.965 209.955 -74.635 210.285 ;
        RECT -74.965 208.595 -74.635 208.925 ;
        RECT -74.965 207.235 -74.635 207.565 ;
        RECT -74.965 205.875 -74.635 206.205 ;
        RECT -74.965 204.515 -74.635 204.845 ;
        RECT -74.965 203.155 -74.635 203.485 ;
        RECT -74.965 201.795 -74.635 202.125 ;
        RECT -74.965 200.435 -74.635 200.765 ;
        RECT -74.965 199.075 -74.635 199.405 ;
        RECT -74.965 197.715 -74.635 198.045 ;
        RECT -74.965 196.355 -74.635 196.685 ;
        RECT -74.965 194.995 -74.635 195.325 ;
        RECT -74.965 193.635 -74.635 193.965 ;
        RECT -74.965 192.275 -74.635 192.605 ;
        RECT -74.965 190.915 -74.635 191.245 ;
        RECT -74.965 189.555 -74.635 189.885 ;
        RECT -74.965 188.195 -74.635 188.525 ;
        RECT -74.965 186.835 -74.635 187.165 ;
        RECT -74.965 185.475 -74.635 185.805 ;
        RECT -74.965 184.115 -74.635 184.445 ;
        RECT -74.965 182.755 -74.635 183.085 ;
        RECT -74.965 181.395 -74.635 181.725 ;
        RECT -74.965 180.035 -74.635 180.365 ;
        RECT -74.965 178.675 -74.635 179.005 ;
        RECT -74.965 177.315 -74.635 177.645 ;
        RECT -74.965 175.955 -74.635 176.285 ;
        RECT -74.965 174.595 -74.635 174.925 ;
        RECT -74.965 173.235 -74.635 173.565 ;
        RECT -74.965 171.875 -74.635 172.205 ;
        RECT -74.965 170.515 -74.635 170.845 ;
        RECT -74.965 169.155 -74.635 169.485 ;
        RECT -74.965 167.795 -74.635 168.125 ;
        RECT -74.965 166.435 -74.635 166.765 ;
        RECT -74.965 165.075 -74.635 165.405 ;
        RECT -74.965 163.715 -74.635 164.045 ;
        RECT -74.965 162.355 -74.635 162.685 ;
        RECT -74.965 160.995 -74.635 161.325 ;
        RECT -74.965 159.635 -74.635 159.965 ;
        RECT -74.965 158.275 -74.635 158.605 ;
        RECT -74.965 156.915 -74.635 157.245 ;
        RECT -74.965 155.555 -74.635 155.885 ;
        RECT -74.965 154.195 -74.635 154.525 ;
        RECT -74.965 152.835 -74.635 153.165 ;
        RECT -74.965 151.475 -74.635 151.805 ;
        RECT -74.965 150.115 -74.635 150.445 ;
        RECT -74.965 148.755 -74.635 149.085 ;
        RECT -74.965 147.395 -74.635 147.725 ;
        RECT -74.965 146.035 -74.635 146.365 ;
        RECT -74.965 144.675 -74.635 145.005 ;
        RECT -74.965 143.315 -74.635 143.645 ;
        RECT -74.965 141.955 -74.635 142.285 ;
        RECT -74.965 140.595 -74.635 140.925 ;
        RECT -74.965 139.235 -74.635 139.565 ;
        RECT -74.965 137.875 -74.635 138.205 ;
        RECT -74.965 136.515 -74.635 136.845 ;
        RECT -74.965 135.155 -74.635 135.485 ;
        RECT -74.965 133.795 -74.635 134.125 ;
        RECT -74.965 132.435 -74.635 132.765 ;
        RECT -74.965 131.075 -74.635 131.405 ;
        RECT -74.965 129.715 -74.635 130.045 ;
        RECT -74.965 128.355 -74.635 128.685 ;
        RECT -74.965 126.995 -74.635 127.325 ;
        RECT -74.965 125.635 -74.635 125.965 ;
        RECT -74.965 124.275 -74.635 124.605 ;
        RECT -74.965 122.915 -74.635 123.245 ;
        RECT -74.965 121.555 -74.635 121.885 ;
        RECT -74.965 120.195 -74.635 120.525 ;
        RECT -74.965 118.835 -74.635 119.165 ;
        RECT -74.965 117.475 -74.635 117.805 ;
        RECT -74.965 116.115 -74.635 116.445 ;
        RECT -74.965 114.755 -74.635 115.085 ;
        RECT -74.965 113.395 -74.635 113.725 ;
        RECT -74.965 112.035 -74.635 112.365 ;
        RECT -74.965 110.675 -74.635 111.005 ;
        RECT -74.965 109.315 -74.635 109.645 ;
        RECT -74.965 107.955 -74.635 108.285 ;
        RECT -74.965 106.595 -74.635 106.925 ;
        RECT -74.965 105.235 -74.635 105.565 ;
        RECT -74.965 103.875 -74.635 104.205 ;
        RECT -74.965 102.515 -74.635 102.845 ;
        RECT -74.965 101.155 -74.635 101.485 ;
        RECT -74.965 99.795 -74.635 100.125 ;
        RECT -74.965 98.435 -74.635 98.765 ;
        RECT -74.965 97.075 -74.635 97.405 ;
        RECT -74.965 95.715 -74.635 96.045 ;
        RECT -74.965 94.355 -74.635 94.685 ;
        RECT -74.965 92.995 -74.635 93.325 ;
        RECT -74.965 91.635 -74.635 91.965 ;
        RECT -74.965 90.275 -74.635 90.605 ;
        RECT -74.965 88.915 -74.635 89.245 ;
        RECT -74.965 87.555 -74.635 87.885 ;
        RECT -74.965 86.195 -74.635 86.525 ;
        RECT -74.965 84.835 -74.635 85.165 ;
        RECT -74.965 83.475 -74.635 83.805 ;
        RECT -74.965 82.115 -74.635 82.445 ;
        RECT -74.965 80.755 -74.635 81.085 ;
        RECT -74.965 79.395 -74.635 79.725 ;
        RECT -74.965 78.035 -74.635 78.365 ;
        RECT -74.965 76.675 -74.635 77.005 ;
        RECT -74.965 75.315 -74.635 75.645 ;
        RECT -74.965 73.955 -74.635 74.285 ;
        RECT -74.965 72.595 -74.635 72.925 ;
        RECT -74.965 71.235 -74.635 71.565 ;
        RECT -74.965 69.875 -74.635 70.205 ;
        RECT -74.965 68.515 -74.635 68.845 ;
        RECT -74.965 67.155 -74.635 67.485 ;
        RECT -74.965 65.795 -74.635 66.125 ;
        RECT -74.965 64.435 -74.635 64.765 ;
        RECT -74.965 63.075 -74.635 63.405 ;
        RECT -74.965 61.715 -74.635 62.045 ;
        RECT -74.965 60.355 -74.635 60.685 ;
        RECT -74.965 58.995 -74.635 59.325 ;
        RECT -74.965 57.635 -74.635 57.965 ;
        RECT -74.965 56.275 -74.635 56.605 ;
        RECT -74.965 54.915 -74.635 55.245 ;
        RECT -74.965 53.555 -74.635 53.885 ;
        RECT -74.965 52.195 -74.635 52.525 ;
        RECT -74.965 50.835 -74.635 51.165 ;
        RECT -74.965 49.475 -74.635 49.805 ;
        RECT -74.965 48.115 -74.635 48.445 ;
        RECT -74.965 46.755 -74.635 47.085 ;
        RECT -74.965 45.395 -74.635 45.725 ;
        RECT -74.965 44.035 -74.635 44.365 ;
        RECT -74.965 42.675 -74.635 43.005 ;
        RECT -74.965 41.315 -74.635 41.645 ;
        RECT -74.965 39.955 -74.635 40.285 ;
        RECT -74.965 38.595 -74.635 38.925 ;
        RECT -74.965 37.235 -74.635 37.565 ;
        RECT -74.965 35.875 -74.635 36.205 ;
        RECT -74.965 34.515 -74.635 34.845 ;
        RECT -74.965 33.155 -74.635 33.485 ;
        RECT -74.965 31.795 -74.635 32.125 ;
        RECT -74.965 30.435 -74.635 30.765 ;
        RECT -74.965 29.075 -74.635 29.405 ;
        RECT -74.965 27.715 -74.635 28.045 ;
        RECT -74.965 26.355 -74.635 26.685 ;
        RECT -74.965 24.995 -74.635 25.325 ;
        RECT -74.965 23.635 -74.635 23.965 ;
        RECT -74.965 22.275 -74.635 22.605 ;
        RECT -74.965 20.915 -74.635 21.245 ;
        RECT -74.965 19.555 -74.635 19.885 ;
        RECT -74.965 18.195 -74.635 18.525 ;
        RECT -74.965 16.835 -74.635 17.165 ;
        RECT -74.965 15.475 -74.635 15.805 ;
        RECT -74.965 14.115 -74.635 14.445 ;
        RECT -74.965 12.755 -74.635 13.085 ;
        RECT -74.965 11.395 -74.635 11.725 ;
        RECT -74.965 10.035 -74.635 10.365 ;
        RECT -74.965 8.675 -74.635 9.005 ;
        RECT -74.965 7.315 -74.635 7.645 ;
        RECT -74.965 5.955 -74.635 6.285 ;
        RECT -74.965 4.595 -74.635 4.925 ;
        RECT -74.965 3.235 -74.635 3.565 ;
        RECT -74.965 1.875 -74.635 2.205 ;
        RECT -74.965 0.515 -74.635 0.845 ;
        RECT -74.965 -0.845 -74.635 -0.515 ;
        RECT -74.965 -2.205 -74.635 -1.875 ;
        RECT -74.965 -3.565 -74.635 -3.235 ;
        RECT -74.965 -4.925 -74.635 -4.595 ;
        RECT -74.965 -6.285 -74.635 -5.955 ;
        RECT -74.965 -7.645 -74.635 -7.315 ;
        RECT -74.965 -9.005 -74.635 -8.675 ;
        RECT -74.965 -10.365 -74.635 -10.035 ;
        RECT -74.965 -11.725 -74.635 -11.395 ;
        RECT -74.965 -13.085 -74.635 -12.755 ;
        RECT -74.965 -14.445 -74.635 -14.115 ;
        RECT -74.965 -15.805 -74.635 -15.475 ;
        RECT -74.965 -17.165 -74.635 -16.835 ;
        RECT -74.965 -18.525 -74.635 -18.195 ;
        RECT -74.965 -19.885 -74.635 -19.555 ;
        RECT -74.965 -21.245 -74.635 -20.915 ;
        RECT -74.965 -22.605 -74.635 -22.275 ;
        RECT -74.965 -23.965 -74.635 -23.635 ;
        RECT -74.965 -25.325 -74.635 -24.995 ;
        RECT -74.965 -26.685 -74.635 -26.355 ;
        RECT -74.965 -28.045 -74.635 -27.715 ;
        RECT -74.965 -29.405 -74.635 -29.075 ;
        RECT -74.965 -30.765 -74.635 -30.435 ;
        RECT -74.965 -32.125 -74.635 -31.795 ;
        RECT -74.965 -33.485 -74.635 -33.155 ;
        RECT -74.965 -34.845 -74.635 -34.515 ;
        RECT -74.965 -36.205 -74.635 -35.875 ;
        RECT -74.965 -37.565 -74.635 -37.235 ;
        RECT -74.965 -38.925 -74.635 -38.595 ;
        RECT -74.965 -40.285 -74.635 -39.955 ;
        RECT -74.965 -41.645 -74.635 -41.315 ;
        RECT -74.965 -43.005 -74.635 -42.675 ;
        RECT -74.965 -44.365 -74.635 -44.035 ;
        RECT -74.965 -45.725 -74.635 -45.395 ;
        RECT -74.965 -47.085 -74.635 -46.755 ;
        RECT -74.965 -48.445 -74.635 -48.115 ;
        RECT -74.965 -49.805 -74.635 -49.475 ;
        RECT -74.965 -51.165 -74.635 -50.835 ;
        RECT -74.965 -52.525 -74.635 -52.195 ;
        RECT -74.965 -53.885 -74.635 -53.555 ;
        RECT -74.965 -55.245 -74.635 -54.915 ;
        RECT -74.965 -56.605 -74.635 -56.275 ;
        RECT -74.965 -57.965 -74.635 -57.635 ;
        RECT -74.965 -59.325 -74.635 -58.995 ;
        RECT -74.965 -60.685 -74.635 -60.355 ;
        RECT -74.965 -62.045 -74.635 -61.715 ;
        RECT -74.965 -63.405 -74.635 -63.075 ;
        RECT -74.965 -64.765 -74.635 -64.435 ;
        RECT -74.965 -66.125 -74.635 -65.795 ;
        RECT -74.965 -67.485 -74.635 -67.155 ;
        RECT -74.965 -68.845 -74.635 -68.515 ;
        RECT -74.965 -70.205 -74.635 -69.875 ;
        RECT -74.965 -71.565 -74.635 -71.235 ;
        RECT -74.965 -72.925 -74.635 -72.595 ;
        RECT -74.965 -74.285 -74.635 -73.955 ;
        RECT -74.965 -75.645 -74.635 -75.315 ;
        RECT -74.965 -77.005 -74.635 -76.675 ;
        RECT -74.965 -78.365 -74.635 -78.035 ;
        RECT -74.965 -79.725 -74.635 -79.395 ;
        RECT -74.965 -81.085 -74.635 -80.755 ;
        RECT -74.965 -82.445 -74.635 -82.115 ;
        RECT -74.965 -83.805 -74.635 -83.475 ;
        RECT -74.965 -85.165 -74.635 -84.835 ;
        RECT -74.965 -86.525 -74.635 -86.195 ;
        RECT -74.965 -87.885 -74.635 -87.555 ;
        RECT -74.965 -89.245 -74.635 -88.915 ;
        RECT -74.965 -90.605 -74.635 -90.275 ;
        RECT -74.965 -91.965 -74.635 -91.635 ;
        RECT -74.965 -93.325 -74.635 -92.995 ;
        RECT -74.965 -94.685 -74.635 -94.355 ;
        RECT -74.965 -96.045 -74.635 -95.715 ;
        RECT -74.965 -97.405 -74.635 -97.075 ;
        RECT -74.965 -98.765 -74.635 -98.435 ;
        RECT -74.965 -100.125 -74.635 -99.795 ;
        RECT -74.965 -101.485 -74.635 -101.155 ;
        RECT -74.965 -102.845 -74.635 -102.515 ;
        RECT -74.965 -104.205 -74.635 -103.875 ;
        RECT -74.965 -105.565 -74.635 -105.235 ;
        RECT -74.965 -106.925 -74.635 -106.595 ;
        RECT -74.965 -108.285 -74.635 -107.955 ;
        RECT -74.965 -109.645 -74.635 -109.315 ;
        RECT -74.965 -111.005 -74.635 -110.675 ;
        RECT -74.965 -112.365 -74.635 -112.035 ;
        RECT -74.965 -113.725 -74.635 -113.395 ;
        RECT -74.965 -115.085 -74.635 -114.755 ;
        RECT -74.965 -116.445 -74.635 -116.115 ;
        RECT -74.965 -117.805 -74.635 -117.475 ;
        RECT -74.965 -119.165 -74.635 -118.835 ;
        RECT -74.965 -120.525 -74.635 -120.195 ;
        RECT -74.965 -121.885 -74.635 -121.555 ;
        RECT -74.965 -123.245 -74.635 -122.915 ;
        RECT -74.965 -124.605 -74.635 -124.275 ;
        RECT -74.965 -125.965 -74.635 -125.635 ;
        RECT -74.965 -127.325 -74.635 -126.995 ;
        RECT -74.965 -128.685 -74.635 -128.355 ;
        RECT -74.965 -130.045 -74.635 -129.715 ;
        RECT -74.965 -131.405 -74.635 -131.075 ;
        RECT -74.965 -132.765 -74.635 -132.435 ;
        RECT -74.965 -134.125 -74.635 -133.795 ;
        RECT -74.965 -135.485 -74.635 -135.155 ;
        RECT -74.965 -136.845 -74.635 -136.515 ;
        RECT -74.965 -138.205 -74.635 -137.875 ;
        RECT -74.965 -139.565 -74.635 -139.235 ;
        RECT -74.965 -140.925 -74.635 -140.595 ;
        RECT -74.965 -142.285 -74.635 -141.955 ;
        RECT -74.965 -143.645 -74.635 -143.315 ;
        RECT -74.965 -145.005 -74.635 -144.675 ;
        RECT -74.965 -146.365 -74.635 -146.035 ;
        RECT -74.965 -147.725 -74.635 -147.395 ;
        RECT -74.965 -149.085 -74.635 -148.755 ;
        RECT -74.965 -150.445 -74.635 -150.115 ;
        RECT -74.965 -151.805 -74.635 -151.475 ;
        RECT -74.965 -153.165 -74.635 -152.835 ;
        RECT -74.965 -154.525 -74.635 -154.195 ;
        RECT -74.965 -155.885 -74.635 -155.555 ;
        RECT -74.965 -157.245 -74.635 -156.915 ;
        RECT -74.965 -158.605 -74.635 -158.275 ;
        RECT -74.965 -159.965 -74.635 -159.635 ;
        RECT -74.965 -161.325 -74.635 -160.995 ;
        RECT -74.965 -162.685 -74.635 -162.355 ;
        RECT -74.965 -164.045 -74.635 -163.715 ;
        RECT -74.965 -165.405 -74.635 -165.075 ;
        RECT -74.965 -166.765 -74.635 -166.435 ;
        RECT -74.965 -168.125 -74.635 -167.795 ;
        RECT -74.965 -169.615 -74.635 -169.285 ;
        RECT -74.965 -170.845 -74.635 -170.515 ;
        RECT -74.965 -172.205 -74.635 -171.875 ;
        RECT -74.965 -173.565 -74.635 -173.235 ;
        RECT -74.965 -174.925 -74.635 -174.595 ;
        RECT -74.965 -177.645 -74.635 -177.315 ;
        RECT -74.965 -179.005 -74.635 -178.675 ;
        RECT -74.965 -184.65 -74.635 -183.52 ;
        RECT -74.96 -184.765 -74.64 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -73.605 200.435 -73.275 200.765 ;
        RECT -73.605 199.075 -73.275 199.405 ;
        RECT -73.605 197.715 -73.275 198.045 ;
        RECT -73.605 196.355 -73.275 196.685 ;
        RECT -73.605 194.995 -73.275 195.325 ;
        RECT -73.605 193.635 -73.275 193.965 ;
        RECT -73.605 192.275 -73.275 192.605 ;
        RECT -73.605 190.915 -73.275 191.245 ;
        RECT -73.605 189.555 -73.275 189.885 ;
        RECT -73.605 188.195 -73.275 188.525 ;
        RECT -73.605 186.835 -73.275 187.165 ;
        RECT -73.605 185.475 -73.275 185.805 ;
        RECT -73.605 184.115 -73.275 184.445 ;
        RECT -73.605 182.755 -73.275 183.085 ;
        RECT -73.605 181.395 -73.275 181.725 ;
        RECT -73.605 180.035 -73.275 180.365 ;
        RECT -73.605 178.675 -73.275 179.005 ;
        RECT -73.605 177.315 -73.275 177.645 ;
        RECT -73.605 175.955 -73.275 176.285 ;
        RECT -73.605 174.595 -73.275 174.925 ;
        RECT -73.605 173.235 -73.275 173.565 ;
        RECT -73.605 171.875 -73.275 172.205 ;
        RECT -73.605 170.515 -73.275 170.845 ;
        RECT -73.605 169.155 -73.275 169.485 ;
        RECT -73.605 167.795 -73.275 168.125 ;
        RECT -73.605 166.435 -73.275 166.765 ;
        RECT -73.605 165.075 -73.275 165.405 ;
        RECT -73.605 163.715 -73.275 164.045 ;
        RECT -73.605 162.355 -73.275 162.685 ;
        RECT -73.605 160.995 -73.275 161.325 ;
        RECT -73.605 159.635 -73.275 159.965 ;
        RECT -73.605 158.275 -73.275 158.605 ;
        RECT -73.605 156.915 -73.275 157.245 ;
        RECT -73.605 155.555 -73.275 155.885 ;
        RECT -73.605 154.195 -73.275 154.525 ;
        RECT -73.605 152.835 -73.275 153.165 ;
        RECT -73.605 151.475 -73.275 151.805 ;
        RECT -73.605 150.115 -73.275 150.445 ;
        RECT -73.605 148.755 -73.275 149.085 ;
        RECT -73.605 147.395 -73.275 147.725 ;
        RECT -73.605 146.035 -73.275 146.365 ;
        RECT -73.605 144.675 -73.275 145.005 ;
        RECT -73.605 143.315 -73.275 143.645 ;
        RECT -73.605 141.955 -73.275 142.285 ;
        RECT -73.605 140.595 -73.275 140.925 ;
        RECT -73.605 139.235 -73.275 139.565 ;
        RECT -73.605 137.875 -73.275 138.205 ;
        RECT -73.605 136.515 -73.275 136.845 ;
        RECT -73.605 135.155 -73.275 135.485 ;
        RECT -73.605 133.795 -73.275 134.125 ;
        RECT -73.605 132.435 -73.275 132.765 ;
        RECT -73.605 131.075 -73.275 131.405 ;
        RECT -73.605 129.715 -73.275 130.045 ;
        RECT -73.605 128.355 -73.275 128.685 ;
        RECT -73.605 126.995 -73.275 127.325 ;
        RECT -73.605 125.635 -73.275 125.965 ;
        RECT -73.605 124.275 -73.275 124.605 ;
        RECT -73.605 122.915 -73.275 123.245 ;
        RECT -73.605 121.555 -73.275 121.885 ;
        RECT -73.605 120.195 -73.275 120.525 ;
        RECT -73.605 118.835 -73.275 119.165 ;
        RECT -73.605 117.475 -73.275 117.805 ;
        RECT -73.605 116.115 -73.275 116.445 ;
        RECT -73.605 114.755 -73.275 115.085 ;
        RECT -73.605 113.395 -73.275 113.725 ;
        RECT -73.605 112.035 -73.275 112.365 ;
        RECT -73.605 110.675 -73.275 111.005 ;
        RECT -73.605 109.315 -73.275 109.645 ;
        RECT -73.605 107.955 -73.275 108.285 ;
        RECT -73.605 106.595 -73.275 106.925 ;
        RECT -73.605 105.235 -73.275 105.565 ;
        RECT -73.605 103.875 -73.275 104.205 ;
        RECT -73.605 102.515 -73.275 102.845 ;
        RECT -73.605 101.155 -73.275 101.485 ;
        RECT -73.605 99.795 -73.275 100.125 ;
        RECT -73.605 98.435 -73.275 98.765 ;
        RECT -73.605 97.075 -73.275 97.405 ;
        RECT -73.605 95.715 -73.275 96.045 ;
        RECT -73.605 94.355 -73.275 94.685 ;
        RECT -73.605 92.995 -73.275 93.325 ;
        RECT -73.605 91.635 -73.275 91.965 ;
        RECT -73.605 90.275 -73.275 90.605 ;
        RECT -73.605 88.915 -73.275 89.245 ;
        RECT -73.605 87.555 -73.275 87.885 ;
        RECT -73.605 86.195 -73.275 86.525 ;
        RECT -73.605 84.835 -73.275 85.165 ;
        RECT -73.605 83.475 -73.275 83.805 ;
        RECT -73.605 82.115 -73.275 82.445 ;
        RECT -73.605 80.755 -73.275 81.085 ;
        RECT -73.605 79.395 -73.275 79.725 ;
        RECT -73.605 78.035 -73.275 78.365 ;
        RECT -73.605 76.675 -73.275 77.005 ;
        RECT -73.605 75.315 -73.275 75.645 ;
        RECT -73.605 73.955 -73.275 74.285 ;
        RECT -73.605 72.595 -73.275 72.925 ;
        RECT -73.605 71.235 -73.275 71.565 ;
        RECT -73.605 69.875 -73.275 70.205 ;
        RECT -73.605 68.515 -73.275 68.845 ;
        RECT -73.605 67.155 -73.275 67.485 ;
        RECT -73.605 65.795 -73.275 66.125 ;
        RECT -73.605 64.435 -73.275 64.765 ;
        RECT -73.605 63.075 -73.275 63.405 ;
        RECT -73.605 61.715 -73.275 62.045 ;
        RECT -73.605 60.355 -73.275 60.685 ;
        RECT -73.605 58.995 -73.275 59.325 ;
        RECT -73.605 57.635 -73.275 57.965 ;
        RECT -73.605 56.275 -73.275 56.605 ;
        RECT -73.605 54.915 -73.275 55.245 ;
        RECT -73.605 53.555 -73.275 53.885 ;
        RECT -73.605 52.195 -73.275 52.525 ;
        RECT -73.605 50.835 -73.275 51.165 ;
        RECT -73.605 49.475 -73.275 49.805 ;
        RECT -73.605 48.115 -73.275 48.445 ;
        RECT -73.605 46.755 -73.275 47.085 ;
        RECT -73.605 45.395 -73.275 45.725 ;
        RECT -73.605 44.035 -73.275 44.365 ;
        RECT -73.605 42.675 -73.275 43.005 ;
        RECT -73.605 41.315 -73.275 41.645 ;
        RECT -73.605 39.955 -73.275 40.285 ;
        RECT -73.605 38.595 -73.275 38.925 ;
        RECT -73.605 37.235 -73.275 37.565 ;
        RECT -73.605 35.875 -73.275 36.205 ;
        RECT -73.605 34.515 -73.275 34.845 ;
        RECT -73.605 33.155 -73.275 33.485 ;
        RECT -73.605 31.795 -73.275 32.125 ;
        RECT -73.605 30.435 -73.275 30.765 ;
        RECT -73.605 29.075 -73.275 29.405 ;
        RECT -73.605 27.715 -73.275 28.045 ;
        RECT -73.605 26.355 -73.275 26.685 ;
        RECT -73.605 24.995 -73.275 25.325 ;
        RECT -73.605 23.635 -73.275 23.965 ;
        RECT -73.605 22.275 -73.275 22.605 ;
        RECT -73.605 20.915 -73.275 21.245 ;
        RECT -73.605 19.555 -73.275 19.885 ;
        RECT -73.605 18.195 -73.275 18.525 ;
        RECT -73.605 16.835 -73.275 17.165 ;
        RECT -73.605 15.475 -73.275 15.805 ;
        RECT -73.605 14.115 -73.275 14.445 ;
        RECT -73.605 12.755 -73.275 13.085 ;
        RECT -73.605 11.395 -73.275 11.725 ;
        RECT -73.605 10.035 -73.275 10.365 ;
        RECT -73.605 8.675 -73.275 9.005 ;
        RECT -73.605 7.315 -73.275 7.645 ;
        RECT -73.605 5.955 -73.275 6.285 ;
        RECT -73.605 4.595 -73.275 4.925 ;
        RECT -73.605 3.235 -73.275 3.565 ;
        RECT -73.605 1.875 -73.275 2.205 ;
        RECT -73.605 0.515 -73.275 0.845 ;
        RECT -73.605 -0.845 -73.275 -0.515 ;
        RECT -73.605 -2.205 -73.275 -1.875 ;
        RECT -73.605 -3.565 -73.275 -3.235 ;
        RECT -73.605 -4.925 -73.275 -4.595 ;
        RECT -73.605 -6.285 -73.275 -5.955 ;
        RECT -73.605 -7.645 -73.275 -7.315 ;
        RECT -73.605 -9.005 -73.275 -8.675 ;
        RECT -73.605 -10.365 -73.275 -10.035 ;
        RECT -73.605 -11.725 -73.275 -11.395 ;
        RECT -73.605 -13.085 -73.275 -12.755 ;
        RECT -73.605 -14.445 -73.275 -14.115 ;
        RECT -73.605 -15.805 -73.275 -15.475 ;
        RECT -73.605 -17.165 -73.275 -16.835 ;
        RECT -73.605 -18.525 -73.275 -18.195 ;
        RECT -73.605 -19.885 -73.275 -19.555 ;
        RECT -73.605 -21.245 -73.275 -20.915 ;
        RECT -73.605 -22.605 -73.275 -22.275 ;
        RECT -73.605 -23.965 -73.275 -23.635 ;
        RECT -73.605 -25.325 -73.275 -24.995 ;
        RECT -73.605 -26.685 -73.275 -26.355 ;
        RECT -73.605 -28.045 -73.275 -27.715 ;
        RECT -73.605 -29.405 -73.275 -29.075 ;
        RECT -73.605 -30.765 -73.275 -30.435 ;
        RECT -73.605 -32.125 -73.275 -31.795 ;
        RECT -73.605 -33.485 -73.275 -33.155 ;
        RECT -73.605 -34.845 -73.275 -34.515 ;
        RECT -73.605 -36.205 -73.275 -35.875 ;
        RECT -73.605 -37.565 -73.275 -37.235 ;
        RECT -73.605 -38.925 -73.275 -38.595 ;
        RECT -73.605 -40.285 -73.275 -39.955 ;
        RECT -73.605 -41.645 -73.275 -41.315 ;
        RECT -73.605 -43.005 -73.275 -42.675 ;
        RECT -73.605 -44.365 -73.275 -44.035 ;
        RECT -73.605 -45.725 -73.275 -45.395 ;
        RECT -73.605 -47.085 -73.275 -46.755 ;
        RECT -73.605 -48.445 -73.275 -48.115 ;
        RECT -73.605 -49.805 -73.275 -49.475 ;
        RECT -73.605 -51.165 -73.275 -50.835 ;
        RECT -73.605 -52.525 -73.275 -52.195 ;
        RECT -73.605 -53.885 -73.275 -53.555 ;
        RECT -73.605 -55.245 -73.275 -54.915 ;
        RECT -73.605 -56.605 -73.275 -56.275 ;
        RECT -73.605 -57.965 -73.275 -57.635 ;
        RECT -73.605 -59.325 -73.275 -58.995 ;
        RECT -73.605 -60.685 -73.275 -60.355 ;
        RECT -73.605 -62.045 -73.275 -61.715 ;
        RECT -73.605 -63.405 -73.275 -63.075 ;
        RECT -73.605 -64.765 -73.275 -64.435 ;
        RECT -73.605 -66.125 -73.275 -65.795 ;
        RECT -73.605 -67.485 -73.275 -67.155 ;
        RECT -73.605 -68.845 -73.275 -68.515 ;
        RECT -73.605 -70.205 -73.275 -69.875 ;
        RECT -73.605 -71.565 -73.275 -71.235 ;
        RECT -73.605 -72.925 -73.275 -72.595 ;
        RECT -73.605 -74.285 -73.275 -73.955 ;
        RECT -73.605 -75.645 -73.275 -75.315 ;
        RECT -73.605 -77.005 -73.275 -76.675 ;
        RECT -73.605 -78.365 -73.275 -78.035 ;
        RECT -73.605 -79.725 -73.275 -79.395 ;
        RECT -73.605 -81.085 -73.275 -80.755 ;
        RECT -73.605 -82.445 -73.275 -82.115 ;
        RECT -73.605 -83.805 -73.275 -83.475 ;
        RECT -73.605 -85.165 -73.275 -84.835 ;
        RECT -73.605 -86.525 -73.275 -86.195 ;
        RECT -73.605 -87.885 -73.275 -87.555 ;
        RECT -73.605 -89.245 -73.275 -88.915 ;
        RECT -73.605 -90.605 -73.275 -90.275 ;
        RECT -73.605 -91.965 -73.275 -91.635 ;
        RECT -73.605 -93.325 -73.275 -92.995 ;
        RECT -73.605 -94.685 -73.275 -94.355 ;
        RECT -73.605 -96.045 -73.275 -95.715 ;
        RECT -73.605 -97.405 -73.275 -97.075 ;
        RECT -73.605 -98.765 -73.275 -98.435 ;
        RECT -73.605 -100.125 -73.275 -99.795 ;
        RECT -73.605 -101.485 -73.275 -101.155 ;
        RECT -73.605 -102.845 -73.275 -102.515 ;
        RECT -73.605 -104.205 -73.275 -103.875 ;
        RECT -73.605 -105.565 -73.275 -105.235 ;
        RECT -73.605 -106.925 -73.275 -106.595 ;
        RECT -73.605 -108.285 -73.275 -107.955 ;
        RECT -73.605 -109.645 -73.275 -109.315 ;
        RECT -73.605 -111.005 -73.275 -110.675 ;
        RECT -73.605 -112.365 -73.275 -112.035 ;
        RECT -73.605 -113.725 -73.275 -113.395 ;
        RECT -73.605 -115.085 -73.275 -114.755 ;
        RECT -73.605 -116.445 -73.275 -116.115 ;
        RECT -73.605 -117.805 -73.275 -117.475 ;
        RECT -73.605 -119.165 -73.275 -118.835 ;
        RECT -73.605 -120.525 -73.275 -120.195 ;
        RECT -73.605 -121.885 -73.275 -121.555 ;
        RECT -73.605 -123.245 -73.275 -122.915 ;
        RECT -73.605 -124.605 -73.275 -124.275 ;
        RECT -73.605 -125.965 -73.275 -125.635 ;
        RECT -73.605 -127.325 -73.275 -126.995 ;
        RECT -73.605 -128.685 -73.275 -128.355 ;
        RECT -73.605 -130.045 -73.275 -129.715 ;
        RECT -73.605 -131.405 -73.275 -131.075 ;
        RECT -73.605 -132.765 -73.275 -132.435 ;
        RECT -73.605 -134.125 -73.275 -133.795 ;
        RECT -73.605 -135.485 -73.275 -135.155 ;
        RECT -73.605 -136.845 -73.275 -136.515 ;
        RECT -73.605 -138.205 -73.275 -137.875 ;
        RECT -73.605 -139.565 -73.275 -139.235 ;
        RECT -73.605 -140.925 -73.275 -140.595 ;
        RECT -73.605 -142.285 -73.275 -141.955 ;
        RECT -73.605 -143.645 -73.275 -143.315 ;
        RECT -73.605 -145.005 -73.275 -144.675 ;
        RECT -73.605 -146.365 -73.275 -146.035 ;
        RECT -73.605 -147.725 -73.275 -147.395 ;
        RECT -73.605 -149.085 -73.275 -148.755 ;
        RECT -73.605 -150.445 -73.275 -150.115 ;
        RECT -73.605 -151.805 -73.275 -151.475 ;
        RECT -73.605 -153.165 -73.275 -152.835 ;
        RECT -73.605 -154.525 -73.275 -154.195 ;
        RECT -73.605 -155.885 -73.275 -155.555 ;
        RECT -73.605 -157.245 -73.275 -156.915 ;
        RECT -73.605 -158.605 -73.275 -158.275 ;
        RECT -73.605 -159.965 -73.275 -159.635 ;
        RECT -73.605 -161.325 -73.275 -160.995 ;
        RECT -73.605 -162.685 -73.275 -162.355 ;
        RECT -73.605 -164.045 -73.275 -163.715 ;
        RECT -73.605 -165.405 -73.275 -165.075 ;
        RECT -73.605 -166.765 -73.275 -166.435 ;
        RECT -73.6 -167.44 -73.28 245.285 ;
        RECT -73.605 244.04 -73.275 245.17 ;
        RECT -73.605 239.875 -73.275 240.205 ;
        RECT -73.605 238.515 -73.275 238.845 ;
        RECT -73.605 237.155 -73.275 237.485 ;
        RECT -73.605 235.795 -73.275 236.125 ;
        RECT -73.605 234.435 -73.275 234.765 ;
        RECT -73.605 233.075 -73.275 233.405 ;
        RECT -73.605 231.715 -73.275 232.045 ;
        RECT -73.605 230.355 -73.275 230.685 ;
        RECT -73.605 228.995 -73.275 229.325 ;
        RECT -73.605 227.635 -73.275 227.965 ;
        RECT -73.605 226.275 -73.275 226.605 ;
        RECT -73.605 224.915 -73.275 225.245 ;
        RECT -73.605 223.555 -73.275 223.885 ;
        RECT -73.605 222.195 -73.275 222.525 ;
        RECT -73.605 220.835 -73.275 221.165 ;
        RECT -73.605 219.475 -73.275 219.805 ;
        RECT -73.605 218.115 -73.275 218.445 ;
        RECT -73.605 216.755 -73.275 217.085 ;
        RECT -73.605 215.395 -73.275 215.725 ;
        RECT -73.605 214.035 -73.275 214.365 ;
        RECT -73.605 212.675 -73.275 213.005 ;
        RECT -73.605 211.315 -73.275 211.645 ;
        RECT -73.605 209.955 -73.275 210.285 ;
        RECT -73.605 208.595 -73.275 208.925 ;
        RECT -73.605 207.235 -73.275 207.565 ;
        RECT -73.605 205.875 -73.275 206.205 ;
        RECT -73.605 204.515 -73.275 204.845 ;
        RECT -73.605 203.155 -73.275 203.485 ;
        RECT -73.605 201.795 -73.275 202.125 ;
    END
    PORT
      LAYER met3 ;
        RECT -80.405 244.04 -80.075 245.17 ;
        RECT -80.405 239.875 -80.075 240.205 ;
        RECT -80.405 238.515 -80.075 238.845 ;
        RECT -80.405 237.155 -80.075 237.485 ;
        RECT -80.405 235.795 -80.075 236.125 ;
        RECT -80.405 234.435 -80.075 234.765 ;
        RECT -80.405 233.075 -80.075 233.405 ;
        RECT -80.405 231.715 -80.075 232.045 ;
        RECT -80.405 230.355 -80.075 230.685 ;
        RECT -80.405 228.995 -80.075 229.325 ;
        RECT -80.405 227.635 -80.075 227.965 ;
        RECT -80.405 226.275 -80.075 226.605 ;
        RECT -80.405 224.915 -80.075 225.245 ;
        RECT -80.405 223.555 -80.075 223.885 ;
        RECT -80.405 222.195 -80.075 222.525 ;
        RECT -80.405 220.835 -80.075 221.165 ;
        RECT -80.405 219.475 -80.075 219.805 ;
        RECT -80.405 218.115 -80.075 218.445 ;
        RECT -80.405 216.755 -80.075 217.085 ;
        RECT -80.405 215.395 -80.075 215.725 ;
        RECT -80.405 214.035 -80.075 214.365 ;
        RECT -80.405 212.675 -80.075 213.005 ;
        RECT -80.405 211.315 -80.075 211.645 ;
        RECT -80.405 209.955 -80.075 210.285 ;
        RECT -80.405 208.595 -80.075 208.925 ;
        RECT -80.405 207.235 -80.075 207.565 ;
        RECT -80.405 205.875 -80.075 206.205 ;
        RECT -80.405 204.515 -80.075 204.845 ;
        RECT -80.405 203.155 -80.075 203.485 ;
        RECT -80.405 201.795 -80.075 202.125 ;
        RECT -80.405 200.435 -80.075 200.765 ;
        RECT -80.405 199.075 -80.075 199.405 ;
        RECT -80.405 197.715 -80.075 198.045 ;
        RECT -80.405 196.355 -80.075 196.685 ;
        RECT -80.405 194.995 -80.075 195.325 ;
        RECT -80.405 193.635 -80.075 193.965 ;
        RECT -80.405 192.275 -80.075 192.605 ;
        RECT -80.405 190.915 -80.075 191.245 ;
        RECT -80.405 189.555 -80.075 189.885 ;
        RECT -80.405 188.195 -80.075 188.525 ;
        RECT -80.405 186.835 -80.075 187.165 ;
        RECT -80.405 185.475 -80.075 185.805 ;
        RECT -80.405 184.115 -80.075 184.445 ;
        RECT -80.405 182.755 -80.075 183.085 ;
        RECT -80.405 181.395 -80.075 181.725 ;
        RECT -80.405 180.035 -80.075 180.365 ;
        RECT -80.405 178.675 -80.075 179.005 ;
        RECT -80.405 177.315 -80.075 177.645 ;
        RECT -80.405 175.955 -80.075 176.285 ;
        RECT -80.405 174.595 -80.075 174.925 ;
        RECT -80.405 173.235 -80.075 173.565 ;
        RECT -80.405 171.875 -80.075 172.205 ;
        RECT -80.405 170.515 -80.075 170.845 ;
        RECT -80.405 169.155 -80.075 169.485 ;
        RECT -80.405 167.795 -80.075 168.125 ;
        RECT -80.405 166.435 -80.075 166.765 ;
        RECT -80.405 165.075 -80.075 165.405 ;
        RECT -80.405 163.715 -80.075 164.045 ;
        RECT -80.405 162.355 -80.075 162.685 ;
        RECT -80.405 160.995 -80.075 161.325 ;
        RECT -80.405 159.635 -80.075 159.965 ;
        RECT -80.405 158.275 -80.075 158.605 ;
        RECT -80.405 156.915 -80.075 157.245 ;
        RECT -80.405 155.555 -80.075 155.885 ;
        RECT -80.405 154.195 -80.075 154.525 ;
        RECT -80.405 152.835 -80.075 153.165 ;
        RECT -80.405 151.475 -80.075 151.805 ;
        RECT -80.405 150.115 -80.075 150.445 ;
        RECT -80.405 148.755 -80.075 149.085 ;
        RECT -80.405 147.395 -80.075 147.725 ;
        RECT -80.405 146.035 -80.075 146.365 ;
        RECT -80.405 144.675 -80.075 145.005 ;
        RECT -80.405 143.315 -80.075 143.645 ;
        RECT -80.405 141.955 -80.075 142.285 ;
        RECT -80.405 140.595 -80.075 140.925 ;
        RECT -80.405 139.235 -80.075 139.565 ;
        RECT -80.405 137.875 -80.075 138.205 ;
        RECT -80.405 136.515 -80.075 136.845 ;
        RECT -80.405 135.155 -80.075 135.485 ;
        RECT -80.405 133.795 -80.075 134.125 ;
        RECT -80.405 132.435 -80.075 132.765 ;
        RECT -80.405 131.075 -80.075 131.405 ;
        RECT -80.405 129.715 -80.075 130.045 ;
        RECT -80.405 128.355 -80.075 128.685 ;
        RECT -80.405 126.995 -80.075 127.325 ;
        RECT -80.405 125.635 -80.075 125.965 ;
        RECT -80.405 124.275 -80.075 124.605 ;
        RECT -80.405 122.915 -80.075 123.245 ;
        RECT -80.405 121.555 -80.075 121.885 ;
        RECT -80.405 120.195 -80.075 120.525 ;
        RECT -80.405 118.835 -80.075 119.165 ;
        RECT -80.405 117.475 -80.075 117.805 ;
        RECT -80.405 116.115 -80.075 116.445 ;
        RECT -80.405 114.755 -80.075 115.085 ;
        RECT -80.405 113.395 -80.075 113.725 ;
        RECT -80.405 112.035 -80.075 112.365 ;
        RECT -80.405 110.675 -80.075 111.005 ;
        RECT -80.405 109.315 -80.075 109.645 ;
        RECT -80.405 107.955 -80.075 108.285 ;
        RECT -80.405 106.595 -80.075 106.925 ;
        RECT -80.405 105.235 -80.075 105.565 ;
        RECT -80.405 103.875 -80.075 104.205 ;
        RECT -80.405 102.515 -80.075 102.845 ;
        RECT -80.405 101.155 -80.075 101.485 ;
        RECT -80.405 99.795 -80.075 100.125 ;
        RECT -80.405 98.435 -80.075 98.765 ;
        RECT -80.405 97.075 -80.075 97.405 ;
        RECT -80.405 95.715 -80.075 96.045 ;
        RECT -80.405 94.355 -80.075 94.685 ;
        RECT -80.405 92.995 -80.075 93.325 ;
        RECT -80.405 91.635 -80.075 91.965 ;
        RECT -80.405 90.275 -80.075 90.605 ;
        RECT -80.405 88.915 -80.075 89.245 ;
        RECT -80.405 87.555 -80.075 87.885 ;
        RECT -80.405 86.195 -80.075 86.525 ;
        RECT -80.405 84.835 -80.075 85.165 ;
        RECT -80.405 83.475 -80.075 83.805 ;
        RECT -80.405 82.115 -80.075 82.445 ;
        RECT -80.405 80.755 -80.075 81.085 ;
        RECT -80.405 79.395 -80.075 79.725 ;
        RECT -80.405 78.035 -80.075 78.365 ;
        RECT -80.405 76.675 -80.075 77.005 ;
        RECT -80.405 75.315 -80.075 75.645 ;
        RECT -80.405 73.955 -80.075 74.285 ;
        RECT -80.405 72.595 -80.075 72.925 ;
        RECT -80.405 71.235 -80.075 71.565 ;
        RECT -80.405 69.875 -80.075 70.205 ;
        RECT -80.405 68.515 -80.075 68.845 ;
        RECT -80.405 67.155 -80.075 67.485 ;
        RECT -80.405 65.795 -80.075 66.125 ;
        RECT -80.405 64.435 -80.075 64.765 ;
        RECT -80.405 63.075 -80.075 63.405 ;
        RECT -80.405 61.715 -80.075 62.045 ;
        RECT -80.405 60.355 -80.075 60.685 ;
        RECT -80.405 58.995 -80.075 59.325 ;
        RECT -80.405 57.635 -80.075 57.965 ;
        RECT -80.405 56.275 -80.075 56.605 ;
        RECT -80.405 54.915 -80.075 55.245 ;
        RECT -80.405 53.555 -80.075 53.885 ;
        RECT -80.405 52.195 -80.075 52.525 ;
        RECT -80.405 50.835 -80.075 51.165 ;
        RECT -80.405 49.475 -80.075 49.805 ;
        RECT -80.405 48.115 -80.075 48.445 ;
        RECT -80.405 46.755 -80.075 47.085 ;
        RECT -80.405 45.395 -80.075 45.725 ;
        RECT -80.405 44.035 -80.075 44.365 ;
        RECT -80.405 42.675 -80.075 43.005 ;
        RECT -80.405 41.315 -80.075 41.645 ;
        RECT -80.405 39.955 -80.075 40.285 ;
        RECT -80.405 38.595 -80.075 38.925 ;
        RECT -80.405 37.235 -80.075 37.565 ;
        RECT -80.405 35.875 -80.075 36.205 ;
        RECT -80.405 34.515 -80.075 34.845 ;
        RECT -80.405 33.155 -80.075 33.485 ;
        RECT -80.405 31.795 -80.075 32.125 ;
        RECT -80.405 30.435 -80.075 30.765 ;
        RECT -80.405 29.075 -80.075 29.405 ;
        RECT -80.405 27.715 -80.075 28.045 ;
        RECT -80.405 26.355 -80.075 26.685 ;
        RECT -80.405 24.995 -80.075 25.325 ;
        RECT -80.405 23.635 -80.075 23.965 ;
        RECT -80.405 22.275 -80.075 22.605 ;
        RECT -80.405 20.915 -80.075 21.245 ;
        RECT -80.405 19.555 -80.075 19.885 ;
        RECT -80.405 18.195 -80.075 18.525 ;
        RECT -80.405 16.835 -80.075 17.165 ;
        RECT -80.405 15.475 -80.075 15.805 ;
        RECT -80.405 14.115 -80.075 14.445 ;
        RECT -80.405 12.755 -80.075 13.085 ;
        RECT -80.405 11.395 -80.075 11.725 ;
        RECT -80.405 10.035 -80.075 10.365 ;
        RECT -80.405 8.675 -80.075 9.005 ;
        RECT -80.405 7.315 -80.075 7.645 ;
        RECT -80.405 5.955 -80.075 6.285 ;
        RECT -80.405 4.595 -80.075 4.925 ;
        RECT -80.405 3.235 -80.075 3.565 ;
        RECT -80.405 1.875 -80.075 2.205 ;
        RECT -80.405 0.515 -80.075 0.845 ;
        RECT -80.405 -0.845 -80.075 -0.515 ;
        RECT -80.405 -2.205 -80.075 -1.875 ;
        RECT -80.405 -3.565 -80.075 -3.235 ;
        RECT -80.405 -4.925 -80.075 -4.595 ;
        RECT -80.405 -6.285 -80.075 -5.955 ;
        RECT -80.405 -7.645 -80.075 -7.315 ;
        RECT -80.405 -9.005 -80.075 -8.675 ;
        RECT -80.405 -10.365 -80.075 -10.035 ;
        RECT -80.405 -11.725 -80.075 -11.395 ;
        RECT -80.405 -13.085 -80.075 -12.755 ;
        RECT -80.405 -14.445 -80.075 -14.115 ;
        RECT -80.405 -15.805 -80.075 -15.475 ;
        RECT -80.405 -17.165 -80.075 -16.835 ;
        RECT -80.405 -18.525 -80.075 -18.195 ;
        RECT -80.405 -19.885 -80.075 -19.555 ;
        RECT -80.405 -21.245 -80.075 -20.915 ;
        RECT -80.405 -22.605 -80.075 -22.275 ;
        RECT -80.405 -23.965 -80.075 -23.635 ;
        RECT -80.405 -25.325 -80.075 -24.995 ;
        RECT -80.405 -26.685 -80.075 -26.355 ;
        RECT -80.405 -28.045 -80.075 -27.715 ;
        RECT -80.405 -29.405 -80.075 -29.075 ;
        RECT -80.405 -30.765 -80.075 -30.435 ;
        RECT -80.405 -32.125 -80.075 -31.795 ;
        RECT -80.405 -33.485 -80.075 -33.155 ;
        RECT -80.405 -34.845 -80.075 -34.515 ;
        RECT -80.405 -36.205 -80.075 -35.875 ;
        RECT -80.405 -37.565 -80.075 -37.235 ;
        RECT -80.405 -38.925 -80.075 -38.595 ;
        RECT -80.405 -40.285 -80.075 -39.955 ;
        RECT -80.405 -41.645 -80.075 -41.315 ;
        RECT -80.405 -43.005 -80.075 -42.675 ;
        RECT -80.405 -44.365 -80.075 -44.035 ;
        RECT -80.405 -45.725 -80.075 -45.395 ;
        RECT -80.405 -47.085 -80.075 -46.755 ;
        RECT -80.405 -48.445 -80.075 -48.115 ;
        RECT -80.405 -49.805 -80.075 -49.475 ;
        RECT -80.405 -51.165 -80.075 -50.835 ;
        RECT -80.405 -52.525 -80.075 -52.195 ;
        RECT -80.405 -53.885 -80.075 -53.555 ;
        RECT -80.405 -55.245 -80.075 -54.915 ;
        RECT -80.405 -56.605 -80.075 -56.275 ;
        RECT -80.405 -57.965 -80.075 -57.635 ;
        RECT -80.405 -59.325 -80.075 -58.995 ;
        RECT -80.405 -60.685 -80.075 -60.355 ;
        RECT -80.405 -62.045 -80.075 -61.715 ;
        RECT -80.405 -63.405 -80.075 -63.075 ;
        RECT -80.405 -64.765 -80.075 -64.435 ;
        RECT -80.405 -66.125 -80.075 -65.795 ;
        RECT -80.405 -67.485 -80.075 -67.155 ;
        RECT -80.405 -68.845 -80.075 -68.515 ;
        RECT -80.405 -70.205 -80.075 -69.875 ;
        RECT -80.405 -71.565 -80.075 -71.235 ;
        RECT -80.405 -72.925 -80.075 -72.595 ;
        RECT -80.405 -74.285 -80.075 -73.955 ;
        RECT -80.405 -75.645 -80.075 -75.315 ;
        RECT -80.405 -77.005 -80.075 -76.675 ;
        RECT -80.405 -78.365 -80.075 -78.035 ;
        RECT -80.405 -79.725 -80.075 -79.395 ;
        RECT -80.405 -81.085 -80.075 -80.755 ;
        RECT -80.405 -82.445 -80.075 -82.115 ;
        RECT -80.405 -83.805 -80.075 -83.475 ;
        RECT -80.405 -85.165 -80.075 -84.835 ;
        RECT -80.405 -86.525 -80.075 -86.195 ;
        RECT -80.405 -87.885 -80.075 -87.555 ;
        RECT -80.405 -89.245 -80.075 -88.915 ;
        RECT -80.405 -90.605 -80.075 -90.275 ;
        RECT -80.405 -91.965 -80.075 -91.635 ;
        RECT -80.405 -93.325 -80.075 -92.995 ;
        RECT -80.405 -94.685 -80.075 -94.355 ;
        RECT -80.405 -96.045 -80.075 -95.715 ;
        RECT -80.405 -97.405 -80.075 -97.075 ;
        RECT -80.405 -98.765 -80.075 -98.435 ;
        RECT -80.405 -100.125 -80.075 -99.795 ;
        RECT -80.405 -101.485 -80.075 -101.155 ;
        RECT -80.405 -102.845 -80.075 -102.515 ;
        RECT -80.405 -104.205 -80.075 -103.875 ;
        RECT -80.405 -105.565 -80.075 -105.235 ;
        RECT -80.405 -106.925 -80.075 -106.595 ;
        RECT -80.405 -108.285 -80.075 -107.955 ;
        RECT -80.405 -109.645 -80.075 -109.315 ;
        RECT -80.405 -111.005 -80.075 -110.675 ;
        RECT -80.405 -112.365 -80.075 -112.035 ;
        RECT -80.405 -113.725 -80.075 -113.395 ;
        RECT -80.405 -115.085 -80.075 -114.755 ;
        RECT -80.405 -116.445 -80.075 -116.115 ;
        RECT -80.405 -117.805 -80.075 -117.475 ;
        RECT -80.405 -119.165 -80.075 -118.835 ;
        RECT -80.405 -120.525 -80.075 -120.195 ;
        RECT -80.405 -121.885 -80.075 -121.555 ;
        RECT -80.405 -123.245 -80.075 -122.915 ;
        RECT -80.405 -124.605 -80.075 -124.275 ;
        RECT -80.405 -125.965 -80.075 -125.635 ;
        RECT -80.405 -127.325 -80.075 -126.995 ;
        RECT -80.405 -128.685 -80.075 -128.355 ;
        RECT -80.405 -130.045 -80.075 -129.715 ;
        RECT -80.405 -131.405 -80.075 -131.075 ;
        RECT -80.405 -132.765 -80.075 -132.435 ;
        RECT -80.405 -134.125 -80.075 -133.795 ;
        RECT -80.405 -135.485 -80.075 -135.155 ;
        RECT -80.405 -136.845 -80.075 -136.515 ;
        RECT -80.405 -138.205 -80.075 -137.875 ;
        RECT -80.405 -139.565 -80.075 -139.235 ;
        RECT -80.405 -140.925 -80.075 -140.595 ;
        RECT -80.405 -142.285 -80.075 -141.955 ;
        RECT -80.405 -143.645 -80.075 -143.315 ;
        RECT -80.405 -145.005 -80.075 -144.675 ;
        RECT -80.405 -146.365 -80.075 -146.035 ;
        RECT -80.405 -147.725 -80.075 -147.395 ;
        RECT -80.405 -149.085 -80.075 -148.755 ;
        RECT -80.405 -150.445 -80.075 -150.115 ;
        RECT -80.405 -151.805 -80.075 -151.475 ;
        RECT -80.405 -153.165 -80.075 -152.835 ;
        RECT -80.405 -154.525 -80.075 -154.195 ;
        RECT -80.405 -155.885 -80.075 -155.555 ;
        RECT -80.405 -157.245 -80.075 -156.915 ;
        RECT -80.405 -158.605 -80.075 -158.275 ;
        RECT -80.405 -159.965 -80.075 -159.635 ;
        RECT -80.405 -161.325 -80.075 -160.995 ;
        RECT -80.405 -162.685 -80.075 -162.355 ;
        RECT -80.405 -164.045 -80.075 -163.715 ;
        RECT -80.405 -165.405 -80.075 -165.075 ;
        RECT -80.405 -166.765 -80.075 -166.435 ;
        RECT -80.405 -168.125 -80.075 -167.795 ;
        RECT -80.405 -169.485 -80.075 -169.155 ;
        RECT -80.405 -170.845 -80.075 -170.515 ;
        RECT -80.405 -172.205 -80.075 -171.875 ;
        RECT -80.405 -173.565 -80.075 -173.235 ;
        RECT -80.405 -174.925 -80.075 -174.595 ;
        RECT -80.405 -176.285 -80.075 -175.955 ;
        RECT -80.405 -177.645 -80.075 -177.315 ;
        RECT -80.405 -179.005 -80.075 -178.675 ;
        RECT -80.405 -184.65 -80.075 -183.52 ;
        RECT -80.4 -184.765 -80.08 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -79.045 244.04 -78.715 245.17 ;
        RECT -79.045 239.875 -78.715 240.205 ;
        RECT -79.045 238.515 -78.715 238.845 ;
        RECT -79.045 237.155 -78.715 237.485 ;
        RECT -79.045 235.795 -78.715 236.125 ;
        RECT -79.045 234.435 -78.715 234.765 ;
        RECT -79.045 233.075 -78.715 233.405 ;
        RECT -79.045 231.715 -78.715 232.045 ;
        RECT -79.045 230.355 -78.715 230.685 ;
        RECT -79.045 228.995 -78.715 229.325 ;
        RECT -79.045 227.635 -78.715 227.965 ;
        RECT -79.045 226.275 -78.715 226.605 ;
        RECT -79.045 224.915 -78.715 225.245 ;
        RECT -79.045 223.555 -78.715 223.885 ;
        RECT -79.045 222.195 -78.715 222.525 ;
        RECT -79.045 220.835 -78.715 221.165 ;
        RECT -79.045 219.475 -78.715 219.805 ;
        RECT -79.045 218.115 -78.715 218.445 ;
        RECT -79.045 216.755 -78.715 217.085 ;
        RECT -79.045 215.395 -78.715 215.725 ;
        RECT -79.045 214.035 -78.715 214.365 ;
        RECT -79.045 212.675 -78.715 213.005 ;
        RECT -79.045 211.315 -78.715 211.645 ;
        RECT -79.045 209.955 -78.715 210.285 ;
        RECT -79.045 208.595 -78.715 208.925 ;
        RECT -79.045 207.235 -78.715 207.565 ;
        RECT -79.045 205.875 -78.715 206.205 ;
        RECT -79.045 204.515 -78.715 204.845 ;
        RECT -79.045 203.155 -78.715 203.485 ;
        RECT -79.045 201.795 -78.715 202.125 ;
        RECT -79.045 200.435 -78.715 200.765 ;
        RECT -79.045 199.075 -78.715 199.405 ;
        RECT -79.045 197.715 -78.715 198.045 ;
        RECT -79.045 196.355 -78.715 196.685 ;
        RECT -79.045 194.995 -78.715 195.325 ;
        RECT -79.045 193.635 -78.715 193.965 ;
        RECT -79.045 192.275 -78.715 192.605 ;
        RECT -79.045 190.915 -78.715 191.245 ;
        RECT -79.045 189.555 -78.715 189.885 ;
        RECT -79.045 188.195 -78.715 188.525 ;
        RECT -79.045 186.835 -78.715 187.165 ;
        RECT -79.045 185.475 -78.715 185.805 ;
        RECT -79.045 184.115 -78.715 184.445 ;
        RECT -79.045 182.755 -78.715 183.085 ;
        RECT -79.045 181.395 -78.715 181.725 ;
        RECT -79.045 180.035 -78.715 180.365 ;
        RECT -79.045 178.675 -78.715 179.005 ;
        RECT -79.045 177.315 -78.715 177.645 ;
        RECT -79.045 175.955 -78.715 176.285 ;
        RECT -79.045 174.595 -78.715 174.925 ;
        RECT -79.045 173.235 -78.715 173.565 ;
        RECT -79.045 171.875 -78.715 172.205 ;
        RECT -79.045 170.515 -78.715 170.845 ;
        RECT -79.045 169.155 -78.715 169.485 ;
        RECT -79.045 167.795 -78.715 168.125 ;
        RECT -79.045 166.435 -78.715 166.765 ;
        RECT -79.045 165.075 -78.715 165.405 ;
        RECT -79.045 163.715 -78.715 164.045 ;
        RECT -79.045 162.355 -78.715 162.685 ;
        RECT -79.045 160.995 -78.715 161.325 ;
        RECT -79.045 159.635 -78.715 159.965 ;
        RECT -79.045 158.275 -78.715 158.605 ;
        RECT -79.045 156.915 -78.715 157.245 ;
        RECT -79.045 155.555 -78.715 155.885 ;
        RECT -79.045 154.195 -78.715 154.525 ;
        RECT -79.045 152.835 -78.715 153.165 ;
        RECT -79.045 151.475 -78.715 151.805 ;
        RECT -79.045 150.115 -78.715 150.445 ;
        RECT -79.045 148.755 -78.715 149.085 ;
        RECT -79.045 147.395 -78.715 147.725 ;
        RECT -79.045 146.035 -78.715 146.365 ;
        RECT -79.045 144.675 -78.715 145.005 ;
        RECT -79.045 143.315 -78.715 143.645 ;
        RECT -79.045 141.955 -78.715 142.285 ;
        RECT -79.045 140.595 -78.715 140.925 ;
        RECT -79.045 139.235 -78.715 139.565 ;
        RECT -79.045 137.875 -78.715 138.205 ;
        RECT -79.045 136.515 -78.715 136.845 ;
        RECT -79.045 135.155 -78.715 135.485 ;
        RECT -79.045 133.795 -78.715 134.125 ;
        RECT -79.045 132.435 -78.715 132.765 ;
        RECT -79.045 131.075 -78.715 131.405 ;
        RECT -79.045 129.715 -78.715 130.045 ;
        RECT -79.045 128.355 -78.715 128.685 ;
        RECT -79.045 126.995 -78.715 127.325 ;
        RECT -79.045 125.635 -78.715 125.965 ;
        RECT -79.045 124.275 -78.715 124.605 ;
        RECT -79.045 122.915 -78.715 123.245 ;
        RECT -79.045 121.555 -78.715 121.885 ;
        RECT -79.045 120.195 -78.715 120.525 ;
        RECT -79.045 118.835 -78.715 119.165 ;
        RECT -79.045 117.475 -78.715 117.805 ;
        RECT -79.045 116.115 -78.715 116.445 ;
        RECT -79.045 114.755 -78.715 115.085 ;
        RECT -79.045 113.395 -78.715 113.725 ;
        RECT -79.045 112.035 -78.715 112.365 ;
        RECT -79.045 110.675 -78.715 111.005 ;
        RECT -79.045 109.315 -78.715 109.645 ;
        RECT -79.045 107.955 -78.715 108.285 ;
        RECT -79.045 106.595 -78.715 106.925 ;
        RECT -79.045 105.235 -78.715 105.565 ;
        RECT -79.045 103.875 -78.715 104.205 ;
        RECT -79.045 102.515 -78.715 102.845 ;
        RECT -79.045 101.155 -78.715 101.485 ;
        RECT -79.045 99.795 -78.715 100.125 ;
        RECT -79.045 98.435 -78.715 98.765 ;
        RECT -79.045 97.075 -78.715 97.405 ;
        RECT -79.045 95.715 -78.715 96.045 ;
        RECT -79.045 94.355 -78.715 94.685 ;
        RECT -79.045 92.995 -78.715 93.325 ;
        RECT -79.045 91.635 -78.715 91.965 ;
        RECT -79.045 90.275 -78.715 90.605 ;
        RECT -79.045 88.915 -78.715 89.245 ;
        RECT -79.045 87.555 -78.715 87.885 ;
        RECT -79.045 86.195 -78.715 86.525 ;
        RECT -79.045 84.835 -78.715 85.165 ;
        RECT -79.045 83.475 -78.715 83.805 ;
        RECT -79.045 82.115 -78.715 82.445 ;
        RECT -79.045 80.755 -78.715 81.085 ;
        RECT -79.045 79.395 -78.715 79.725 ;
        RECT -79.045 78.035 -78.715 78.365 ;
        RECT -79.045 76.675 -78.715 77.005 ;
        RECT -79.045 75.315 -78.715 75.645 ;
        RECT -79.045 73.955 -78.715 74.285 ;
        RECT -79.045 72.595 -78.715 72.925 ;
        RECT -79.045 71.235 -78.715 71.565 ;
        RECT -79.045 69.875 -78.715 70.205 ;
        RECT -79.045 68.515 -78.715 68.845 ;
        RECT -79.045 67.155 -78.715 67.485 ;
        RECT -79.045 65.795 -78.715 66.125 ;
        RECT -79.045 64.435 -78.715 64.765 ;
        RECT -79.045 63.075 -78.715 63.405 ;
        RECT -79.045 61.715 -78.715 62.045 ;
        RECT -79.045 60.355 -78.715 60.685 ;
        RECT -79.045 58.995 -78.715 59.325 ;
        RECT -79.045 57.635 -78.715 57.965 ;
        RECT -79.045 56.275 -78.715 56.605 ;
        RECT -79.045 54.915 -78.715 55.245 ;
        RECT -79.045 53.555 -78.715 53.885 ;
        RECT -79.045 52.195 -78.715 52.525 ;
        RECT -79.045 50.835 -78.715 51.165 ;
        RECT -79.045 49.475 -78.715 49.805 ;
        RECT -79.045 48.115 -78.715 48.445 ;
        RECT -79.045 46.755 -78.715 47.085 ;
        RECT -79.045 45.395 -78.715 45.725 ;
        RECT -79.045 44.035 -78.715 44.365 ;
        RECT -79.045 42.675 -78.715 43.005 ;
        RECT -79.045 41.315 -78.715 41.645 ;
        RECT -79.045 39.955 -78.715 40.285 ;
        RECT -79.045 38.595 -78.715 38.925 ;
        RECT -79.045 37.235 -78.715 37.565 ;
        RECT -79.045 35.875 -78.715 36.205 ;
        RECT -79.045 34.515 -78.715 34.845 ;
        RECT -79.045 33.155 -78.715 33.485 ;
        RECT -79.045 31.795 -78.715 32.125 ;
        RECT -79.045 30.435 -78.715 30.765 ;
        RECT -79.045 29.075 -78.715 29.405 ;
        RECT -79.045 27.715 -78.715 28.045 ;
        RECT -79.045 26.355 -78.715 26.685 ;
        RECT -79.045 24.995 -78.715 25.325 ;
        RECT -79.045 23.635 -78.715 23.965 ;
        RECT -79.045 22.275 -78.715 22.605 ;
        RECT -79.045 20.915 -78.715 21.245 ;
        RECT -79.045 19.555 -78.715 19.885 ;
        RECT -79.045 18.195 -78.715 18.525 ;
        RECT -79.045 16.835 -78.715 17.165 ;
        RECT -79.045 15.475 -78.715 15.805 ;
        RECT -79.045 14.115 -78.715 14.445 ;
        RECT -79.045 12.755 -78.715 13.085 ;
        RECT -79.045 11.395 -78.715 11.725 ;
        RECT -79.045 10.035 -78.715 10.365 ;
        RECT -79.045 8.675 -78.715 9.005 ;
        RECT -79.045 7.315 -78.715 7.645 ;
        RECT -79.045 5.955 -78.715 6.285 ;
        RECT -79.045 4.595 -78.715 4.925 ;
        RECT -79.045 3.235 -78.715 3.565 ;
        RECT -79.045 1.875 -78.715 2.205 ;
        RECT -79.045 0.515 -78.715 0.845 ;
        RECT -79.045 -0.845 -78.715 -0.515 ;
        RECT -79.045 -2.205 -78.715 -1.875 ;
        RECT -79.045 -3.565 -78.715 -3.235 ;
        RECT -79.045 -4.925 -78.715 -4.595 ;
        RECT -79.045 -6.285 -78.715 -5.955 ;
        RECT -79.045 -7.645 -78.715 -7.315 ;
        RECT -79.045 -9.005 -78.715 -8.675 ;
        RECT -79.045 -10.365 -78.715 -10.035 ;
        RECT -79.045 -11.725 -78.715 -11.395 ;
        RECT -79.045 -13.085 -78.715 -12.755 ;
        RECT -79.045 -14.445 -78.715 -14.115 ;
        RECT -79.045 -15.805 -78.715 -15.475 ;
        RECT -79.045 -17.165 -78.715 -16.835 ;
        RECT -79.045 -18.525 -78.715 -18.195 ;
        RECT -79.045 -19.885 -78.715 -19.555 ;
        RECT -79.045 -21.245 -78.715 -20.915 ;
        RECT -79.045 -22.605 -78.715 -22.275 ;
        RECT -79.045 -23.965 -78.715 -23.635 ;
        RECT -79.045 -25.325 -78.715 -24.995 ;
        RECT -79.045 -26.685 -78.715 -26.355 ;
        RECT -79.045 -28.045 -78.715 -27.715 ;
        RECT -79.045 -29.405 -78.715 -29.075 ;
        RECT -79.045 -30.765 -78.715 -30.435 ;
        RECT -79.045 -32.125 -78.715 -31.795 ;
        RECT -79.045 -33.485 -78.715 -33.155 ;
        RECT -79.045 -34.845 -78.715 -34.515 ;
        RECT -79.045 -36.205 -78.715 -35.875 ;
        RECT -79.045 -37.565 -78.715 -37.235 ;
        RECT -79.045 -38.925 -78.715 -38.595 ;
        RECT -79.045 -40.285 -78.715 -39.955 ;
        RECT -79.045 -41.645 -78.715 -41.315 ;
        RECT -79.045 -43.005 -78.715 -42.675 ;
        RECT -79.045 -44.365 -78.715 -44.035 ;
        RECT -79.045 -45.725 -78.715 -45.395 ;
        RECT -79.045 -47.085 -78.715 -46.755 ;
        RECT -79.045 -48.445 -78.715 -48.115 ;
        RECT -79.045 -49.805 -78.715 -49.475 ;
        RECT -79.045 -51.165 -78.715 -50.835 ;
        RECT -79.045 -52.525 -78.715 -52.195 ;
        RECT -79.045 -53.885 -78.715 -53.555 ;
        RECT -79.045 -55.245 -78.715 -54.915 ;
        RECT -79.045 -56.605 -78.715 -56.275 ;
        RECT -79.045 -57.965 -78.715 -57.635 ;
        RECT -79.045 -59.325 -78.715 -58.995 ;
        RECT -79.045 -60.685 -78.715 -60.355 ;
        RECT -79.045 -62.045 -78.715 -61.715 ;
        RECT -79.045 -63.405 -78.715 -63.075 ;
        RECT -79.045 -64.765 -78.715 -64.435 ;
        RECT -79.045 -66.125 -78.715 -65.795 ;
        RECT -79.045 -67.485 -78.715 -67.155 ;
        RECT -79.045 -68.845 -78.715 -68.515 ;
        RECT -79.045 -70.205 -78.715 -69.875 ;
        RECT -79.045 -71.565 -78.715 -71.235 ;
        RECT -79.045 -72.925 -78.715 -72.595 ;
        RECT -79.045 -74.285 -78.715 -73.955 ;
        RECT -79.045 -75.645 -78.715 -75.315 ;
        RECT -79.045 -77.005 -78.715 -76.675 ;
        RECT -79.045 -78.365 -78.715 -78.035 ;
        RECT -79.045 -79.725 -78.715 -79.395 ;
        RECT -79.045 -81.085 -78.715 -80.755 ;
        RECT -79.045 -82.445 -78.715 -82.115 ;
        RECT -79.045 -83.805 -78.715 -83.475 ;
        RECT -79.045 -85.165 -78.715 -84.835 ;
        RECT -79.045 -86.525 -78.715 -86.195 ;
        RECT -79.045 -87.885 -78.715 -87.555 ;
        RECT -79.045 -89.245 -78.715 -88.915 ;
        RECT -79.045 -90.605 -78.715 -90.275 ;
        RECT -79.045 -91.965 -78.715 -91.635 ;
        RECT -79.045 -93.325 -78.715 -92.995 ;
        RECT -79.045 -94.685 -78.715 -94.355 ;
        RECT -79.045 -96.045 -78.715 -95.715 ;
        RECT -79.045 -97.405 -78.715 -97.075 ;
        RECT -79.045 -98.765 -78.715 -98.435 ;
        RECT -79.045 -100.125 -78.715 -99.795 ;
        RECT -79.045 -101.485 -78.715 -101.155 ;
        RECT -79.045 -102.845 -78.715 -102.515 ;
        RECT -79.045 -104.205 -78.715 -103.875 ;
        RECT -79.045 -105.565 -78.715 -105.235 ;
        RECT -79.045 -106.925 -78.715 -106.595 ;
        RECT -79.045 -108.285 -78.715 -107.955 ;
        RECT -79.045 -109.645 -78.715 -109.315 ;
        RECT -79.045 -111.005 -78.715 -110.675 ;
        RECT -79.045 -112.365 -78.715 -112.035 ;
        RECT -79.045 -113.725 -78.715 -113.395 ;
        RECT -79.045 -115.085 -78.715 -114.755 ;
        RECT -79.045 -116.445 -78.715 -116.115 ;
        RECT -79.045 -117.805 -78.715 -117.475 ;
        RECT -79.045 -119.165 -78.715 -118.835 ;
        RECT -79.045 -120.525 -78.715 -120.195 ;
        RECT -79.045 -121.885 -78.715 -121.555 ;
        RECT -79.045 -123.245 -78.715 -122.915 ;
        RECT -79.045 -124.605 -78.715 -124.275 ;
        RECT -79.045 -125.965 -78.715 -125.635 ;
        RECT -79.045 -127.325 -78.715 -126.995 ;
        RECT -79.045 -128.685 -78.715 -128.355 ;
        RECT -79.045 -130.045 -78.715 -129.715 ;
        RECT -79.045 -131.405 -78.715 -131.075 ;
        RECT -79.045 -132.765 -78.715 -132.435 ;
        RECT -79.045 -134.125 -78.715 -133.795 ;
        RECT -79.045 -135.485 -78.715 -135.155 ;
        RECT -79.045 -136.845 -78.715 -136.515 ;
        RECT -79.045 -138.205 -78.715 -137.875 ;
        RECT -79.045 -139.565 -78.715 -139.235 ;
        RECT -79.045 -140.925 -78.715 -140.595 ;
        RECT -79.045 -142.285 -78.715 -141.955 ;
        RECT -79.045 -143.645 -78.715 -143.315 ;
        RECT -79.045 -145.005 -78.715 -144.675 ;
        RECT -79.045 -146.365 -78.715 -146.035 ;
        RECT -79.045 -147.725 -78.715 -147.395 ;
        RECT -79.045 -149.085 -78.715 -148.755 ;
        RECT -79.045 -150.445 -78.715 -150.115 ;
        RECT -79.045 -151.805 -78.715 -151.475 ;
        RECT -79.045 -153.165 -78.715 -152.835 ;
        RECT -79.045 -154.525 -78.715 -154.195 ;
        RECT -79.045 -155.885 -78.715 -155.555 ;
        RECT -79.045 -157.245 -78.715 -156.915 ;
        RECT -79.045 -158.605 -78.715 -158.275 ;
        RECT -79.045 -159.965 -78.715 -159.635 ;
        RECT -79.045 -161.325 -78.715 -160.995 ;
        RECT -79.045 -162.685 -78.715 -162.355 ;
        RECT -79.045 -164.045 -78.715 -163.715 ;
        RECT -79.045 -165.405 -78.715 -165.075 ;
        RECT -79.045 -166.765 -78.715 -166.435 ;
        RECT -79.045 -168.125 -78.715 -167.795 ;
        RECT -79.045 -169.485 -78.715 -169.155 ;
        RECT -79.045 -170.845 -78.715 -170.515 ;
        RECT -79.045 -172.205 -78.715 -171.875 ;
        RECT -79.045 -173.565 -78.715 -173.235 ;
        RECT -79.045 -174.925 -78.715 -174.595 ;
        RECT -79.045 -176.285 -78.715 -175.955 ;
        RECT -79.045 -177.645 -78.715 -177.315 ;
        RECT -79.045 -179.005 -78.715 -178.675 ;
        RECT -79.045 -184.65 -78.715 -183.52 ;
        RECT -79.04 -184.765 -78.72 245.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -77.685 95.715 -77.355 96.045 ;
        RECT -77.685 94.355 -77.355 94.685 ;
        RECT -77.685 92.995 -77.355 93.325 ;
        RECT -77.685 91.635 -77.355 91.965 ;
        RECT -77.685 90.275 -77.355 90.605 ;
        RECT -77.685 88.915 -77.355 89.245 ;
        RECT -77.685 87.555 -77.355 87.885 ;
        RECT -77.685 86.195 -77.355 86.525 ;
        RECT -77.685 84.835 -77.355 85.165 ;
        RECT -77.685 83.475 -77.355 83.805 ;
        RECT -77.685 82.115 -77.355 82.445 ;
        RECT -77.685 80.755 -77.355 81.085 ;
        RECT -77.685 79.395 -77.355 79.725 ;
        RECT -77.685 78.035 -77.355 78.365 ;
        RECT -77.685 76.675 -77.355 77.005 ;
        RECT -77.685 75.315 -77.355 75.645 ;
        RECT -77.685 73.955 -77.355 74.285 ;
        RECT -77.685 72.595 -77.355 72.925 ;
        RECT -77.685 71.235 -77.355 71.565 ;
        RECT -77.685 69.875 -77.355 70.205 ;
        RECT -77.685 68.515 -77.355 68.845 ;
        RECT -77.685 67.155 -77.355 67.485 ;
        RECT -77.685 65.795 -77.355 66.125 ;
        RECT -77.685 64.435 -77.355 64.765 ;
        RECT -77.685 63.075 -77.355 63.405 ;
        RECT -77.685 61.715 -77.355 62.045 ;
        RECT -77.685 60.355 -77.355 60.685 ;
        RECT -77.685 58.995 -77.355 59.325 ;
        RECT -77.685 57.635 -77.355 57.965 ;
        RECT -77.685 56.275 -77.355 56.605 ;
        RECT -77.685 54.915 -77.355 55.245 ;
        RECT -77.685 53.555 -77.355 53.885 ;
        RECT -77.685 52.195 -77.355 52.525 ;
        RECT -77.685 50.835 -77.355 51.165 ;
        RECT -77.685 49.475 -77.355 49.805 ;
        RECT -77.685 48.115 -77.355 48.445 ;
        RECT -77.685 46.755 -77.355 47.085 ;
        RECT -77.685 45.395 -77.355 45.725 ;
        RECT -77.685 44.035 -77.355 44.365 ;
        RECT -77.685 42.675 -77.355 43.005 ;
        RECT -77.685 41.315 -77.355 41.645 ;
        RECT -77.685 39.955 -77.355 40.285 ;
        RECT -77.685 38.595 -77.355 38.925 ;
        RECT -77.685 37.235 -77.355 37.565 ;
        RECT -77.685 35.875 -77.355 36.205 ;
        RECT -77.685 34.515 -77.355 34.845 ;
        RECT -77.685 33.155 -77.355 33.485 ;
        RECT -77.685 31.795 -77.355 32.125 ;
        RECT -77.685 30.435 -77.355 30.765 ;
        RECT -77.685 29.075 -77.355 29.405 ;
        RECT -77.685 27.715 -77.355 28.045 ;
        RECT -77.685 26.355 -77.355 26.685 ;
        RECT -77.685 24.995 -77.355 25.325 ;
        RECT -77.685 23.635 -77.355 23.965 ;
        RECT -77.685 22.275 -77.355 22.605 ;
        RECT -77.685 20.915 -77.355 21.245 ;
        RECT -77.685 19.555 -77.355 19.885 ;
        RECT -77.685 18.195 -77.355 18.525 ;
        RECT -77.685 16.835 -77.355 17.165 ;
        RECT -77.685 15.475 -77.355 15.805 ;
        RECT -77.685 14.115 -77.355 14.445 ;
        RECT -77.685 12.755 -77.355 13.085 ;
        RECT -77.685 11.395 -77.355 11.725 ;
        RECT -77.685 10.035 -77.355 10.365 ;
        RECT -77.685 8.675 -77.355 9.005 ;
        RECT -77.685 7.315 -77.355 7.645 ;
        RECT -77.685 5.955 -77.355 6.285 ;
        RECT -77.685 4.595 -77.355 4.925 ;
        RECT -77.685 3.235 -77.355 3.565 ;
        RECT -77.685 1.875 -77.355 2.205 ;
        RECT -77.685 0.515 -77.355 0.845 ;
        RECT -77.685 -0.845 -77.355 -0.515 ;
        RECT -77.685 -2.205 -77.355 -1.875 ;
        RECT -77.685 -3.565 -77.355 -3.235 ;
        RECT -77.685 -4.925 -77.355 -4.595 ;
        RECT -77.685 -6.285 -77.355 -5.955 ;
        RECT -77.685 -7.645 -77.355 -7.315 ;
        RECT -77.685 -9.005 -77.355 -8.675 ;
        RECT -77.685 -10.365 -77.355 -10.035 ;
        RECT -77.685 -11.725 -77.355 -11.395 ;
        RECT -77.685 -13.085 -77.355 -12.755 ;
        RECT -77.685 -14.445 -77.355 -14.115 ;
        RECT -77.685 -15.805 -77.355 -15.475 ;
        RECT -77.685 -17.165 -77.355 -16.835 ;
        RECT -77.685 -18.525 -77.355 -18.195 ;
        RECT -77.685 -19.885 -77.355 -19.555 ;
        RECT -77.685 -21.245 -77.355 -20.915 ;
        RECT -77.685 -22.605 -77.355 -22.275 ;
        RECT -77.685 -23.965 -77.355 -23.635 ;
        RECT -77.685 -25.325 -77.355 -24.995 ;
        RECT -77.685 -26.685 -77.355 -26.355 ;
        RECT -77.685 -28.045 -77.355 -27.715 ;
        RECT -77.685 -29.405 -77.355 -29.075 ;
        RECT -77.685 -30.765 -77.355 -30.435 ;
        RECT -77.685 -32.125 -77.355 -31.795 ;
        RECT -77.685 -33.485 -77.355 -33.155 ;
        RECT -77.685 -34.845 -77.355 -34.515 ;
        RECT -77.685 -36.205 -77.355 -35.875 ;
        RECT -77.685 -37.565 -77.355 -37.235 ;
        RECT -77.685 -38.925 -77.355 -38.595 ;
        RECT -77.685 -40.285 -77.355 -39.955 ;
        RECT -77.685 -41.645 -77.355 -41.315 ;
        RECT -77.685 -43.005 -77.355 -42.675 ;
        RECT -77.685 -44.365 -77.355 -44.035 ;
        RECT -77.685 -45.725 -77.355 -45.395 ;
        RECT -77.685 -47.085 -77.355 -46.755 ;
        RECT -77.685 -48.445 -77.355 -48.115 ;
        RECT -77.685 -49.805 -77.355 -49.475 ;
        RECT -77.685 -51.165 -77.355 -50.835 ;
        RECT -77.685 -52.525 -77.355 -52.195 ;
        RECT -77.685 -53.885 -77.355 -53.555 ;
        RECT -77.685 -55.245 -77.355 -54.915 ;
        RECT -77.685 -56.605 -77.355 -56.275 ;
        RECT -77.685 -57.965 -77.355 -57.635 ;
        RECT -77.685 -59.325 -77.355 -58.995 ;
        RECT -77.685 -60.685 -77.355 -60.355 ;
        RECT -77.685 -62.045 -77.355 -61.715 ;
        RECT -77.685 -63.405 -77.355 -63.075 ;
        RECT -77.685 -64.765 -77.355 -64.435 ;
        RECT -77.685 -66.125 -77.355 -65.795 ;
        RECT -77.685 -67.485 -77.355 -67.155 ;
        RECT -77.685 -68.845 -77.355 -68.515 ;
        RECT -77.685 -70.205 -77.355 -69.875 ;
        RECT -77.685 -71.565 -77.355 -71.235 ;
        RECT -77.685 -72.925 -77.355 -72.595 ;
        RECT -77.685 -74.285 -77.355 -73.955 ;
        RECT -77.685 -75.645 -77.355 -75.315 ;
        RECT -77.685 -77.005 -77.355 -76.675 ;
        RECT -77.685 -78.365 -77.355 -78.035 ;
        RECT -77.685 -79.725 -77.355 -79.395 ;
        RECT -77.685 -81.085 -77.355 -80.755 ;
        RECT -77.685 -82.445 -77.355 -82.115 ;
        RECT -77.685 -83.805 -77.355 -83.475 ;
        RECT -77.685 -85.165 -77.355 -84.835 ;
        RECT -77.685 -86.525 -77.355 -86.195 ;
        RECT -77.685 -87.885 -77.355 -87.555 ;
        RECT -77.685 -89.245 -77.355 -88.915 ;
        RECT -77.685 -90.605 -77.355 -90.275 ;
        RECT -77.685 -91.965 -77.355 -91.635 ;
        RECT -77.685 -93.325 -77.355 -92.995 ;
        RECT -77.685 -94.685 -77.355 -94.355 ;
        RECT -77.685 -96.045 -77.355 -95.715 ;
        RECT -77.685 -97.405 -77.355 -97.075 ;
        RECT -77.685 -98.765 -77.355 -98.435 ;
        RECT -77.685 -100.125 -77.355 -99.795 ;
        RECT -77.685 -101.485 -77.355 -101.155 ;
        RECT -77.685 -102.845 -77.355 -102.515 ;
        RECT -77.685 -104.205 -77.355 -103.875 ;
        RECT -77.685 -105.565 -77.355 -105.235 ;
        RECT -77.685 -106.925 -77.355 -106.595 ;
        RECT -77.685 -108.285 -77.355 -107.955 ;
        RECT -77.685 -109.645 -77.355 -109.315 ;
        RECT -77.685 -111.005 -77.355 -110.675 ;
        RECT -77.685 -112.365 -77.355 -112.035 ;
        RECT -77.685 -113.725 -77.355 -113.395 ;
        RECT -77.685 -115.085 -77.355 -114.755 ;
        RECT -77.685 -116.445 -77.355 -116.115 ;
        RECT -77.685 -117.805 -77.355 -117.475 ;
        RECT -77.685 -119.165 -77.355 -118.835 ;
        RECT -77.685 -120.525 -77.355 -120.195 ;
        RECT -77.685 -121.885 -77.355 -121.555 ;
        RECT -77.685 -123.245 -77.355 -122.915 ;
        RECT -77.685 -124.605 -77.355 -124.275 ;
        RECT -77.685 -125.965 -77.355 -125.635 ;
        RECT -77.685 -127.325 -77.355 -126.995 ;
        RECT -77.685 -128.685 -77.355 -128.355 ;
        RECT -77.685 -130.045 -77.355 -129.715 ;
        RECT -77.685 -131.405 -77.355 -131.075 ;
        RECT -77.685 -132.765 -77.355 -132.435 ;
        RECT -77.685 -134.125 -77.355 -133.795 ;
        RECT -77.685 -135.485 -77.355 -135.155 ;
        RECT -77.685 -136.845 -77.355 -136.515 ;
        RECT -77.685 -138.205 -77.355 -137.875 ;
        RECT -77.685 -139.565 -77.355 -139.235 ;
        RECT -77.685 -140.925 -77.355 -140.595 ;
        RECT -77.685 -142.285 -77.355 -141.955 ;
        RECT -77.685 -143.645 -77.355 -143.315 ;
        RECT -77.685 -145.005 -77.355 -144.675 ;
        RECT -77.685 -146.365 -77.355 -146.035 ;
        RECT -77.685 -147.725 -77.355 -147.395 ;
        RECT -77.685 -149.085 -77.355 -148.755 ;
        RECT -77.685 -150.445 -77.355 -150.115 ;
        RECT -77.685 -151.805 -77.355 -151.475 ;
        RECT -77.685 -153.165 -77.355 -152.835 ;
        RECT -77.685 -154.525 -77.355 -154.195 ;
        RECT -77.685 -155.885 -77.355 -155.555 ;
        RECT -77.685 -157.245 -77.355 -156.915 ;
        RECT -77.685 -158.605 -77.355 -158.275 ;
        RECT -77.685 -159.965 -77.355 -159.635 ;
        RECT -77.685 -161.325 -77.355 -160.995 ;
        RECT -77.685 -162.685 -77.355 -162.355 ;
        RECT -77.685 -164.045 -77.355 -163.715 ;
        RECT -77.685 -165.405 -77.355 -165.075 ;
        RECT -77.685 -166.765 -77.355 -166.435 ;
        RECT -77.685 -168.125 -77.355 -167.795 ;
        RECT -77.685 -169.615 -77.355 -169.285 ;
        RECT -77.685 -170.845 -77.355 -170.515 ;
        RECT -77.685 -172.205 -77.355 -171.875 ;
        RECT -77.68 -172.88 -77.36 245.285 ;
        RECT -77.685 244.04 -77.355 245.17 ;
        RECT -77.685 239.875 -77.355 240.205 ;
        RECT -77.685 238.515 -77.355 238.845 ;
        RECT -77.685 237.155 -77.355 237.485 ;
        RECT -77.685 235.795 -77.355 236.125 ;
        RECT -77.685 234.435 -77.355 234.765 ;
        RECT -77.685 233.075 -77.355 233.405 ;
        RECT -77.685 231.715 -77.355 232.045 ;
        RECT -77.685 230.355 -77.355 230.685 ;
        RECT -77.685 228.995 -77.355 229.325 ;
        RECT -77.685 227.635 -77.355 227.965 ;
        RECT -77.685 226.275 -77.355 226.605 ;
        RECT -77.685 224.915 -77.355 225.245 ;
        RECT -77.685 223.555 -77.355 223.885 ;
        RECT -77.685 222.195 -77.355 222.525 ;
        RECT -77.685 220.835 -77.355 221.165 ;
        RECT -77.685 219.475 -77.355 219.805 ;
        RECT -77.685 218.115 -77.355 218.445 ;
        RECT -77.685 216.755 -77.355 217.085 ;
        RECT -77.685 215.395 -77.355 215.725 ;
        RECT -77.685 214.035 -77.355 214.365 ;
        RECT -77.685 212.675 -77.355 213.005 ;
        RECT -77.685 211.315 -77.355 211.645 ;
        RECT -77.685 209.955 -77.355 210.285 ;
        RECT -77.685 208.595 -77.355 208.925 ;
        RECT -77.685 207.235 -77.355 207.565 ;
        RECT -77.685 205.875 -77.355 206.205 ;
        RECT -77.685 204.515 -77.355 204.845 ;
        RECT -77.685 203.155 -77.355 203.485 ;
        RECT -77.685 201.795 -77.355 202.125 ;
        RECT -77.685 200.435 -77.355 200.765 ;
        RECT -77.685 199.075 -77.355 199.405 ;
        RECT -77.685 197.715 -77.355 198.045 ;
        RECT -77.685 196.355 -77.355 196.685 ;
        RECT -77.685 194.995 -77.355 195.325 ;
        RECT -77.685 193.635 -77.355 193.965 ;
        RECT -77.685 192.275 -77.355 192.605 ;
        RECT -77.685 190.915 -77.355 191.245 ;
        RECT -77.685 189.555 -77.355 189.885 ;
        RECT -77.685 188.195 -77.355 188.525 ;
        RECT -77.685 186.835 -77.355 187.165 ;
        RECT -77.685 185.475 -77.355 185.805 ;
        RECT -77.685 184.115 -77.355 184.445 ;
        RECT -77.685 182.755 -77.355 183.085 ;
        RECT -77.685 181.395 -77.355 181.725 ;
        RECT -77.685 180.035 -77.355 180.365 ;
        RECT -77.685 178.675 -77.355 179.005 ;
        RECT -77.685 177.315 -77.355 177.645 ;
        RECT -77.685 175.955 -77.355 176.285 ;
        RECT -77.685 174.595 -77.355 174.925 ;
        RECT -77.685 173.235 -77.355 173.565 ;
        RECT -77.685 171.875 -77.355 172.205 ;
        RECT -77.685 170.515 -77.355 170.845 ;
        RECT -77.685 169.155 -77.355 169.485 ;
        RECT -77.685 167.795 -77.355 168.125 ;
        RECT -77.685 166.435 -77.355 166.765 ;
        RECT -77.685 165.075 -77.355 165.405 ;
        RECT -77.685 163.715 -77.355 164.045 ;
        RECT -77.685 162.355 -77.355 162.685 ;
        RECT -77.685 160.995 -77.355 161.325 ;
        RECT -77.685 159.635 -77.355 159.965 ;
        RECT -77.685 158.275 -77.355 158.605 ;
        RECT -77.685 156.915 -77.355 157.245 ;
        RECT -77.685 155.555 -77.355 155.885 ;
        RECT -77.685 154.195 -77.355 154.525 ;
        RECT -77.685 152.835 -77.355 153.165 ;
        RECT -77.685 151.475 -77.355 151.805 ;
        RECT -77.685 150.115 -77.355 150.445 ;
        RECT -77.685 148.755 -77.355 149.085 ;
        RECT -77.685 147.395 -77.355 147.725 ;
        RECT -77.685 146.035 -77.355 146.365 ;
        RECT -77.685 144.675 -77.355 145.005 ;
        RECT -77.685 143.315 -77.355 143.645 ;
        RECT -77.685 141.955 -77.355 142.285 ;
        RECT -77.685 140.595 -77.355 140.925 ;
        RECT -77.685 139.235 -77.355 139.565 ;
        RECT -77.685 137.875 -77.355 138.205 ;
        RECT -77.685 136.515 -77.355 136.845 ;
        RECT -77.685 135.155 -77.355 135.485 ;
        RECT -77.685 133.795 -77.355 134.125 ;
        RECT -77.685 132.435 -77.355 132.765 ;
        RECT -77.685 131.075 -77.355 131.405 ;
        RECT -77.685 129.715 -77.355 130.045 ;
        RECT -77.685 128.355 -77.355 128.685 ;
        RECT -77.685 126.995 -77.355 127.325 ;
        RECT -77.685 125.635 -77.355 125.965 ;
        RECT -77.685 124.275 -77.355 124.605 ;
        RECT -77.685 122.915 -77.355 123.245 ;
        RECT -77.685 121.555 -77.355 121.885 ;
        RECT -77.685 120.195 -77.355 120.525 ;
        RECT -77.685 118.835 -77.355 119.165 ;
        RECT -77.685 117.475 -77.355 117.805 ;
        RECT -77.685 116.115 -77.355 116.445 ;
        RECT -77.685 114.755 -77.355 115.085 ;
        RECT -77.685 113.395 -77.355 113.725 ;
        RECT -77.685 112.035 -77.355 112.365 ;
        RECT -77.685 110.675 -77.355 111.005 ;
        RECT -77.685 109.315 -77.355 109.645 ;
        RECT -77.685 107.955 -77.355 108.285 ;
        RECT -77.685 106.595 -77.355 106.925 ;
        RECT -77.685 105.235 -77.355 105.565 ;
        RECT -77.685 103.875 -77.355 104.205 ;
        RECT -77.685 102.515 -77.355 102.845 ;
        RECT -77.685 101.155 -77.355 101.485 ;
        RECT -77.685 99.795 -77.355 100.125 ;
        RECT -77.685 98.435 -77.355 98.765 ;
        RECT -77.685 97.075 -77.355 97.405 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 356.835 241.32 357.165 242.45 ;
        RECT 356.835 239.195 357.165 239.525 ;
        RECT 356.835 237.835 357.165 238.165 ;
        RECT 356.835 235.975 357.165 236.305 ;
        RECT 356.835 233.925 357.165 234.255 ;
        RECT 356.835 231.995 357.165 232.325 ;
        RECT 356.835 230.155 357.165 230.485 ;
        RECT 356.835 228.665 357.165 228.995 ;
        RECT 356.835 226.995 357.165 227.325 ;
        RECT 356.835 225.505 357.165 225.835 ;
        RECT 356.835 223.835 357.165 224.165 ;
        RECT 356.835 222.345 357.165 222.675 ;
        RECT 356.835 220.675 357.165 221.005 ;
        RECT 356.835 219.185 357.165 219.515 ;
        RECT 356.835 217.775 357.165 218.105 ;
        RECT 356.835 215.935 357.165 216.265 ;
        RECT 356.835 214.445 357.165 214.775 ;
        RECT 356.835 212.775 357.165 213.105 ;
        RECT 356.835 211.285 357.165 211.615 ;
        RECT 356.835 209.615 357.165 209.945 ;
        RECT 356.835 208.125 357.165 208.455 ;
        RECT 356.835 206.455 357.165 206.785 ;
        RECT 356.835 204.965 357.165 205.295 ;
        RECT 356.835 203.555 357.165 203.885 ;
        RECT 356.835 201.715 357.165 202.045 ;
        RECT 356.835 200.225 357.165 200.555 ;
        RECT 356.835 198.555 357.165 198.885 ;
        RECT 356.835 197.065 357.165 197.395 ;
        RECT 356.835 195.395 357.165 195.725 ;
        RECT 356.835 193.905 357.165 194.235 ;
        RECT 356.835 192.235 357.165 192.565 ;
        RECT 356.835 190.745 357.165 191.075 ;
        RECT 356.835 189.335 357.165 189.665 ;
        RECT 356.835 187.495 357.165 187.825 ;
        RECT 356.835 186.005 357.165 186.335 ;
        RECT 356.835 184.335 357.165 184.665 ;
        RECT 356.835 182.845 357.165 183.175 ;
        RECT 356.835 181.175 357.165 181.505 ;
        RECT 356.835 179.685 357.165 180.015 ;
        RECT 356.835 178.015 357.165 178.345 ;
        RECT 356.835 176.525 357.165 176.855 ;
        RECT 356.835 175.115 357.165 175.445 ;
        RECT 356.835 173.275 357.165 173.605 ;
        RECT 356.835 171.785 357.165 172.115 ;
        RECT 356.835 170.115 357.165 170.445 ;
        RECT 356.835 168.625 357.165 168.955 ;
        RECT 356.835 166.955 357.165 167.285 ;
        RECT 356.835 165.465 357.165 165.795 ;
        RECT 356.835 163.795 357.165 164.125 ;
        RECT 356.835 162.305 357.165 162.635 ;
        RECT 356.835 160.895 357.165 161.225 ;
        RECT 356.835 159.055 357.165 159.385 ;
        RECT 356.835 157.565 357.165 157.895 ;
        RECT 356.835 155.895 357.165 156.225 ;
        RECT 356.835 154.405 357.165 154.735 ;
        RECT 356.835 152.735 357.165 153.065 ;
        RECT 356.835 151.245 357.165 151.575 ;
        RECT 356.835 149.575 357.165 149.905 ;
        RECT 356.835 148.085 357.165 148.415 ;
        RECT 356.835 146.675 357.165 147.005 ;
        RECT 356.835 144.835 357.165 145.165 ;
        RECT 356.835 143.345 357.165 143.675 ;
        RECT 356.835 141.675 357.165 142.005 ;
        RECT 356.835 140.185 357.165 140.515 ;
        RECT 356.835 138.515 357.165 138.845 ;
        RECT 356.835 137.025 357.165 137.355 ;
        RECT 356.835 135.355 357.165 135.685 ;
        RECT 356.835 133.865 357.165 134.195 ;
        RECT 356.835 132.455 357.165 132.785 ;
        RECT 356.835 130.615 357.165 130.945 ;
        RECT 356.835 129.125 357.165 129.455 ;
        RECT 356.835 127.455 357.165 127.785 ;
        RECT 356.835 125.965 357.165 126.295 ;
        RECT 356.835 124.295 357.165 124.625 ;
        RECT 356.835 122.805 357.165 123.135 ;
        RECT 356.835 121.135 357.165 121.465 ;
        RECT 356.835 119.645 357.165 119.975 ;
        RECT 356.835 118.235 357.165 118.565 ;
        RECT 356.835 116.395 357.165 116.725 ;
        RECT 356.835 114.905 357.165 115.235 ;
        RECT 356.835 113.235 357.165 113.565 ;
        RECT 356.835 111.745 357.165 112.075 ;
        RECT 356.835 110.075 357.165 110.405 ;
        RECT 356.835 108.585 357.165 108.915 ;
        RECT 356.835 106.915 357.165 107.245 ;
        RECT 356.835 105.425 357.165 105.755 ;
        RECT 356.835 104.015 357.165 104.345 ;
        RECT 356.835 102.175 357.165 102.505 ;
        RECT 356.835 100.685 357.165 101.015 ;
        RECT 356.835 99.015 357.165 99.345 ;
        RECT 356.835 97.525 357.165 97.855 ;
        RECT 356.835 95.855 357.165 96.185 ;
        RECT 356.835 94.365 357.165 94.695 ;
        RECT 356.835 92.695 357.165 93.025 ;
        RECT 356.835 91.205 357.165 91.535 ;
        RECT 356.835 89.795 357.165 90.125 ;
        RECT 356.835 87.955 357.165 88.285 ;
        RECT 356.835 86.465 357.165 86.795 ;
        RECT 356.835 84.795 357.165 85.125 ;
        RECT 356.835 83.305 357.165 83.635 ;
        RECT 356.835 81.635 357.165 81.965 ;
        RECT 356.835 80.145 357.165 80.475 ;
        RECT 356.835 78.475 357.165 78.805 ;
        RECT 356.835 76.985 357.165 77.315 ;
        RECT 356.835 75.575 357.165 75.905 ;
        RECT 356.835 73.735 357.165 74.065 ;
        RECT 356.835 72.245 357.165 72.575 ;
        RECT 356.835 70.575 357.165 70.905 ;
        RECT 356.835 69.085 357.165 69.415 ;
        RECT 356.835 67.415 357.165 67.745 ;
        RECT 356.835 65.925 357.165 66.255 ;
        RECT 356.835 64.255 357.165 64.585 ;
        RECT 356.835 62.765 357.165 63.095 ;
        RECT 356.835 61.355 357.165 61.685 ;
        RECT 356.835 59.515 357.165 59.845 ;
        RECT 356.835 58.025 357.165 58.355 ;
        RECT 356.835 56.355 357.165 56.685 ;
        RECT 356.835 54.865 357.165 55.195 ;
        RECT 356.835 53.195 357.165 53.525 ;
        RECT 356.835 51.705 357.165 52.035 ;
        RECT 356.835 50.035 357.165 50.365 ;
        RECT 356.835 48.545 357.165 48.875 ;
        RECT 356.835 47.135 357.165 47.465 ;
        RECT 356.835 45.295 357.165 45.625 ;
        RECT 356.835 43.805 357.165 44.135 ;
        RECT 356.835 42.135 357.165 42.465 ;
        RECT 356.835 40.645 357.165 40.975 ;
        RECT 356.835 38.975 357.165 39.305 ;
        RECT 356.835 37.485 357.165 37.815 ;
        RECT 356.835 35.815 357.165 36.145 ;
        RECT 356.835 34.325 357.165 34.655 ;
        RECT 356.835 32.915 357.165 33.245 ;
        RECT 356.835 31.075 357.165 31.405 ;
        RECT 356.835 29.585 357.165 29.915 ;
        RECT 356.835 27.915 357.165 28.245 ;
        RECT 356.835 26.425 357.165 26.755 ;
        RECT 356.835 24.755 357.165 25.085 ;
        RECT 356.835 23.265 357.165 23.595 ;
        RECT 356.835 21.595 357.165 21.925 ;
        RECT 356.835 20.105 357.165 20.435 ;
        RECT 356.835 18.695 357.165 19.025 ;
        RECT 356.835 16.855 357.165 17.185 ;
        RECT 356.835 15.365 357.165 15.695 ;
        RECT 356.835 13.695 357.165 14.025 ;
        RECT 356.835 12.205 357.165 12.535 ;
        RECT 356.835 10.535 357.165 10.865 ;
        RECT 356.835 9.045 357.165 9.375 ;
        RECT 356.835 7.375 357.165 7.705 ;
        RECT 356.835 5.885 357.165 6.215 ;
        RECT 356.835 4.475 357.165 4.805 ;
        RECT 356.835 2.115 357.165 2.445 ;
        RECT 356.835 0.06 357.165 0.39 ;
        RECT 356.835 -1.525 357.165 -1.195 ;
        RECT 356.835 -2.885 357.165 -2.555 ;
        RECT 356.835 -4.245 357.165 -3.915 ;
        RECT 356.835 -5.605 357.165 -5.275 ;
        RECT 356.835 -6.965 357.165 -6.635 ;
        RECT 356.835 -8.325 357.165 -7.995 ;
        RECT 356.835 -9.685 357.165 -9.355 ;
        RECT 356.835 -11.045 357.165 -10.715 ;
        RECT 356.835 -12.405 357.165 -12.075 ;
        RECT 356.835 -13.765 357.165 -13.435 ;
        RECT 356.835 -15.125 357.165 -14.795 ;
        RECT 356.835 -16.485 357.165 -16.155 ;
        RECT 356.835 -17.845 357.165 -17.515 ;
        RECT 356.835 -19.205 357.165 -18.875 ;
        RECT 356.835 -20.565 357.165 -20.235 ;
        RECT 356.835 -21.925 357.165 -21.595 ;
        RECT 356.835 -23.285 357.165 -22.955 ;
        RECT 356.835 -24.645 357.165 -24.315 ;
        RECT 356.835 -26.005 357.165 -25.675 ;
        RECT 356.835 -27.365 357.165 -27.035 ;
        RECT 356.835 -28.725 357.165 -28.395 ;
        RECT 356.835 -30.085 357.165 -29.755 ;
        RECT 356.835 -31.445 357.165 -31.115 ;
        RECT 356.835 -32.805 357.165 -32.475 ;
        RECT 356.835 -34.165 357.165 -33.835 ;
        RECT 356.835 -35.525 357.165 -35.195 ;
        RECT 356.835 -36.885 357.165 -36.555 ;
        RECT 356.835 -38.245 357.165 -37.915 ;
        RECT 356.835 -39.605 357.165 -39.275 ;
        RECT 356.835 -40.965 357.165 -40.635 ;
        RECT 356.835 -42.325 357.165 -41.995 ;
        RECT 356.835 -43.685 357.165 -43.355 ;
        RECT 356.835 -45.045 357.165 -44.715 ;
        RECT 356.835 -46.405 357.165 -46.075 ;
        RECT 356.835 -47.765 357.165 -47.435 ;
        RECT 356.835 -49.125 357.165 -48.795 ;
        RECT 356.835 -50.485 357.165 -50.155 ;
        RECT 356.835 -51.845 357.165 -51.515 ;
        RECT 356.835 -53.205 357.165 -52.875 ;
        RECT 356.835 -54.565 357.165 -54.235 ;
        RECT 356.835 -55.925 357.165 -55.595 ;
        RECT 356.835 -57.285 357.165 -56.955 ;
        RECT 356.835 -58.645 357.165 -58.315 ;
        RECT 356.835 -60.005 357.165 -59.675 ;
        RECT 356.835 -61.365 357.165 -61.035 ;
        RECT 356.835 -62.725 357.165 -62.395 ;
        RECT 356.835 -64.085 357.165 -63.755 ;
        RECT 356.835 -65.445 357.165 -65.115 ;
        RECT 356.835 -66.805 357.165 -66.475 ;
        RECT 356.835 -68.165 357.165 -67.835 ;
        RECT 356.835 -69.525 357.165 -69.195 ;
        RECT 356.835 -70.885 357.165 -70.555 ;
        RECT 356.835 -72.245 357.165 -71.915 ;
        RECT 356.835 -73.605 357.165 -73.275 ;
        RECT 356.835 -74.965 357.165 -74.635 ;
        RECT 356.835 -76.325 357.165 -75.995 ;
        RECT 356.835 -77.685 357.165 -77.355 ;
        RECT 356.835 -79.045 357.165 -78.715 ;
        RECT 356.835 -80.405 357.165 -80.075 ;
        RECT 356.835 -81.765 357.165 -81.435 ;
        RECT 356.835 -83.125 357.165 -82.795 ;
        RECT 356.835 -84.485 357.165 -84.155 ;
        RECT 356.835 -85.845 357.165 -85.515 ;
        RECT 356.835 -87.205 357.165 -86.875 ;
        RECT 356.835 -88.565 357.165 -88.235 ;
        RECT 356.835 -89.925 357.165 -89.595 ;
        RECT 356.835 -91.285 357.165 -90.955 ;
        RECT 356.835 -92.645 357.165 -92.315 ;
        RECT 356.835 -94.005 357.165 -93.675 ;
        RECT 356.835 -95.365 357.165 -95.035 ;
        RECT 356.835 -96.725 357.165 -96.395 ;
        RECT 356.835 -98.085 357.165 -97.755 ;
        RECT 356.835 -99.445 357.165 -99.115 ;
        RECT 356.835 -100.805 357.165 -100.475 ;
        RECT 356.835 -102.165 357.165 -101.835 ;
        RECT 356.835 -103.525 357.165 -103.195 ;
        RECT 356.835 -104.885 357.165 -104.555 ;
        RECT 356.835 -106.245 357.165 -105.915 ;
        RECT 356.835 -107.605 357.165 -107.275 ;
        RECT 356.835 -108.965 357.165 -108.635 ;
        RECT 356.835 -110.325 357.165 -109.995 ;
        RECT 356.835 -111.685 357.165 -111.355 ;
        RECT 356.835 -113.045 357.165 -112.715 ;
        RECT 356.835 -114.405 357.165 -114.075 ;
        RECT 356.835 -115.765 357.165 -115.435 ;
        RECT 356.835 -117.125 357.165 -116.795 ;
        RECT 356.835 -118.485 357.165 -118.155 ;
        RECT 356.835 -119.845 357.165 -119.515 ;
        RECT 356.835 -121.205 357.165 -120.875 ;
        RECT 356.835 -122.565 357.165 -122.235 ;
        RECT 356.835 -123.925 357.165 -123.595 ;
        RECT 356.835 -125.285 357.165 -124.955 ;
        RECT 356.835 -126.645 357.165 -126.315 ;
        RECT 356.835 -128.005 357.165 -127.675 ;
        RECT 356.835 -129.365 357.165 -129.035 ;
        RECT 356.835 -130.725 357.165 -130.395 ;
        RECT 356.835 -132.085 357.165 -131.755 ;
        RECT 356.835 -133.445 357.165 -133.115 ;
        RECT 356.835 -134.805 357.165 -134.475 ;
        RECT 356.835 -136.165 357.165 -135.835 ;
        RECT 356.835 -137.525 357.165 -137.195 ;
        RECT 356.835 -138.885 357.165 -138.555 ;
        RECT 356.835 -140.245 357.165 -139.915 ;
        RECT 356.835 -141.605 357.165 -141.275 ;
        RECT 356.835 -142.965 357.165 -142.635 ;
        RECT 356.835 -144.325 357.165 -143.995 ;
        RECT 356.835 -145.685 357.165 -145.355 ;
        RECT 356.835 -147.045 357.165 -146.715 ;
        RECT 356.835 -148.405 357.165 -148.075 ;
        RECT 356.835 -149.765 357.165 -149.435 ;
        RECT 356.835 -151.125 357.165 -150.795 ;
        RECT 356.835 -152.485 357.165 -152.155 ;
        RECT 356.835 -153.845 357.165 -153.515 ;
        RECT 356.835 -155.205 357.165 -154.875 ;
        RECT 356.835 -156.565 357.165 -156.235 ;
        RECT 356.835 -157.925 357.165 -157.595 ;
        RECT 356.835 -159.285 357.165 -158.955 ;
        RECT 356.835 -160.645 357.165 -160.315 ;
        RECT 356.835 -162.005 357.165 -161.675 ;
        RECT 356.835 -163.365 357.165 -163.035 ;
        RECT 356.835 -164.725 357.165 -164.395 ;
        RECT 356.835 -166.085 357.165 -165.755 ;
        RECT 356.835 -167.445 357.165 -167.115 ;
        RECT 356.835 -168.805 357.165 -168.475 ;
        RECT 356.835 -170.165 357.165 -169.835 ;
        RECT 356.835 -171.525 357.165 -171.195 ;
        RECT 356.835 -172.885 357.165 -172.555 ;
        RECT 356.835 -174.245 357.165 -173.915 ;
        RECT 356.835 -175.605 357.165 -175.275 ;
        RECT 356.835 -176.965 357.165 -176.635 ;
        RECT 356.835 -178.325 357.165 -177.995 ;
        RECT 356.835 -179.685 357.165 -179.355 ;
        RECT 356.835 -181.93 357.165 -180.8 ;
        RECT 356.84 -182.045 357.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 358.195 241.32 358.525 242.45 ;
        RECT 358.195 239.195 358.525 239.525 ;
        RECT 358.195 237.835 358.525 238.165 ;
        RECT 358.195 235.975 358.525 236.305 ;
        RECT 358.195 233.925 358.525 234.255 ;
        RECT 358.195 231.995 358.525 232.325 ;
        RECT 358.195 230.155 358.525 230.485 ;
        RECT 358.195 228.665 358.525 228.995 ;
        RECT 358.195 226.995 358.525 227.325 ;
        RECT 358.195 225.505 358.525 225.835 ;
        RECT 358.195 223.835 358.525 224.165 ;
        RECT 358.195 222.345 358.525 222.675 ;
        RECT 358.195 220.675 358.525 221.005 ;
        RECT 358.195 219.185 358.525 219.515 ;
        RECT 358.195 217.775 358.525 218.105 ;
        RECT 358.195 215.935 358.525 216.265 ;
        RECT 358.195 214.445 358.525 214.775 ;
        RECT 358.195 212.775 358.525 213.105 ;
        RECT 358.195 211.285 358.525 211.615 ;
        RECT 358.195 209.615 358.525 209.945 ;
        RECT 358.195 208.125 358.525 208.455 ;
        RECT 358.195 206.455 358.525 206.785 ;
        RECT 358.195 204.965 358.525 205.295 ;
        RECT 358.195 203.555 358.525 203.885 ;
        RECT 358.195 201.715 358.525 202.045 ;
        RECT 358.195 200.225 358.525 200.555 ;
        RECT 358.195 198.555 358.525 198.885 ;
        RECT 358.195 197.065 358.525 197.395 ;
        RECT 358.195 195.395 358.525 195.725 ;
        RECT 358.195 193.905 358.525 194.235 ;
        RECT 358.195 192.235 358.525 192.565 ;
        RECT 358.195 190.745 358.525 191.075 ;
        RECT 358.195 189.335 358.525 189.665 ;
        RECT 358.195 187.495 358.525 187.825 ;
        RECT 358.195 186.005 358.525 186.335 ;
        RECT 358.195 184.335 358.525 184.665 ;
        RECT 358.195 182.845 358.525 183.175 ;
        RECT 358.195 181.175 358.525 181.505 ;
        RECT 358.195 179.685 358.525 180.015 ;
        RECT 358.195 178.015 358.525 178.345 ;
        RECT 358.195 176.525 358.525 176.855 ;
        RECT 358.195 175.115 358.525 175.445 ;
        RECT 358.195 173.275 358.525 173.605 ;
        RECT 358.195 171.785 358.525 172.115 ;
        RECT 358.195 170.115 358.525 170.445 ;
        RECT 358.195 168.625 358.525 168.955 ;
        RECT 358.195 166.955 358.525 167.285 ;
        RECT 358.195 165.465 358.525 165.795 ;
        RECT 358.195 163.795 358.525 164.125 ;
        RECT 358.195 162.305 358.525 162.635 ;
        RECT 358.195 160.895 358.525 161.225 ;
        RECT 358.195 159.055 358.525 159.385 ;
        RECT 358.195 157.565 358.525 157.895 ;
        RECT 358.195 155.895 358.525 156.225 ;
        RECT 358.195 154.405 358.525 154.735 ;
        RECT 358.195 152.735 358.525 153.065 ;
        RECT 358.195 151.245 358.525 151.575 ;
        RECT 358.195 149.575 358.525 149.905 ;
        RECT 358.195 148.085 358.525 148.415 ;
        RECT 358.195 146.675 358.525 147.005 ;
        RECT 358.195 144.835 358.525 145.165 ;
        RECT 358.195 143.345 358.525 143.675 ;
        RECT 358.195 141.675 358.525 142.005 ;
        RECT 358.195 140.185 358.525 140.515 ;
        RECT 358.195 138.515 358.525 138.845 ;
        RECT 358.195 137.025 358.525 137.355 ;
        RECT 358.195 135.355 358.525 135.685 ;
        RECT 358.195 133.865 358.525 134.195 ;
        RECT 358.195 132.455 358.525 132.785 ;
        RECT 358.195 130.615 358.525 130.945 ;
        RECT 358.195 129.125 358.525 129.455 ;
        RECT 358.195 127.455 358.525 127.785 ;
        RECT 358.195 125.965 358.525 126.295 ;
        RECT 358.195 124.295 358.525 124.625 ;
        RECT 358.195 122.805 358.525 123.135 ;
        RECT 358.195 121.135 358.525 121.465 ;
        RECT 358.195 119.645 358.525 119.975 ;
        RECT 358.195 118.235 358.525 118.565 ;
        RECT 358.195 116.395 358.525 116.725 ;
        RECT 358.195 114.905 358.525 115.235 ;
        RECT 358.195 113.235 358.525 113.565 ;
        RECT 358.195 111.745 358.525 112.075 ;
        RECT 358.195 110.075 358.525 110.405 ;
        RECT 358.195 108.585 358.525 108.915 ;
        RECT 358.195 106.915 358.525 107.245 ;
        RECT 358.195 105.425 358.525 105.755 ;
        RECT 358.195 104.015 358.525 104.345 ;
        RECT 358.195 102.175 358.525 102.505 ;
        RECT 358.195 100.685 358.525 101.015 ;
        RECT 358.195 99.015 358.525 99.345 ;
        RECT 358.195 97.525 358.525 97.855 ;
        RECT 358.195 95.855 358.525 96.185 ;
        RECT 358.195 94.365 358.525 94.695 ;
        RECT 358.195 92.695 358.525 93.025 ;
        RECT 358.195 91.205 358.525 91.535 ;
        RECT 358.195 89.795 358.525 90.125 ;
        RECT 358.195 87.955 358.525 88.285 ;
        RECT 358.195 86.465 358.525 86.795 ;
        RECT 358.195 84.795 358.525 85.125 ;
        RECT 358.195 83.305 358.525 83.635 ;
        RECT 358.195 81.635 358.525 81.965 ;
        RECT 358.195 80.145 358.525 80.475 ;
        RECT 358.195 78.475 358.525 78.805 ;
        RECT 358.195 76.985 358.525 77.315 ;
        RECT 358.195 75.575 358.525 75.905 ;
        RECT 358.195 73.735 358.525 74.065 ;
        RECT 358.195 72.245 358.525 72.575 ;
        RECT 358.195 70.575 358.525 70.905 ;
        RECT 358.195 69.085 358.525 69.415 ;
        RECT 358.195 67.415 358.525 67.745 ;
        RECT 358.195 65.925 358.525 66.255 ;
        RECT 358.195 64.255 358.525 64.585 ;
        RECT 358.195 62.765 358.525 63.095 ;
        RECT 358.195 61.355 358.525 61.685 ;
        RECT 358.195 59.515 358.525 59.845 ;
        RECT 358.195 58.025 358.525 58.355 ;
        RECT 358.195 56.355 358.525 56.685 ;
        RECT 358.195 54.865 358.525 55.195 ;
        RECT 358.195 53.195 358.525 53.525 ;
        RECT 358.195 51.705 358.525 52.035 ;
        RECT 358.195 50.035 358.525 50.365 ;
        RECT 358.195 48.545 358.525 48.875 ;
        RECT 358.195 47.135 358.525 47.465 ;
        RECT 358.195 45.295 358.525 45.625 ;
        RECT 358.195 43.805 358.525 44.135 ;
        RECT 358.195 42.135 358.525 42.465 ;
        RECT 358.195 40.645 358.525 40.975 ;
        RECT 358.195 38.975 358.525 39.305 ;
        RECT 358.195 37.485 358.525 37.815 ;
        RECT 358.195 35.815 358.525 36.145 ;
        RECT 358.195 34.325 358.525 34.655 ;
        RECT 358.195 32.915 358.525 33.245 ;
        RECT 358.195 31.075 358.525 31.405 ;
        RECT 358.195 29.585 358.525 29.915 ;
        RECT 358.195 27.915 358.525 28.245 ;
        RECT 358.195 26.425 358.525 26.755 ;
        RECT 358.195 24.755 358.525 25.085 ;
        RECT 358.195 23.265 358.525 23.595 ;
        RECT 358.195 21.595 358.525 21.925 ;
        RECT 358.195 20.105 358.525 20.435 ;
        RECT 358.195 18.695 358.525 19.025 ;
        RECT 358.195 16.855 358.525 17.185 ;
        RECT 358.195 15.365 358.525 15.695 ;
        RECT 358.195 13.695 358.525 14.025 ;
        RECT 358.195 12.205 358.525 12.535 ;
        RECT 358.195 10.535 358.525 10.865 ;
        RECT 358.195 9.045 358.525 9.375 ;
        RECT 358.195 7.375 358.525 7.705 ;
        RECT 358.195 5.885 358.525 6.215 ;
        RECT 358.195 4.475 358.525 4.805 ;
        RECT 358.195 2.115 358.525 2.445 ;
        RECT 358.195 0.06 358.525 0.39 ;
        RECT 358.195 -1.525 358.525 -1.195 ;
        RECT 358.195 -2.885 358.525 -2.555 ;
        RECT 358.195 -4.245 358.525 -3.915 ;
        RECT 358.195 -5.605 358.525 -5.275 ;
        RECT 358.195 -6.965 358.525 -6.635 ;
        RECT 358.195 -8.325 358.525 -7.995 ;
        RECT 358.195 -9.685 358.525 -9.355 ;
        RECT 358.195 -11.045 358.525 -10.715 ;
        RECT 358.195 -12.405 358.525 -12.075 ;
        RECT 358.195 -13.765 358.525 -13.435 ;
        RECT 358.195 -15.125 358.525 -14.795 ;
        RECT 358.195 -16.485 358.525 -16.155 ;
        RECT 358.195 -17.845 358.525 -17.515 ;
        RECT 358.195 -19.205 358.525 -18.875 ;
        RECT 358.195 -20.565 358.525 -20.235 ;
        RECT 358.195 -21.925 358.525 -21.595 ;
        RECT 358.195 -23.285 358.525 -22.955 ;
        RECT 358.195 -24.645 358.525 -24.315 ;
        RECT 358.195 -26.005 358.525 -25.675 ;
        RECT 358.195 -27.365 358.525 -27.035 ;
        RECT 358.195 -28.725 358.525 -28.395 ;
        RECT 358.195 -30.085 358.525 -29.755 ;
        RECT 358.195 -31.445 358.525 -31.115 ;
        RECT 358.195 -32.805 358.525 -32.475 ;
        RECT 358.195 -34.165 358.525 -33.835 ;
        RECT 358.195 -35.525 358.525 -35.195 ;
        RECT 358.195 -36.885 358.525 -36.555 ;
        RECT 358.195 -38.245 358.525 -37.915 ;
        RECT 358.195 -39.605 358.525 -39.275 ;
        RECT 358.195 -40.965 358.525 -40.635 ;
        RECT 358.195 -42.325 358.525 -41.995 ;
        RECT 358.195 -43.685 358.525 -43.355 ;
        RECT 358.195 -45.045 358.525 -44.715 ;
        RECT 358.195 -46.405 358.525 -46.075 ;
        RECT 358.195 -47.765 358.525 -47.435 ;
        RECT 358.195 -49.125 358.525 -48.795 ;
        RECT 358.195 -50.485 358.525 -50.155 ;
        RECT 358.195 -51.845 358.525 -51.515 ;
        RECT 358.195 -53.205 358.525 -52.875 ;
        RECT 358.195 -54.565 358.525 -54.235 ;
        RECT 358.195 -55.925 358.525 -55.595 ;
        RECT 358.195 -57.285 358.525 -56.955 ;
        RECT 358.195 -58.645 358.525 -58.315 ;
        RECT 358.195 -60.005 358.525 -59.675 ;
        RECT 358.195 -61.365 358.525 -61.035 ;
        RECT 358.195 -62.725 358.525 -62.395 ;
        RECT 358.195 -64.085 358.525 -63.755 ;
        RECT 358.195 -65.445 358.525 -65.115 ;
        RECT 358.195 -66.805 358.525 -66.475 ;
        RECT 358.195 -68.165 358.525 -67.835 ;
        RECT 358.195 -69.525 358.525 -69.195 ;
        RECT 358.195 -70.885 358.525 -70.555 ;
        RECT 358.195 -72.245 358.525 -71.915 ;
        RECT 358.195 -73.605 358.525 -73.275 ;
        RECT 358.195 -74.965 358.525 -74.635 ;
        RECT 358.195 -76.325 358.525 -75.995 ;
        RECT 358.195 -77.685 358.525 -77.355 ;
        RECT 358.195 -79.045 358.525 -78.715 ;
        RECT 358.195 -80.405 358.525 -80.075 ;
        RECT 358.195 -81.765 358.525 -81.435 ;
        RECT 358.195 -83.125 358.525 -82.795 ;
        RECT 358.195 -84.485 358.525 -84.155 ;
        RECT 358.195 -85.845 358.525 -85.515 ;
        RECT 358.195 -87.205 358.525 -86.875 ;
        RECT 358.195 -88.565 358.525 -88.235 ;
        RECT 358.195 -89.925 358.525 -89.595 ;
        RECT 358.195 -91.285 358.525 -90.955 ;
        RECT 358.195 -92.645 358.525 -92.315 ;
        RECT 358.195 -94.005 358.525 -93.675 ;
        RECT 358.195 -95.365 358.525 -95.035 ;
        RECT 358.195 -96.725 358.525 -96.395 ;
        RECT 358.195 -98.085 358.525 -97.755 ;
        RECT 358.195 -99.445 358.525 -99.115 ;
        RECT 358.195 -100.805 358.525 -100.475 ;
        RECT 358.195 -102.165 358.525 -101.835 ;
        RECT 358.195 -103.525 358.525 -103.195 ;
        RECT 358.195 -104.885 358.525 -104.555 ;
        RECT 358.195 -106.245 358.525 -105.915 ;
        RECT 358.195 -107.605 358.525 -107.275 ;
        RECT 358.195 -108.965 358.525 -108.635 ;
        RECT 358.195 -110.325 358.525 -109.995 ;
        RECT 358.195 -111.685 358.525 -111.355 ;
        RECT 358.195 -113.045 358.525 -112.715 ;
        RECT 358.195 -114.405 358.525 -114.075 ;
        RECT 358.195 -115.765 358.525 -115.435 ;
        RECT 358.195 -117.125 358.525 -116.795 ;
        RECT 358.195 -118.485 358.525 -118.155 ;
        RECT 358.195 -119.845 358.525 -119.515 ;
        RECT 358.195 -121.205 358.525 -120.875 ;
        RECT 358.195 -122.565 358.525 -122.235 ;
        RECT 358.195 -123.925 358.525 -123.595 ;
        RECT 358.195 -125.285 358.525 -124.955 ;
        RECT 358.195 -126.645 358.525 -126.315 ;
        RECT 358.195 -128.005 358.525 -127.675 ;
        RECT 358.195 -129.365 358.525 -129.035 ;
        RECT 358.195 -130.725 358.525 -130.395 ;
        RECT 358.195 -132.085 358.525 -131.755 ;
        RECT 358.195 -133.445 358.525 -133.115 ;
        RECT 358.195 -134.805 358.525 -134.475 ;
        RECT 358.195 -136.165 358.525 -135.835 ;
        RECT 358.195 -137.525 358.525 -137.195 ;
        RECT 358.195 -138.885 358.525 -138.555 ;
        RECT 358.195 -140.245 358.525 -139.915 ;
        RECT 358.195 -141.605 358.525 -141.275 ;
        RECT 358.195 -142.965 358.525 -142.635 ;
        RECT 358.195 -144.325 358.525 -143.995 ;
        RECT 358.195 -145.685 358.525 -145.355 ;
        RECT 358.195 -147.045 358.525 -146.715 ;
        RECT 358.195 -148.405 358.525 -148.075 ;
        RECT 358.195 -149.765 358.525 -149.435 ;
        RECT 358.195 -151.125 358.525 -150.795 ;
        RECT 358.195 -152.485 358.525 -152.155 ;
        RECT 358.195 -153.845 358.525 -153.515 ;
        RECT 358.195 -155.205 358.525 -154.875 ;
        RECT 358.195 -156.565 358.525 -156.235 ;
        RECT 358.195 -157.925 358.525 -157.595 ;
        RECT 358.195 -159.285 358.525 -158.955 ;
        RECT 358.195 -160.645 358.525 -160.315 ;
        RECT 358.195 -162.005 358.525 -161.675 ;
        RECT 358.195 -163.365 358.525 -163.035 ;
        RECT 358.195 -164.725 358.525 -164.395 ;
        RECT 358.195 -166.085 358.525 -165.755 ;
        RECT 358.195 -167.445 358.525 -167.115 ;
        RECT 358.195 -168.805 358.525 -168.475 ;
        RECT 358.195 -170.165 358.525 -169.835 ;
        RECT 358.195 -171.525 358.525 -171.195 ;
        RECT 358.195 -172.885 358.525 -172.555 ;
        RECT 358.195 -174.245 358.525 -173.915 ;
        RECT 358.195 -175.605 358.525 -175.275 ;
        RECT 358.195 -176.965 358.525 -176.635 ;
        RECT 358.195 -178.325 358.525 -177.995 ;
        RECT 358.195 -179.685 358.525 -179.355 ;
        RECT 358.195 -181.93 358.525 -180.8 ;
        RECT 358.2 -182.045 358.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 359.555 241.32 359.885 242.45 ;
        RECT 359.555 239.195 359.885 239.525 ;
        RECT 359.555 237.835 359.885 238.165 ;
        RECT 359.555 235.975 359.885 236.305 ;
        RECT 359.555 233.925 359.885 234.255 ;
        RECT 359.555 231.995 359.885 232.325 ;
        RECT 359.555 230.155 359.885 230.485 ;
        RECT 359.555 228.665 359.885 228.995 ;
        RECT 359.555 226.995 359.885 227.325 ;
        RECT 359.555 225.505 359.885 225.835 ;
        RECT 359.555 223.835 359.885 224.165 ;
        RECT 359.555 222.345 359.885 222.675 ;
        RECT 359.555 220.675 359.885 221.005 ;
        RECT 359.555 219.185 359.885 219.515 ;
        RECT 359.555 217.775 359.885 218.105 ;
        RECT 359.555 215.935 359.885 216.265 ;
        RECT 359.555 214.445 359.885 214.775 ;
        RECT 359.555 212.775 359.885 213.105 ;
        RECT 359.555 211.285 359.885 211.615 ;
        RECT 359.555 209.615 359.885 209.945 ;
        RECT 359.555 208.125 359.885 208.455 ;
        RECT 359.555 206.455 359.885 206.785 ;
        RECT 359.555 204.965 359.885 205.295 ;
        RECT 359.555 203.555 359.885 203.885 ;
        RECT 359.555 201.715 359.885 202.045 ;
        RECT 359.555 200.225 359.885 200.555 ;
        RECT 359.555 198.555 359.885 198.885 ;
        RECT 359.555 197.065 359.885 197.395 ;
        RECT 359.555 195.395 359.885 195.725 ;
        RECT 359.555 193.905 359.885 194.235 ;
        RECT 359.555 192.235 359.885 192.565 ;
        RECT 359.555 190.745 359.885 191.075 ;
        RECT 359.555 189.335 359.885 189.665 ;
        RECT 359.555 187.495 359.885 187.825 ;
        RECT 359.555 186.005 359.885 186.335 ;
        RECT 359.555 184.335 359.885 184.665 ;
        RECT 359.555 182.845 359.885 183.175 ;
        RECT 359.555 181.175 359.885 181.505 ;
        RECT 359.555 179.685 359.885 180.015 ;
        RECT 359.555 178.015 359.885 178.345 ;
        RECT 359.555 176.525 359.885 176.855 ;
        RECT 359.555 175.115 359.885 175.445 ;
        RECT 359.555 173.275 359.885 173.605 ;
        RECT 359.555 171.785 359.885 172.115 ;
        RECT 359.555 170.115 359.885 170.445 ;
        RECT 359.555 168.625 359.885 168.955 ;
        RECT 359.555 166.955 359.885 167.285 ;
        RECT 359.555 165.465 359.885 165.795 ;
        RECT 359.555 163.795 359.885 164.125 ;
        RECT 359.555 162.305 359.885 162.635 ;
        RECT 359.555 160.895 359.885 161.225 ;
        RECT 359.555 159.055 359.885 159.385 ;
        RECT 359.555 157.565 359.885 157.895 ;
        RECT 359.555 155.895 359.885 156.225 ;
        RECT 359.555 154.405 359.885 154.735 ;
        RECT 359.555 152.735 359.885 153.065 ;
        RECT 359.555 151.245 359.885 151.575 ;
        RECT 359.555 149.575 359.885 149.905 ;
        RECT 359.555 148.085 359.885 148.415 ;
        RECT 359.555 146.675 359.885 147.005 ;
        RECT 359.555 144.835 359.885 145.165 ;
        RECT 359.555 143.345 359.885 143.675 ;
        RECT 359.555 141.675 359.885 142.005 ;
        RECT 359.555 140.185 359.885 140.515 ;
        RECT 359.555 138.515 359.885 138.845 ;
        RECT 359.555 137.025 359.885 137.355 ;
        RECT 359.555 135.355 359.885 135.685 ;
        RECT 359.555 133.865 359.885 134.195 ;
        RECT 359.555 132.455 359.885 132.785 ;
        RECT 359.555 130.615 359.885 130.945 ;
        RECT 359.555 129.125 359.885 129.455 ;
        RECT 359.555 127.455 359.885 127.785 ;
        RECT 359.555 125.965 359.885 126.295 ;
        RECT 359.555 124.295 359.885 124.625 ;
        RECT 359.555 122.805 359.885 123.135 ;
        RECT 359.555 121.135 359.885 121.465 ;
        RECT 359.555 119.645 359.885 119.975 ;
        RECT 359.555 118.235 359.885 118.565 ;
        RECT 359.555 116.395 359.885 116.725 ;
        RECT 359.555 114.905 359.885 115.235 ;
        RECT 359.555 113.235 359.885 113.565 ;
        RECT 359.555 111.745 359.885 112.075 ;
        RECT 359.555 110.075 359.885 110.405 ;
        RECT 359.555 108.585 359.885 108.915 ;
        RECT 359.555 106.915 359.885 107.245 ;
        RECT 359.555 105.425 359.885 105.755 ;
        RECT 359.555 104.015 359.885 104.345 ;
        RECT 359.555 102.175 359.885 102.505 ;
        RECT 359.555 100.685 359.885 101.015 ;
        RECT 359.555 99.015 359.885 99.345 ;
        RECT 359.555 97.525 359.885 97.855 ;
        RECT 359.555 95.855 359.885 96.185 ;
        RECT 359.555 94.365 359.885 94.695 ;
        RECT 359.555 92.695 359.885 93.025 ;
        RECT 359.555 91.205 359.885 91.535 ;
        RECT 359.555 89.795 359.885 90.125 ;
        RECT 359.555 87.955 359.885 88.285 ;
        RECT 359.555 86.465 359.885 86.795 ;
        RECT 359.555 84.795 359.885 85.125 ;
        RECT 359.555 83.305 359.885 83.635 ;
        RECT 359.555 81.635 359.885 81.965 ;
        RECT 359.555 80.145 359.885 80.475 ;
        RECT 359.555 78.475 359.885 78.805 ;
        RECT 359.555 76.985 359.885 77.315 ;
        RECT 359.555 75.575 359.885 75.905 ;
        RECT 359.555 73.735 359.885 74.065 ;
        RECT 359.555 72.245 359.885 72.575 ;
        RECT 359.555 70.575 359.885 70.905 ;
        RECT 359.555 69.085 359.885 69.415 ;
        RECT 359.555 67.415 359.885 67.745 ;
        RECT 359.555 65.925 359.885 66.255 ;
        RECT 359.555 64.255 359.885 64.585 ;
        RECT 359.555 62.765 359.885 63.095 ;
        RECT 359.555 61.355 359.885 61.685 ;
        RECT 359.555 59.515 359.885 59.845 ;
        RECT 359.555 58.025 359.885 58.355 ;
        RECT 359.555 56.355 359.885 56.685 ;
        RECT 359.555 54.865 359.885 55.195 ;
        RECT 359.555 53.195 359.885 53.525 ;
        RECT 359.555 51.705 359.885 52.035 ;
        RECT 359.555 50.035 359.885 50.365 ;
        RECT 359.555 48.545 359.885 48.875 ;
        RECT 359.555 47.135 359.885 47.465 ;
        RECT 359.555 45.295 359.885 45.625 ;
        RECT 359.555 43.805 359.885 44.135 ;
        RECT 359.555 42.135 359.885 42.465 ;
        RECT 359.555 40.645 359.885 40.975 ;
        RECT 359.555 38.975 359.885 39.305 ;
        RECT 359.555 37.485 359.885 37.815 ;
        RECT 359.555 35.815 359.885 36.145 ;
        RECT 359.555 34.325 359.885 34.655 ;
        RECT 359.555 32.915 359.885 33.245 ;
        RECT 359.555 31.075 359.885 31.405 ;
        RECT 359.555 29.585 359.885 29.915 ;
        RECT 359.555 27.915 359.885 28.245 ;
        RECT 359.555 26.425 359.885 26.755 ;
        RECT 359.555 24.755 359.885 25.085 ;
        RECT 359.555 23.265 359.885 23.595 ;
        RECT 359.555 21.595 359.885 21.925 ;
        RECT 359.555 20.105 359.885 20.435 ;
        RECT 359.555 18.695 359.885 19.025 ;
        RECT 359.555 16.855 359.885 17.185 ;
        RECT 359.555 15.365 359.885 15.695 ;
        RECT 359.555 13.695 359.885 14.025 ;
        RECT 359.555 12.205 359.885 12.535 ;
        RECT 359.555 10.535 359.885 10.865 ;
        RECT 359.555 9.045 359.885 9.375 ;
        RECT 359.555 7.375 359.885 7.705 ;
        RECT 359.555 5.885 359.885 6.215 ;
        RECT 359.555 4.475 359.885 4.805 ;
        RECT 359.555 2.115 359.885 2.445 ;
        RECT 359.555 0.06 359.885 0.39 ;
        RECT 359.555 -1.525 359.885 -1.195 ;
        RECT 359.555 -2.885 359.885 -2.555 ;
        RECT 359.555 -4.245 359.885 -3.915 ;
        RECT 359.555 -5.605 359.885 -5.275 ;
        RECT 359.555 -6.965 359.885 -6.635 ;
        RECT 359.555 -8.325 359.885 -7.995 ;
        RECT 359.555 -9.685 359.885 -9.355 ;
        RECT 359.555 -11.045 359.885 -10.715 ;
        RECT 359.555 -12.405 359.885 -12.075 ;
        RECT 359.555 -13.765 359.885 -13.435 ;
        RECT 359.555 -15.125 359.885 -14.795 ;
        RECT 359.555 -16.485 359.885 -16.155 ;
        RECT 359.555 -17.845 359.885 -17.515 ;
        RECT 359.555 -19.205 359.885 -18.875 ;
        RECT 359.555 -20.565 359.885 -20.235 ;
        RECT 359.555 -21.925 359.885 -21.595 ;
        RECT 359.555 -23.285 359.885 -22.955 ;
        RECT 359.555 -24.645 359.885 -24.315 ;
        RECT 359.555 -26.005 359.885 -25.675 ;
        RECT 359.555 -27.365 359.885 -27.035 ;
        RECT 359.555 -28.725 359.885 -28.395 ;
        RECT 359.555 -30.085 359.885 -29.755 ;
        RECT 359.555 -31.445 359.885 -31.115 ;
        RECT 359.555 -32.805 359.885 -32.475 ;
        RECT 359.555 -34.165 359.885 -33.835 ;
        RECT 359.555 -35.525 359.885 -35.195 ;
        RECT 359.555 -36.885 359.885 -36.555 ;
        RECT 359.555 -38.245 359.885 -37.915 ;
        RECT 359.555 -39.605 359.885 -39.275 ;
        RECT 359.555 -40.965 359.885 -40.635 ;
        RECT 359.555 -42.325 359.885 -41.995 ;
        RECT 359.555 -43.685 359.885 -43.355 ;
        RECT 359.555 -45.045 359.885 -44.715 ;
        RECT 359.555 -46.405 359.885 -46.075 ;
        RECT 359.555 -47.765 359.885 -47.435 ;
        RECT 359.555 -49.125 359.885 -48.795 ;
        RECT 359.555 -50.485 359.885 -50.155 ;
        RECT 359.555 -51.845 359.885 -51.515 ;
        RECT 359.555 -53.205 359.885 -52.875 ;
        RECT 359.555 -54.565 359.885 -54.235 ;
        RECT 359.555 -55.925 359.885 -55.595 ;
        RECT 359.555 -57.285 359.885 -56.955 ;
        RECT 359.555 -58.645 359.885 -58.315 ;
        RECT 359.555 -60.005 359.885 -59.675 ;
        RECT 359.555 -61.365 359.885 -61.035 ;
        RECT 359.555 -62.725 359.885 -62.395 ;
        RECT 359.555 -64.085 359.885 -63.755 ;
        RECT 359.555 -65.445 359.885 -65.115 ;
        RECT 359.555 -66.805 359.885 -66.475 ;
        RECT 359.555 -68.165 359.885 -67.835 ;
        RECT 359.555 -69.525 359.885 -69.195 ;
        RECT 359.555 -70.885 359.885 -70.555 ;
        RECT 359.555 -72.245 359.885 -71.915 ;
        RECT 359.555 -73.605 359.885 -73.275 ;
        RECT 359.555 -74.965 359.885 -74.635 ;
        RECT 359.555 -76.325 359.885 -75.995 ;
        RECT 359.555 -77.685 359.885 -77.355 ;
        RECT 359.555 -79.045 359.885 -78.715 ;
        RECT 359.555 -80.405 359.885 -80.075 ;
        RECT 359.555 -81.765 359.885 -81.435 ;
        RECT 359.555 -83.125 359.885 -82.795 ;
        RECT 359.555 -84.485 359.885 -84.155 ;
        RECT 359.555 -85.845 359.885 -85.515 ;
        RECT 359.555 -87.205 359.885 -86.875 ;
        RECT 359.555 -88.565 359.885 -88.235 ;
        RECT 359.555 -89.925 359.885 -89.595 ;
        RECT 359.555 -91.285 359.885 -90.955 ;
        RECT 359.555 -92.645 359.885 -92.315 ;
        RECT 359.555 -94.005 359.885 -93.675 ;
        RECT 359.555 -95.365 359.885 -95.035 ;
        RECT 359.555 -96.725 359.885 -96.395 ;
        RECT 359.555 -98.085 359.885 -97.755 ;
        RECT 359.555 -99.445 359.885 -99.115 ;
        RECT 359.555 -100.805 359.885 -100.475 ;
        RECT 359.555 -102.165 359.885 -101.835 ;
        RECT 359.555 -103.525 359.885 -103.195 ;
        RECT 359.555 -104.885 359.885 -104.555 ;
        RECT 359.555 -106.245 359.885 -105.915 ;
        RECT 359.555 -107.605 359.885 -107.275 ;
        RECT 359.555 -108.965 359.885 -108.635 ;
        RECT 359.555 -110.325 359.885 -109.995 ;
        RECT 359.555 -111.685 359.885 -111.355 ;
        RECT 359.555 -113.045 359.885 -112.715 ;
        RECT 359.555 -114.405 359.885 -114.075 ;
        RECT 359.555 -115.765 359.885 -115.435 ;
        RECT 359.555 -117.125 359.885 -116.795 ;
        RECT 359.555 -118.485 359.885 -118.155 ;
        RECT 359.555 -119.845 359.885 -119.515 ;
        RECT 359.555 -121.205 359.885 -120.875 ;
        RECT 359.555 -122.565 359.885 -122.235 ;
        RECT 359.555 -123.925 359.885 -123.595 ;
        RECT 359.555 -125.285 359.885 -124.955 ;
        RECT 359.555 -126.645 359.885 -126.315 ;
        RECT 359.555 -128.005 359.885 -127.675 ;
        RECT 359.555 -129.365 359.885 -129.035 ;
        RECT 359.555 -130.725 359.885 -130.395 ;
        RECT 359.555 -132.085 359.885 -131.755 ;
        RECT 359.555 -133.445 359.885 -133.115 ;
        RECT 359.555 -134.805 359.885 -134.475 ;
        RECT 359.555 -136.165 359.885 -135.835 ;
        RECT 359.555 -137.525 359.885 -137.195 ;
        RECT 359.555 -138.885 359.885 -138.555 ;
        RECT 359.555 -140.245 359.885 -139.915 ;
        RECT 359.555 -141.605 359.885 -141.275 ;
        RECT 359.555 -142.965 359.885 -142.635 ;
        RECT 359.555 -144.325 359.885 -143.995 ;
        RECT 359.555 -145.685 359.885 -145.355 ;
        RECT 359.555 -147.045 359.885 -146.715 ;
        RECT 359.555 -148.405 359.885 -148.075 ;
        RECT 359.555 -149.765 359.885 -149.435 ;
        RECT 359.555 -151.125 359.885 -150.795 ;
        RECT 359.555 -152.485 359.885 -152.155 ;
        RECT 359.555 -153.845 359.885 -153.515 ;
        RECT 359.555 -155.205 359.885 -154.875 ;
        RECT 359.555 -156.565 359.885 -156.235 ;
        RECT 359.555 -157.925 359.885 -157.595 ;
        RECT 359.555 -159.285 359.885 -158.955 ;
        RECT 359.555 -160.645 359.885 -160.315 ;
        RECT 359.555 -162.005 359.885 -161.675 ;
        RECT 359.555 -163.365 359.885 -163.035 ;
        RECT 359.555 -164.725 359.885 -164.395 ;
        RECT 359.555 -166.085 359.885 -165.755 ;
        RECT 359.555 -167.445 359.885 -167.115 ;
        RECT 359.555 -168.805 359.885 -168.475 ;
        RECT 359.555 -170.165 359.885 -169.835 ;
        RECT 359.555 -171.525 359.885 -171.195 ;
        RECT 359.555 -172.885 359.885 -172.555 ;
        RECT 359.555 -174.245 359.885 -173.915 ;
        RECT 359.555 -175.605 359.885 -175.275 ;
        RECT 359.555 -176.965 359.885 -176.635 ;
        RECT 359.555 -178.325 359.885 -177.995 ;
        RECT 359.555 -179.685 359.885 -179.355 ;
        RECT 359.555 -181.93 359.885 -180.8 ;
        RECT 359.56 -182.045 359.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 360.915 241.32 361.245 242.45 ;
        RECT 360.915 239.195 361.245 239.525 ;
        RECT 360.915 237.835 361.245 238.165 ;
        RECT 360.915 -1.525 361.245 -1.195 ;
        RECT 360.915 -2.885 361.245 -2.555 ;
        RECT 360.915 -4.245 361.245 -3.915 ;
        RECT 360.915 -5.605 361.245 -5.275 ;
        RECT 360.915 -6.965 361.245 -6.635 ;
        RECT 360.915 -8.325 361.245 -7.995 ;
        RECT 360.915 -9.685 361.245 -9.355 ;
        RECT 360.915 -11.045 361.245 -10.715 ;
        RECT 360.915 -12.405 361.245 -12.075 ;
        RECT 360.915 -13.765 361.245 -13.435 ;
        RECT 360.915 -15.125 361.245 -14.795 ;
        RECT 360.915 -16.485 361.245 -16.155 ;
        RECT 360.915 -17.845 361.245 -17.515 ;
        RECT 360.915 -19.205 361.245 -18.875 ;
        RECT 360.915 -20.565 361.245 -20.235 ;
        RECT 360.915 -21.925 361.245 -21.595 ;
        RECT 360.915 -23.285 361.245 -22.955 ;
        RECT 360.915 -24.645 361.245 -24.315 ;
        RECT 360.915 -26.005 361.245 -25.675 ;
        RECT 360.915 -27.365 361.245 -27.035 ;
        RECT 360.915 -28.725 361.245 -28.395 ;
        RECT 360.915 -30.085 361.245 -29.755 ;
        RECT 360.915 -31.445 361.245 -31.115 ;
        RECT 360.915 -32.805 361.245 -32.475 ;
        RECT 360.915 -34.165 361.245 -33.835 ;
        RECT 360.915 -35.525 361.245 -35.195 ;
        RECT 360.915 -36.885 361.245 -36.555 ;
        RECT 360.915 -38.245 361.245 -37.915 ;
        RECT 360.915 -39.605 361.245 -39.275 ;
        RECT 360.915 -40.965 361.245 -40.635 ;
        RECT 360.915 -42.325 361.245 -41.995 ;
        RECT 360.915 -43.685 361.245 -43.355 ;
        RECT 360.915 -45.045 361.245 -44.715 ;
        RECT 360.915 -46.405 361.245 -46.075 ;
        RECT 360.915 -47.765 361.245 -47.435 ;
        RECT 360.915 -49.125 361.245 -48.795 ;
        RECT 360.915 -50.485 361.245 -50.155 ;
        RECT 360.915 -51.845 361.245 -51.515 ;
        RECT 360.915 -53.205 361.245 -52.875 ;
        RECT 360.915 -54.565 361.245 -54.235 ;
        RECT 360.915 -55.925 361.245 -55.595 ;
        RECT 360.915 -57.285 361.245 -56.955 ;
        RECT 360.915 -58.645 361.245 -58.315 ;
        RECT 360.915 -60.005 361.245 -59.675 ;
        RECT 360.915 -61.365 361.245 -61.035 ;
        RECT 360.915 -62.725 361.245 -62.395 ;
        RECT 360.915 -64.085 361.245 -63.755 ;
        RECT 360.915 -65.445 361.245 -65.115 ;
        RECT 360.915 -66.805 361.245 -66.475 ;
        RECT 360.915 -68.165 361.245 -67.835 ;
        RECT 360.915 -69.525 361.245 -69.195 ;
        RECT 360.915 -70.885 361.245 -70.555 ;
        RECT 360.915 -72.245 361.245 -71.915 ;
        RECT 360.915 -73.605 361.245 -73.275 ;
        RECT 360.915 -74.965 361.245 -74.635 ;
        RECT 360.915 -76.325 361.245 -75.995 ;
        RECT 360.915 -77.685 361.245 -77.355 ;
        RECT 360.915 -79.045 361.245 -78.715 ;
        RECT 360.915 -80.405 361.245 -80.075 ;
        RECT 360.915 -81.765 361.245 -81.435 ;
        RECT 360.915 -83.125 361.245 -82.795 ;
        RECT 360.915 -84.485 361.245 -84.155 ;
        RECT 360.915 -85.845 361.245 -85.515 ;
        RECT 360.915 -87.205 361.245 -86.875 ;
        RECT 360.915 -88.565 361.245 -88.235 ;
        RECT 360.915 -89.925 361.245 -89.595 ;
        RECT 360.915 -91.285 361.245 -90.955 ;
        RECT 360.915 -92.645 361.245 -92.315 ;
        RECT 360.915 -94.005 361.245 -93.675 ;
        RECT 360.915 -95.365 361.245 -95.035 ;
        RECT 360.915 -96.725 361.245 -96.395 ;
        RECT 360.915 -98.085 361.245 -97.755 ;
        RECT 360.915 -99.445 361.245 -99.115 ;
        RECT 360.915 -100.805 361.245 -100.475 ;
        RECT 360.915 -102.165 361.245 -101.835 ;
        RECT 360.915 -103.525 361.245 -103.195 ;
        RECT 360.915 -104.885 361.245 -104.555 ;
        RECT 360.915 -106.245 361.245 -105.915 ;
        RECT 360.915 -107.605 361.245 -107.275 ;
        RECT 360.915 -108.965 361.245 -108.635 ;
        RECT 360.915 -110.325 361.245 -109.995 ;
        RECT 360.915 -111.685 361.245 -111.355 ;
        RECT 360.915 -113.045 361.245 -112.715 ;
        RECT 360.915 -114.405 361.245 -114.075 ;
        RECT 360.915 -115.765 361.245 -115.435 ;
        RECT 360.915 -117.125 361.245 -116.795 ;
        RECT 360.915 -118.485 361.245 -118.155 ;
        RECT 360.915 -119.845 361.245 -119.515 ;
        RECT 360.915 -121.205 361.245 -120.875 ;
        RECT 360.915 -122.565 361.245 -122.235 ;
        RECT 360.915 -123.925 361.245 -123.595 ;
        RECT 360.915 -125.285 361.245 -124.955 ;
        RECT 360.915 -126.645 361.245 -126.315 ;
        RECT 360.915 -128.005 361.245 -127.675 ;
        RECT 360.915 -129.365 361.245 -129.035 ;
        RECT 360.915 -130.725 361.245 -130.395 ;
        RECT 360.915 -132.085 361.245 -131.755 ;
        RECT 360.915 -133.445 361.245 -133.115 ;
        RECT 360.915 -134.805 361.245 -134.475 ;
        RECT 360.915 -136.165 361.245 -135.835 ;
        RECT 360.915 -137.525 361.245 -137.195 ;
        RECT 360.915 -138.885 361.245 -138.555 ;
        RECT 360.915 -140.245 361.245 -139.915 ;
        RECT 360.915 -141.605 361.245 -141.275 ;
        RECT 360.915 -142.965 361.245 -142.635 ;
        RECT 360.915 -144.325 361.245 -143.995 ;
        RECT 360.915 -145.685 361.245 -145.355 ;
        RECT 360.915 -147.045 361.245 -146.715 ;
        RECT 360.915 -148.405 361.245 -148.075 ;
        RECT 360.915 -149.765 361.245 -149.435 ;
        RECT 360.915 -151.125 361.245 -150.795 ;
        RECT 360.915 -152.485 361.245 -152.155 ;
        RECT 360.915 -153.845 361.245 -153.515 ;
        RECT 360.915 -155.205 361.245 -154.875 ;
        RECT 360.915 -156.565 361.245 -156.235 ;
        RECT 360.915 -157.925 361.245 -157.595 ;
        RECT 360.915 -159.285 361.245 -158.955 ;
        RECT 360.915 -160.645 361.245 -160.315 ;
        RECT 360.915 -162.005 361.245 -161.675 ;
        RECT 360.915 -163.365 361.245 -163.035 ;
        RECT 360.915 -164.725 361.245 -164.395 ;
        RECT 360.915 -166.085 361.245 -165.755 ;
        RECT 360.915 -167.445 361.245 -167.115 ;
        RECT 360.915 -168.805 361.245 -168.475 ;
        RECT 360.915 -170.165 361.245 -169.835 ;
        RECT 360.915 -171.525 361.245 -171.195 ;
        RECT 360.915 -172.885 361.245 -172.555 ;
        RECT 360.915 -174.245 361.245 -173.915 ;
        RECT 360.915 -175.605 361.245 -175.275 ;
        RECT 360.915 -176.965 361.245 -176.635 ;
        RECT 360.915 -178.325 361.245 -177.995 ;
        RECT 360.915 -179.685 361.245 -179.355 ;
        RECT 360.915 -181.93 361.245 -180.8 ;
        RECT 360.92 -182.045 361.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 241.32 339.485 242.45 ;
        RECT 339.155 239.195 339.485 239.525 ;
        RECT 339.155 237.835 339.485 238.165 ;
        RECT 339.16 237.16 339.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 -1.525 339.485 -1.195 ;
        RECT 339.155 -2.885 339.485 -2.555 ;
        RECT 339.16 -3.56 339.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 339.155 -95.365 339.485 -95.035 ;
        RECT 339.155 -96.725 339.485 -96.395 ;
        RECT 339.155 -98.085 339.485 -97.755 ;
        RECT 339.155 -99.445 339.485 -99.115 ;
        RECT 339.155 -100.805 339.485 -100.475 ;
        RECT 339.155 -102.165 339.485 -101.835 ;
        RECT 339.155 -103.525 339.485 -103.195 ;
        RECT 339.155 -104.885 339.485 -104.555 ;
        RECT 339.155 -106.245 339.485 -105.915 ;
        RECT 339.155 -107.605 339.485 -107.275 ;
        RECT 339.155 -108.965 339.485 -108.635 ;
        RECT 339.155 -110.325 339.485 -109.995 ;
        RECT 339.155 -111.685 339.485 -111.355 ;
        RECT 339.155 -113.045 339.485 -112.715 ;
        RECT 339.155 -114.405 339.485 -114.075 ;
        RECT 339.155 -115.765 339.485 -115.435 ;
        RECT 339.155 -117.125 339.485 -116.795 ;
        RECT 339.155 -118.485 339.485 -118.155 ;
        RECT 339.155 -119.845 339.485 -119.515 ;
        RECT 339.155 -121.205 339.485 -120.875 ;
        RECT 339.155 -122.565 339.485 -122.235 ;
        RECT 339.155 -123.925 339.485 -123.595 ;
        RECT 339.155 -125.285 339.485 -124.955 ;
        RECT 339.155 -126.645 339.485 -126.315 ;
        RECT 339.155 -128.005 339.485 -127.675 ;
        RECT 339.155 -129.365 339.485 -129.035 ;
        RECT 339.155 -130.725 339.485 -130.395 ;
        RECT 339.155 -132.085 339.485 -131.755 ;
        RECT 339.155 -133.445 339.485 -133.115 ;
        RECT 339.155 -134.805 339.485 -134.475 ;
        RECT 339.155 -136.165 339.485 -135.835 ;
        RECT 339.155 -137.525 339.485 -137.195 ;
        RECT 339.155 -138.885 339.485 -138.555 ;
        RECT 339.155 -140.245 339.485 -139.915 ;
        RECT 339.155 -141.605 339.485 -141.275 ;
        RECT 339.155 -142.965 339.485 -142.635 ;
        RECT 339.155 -144.325 339.485 -143.995 ;
        RECT 339.155 -145.685 339.485 -145.355 ;
        RECT 339.155 -147.045 339.485 -146.715 ;
        RECT 339.155 -148.405 339.485 -148.075 ;
        RECT 339.155 -149.765 339.485 -149.435 ;
        RECT 339.155 -151.125 339.485 -150.795 ;
        RECT 339.155 -152.485 339.485 -152.155 ;
        RECT 339.155 -153.845 339.485 -153.515 ;
        RECT 339.155 -155.205 339.485 -154.875 ;
        RECT 339.155 -156.565 339.485 -156.235 ;
        RECT 339.155 -157.925 339.485 -157.595 ;
        RECT 339.155 -159.285 339.485 -158.955 ;
        RECT 339.155 -160.645 339.485 -160.315 ;
        RECT 339.155 -162.005 339.485 -161.675 ;
        RECT 339.155 -163.365 339.485 -163.035 ;
        RECT 339.155 -164.725 339.485 -164.395 ;
        RECT 339.155 -166.085 339.485 -165.755 ;
        RECT 339.155 -167.445 339.485 -167.115 ;
        RECT 339.155 -168.805 339.485 -168.475 ;
        RECT 339.155 -170.165 339.485 -169.835 ;
        RECT 339.155 -171.525 339.485 -171.195 ;
        RECT 339.155 -172.885 339.485 -172.555 ;
        RECT 339.155 -174.245 339.485 -173.915 ;
        RECT 339.155 -175.605 339.485 -175.275 ;
        RECT 339.155 -176.965 339.485 -176.635 ;
        RECT 339.155 -178.325 339.485 -177.995 ;
        RECT 339.155 -179.685 339.485 -179.355 ;
        RECT 339.155 -181.93 339.485 -180.8 ;
        RECT 339.16 -182.045 339.48 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.515 241.32 340.845 242.45 ;
        RECT 340.515 239.195 340.845 239.525 ;
        RECT 340.515 237.835 340.845 238.165 ;
        RECT 340.52 237.16 340.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 340.515 -99.445 340.845 -99.115 ;
        RECT 340.515 -100.805 340.845 -100.475 ;
        RECT 340.515 -102.165 340.845 -101.835 ;
        RECT 340.515 -103.525 340.845 -103.195 ;
        RECT 340.515 -104.885 340.845 -104.555 ;
        RECT 340.515 -106.245 340.845 -105.915 ;
        RECT 340.515 -107.605 340.845 -107.275 ;
        RECT 340.515 -108.965 340.845 -108.635 ;
        RECT 340.515 -110.325 340.845 -109.995 ;
        RECT 340.515 -111.685 340.845 -111.355 ;
        RECT 340.515 -113.045 340.845 -112.715 ;
        RECT 340.515 -114.405 340.845 -114.075 ;
        RECT 340.515 -115.765 340.845 -115.435 ;
        RECT 340.515 -117.125 340.845 -116.795 ;
        RECT 340.515 -118.485 340.845 -118.155 ;
        RECT 340.515 -119.845 340.845 -119.515 ;
        RECT 340.515 -121.205 340.845 -120.875 ;
        RECT 340.515 -122.565 340.845 -122.235 ;
        RECT 340.515 -123.925 340.845 -123.595 ;
        RECT 340.515 -125.285 340.845 -124.955 ;
        RECT 340.515 -126.645 340.845 -126.315 ;
        RECT 340.515 -128.005 340.845 -127.675 ;
        RECT 340.515 -129.365 340.845 -129.035 ;
        RECT 340.515 -130.725 340.845 -130.395 ;
        RECT 340.515 -132.085 340.845 -131.755 ;
        RECT 340.515 -133.445 340.845 -133.115 ;
        RECT 340.515 -134.805 340.845 -134.475 ;
        RECT 340.515 -136.165 340.845 -135.835 ;
        RECT 340.515 -137.525 340.845 -137.195 ;
        RECT 340.515 -138.885 340.845 -138.555 ;
        RECT 340.515 -140.245 340.845 -139.915 ;
        RECT 340.515 -141.605 340.845 -141.275 ;
        RECT 340.515 -142.965 340.845 -142.635 ;
        RECT 340.515 -144.325 340.845 -143.995 ;
        RECT 340.515 -145.685 340.845 -145.355 ;
        RECT 340.515 -147.045 340.845 -146.715 ;
        RECT 340.515 -148.405 340.845 -148.075 ;
        RECT 340.515 -149.765 340.845 -149.435 ;
        RECT 340.515 -151.125 340.845 -150.795 ;
        RECT 340.515 -152.485 340.845 -152.155 ;
        RECT 340.515 -153.845 340.845 -153.515 ;
        RECT 340.515 -155.205 340.845 -154.875 ;
        RECT 340.515 -156.565 340.845 -156.235 ;
        RECT 340.515 -157.925 340.845 -157.595 ;
        RECT 340.515 -159.285 340.845 -158.955 ;
        RECT 340.515 -160.645 340.845 -160.315 ;
        RECT 340.515 -162.005 340.845 -161.675 ;
        RECT 340.515 -163.365 340.845 -163.035 ;
        RECT 340.515 -164.725 340.845 -164.395 ;
        RECT 340.515 -166.085 340.845 -165.755 ;
        RECT 340.515 -167.445 340.845 -167.115 ;
        RECT 340.515 -168.805 340.845 -168.475 ;
        RECT 340.515 -170.165 340.845 -169.835 ;
        RECT 340.515 -171.525 340.845 -171.195 ;
        RECT 340.515 -172.885 340.845 -172.555 ;
        RECT 340.515 -174.245 340.845 -173.915 ;
        RECT 340.515 -175.605 340.845 -175.275 ;
        RECT 340.515 -176.965 340.845 -176.635 ;
        RECT 340.515 -178.325 340.845 -177.995 ;
        RECT 340.515 -179.685 340.845 -179.355 ;
        RECT 340.515 -181.93 340.845 -180.8 ;
        RECT 340.52 -182.045 340.84 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.21 -98.075 341.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 341.875 241.32 342.205 242.45 ;
        RECT 341.875 239.195 342.205 239.525 ;
        RECT 341.875 237.835 342.205 238.165 ;
        RECT 341.88 237.16 342.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.235 241.32 343.565 242.45 ;
        RECT 343.235 239.195 343.565 239.525 ;
        RECT 343.235 237.835 343.565 238.165 ;
        RECT 343.24 237.16 343.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 343.235 -1.525 343.565 -1.195 ;
        RECT 343.235 -2.885 343.565 -2.555 ;
        RECT 343.24 -3.56 343.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.595 241.32 344.925 242.45 ;
        RECT 344.595 239.195 344.925 239.525 ;
        RECT 344.595 237.835 344.925 238.165 ;
        RECT 344.6 237.16 344.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.595 -1.525 344.925 -1.195 ;
        RECT 344.595 -2.885 344.925 -2.555 ;
        RECT 344.6 -3.56 344.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 344.595 -95.365 344.925 -95.035 ;
        RECT 344.595 -96.725 344.925 -96.395 ;
        RECT 344.595 -98.085 344.925 -97.755 ;
        RECT 344.595 -99.445 344.925 -99.115 ;
        RECT 344.595 -100.805 344.925 -100.475 ;
        RECT 344.595 -102.165 344.925 -101.835 ;
        RECT 344.595 -103.525 344.925 -103.195 ;
        RECT 344.595 -104.885 344.925 -104.555 ;
        RECT 344.595 -106.245 344.925 -105.915 ;
        RECT 344.595 -107.605 344.925 -107.275 ;
        RECT 344.595 -108.965 344.925 -108.635 ;
        RECT 344.595 -110.325 344.925 -109.995 ;
        RECT 344.595 -111.685 344.925 -111.355 ;
        RECT 344.595 -113.045 344.925 -112.715 ;
        RECT 344.595 -114.405 344.925 -114.075 ;
        RECT 344.595 -115.765 344.925 -115.435 ;
        RECT 344.595 -117.125 344.925 -116.795 ;
        RECT 344.595 -118.485 344.925 -118.155 ;
        RECT 344.595 -119.845 344.925 -119.515 ;
        RECT 344.595 -121.205 344.925 -120.875 ;
        RECT 344.595 -122.565 344.925 -122.235 ;
        RECT 344.595 -123.925 344.925 -123.595 ;
        RECT 344.595 -125.285 344.925 -124.955 ;
        RECT 344.595 -126.645 344.925 -126.315 ;
        RECT 344.595 -128.005 344.925 -127.675 ;
        RECT 344.595 -129.365 344.925 -129.035 ;
        RECT 344.595 -130.725 344.925 -130.395 ;
        RECT 344.595 -132.085 344.925 -131.755 ;
        RECT 344.595 -133.445 344.925 -133.115 ;
        RECT 344.595 -134.805 344.925 -134.475 ;
        RECT 344.595 -136.165 344.925 -135.835 ;
        RECT 344.595 -137.525 344.925 -137.195 ;
        RECT 344.595 -138.885 344.925 -138.555 ;
        RECT 344.595 -140.245 344.925 -139.915 ;
        RECT 344.595 -141.605 344.925 -141.275 ;
        RECT 344.595 -142.965 344.925 -142.635 ;
        RECT 344.595 -144.325 344.925 -143.995 ;
        RECT 344.595 -145.685 344.925 -145.355 ;
        RECT 344.595 -147.045 344.925 -146.715 ;
        RECT 344.595 -148.405 344.925 -148.075 ;
        RECT 344.595 -149.765 344.925 -149.435 ;
        RECT 344.595 -151.125 344.925 -150.795 ;
        RECT 344.595 -152.485 344.925 -152.155 ;
        RECT 344.595 -153.845 344.925 -153.515 ;
        RECT 344.595 -155.205 344.925 -154.875 ;
        RECT 344.595 -156.565 344.925 -156.235 ;
        RECT 344.595 -157.925 344.925 -157.595 ;
        RECT 344.595 -159.285 344.925 -158.955 ;
        RECT 344.595 -160.645 344.925 -160.315 ;
        RECT 344.595 -162.005 344.925 -161.675 ;
        RECT 344.595 -163.365 344.925 -163.035 ;
        RECT 344.595 -164.725 344.925 -164.395 ;
        RECT 344.595 -166.085 344.925 -165.755 ;
        RECT 344.595 -167.445 344.925 -167.115 ;
        RECT 344.595 -168.805 344.925 -168.475 ;
        RECT 344.595 -170.165 344.925 -169.835 ;
        RECT 344.595 -171.525 344.925 -171.195 ;
        RECT 344.595 -172.885 344.925 -172.555 ;
        RECT 344.595 -174.245 344.925 -173.915 ;
        RECT 344.595 -175.605 344.925 -175.275 ;
        RECT 344.595 -176.965 344.925 -176.635 ;
        RECT 344.595 -178.325 344.925 -177.995 ;
        RECT 344.595 -179.685 344.925 -179.355 ;
        RECT 344.595 -181.93 344.925 -180.8 ;
        RECT 344.6 -182.045 344.92 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.955 241.32 346.285 242.45 ;
        RECT 345.955 239.195 346.285 239.525 ;
        RECT 345.955 237.835 346.285 238.165 ;
        RECT 345.96 237.16 346.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.955 -1.525 346.285 -1.195 ;
        RECT 345.955 -2.885 346.285 -2.555 ;
        RECT 345.96 -3.56 346.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 345.955 -95.365 346.285 -95.035 ;
        RECT 345.955 -96.725 346.285 -96.395 ;
        RECT 345.955 -98.085 346.285 -97.755 ;
        RECT 345.955 -99.445 346.285 -99.115 ;
        RECT 345.955 -100.805 346.285 -100.475 ;
        RECT 345.955 -102.165 346.285 -101.835 ;
        RECT 345.955 -103.525 346.285 -103.195 ;
        RECT 345.955 -104.885 346.285 -104.555 ;
        RECT 345.955 -106.245 346.285 -105.915 ;
        RECT 345.955 -107.605 346.285 -107.275 ;
        RECT 345.955 -108.965 346.285 -108.635 ;
        RECT 345.955 -110.325 346.285 -109.995 ;
        RECT 345.955 -111.685 346.285 -111.355 ;
        RECT 345.955 -113.045 346.285 -112.715 ;
        RECT 345.955 -114.405 346.285 -114.075 ;
        RECT 345.955 -115.765 346.285 -115.435 ;
        RECT 345.955 -117.125 346.285 -116.795 ;
        RECT 345.955 -118.485 346.285 -118.155 ;
        RECT 345.955 -119.845 346.285 -119.515 ;
        RECT 345.955 -121.205 346.285 -120.875 ;
        RECT 345.955 -122.565 346.285 -122.235 ;
        RECT 345.955 -123.925 346.285 -123.595 ;
        RECT 345.955 -125.285 346.285 -124.955 ;
        RECT 345.955 -126.645 346.285 -126.315 ;
        RECT 345.955 -128.005 346.285 -127.675 ;
        RECT 345.955 -129.365 346.285 -129.035 ;
        RECT 345.955 -130.725 346.285 -130.395 ;
        RECT 345.955 -132.085 346.285 -131.755 ;
        RECT 345.955 -133.445 346.285 -133.115 ;
        RECT 345.955 -134.805 346.285 -134.475 ;
        RECT 345.955 -136.165 346.285 -135.835 ;
        RECT 345.955 -137.525 346.285 -137.195 ;
        RECT 345.955 -138.885 346.285 -138.555 ;
        RECT 345.955 -140.245 346.285 -139.915 ;
        RECT 345.955 -141.605 346.285 -141.275 ;
        RECT 345.955 -142.965 346.285 -142.635 ;
        RECT 345.955 -144.325 346.285 -143.995 ;
        RECT 345.955 -145.685 346.285 -145.355 ;
        RECT 345.955 -147.045 346.285 -146.715 ;
        RECT 345.955 -148.405 346.285 -148.075 ;
        RECT 345.955 -149.765 346.285 -149.435 ;
        RECT 345.955 -151.125 346.285 -150.795 ;
        RECT 345.955 -152.485 346.285 -152.155 ;
        RECT 345.955 -153.845 346.285 -153.515 ;
        RECT 345.955 -155.205 346.285 -154.875 ;
        RECT 345.955 -156.565 346.285 -156.235 ;
        RECT 345.955 -157.925 346.285 -157.595 ;
        RECT 345.955 -159.285 346.285 -158.955 ;
        RECT 345.955 -160.645 346.285 -160.315 ;
        RECT 345.955 -162.005 346.285 -161.675 ;
        RECT 345.955 -163.365 346.285 -163.035 ;
        RECT 345.955 -164.725 346.285 -164.395 ;
        RECT 345.955 -166.085 346.285 -165.755 ;
        RECT 345.955 -167.445 346.285 -167.115 ;
        RECT 345.955 -168.805 346.285 -168.475 ;
        RECT 345.955 -170.165 346.285 -169.835 ;
        RECT 345.955 -171.525 346.285 -171.195 ;
        RECT 345.955 -172.885 346.285 -172.555 ;
        RECT 345.955 -174.245 346.285 -173.915 ;
        RECT 345.955 -175.605 346.285 -175.275 ;
        RECT 345.955 -176.965 346.285 -176.635 ;
        RECT 345.955 -178.325 346.285 -177.995 ;
        RECT 345.955 -179.685 346.285 -179.355 ;
        RECT 345.955 -181.93 346.285 -180.8 ;
        RECT 345.96 -182.045 346.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.315 241.32 347.645 242.45 ;
        RECT 347.315 239.195 347.645 239.525 ;
        RECT 347.315 237.835 347.645 238.165 ;
        RECT 347.32 237.16 347.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.315 -1.525 347.645 -1.195 ;
        RECT 347.315 -2.885 347.645 -2.555 ;
        RECT 347.32 -3.56 347.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 347.315 -95.365 347.645 -95.035 ;
        RECT 347.315 -96.725 347.645 -96.395 ;
        RECT 347.315 -98.085 347.645 -97.755 ;
        RECT 347.315 -99.445 347.645 -99.115 ;
        RECT 347.315 -100.805 347.645 -100.475 ;
        RECT 347.315 -102.165 347.645 -101.835 ;
        RECT 347.315 -103.525 347.645 -103.195 ;
        RECT 347.315 -104.885 347.645 -104.555 ;
        RECT 347.315 -106.245 347.645 -105.915 ;
        RECT 347.315 -107.605 347.645 -107.275 ;
        RECT 347.315 -108.965 347.645 -108.635 ;
        RECT 347.315 -110.325 347.645 -109.995 ;
        RECT 347.315 -111.685 347.645 -111.355 ;
        RECT 347.315 -113.045 347.645 -112.715 ;
        RECT 347.315 -114.405 347.645 -114.075 ;
        RECT 347.315 -115.765 347.645 -115.435 ;
        RECT 347.315 -117.125 347.645 -116.795 ;
        RECT 347.315 -118.485 347.645 -118.155 ;
        RECT 347.315 -119.845 347.645 -119.515 ;
        RECT 347.315 -121.205 347.645 -120.875 ;
        RECT 347.315 -122.565 347.645 -122.235 ;
        RECT 347.315 -123.925 347.645 -123.595 ;
        RECT 347.315 -125.285 347.645 -124.955 ;
        RECT 347.315 -126.645 347.645 -126.315 ;
        RECT 347.315 -128.005 347.645 -127.675 ;
        RECT 347.315 -129.365 347.645 -129.035 ;
        RECT 347.315 -130.725 347.645 -130.395 ;
        RECT 347.315 -132.085 347.645 -131.755 ;
        RECT 347.315 -133.445 347.645 -133.115 ;
        RECT 347.315 -134.805 347.645 -134.475 ;
        RECT 347.315 -136.165 347.645 -135.835 ;
        RECT 347.315 -137.525 347.645 -137.195 ;
        RECT 347.315 -138.885 347.645 -138.555 ;
        RECT 347.315 -140.245 347.645 -139.915 ;
        RECT 347.315 -141.605 347.645 -141.275 ;
        RECT 347.315 -142.965 347.645 -142.635 ;
        RECT 347.315 -144.325 347.645 -143.995 ;
        RECT 347.315 -145.685 347.645 -145.355 ;
        RECT 347.315 -147.045 347.645 -146.715 ;
        RECT 347.315 -148.405 347.645 -148.075 ;
        RECT 347.315 -149.765 347.645 -149.435 ;
        RECT 347.315 -151.125 347.645 -150.795 ;
        RECT 347.315 -152.485 347.645 -152.155 ;
        RECT 347.315 -153.845 347.645 -153.515 ;
        RECT 347.315 -155.205 347.645 -154.875 ;
        RECT 347.315 -156.565 347.645 -156.235 ;
        RECT 347.315 -157.925 347.645 -157.595 ;
        RECT 347.315 -159.285 347.645 -158.955 ;
        RECT 347.315 -160.645 347.645 -160.315 ;
        RECT 347.315 -162.005 347.645 -161.675 ;
        RECT 347.315 -163.365 347.645 -163.035 ;
        RECT 347.315 -164.725 347.645 -164.395 ;
        RECT 347.315 -166.085 347.645 -165.755 ;
        RECT 347.315 -167.445 347.645 -167.115 ;
        RECT 347.315 -168.805 347.645 -168.475 ;
        RECT 347.315 -170.165 347.645 -169.835 ;
        RECT 347.315 -171.525 347.645 -171.195 ;
        RECT 347.315 -172.885 347.645 -172.555 ;
        RECT 347.315 -174.245 347.645 -173.915 ;
        RECT 347.315 -175.605 347.645 -175.275 ;
        RECT 347.315 -176.965 347.645 -176.635 ;
        RECT 347.315 -178.325 347.645 -177.995 ;
        RECT 347.315 -179.685 347.645 -179.355 ;
        RECT 347.315 -181.93 347.645 -180.8 ;
        RECT 347.32 -182.045 347.64 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.675 241.32 349.005 242.45 ;
        RECT 348.675 239.195 349.005 239.525 ;
        RECT 348.675 237.835 349.005 238.165 ;
        RECT 348.68 237.16 349 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.675 -1.525 349.005 -1.195 ;
        RECT 348.675 -2.885 349.005 -2.555 ;
        RECT 348.68 -3.56 349 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 348.675 -95.365 349.005 -95.035 ;
        RECT 348.675 -96.725 349.005 -96.395 ;
        RECT 348.675 -98.085 349.005 -97.755 ;
        RECT 348.675 -99.445 349.005 -99.115 ;
        RECT 348.675 -100.805 349.005 -100.475 ;
        RECT 348.675 -102.165 349.005 -101.835 ;
        RECT 348.675 -103.525 349.005 -103.195 ;
        RECT 348.675 -104.885 349.005 -104.555 ;
        RECT 348.675 -106.245 349.005 -105.915 ;
        RECT 348.675 -107.605 349.005 -107.275 ;
        RECT 348.675 -108.965 349.005 -108.635 ;
        RECT 348.675 -110.325 349.005 -109.995 ;
        RECT 348.675 -111.685 349.005 -111.355 ;
        RECT 348.675 -113.045 349.005 -112.715 ;
        RECT 348.675 -114.405 349.005 -114.075 ;
        RECT 348.675 -115.765 349.005 -115.435 ;
        RECT 348.675 -117.125 349.005 -116.795 ;
        RECT 348.675 -118.485 349.005 -118.155 ;
        RECT 348.675 -119.845 349.005 -119.515 ;
        RECT 348.675 -121.205 349.005 -120.875 ;
        RECT 348.675 -122.565 349.005 -122.235 ;
        RECT 348.675 -123.925 349.005 -123.595 ;
        RECT 348.675 -125.285 349.005 -124.955 ;
        RECT 348.675 -126.645 349.005 -126.315 ;
        RECT 348.675 -128.005 349.005 -127.675 ;
        RECT 348.675 -129.365 349.005 -129.035 ;
        RECT 348.675 -130.725 349.005 -130.395 ;
        RECT 348.675 -132.085 349.005 -131.755 ;
        RECT 348.675 -133.445 349.005 -133.115 ;
        RECT 348.675 -134.805 349.005 -134.475 ;
        RECT 348.675 -136.165 349.005 -135.835 ;
        RECT 348.675 -137.525 349.005 -137.195 ;
        RECT 348.675 -138.885 349.005 -138.555 ;
        RECT 348.675 -140.245 349.005 -139.915 ;
        RECT 348.675 -141.605 349.005 -141.275 ;
        RECT 348.675 -142.965 349.005 -142.635 ;
        RECT 348.675 -144.325 349.005 -143.995 ;
        RECT 348.675 -145.685 349.005 -145.355 ;
        RECT 348.675 -147.045 349.005 -146.715 ;
        RECT 348.675 -148.405 349.005 -148.075 ;
        RECT 348.675 -149.765 349.005 -149.435 ;
        RECT 348.675 -151.125 349.005 -150.795 ;
        RECT 348.675 -152.485 349.005 -152.155 ;
        RECT 348.675 -153.845 349.005 -153.515 ;
        RECT 348.675 -155.205 349.005 -154.875 ;
        RECT 348.675 -156.565 349.005 -156.235 ;
        RECT 348.675 -157.925 349.005 -157.595 ;
        RECT 348.675 -159.285 349.005 -158.955 ;
        RECT 348.675 -160.645 349.005 -160.315 ;
        RECT 348.675 -162.005 349.005 -161.675 ;
        RECT 348.675 -163.365 349.005 -163.035 ;
        RECT 348.675 -164.725 349.005 -164.395 ;
        RECT 348.675 -166.085 349.005 -165.755 ;
        RECT 348.675 -167.445 349.005 -167.115 ;
        RECT 348.675 -168.805 349.005 -168.475 ;
        RECT 348.675 -170.165 349.005 -169.835 ;
        RECT 348.675 -171.525 349.005 -171.195 ;
        RECT 348.675 -172.885 349.005 -172.555 ;
        RECT 348.675 -174.245 349.005 -173.915 ;
        RECT 348.675 -175.605 349.005 -175.275 ;
        RECT 348.675 -176.965 349.005 -176.635 ;
        RECT 348.675 -178.325 349.005 -177.995 ;
        RECT 348.675 -179.685 349.005 -179.355 ;
        RECT 348.675 -181.93 349.005 -180.8 ;
        RECT 348.68 -182.045 349 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.035 241.32 350.365 242.45 ;
        RECT 350.035 239.195 350.365 239.525 ;
        RECT 350.035 237.835 350.365 238.165 ;
        RECT 350.04 237.16 350.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.035 -1.525 350.365 -1.195 ;
        RECT 350.035 -2.885 350.365 -2.555 ;
        RECT 350.04 -3.56 350.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 350.035 -95.365 350.365 -95.035 ;
        RECT 350.035 -96.725 350.365 -96.395 ;
        RECT 350.035 -98.085 350.365 -97.755 ;
        RECT 350.035 -99.445 350.365 -99.115 ;
        RECT 350.035 -100.805 350.365 -100.475 ;
        RECT 350.035 -102.165 350.365 -101.835 ;
        RECT 350.035 -103.525 350.365 -103.195 ;
        RECT 350.035 -104.885 350.365 -104.555 ;
        RECT 350.035 -106.245 350.365 -105.915 ;
        RECT 350.035 -107.605 350.365 -107.275 ;
        RECT 350.035 -108.965 350.365 -108.635 ;
        RECT 350.035 -110.325 350.365 -109.995 ;
        RECT 350.035 -111.685 350.365 -111.355 ;
        RECT 350.035 -113.045 350.365 -112.715 ;
        RECT 350.035 -114.405 350.365 -114.075 ;
        RECT 350.035 -115.765 350.365 -115.435 ;
        RECT 350.035 -117.125 350.365 -116.795 ;
        RECT 350.035 -118.485 350.365 -118.155 ;
        RECT 350.035 -119.845 350.365 -119.515 ;
        RECT 350.035 -121.205 350.365 -120.875 ;
        RECT 350.035 -122.565 350.365 -122.235 ;
        RECT 350.035 -123.925 350.365 -123.595 ;
        RECT 350.035 -125.285 350.365 -124.955 ;
        RECT 350.035 -126.645 350.365 -126.315 ;
        RECT 350.035 -128.005 350.365 -127.675 ;
        RECT 350.035 -129.365 350.365 -129.035 ;
        RECT 350.035 -130.725 350.365 -130.395 ;
        RECT 350.035 -132.085 350.365 -131.755 ;
        RECT 350.035 -133.445 350.365 -133.115 ;
        RECT 350.035 -134.805 350.365 -134.475 ;
        RECT 350.035 -136.165 350.365 -135.835 ;
        RECT 350.035 -137.525 350.365 -137.195 ;
        RECT 350.035 -138.885 350.365 -138.555 ;
        RECT 350.035 -140.245 350.365 -139.915 ;
        RECT 350.035 -141.605 350.365 -141.275 ;
        RECT 350.035 -142.965 350.365 -142.635 ;
        RECT 350.035 -144.325 350.365 -143.995 ;
        RECT 350.035 -145.685 350.365 -145.355 ;
        RECT 350.035 -147.045 350.365 -146.715 ;
        RECT 350.035 -148.405 350.365 -148.075 ;
        RECT 350.035 -149.765 350.365 -149.435 ;
        RECT 350.035 -151.125 350.365 -150.795 ;
        RECT 350.035 -152.485 350.365 -152.155 ;
        RECT 350.035 -153.845 350.365 -153.515 ;
        RECT 350.035 -155.205 350.365 -154.875 ;
        RECT 350.035 -156.565 350.365 -156.235 ;
        RECT 350.035 -157.925 350.365 -157.595 ;
        RECT 350.035 -159.285 350.365 -158.955 ;
        RECT 350.035 -160.645 350.365 -160.315 ;
        RECT 350.035 -162.005 350.365 -161.675 ;
        RECT 350.035 -163.365 350.365 -163.035 ;
        RECT 350.035 -164.725 350.365 -164.395 ;
        RECT 350.035 -166.085 350.365 -165.755 ;
        RECT 350.035 -167.445 350.365 -167.115 ;
        RECT 350.035 -168.805 350.365 -168.475 ;
        RECT 350.035 -170.165 350.365 -169.835 ;
        RECT 350.035 -171.525 350.365 -171.195 ;
        RECT 350.035 -172.885 350.365 -172.555 ;
        RECT 350.035 -174.245 350.365 -173.915 ;
        RECT 350.035 -175.605 350.365 -175.275 ;
        RECT 350.035 -176.965 350.365 -176.635 ;
        RECT 350.035 -178.325 350.365 -177.995 ;
        RECT 350.035 -179.685 350.365 -179.355 ;
        RECT 350.035 -181.93 350.365 -180.8 ;
        RECT 350.04 -182.045 350.36 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.395 241.32 351.725 242.45 ;
        RECT 351.395 239.195 351.725 239.525 ;
        RECT 351.395 237.835 351.725 238.165 ;
        RECT 351.4 237.16 351.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.395 -99.445 351.725 -99.115 ;
        RECT 351.395 -100.805 351.725 -100.475 ;
        RECT 351.395 -102.165 351.725 -101.835 ;
        RECT 351.395 -103.525 351.725 -103.195 ;
        RECT 351.395 -104.885 351.725 -104.555 ;
        RECT 351.395 -106.245 351.725 -105.915 ;
        RECT 351.395 -107.605 351.725 -107.275 ;
        RECT 351.395 -108.965 351.725 -108.635 ;
        RECT 351.395 -110.325 351.725 -109.995 ;
        RECT 351.395 -111.685 351.725 -111.355 ;
        RECT 351.395 -113.045 351.725 -112.715 ;
        RECT 351.395 -114.405 351.725 -114.075 ;
        RECT 351.395 -115.765 351.725 -115.435 ;
        RECT 351.395 -117.125 351.725 -116.795 ;
        RECT 351.395 -118.485 351.725 -118.155 ;
        RECT 351.395 -119.845 351.725 -119.515 ;
        RECT 351.395 -121.205 351.725 -120.875 ;
        RECT 351.395 -122.565 351.725 -122.235 ;
        RECT 351.395 -123.925 351.725 -123.595 ;
        RECT 351.395 -125.285 351.725 -124.955 ;
        RECT 351.395 -126.645 351.725 -126.315 ;
        RECT 351.395 -128.005 351.725 -127.675 ;
        RECT 351.395 -129.365 351.725 -129.035 ;
        RECT 351.395 -130.725 351.725 -130.395 ;
        RECT 351.395 -132.085 351.725 -131.755 ;
        RECT 351.395 -133.445 351.725 -133.115 ;
        RECT 351.395 -134.805 351.725 -134.475 ;
        RECT 351.395 -136.165 351.725 -135.835 ;
        RECT 351.395 -137.525 351.725 -137.195 ;
        RECT 351.395 -138.885 351.725 -138.555 ;
        RECT 351.395 -140.245 351.725 -139.915 ;
        RECT 351.395 -141.605 351.725 -141.275 ;
        RECT 351.395 -142.965 351.725 -142.635 ;
        RECT 351.395 -144.325 351.725 -143.995 ;
        RECT 351.395 -145.685 351.725 -145.355 ;
        RECT 351.395 -147.045 351.725 -146.715 ;
        RECT 351.395 -148.405 351.725 -148.075 ;
        RECT 351.395 -149.765 351.725 -149.435 ;
        RECT 351.395 -151.125 351.725 -150.795 ;
        RECT 351.395 -152.485 351.725 -152.155 ;
        RECT 351.395 -153.845 351.725 -153.515 ;
        RECT 351.395 -155.205 351.725 -154.875 ;
        RECT 351.395 -156.565 351.725 -156.235 ;
        RECT 351.395 -157.925 351.725 -157.595 ;
        RECT 351.395 -159.285 351.725 -158.955 ;
        RECT 351.395 -160.645 351.725 -160.315 ;
        RECT 351.395 -162.005 351.725 -161.675 ;
        RECT 351.395 -163.365 351.725 -163.035 ;
        RECT 351.395 -164.725 351.725 -164.395 ;
        RECT 351.395 -166.085 351.725 -165.755 ;
        RECT 351.395 -167.445 351.725 -167.115 ;
        RECT 351.395 -168.805 351.725 -168.475 ;
        RECT 351.395 -170.165 351.725 -169.835 ;
        RECT 351.395 -171.525 351.725 -171.195 ;
        RECT 351.395 -172.885 351.725 -172.555 ;
        RECT 351.395 -174.245 351.725 -173.915 ;
        RECT 351.395 -175.605 351.725 -175.275 ;
        RECT 351.395 -176.965 351.725 -176.635 ;
        RECT 351.395 -178.325 351.725 -177.995 ;
        RECT 351.395 -179.685 351.725 -179.355 ;
        RECT 351.395 -181.93 351.725 -180.8 ;
        RECT 351.4 -182.045 351.72 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 351.46 -98.075 351.79 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.755 241.32 353.085 242.45 ;
        RECT 352.755 239.195 353.085 239.525 ;
        RECT 352.755 237.835 353.085 238.165 ;
        RECT 352.76 237.16 353.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 352.755 -99.445 353.085 -99.115 ;
        RECT 352.755 -100.805 353.085 -100.475 ;
        RECT 352.755 -102.165 353.085 -101.835 ;
        RECT 352.755 -103.525 353.085 -103.195 ;
        RECT 352.755 -104.885 353.085 -104.555 ;
        RECT 352.755 -106.245 353.085 -105.915 ;
        RECT 352.755 -107.605 353.085 -107.275 ;
        RECT 352.755 -108.965 353.085 -108.635 ;
        RECT 352.755 -110.325 353.085 -109.995 ;
        RECT 352.755 -111.685 353.085 -111.355 ;
        RECT 352.755 -113.045 353.085 -112.715 ;
        RECT 352.755 -114.405 353.085 -114.075 ;
        RECT 352.755 -115.765 353.085 -115.435 ;
        RECT 352.755 -117.125 353.085 -116.795 ;
        RECT 352.755 -118.485 353.085 -118.155 ;
        RECT 352.755 -119.845 353.085 -119.515 ;
        RECT 352.755 -121.205 353.085 -120.875 ;
        RECT 352.755 -122.565 353.085 -122.235 ;
        RECT 352.755 -123.925 353.085 -123.595 ;
        RECT 352.755 -125.285 353.085 -124.955 ;
        RECT 352.755 -126.645 353.085 -126.315 ;
        RECT 352.755 -128.005 353.085 -127.675 ;
        RECT 352.755 -129.365 353.085 -129.035 ;
        RECT 352.755 -130.725 353.085 -130.395 ;
        RECT 352.755 -132.085 353.085 -131.755 ;
        RECT 352.755 -133.445 353.085 -133.115 ;
        RECT 352.755 -134.805 353.085 -134.475 ;
        RECT 352.755 -136.165 353.085 -135.835 ;
        RECT 352.755 -137.525 353.085 -137.195 ;
        RECT 352.755 -138.885 353.085 -138.555 ;
        RECT 352.755 -140.245 353.085 -139.915 ;
        RECT 352.755 -141.605 353.085 -141.275 ;
        RECT 352.755 -142.965 353.085 -142.635 ;
        RECT 352.755 -144.325 353.085 -143.995 ;
        RECT 352.755 -145.685 353.085 -145.355 ;
        RECT 352.755 -147.045 353.085 -146.715 ;
        RECT 352.755 -148.405 353.085 -148.075 ;
        RECT 352.755 -149.765 353.085 -149.435 ;
        RECT 352.755 -151.125 353.085 -150.795 ;
        RECT 352.755 -152.485 353.085 -152.155 ;
        RECT 352.755 -153.845 353.085 -153.515 ;
        RECT 352.755 -155.205 353.085 -154.875 ;
        RECT 352.755 -156.565 353.085 -156.235 ;
        RECT 352.755 -157.925 353.085 -157.595 ;
        RECT 352.755 -159.285 353.085 -158.955 ;
        RECT 352.755 -160.645 353.085 -160.315 ;
        RECT 352.755 -162.005 353.085 -161.675 ;
        RECT 352.755 -163.365 353.085 -163.035 ;
        RECT 352.755 -164.725 353.085 -164.395 ;
        RECT 352.755 -166.085 353.085 -165.755 ;
        RECT 352.755 -167.445 353.085 -167.115 ;
        RECT 352.755 -168.805 353.085 -168.475 ;
        RECT 352.755 -170.165 353.085 -169.835 ;
        RECT 352.755 -171.525 353.085 -171.195 ;
        RECT 352.755 -172.885 353.085 -172.555 ;
        RECT 352.755 -174.245 353.085 -173.915 ;
        RECT 352.755 -175.605 353.085 -175.275 ;
        RECT 352.755 -176.965 353.085 -176.635 ;
        RECT 352.755 -178.325 353.085 -177.995 ;
        RECT 352.755 -179.685 353.085 -179.355 ;
        RECT 352.755 -181.93 353.085 -180.8 ;
        RECT 352.76 -182.045 353.08 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.115 241.32 354.445 242.45 ;
        RECT 354.115 239.195 354.445 239.525 ;
        RECT 354.115 237.835 354.445 238.165 ;
        RECT 354.12 237.16 354.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.115 -1.525 354.445 -1.195 ;
        RECT 354.115 -2.885 354.445 -2.555 ;
        RECT 354.12 -3.56 354.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 354.115 -95.365 354.445 -95.035 ;
        RECT 354.115 -96.725 354.445 -96.395 ;
        RECT 354.115 -98.085 354.445 -97.755 ;
        RECT 354.115 -99.445 354.445 -99.115 ;
        RECT 354.115 -100.805 354.445 -100.475 ;
        RECT 354.115 -102.165 354.445 -101.835 ;
        RECT 354.115 -103.525 354.445 -103.195 ;
        RECT 354.115 -104.885 354.445 -104.555 ;
        RECT 354.115 -106.245 354.445 -105.915 ;
        RECT 354.115 -107.605 354.445 -107.275 ;
        RECT 354.115 -108.965 354.445 -108.635 ;
        RECT 354.115 -110.325 354.445 -109.995 ;
        RECT 354.115 -111.685 354.445 -111.355 ;
        RECT 354.115 -113.045 354.445 -112.715 ;
        RECT 354.115 -114.405 354.445 -114.075 ;
        RECT 354.115 -115.765 354.445 -115.435 ;
        RECT 354.115 -117.125 354.445 -116.795 ;
        RECT 354.115 -118.485 354.445 -118.155 ;
        RECT 354.115 -119.845 354.445 -119.515 ;
        RECT 354.115 -121.205 354.445 -120.875 ;
        RECT 354.115 -122.565 354.445 -122.235 ;
        RECT 354.115 -123.925 354.445 -123.595 ;
        RECT 354.115 -125.285 354.445 -124.955 ;
        RECT 354.115 -126.645 354.445 -126.315 ;
        RECT 354.115 -128.005 354.445 -127.675 ;
        RECT 354.115 -129.365 354.445 -129.035 ;
        RECT 354.115 -130.725 354.445 -130.395 ;
        RECT 354.115 -132.085 354.445 -131.755 ;
        RECT 354.115 -133.445 354.445 -133.115 ;
        RECT 354.115 -134.805 354.445 -134.475 ;
        RECT 354.115 -136.165 354.445 -135.835 ;
        RECT 354.115 -137.525 354.445 -137.195 ;
        RECT 354.115 -138.885 354.445 -138.555 ;
        RECT 354.115 -140.245 354.445 -139.915 ;
        RECT 354.115 -141.605 354.445 -141.275 ;
        RECT 354.115 -142.965 354.445 -142.635 ;
        RECT 354.115 -144.325 354.445 -143.995 ;
        RECT 354.115 -145.685 354.445 -145.355 ;
        RECT 354.115 -147.045 354.445 -146.715 ;
        RECT 354.115 -148.405 354.445 -148.075 ;
        RECT 354.115 -149.765 354.445 -149.435 ;
        RECT 354.115 -151.125 354.445 -150.795 ;
        RECT 354.115 -152.485 354.445 -152.155 ;
        RECT 354.115 -153.845 354.445 -153.515 ;
        RECT 354.115 -155.205 354.445 -154.875 ;
        RECT 354.115 -156.565 354.445 -156.235 ;
        RECT 354.115 -157.925 354.445 -157.595 ;
        RECT 354.115 -159.285 354.445 -158.955 ;
        RECT 354.115 -160.645 354.445 -160.315 ;
        RECT 354.115 -162.005 354.445 -161.675 ;
        RECT 354.115 -163.365 354.445 -163.035 ;
        RECT 354.115 -164.725 354.445 -164.395 ;
        RECT 354.115 -166.085 354.445 -165.755 ;
        RECT 354.115 -167.445 354.445 -167.115 ;
        RECT 354.115 -168.805 354.445 -168.475 ;
        RECT 354.115 -170.165 354.445 -169.835 ;
        RECT 354.115 -171.525 354.445 -171.195 ;
        RECT 354.115 -172.885 354.445 -172.555 ;
        RECT 354.115 -174.245 354.445 -173.915 ;
        RECT 354.115 -175.605 354.445 -175.275 ;
        RECT 354.115 -176.965 354.445 -176.635 ;
        RECT 354.115 -178.325 354.445 -177.995 ;
        RECT 354.115 -179.685 354.445 -179.355 ;
        RECT 354.115 -181.93 354.445 -180.8 ;
        RECT 354.12 -182.045 354.44 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 355.475 231.995 355.805 232.325 ;
        RECT 355.475 230.155 355.805 230.485 ;
        RECT 355.475 228.665 355.805 228.995 ;
        RECT 355.475 226.995 355.805 227.325 ;
        RECT 355.475 225.505 355.805 225.835 ;
        RECT 355.475 223.835 355.805 224.165 ;
        RECT 355.475 222.345 355.805 222.675 ;
        RECT 355.475 220.675 355.805 221.005 ;
        RECT 355.475 219.185 355.805 219.515 ;
        RECT 355.475 217.775 355.805 218.105 ;
        RECT 355.475 215.935 355.805 216.265 ;
        RECT 355.475 214.445 355.805 214.775 ;
        RECT 355.475 212.775 355.805 213.105 ;
        RECT 355.475 211.285 355.805 211.615 ;
        RECT 355.475 209.615 355.805 209.945 ;
        RECT 355.475 208.125 355.805 208.455 ;
        RECT 355.475 206.455 355.805 206.785 ;
        RECT 355.475 204.965 355.805 205.295 ;
        RECT 355.475 203.555 355.805 203.885 ;
        RECT 355.475 201.715 355.805 202.045 ;
        RECT 355.475 200.225 355.805 200.555 ;
        RECT 355.475 198.555 355.805 198.885 ;
        RECT 355.475 197.065 355.805 197.395 ;
        RECT 355.475 195.395 355.805 195.725 ;
        RECT 355.475 193.905 355.805 194.235 ;
        RECT 355.475 192.235 355.805 192.565 ;
        RECT 355.475 190.745 355.805 191.075 ;
        RECT 355.475 189.335 355.805 189.665 ;
        RECT 355.475 187.495 355.805 187.825 ;
        RECT 355.475 186.005 355.805 186.335 ;
        RECT 355.475 184.335 355.805 184.665 ;
        RECT 355.475 182.845 355.805 183.175 ;
        RECT 355.475 181.175 355.805 181.505 ;
        RECT 355.475 179.685 355.805 180.015 ;
        RECT 355.475 178.015 355.805 178.345 ;
        RECT 355.475 176.525 355.805 176.855 ;
        RECT 355.475 175.115 355.805 175.445 ;
        RECT 355.475 173.275 355.805 173.605 ;
        RECT 355.475 171.785 355.805 172.115 ;
        RECT 355.475 170.115 355.805 170.445 ;
        RECT 355.475 168.625 355.805 168.955 ;
        RECT 355.475 166.955 355.805 167.285 ;
        RECT 355.475 165.465 355.805 165.795 ;
        RECT 355.475 163.795 355.805 164.125 ;
        RECT 355.475 162.305 355.805 162.635 ;
        RECT 355.475 160.895 355.805 161.225 ;
        RECT 355.475 159.055 355.805 159.385 ;
        RECT 355.475 157.565 355.805 157.895 ;
        RECT 355.475 155.895 355.805 156.225 ;
        RECT 355.475 154.405 355.805 154.735 ;
        RECT 355.475 152.735 355.805 153.065 ;
        RECT 355.475 151.245 355.805 151.575 ;
        RECT 355.475 149.575 355.805 149.905 ;
        RECT 355.475 148.085 355.805 148.415 ;
        RECT 355.475 146.675 355.805 147.005 ;
        RECT 355.475 144.835 355.805 145.165 ;
        RECT 355.475 143.345 355.805 143.675 ;
        RECT 355.475 141.675 355.805 142.005 ;
        RECT 355.475 140.185 355.805 140.515 ;
        RECT 355.475 138.515 355.805 138.845 ;
        RECT 355.475 137.025 355.805 137.355 ;
        RECT 355.475 135.355 355.805 135.685 ;
        RECT 355.475 133.865 355.805 134.195 ;
        RECT 355.475 132.455 355.805 132.785 ;
        RECT 355.475 130.615 355.805 130.945 ;
        RECT 355.475 129.125 355.805 129.455 ;
        RECT 355.475 127.455 355.805 127.785 ;
        RECT 355.475 125.965 355.805 126.295 ;
        RECT 355.475 124.295 355.805 124.625 ;
        RECT 355.475 122.805 355.805 123.135 ;
        RECT 355.475 121.135 355.805 121.465 ;
        RECT 355.475 119.645 355.805 119.975 ;
        RECT 355.475 118.235 355.805 118.565 ;
        RECT 355.475 116.395 355.805 116.725 ;
        RECT 355.475 114.905 355.805 115.235 ;
        RECT 355.475 113.235 355.805 113.565 ;
        RECT 355.475 111.745 355.805 112.075 ;
        RECT 355.475 110.075 355.805 110.405 ;
        RECT 355.475 108.585 355.805 108.915 ;
        RECT 355.475 106.915 355.805 107.245 ;
        RECT 355.475 105.425 355.805 105.755 ;
        RECT 355.475 104.015 355.805 104.345 ;
        RECT 355.475 102.175 355.805 102.505 ;
        RECT 355.475 100.685 355.805 101.015 ;
        RECT 355.475 99.015 355.805 99.345 ;
        RECT 355.475 97.525 355.805 97.855 ;
        RECT 355.475 95.855 355.805 96.185 ;
        RECT 355.475 94.365 355.805 94.695 ;
        RECT 355.475 92.695 355.805 93.025 ;
        RECT 355.475 91.205 355.805 91.535 ;
        RECT 355.475 89.795 355.805 90.125 ;
        RECT 355.475 87.955 355.805 88.285 ;
        RECT 355.475 86.465 355.805 86.795 ;
        RECT 355.475 84.795 355.805 85.125 ;
        RECT 355.475 83.305 355.805 83.635 ;
        RECT 355.475 81.635 355.805 81.965 ;
        RECT 355.475 80.145 355.805 80.475 ;
        RECT 355.475 78.475 355.805 78.805 ;
        RECT 355.475 76.985 355.805 77.315 ;
        RECT 355.475 75.575 355.805 75.905 ;
        RECT 355.475 73.735 355.805 74.065 ;
        RECT 355.475 72.245 355.805 72.575 ;
        RECT 355.475 70.575 355.805 70.905 ;
        RECT 355.475 69.085 355.805 69.415 ;
        RECT 355.475 67.415 355.805 67.745 ;
        RECT 355.475 65.925 355.805 66.255 ;
        RECT 355.475 64.255 355.805 64.585 ;
        RECT 355.475 62.765 355.805 63.095 ;
        RECT 355.475 61.355 355.805 61.685 ;
        RECT 355.475 59.515 355.805 59.845 ;
        RECT 355.475 58.025 355.805 58.355 ;
        RECT 355.475 56.355 355.805 56.685 ;
        RECT 355.475 54.865 355.805 55.195 ;
        RECT 355.475 53.195 355.805 53.525 ;
        RECT 355.475 51.705 355.805 52.035 ;
        RECT 355.475 50.035 355.805 50.365 ;
        RECT 355.475 48.545 355.805 48.875 ;
        RECT 355.475 47.135 355.805 47.465 ;
        RECT 355.475 45.295 355.805 45.625 ;
        RECT 355.475 43.805 355.805 44.135 ;
        RECT 355.475 42.135 355.805 42.465 ;
        RECT 355.475 40.645 355.805 40.975 ;
        RECT 355.475 38.975 355.805 39.305 ;
        RECT 355.475 37.485 355.805 37.815 ;
        RECT 355.475 35.815 355.805 36.145 ;
        RECT 355.475 34.325 355.805 34.655 ;
        RECT 355.475 32.915 355.805 33.245 ;
        RECT 355.475 31.075 355.805 31.405 ;
        RECT 355.475 29.585 355.805 29.915 ;
        RECT 355.475 27.915 355.805 28.245 ;
        RECT 355.475 26.425 355.805 26.755 ;
        RECT 355.475 24.755 355.805 25.085 ;
        RECT 355.475 23.265 355.805 23.595 ;
        RECT 355.475 21.595 355.805 21.925 ;
        RECT 355.475 20.105 355.805 20.435 ;
        RECT 355.475 18.695 355.805 19.025 ;
        RECT 355.475 16.855 355.805 17.185 ;
        RECT 355.475 15.365 355.805 15.695 ;
        RECT 355.475 13.695 355.805 14.025 ;
        RECT 355.475 12.205 355.805 12.535 ;
        RECT 355.475 10.535 355.805 10.865 ;
        RECT 355.475 9.045 355.805 9.375 ;
        RECT 355.475 7.375 355.805 7.705 ;
        RECT 355.475 5.885 355.805 6.215 ;
        RECT 355.475 4.475 355.805 4.805 ;
        RECT 355.475 2.115 355.805 2.445 ;
        RECT 355.475 0.06 355.805 0.39 ;
        RECT 355.475 -1.525 355.805 -1.195 ;
        RECT 355.475 -2.885 355.805 -2.555 ;
        RECT 355.475 -4.245 355.805 -3.915 ;
        RECT 355.475 -5.605 355.805 -5.275 ;
        RECT 355.475 -6.965 355.805 -6.635 ;
        RECT 355.475 -8.325 355.805 -7.995 ;
        RECT 355.475 -9.685 355.805 -9.355 ;
        RECT 355.475 -11.045 355.805 -10.715 ;
        RECT 355.475 -12.405 355.805 -12.075 ;
        RECT 355.475 -13.765 355.805 -13.435 ;
        RECT 355.475 -15.125 355.805 -14.795 ;
        RECT 355.475 -16.485 355.805 -16.155 ;
        RECT 355.475 -17.845 355.805 -17.515 ;
        RECT 355.475 -19.205 355.805 -18.875 ;
        RECT 355.475 -20.565 355.805 -20.235 ;
        RECT 355.475 -21.925 355.805 -21.595 ;
        RECT 355.475 -23.285 355.805 -22.955 ;
        RECT 355.475 -24.645 355.805 -24.315 ;
        RECT 355.475 -26.005 355.805 -25.675 ;
        RECT 355.475 -27.365 355.805 -27.035 ;
        RECT 355.475 -28.725 355.805 -28.395 ;
        RECT 355.475 -30.085 355.805 -29.755 ;
        RECT 355.475 -31.445 355.805 -31.115 ;
        RECT 355.475 -32.805 355.805 -32.475 ;
        RECT 355.475 -34.165 355.805 -33.835 ;
        RECT 355.475 -35.525 355.805 -35.195 ;
        RECT 355.475 -36.885 355.805 -36.555 ;
        RECT 355.475 -38.245 355.805 -37.915 ;
        RECT 355.475 -39.605 355.805 -39.275 ;
        RECT 355.475 -40.965 355.805 -40.635 ;
        RECT 355.475 -42.325 355.805 -41.995 ;
        RECT 355.475 -43.685 355.805 -43.355 ;
        RECT 355.475 -45.045 355.805 -44.715 ;
        RECT 355.475 -46.405 355.805 -46.075 ;
        RECT 355.475 -47.765 355.805 -47.435 ;
        RECT 355.475 -49.125 355.805 -48.795 ;
        RECT 355.475 -50.485 355.805 -50.155 ;
        RECT 355.475 -51.845 355.805 -51.515 ;
        RECT 355.475 -53.205 355.805 -52.875 ;
        RECT 355.475 -54.565 355.805 -54.235 ;
        RECT 355.475 -55.925 355.805 -55.595 ;
        RECT 355.475 -57.285 355.805 -56.955 ;
        RECT 355.475 -58.645 355.805 -58.315 ;
        RECT 355.475 -60.005 355.805 -59.675 ;
        RECT 355.475 -61.365 355.805 -61.035 ;
        RECT 355.475 -62.725 355.805 -62.395 ;
        RECT 355.475 -64.085 355.805 -63.755 ;
        RECT 355.475 -65.445 355.805 -65.115 ;
        RECT 355.475 -66.805 355.805 -66.475 ;
        RECT 355.475 -68.165 355.805 -67.835 ;
        RECT 355.475 -69.525 355.805 -69.195 ;
        RECT 355.475 -70.885 355.805 -70.555 ;
        RECT 355.475 -72.245 355.805 -71.915 ;
        RECT 355.475 -73.605 355.805 -73.275 ;
        RECT 355.475 -74.965 355.805 -74.635 ;
        RECT 355.475 -76.325 355.805 -75.995 ;
        RECT 355.475 -77.685 355.805 -77.355 ;
        RECT 355.475 -79.045 355.805 -78.715 ;
        RECT 355.475 -80.405 355.805 -80.075 ;
        RECT 355.475 -81.765 355.805 -81.435 ;
        RECT 355.475 -83.125 355.805 -82.795 ;
        RECT 355.475 -84.485 355.805 -84.155 ;
        RECT 355.475 -85.845 355.805 -85.515 ;
        RECT 355.475 -87.205 355.805 -86.875 ;
        RECT 355.475 -88.565 355.805 -88.235 ;
        RECT 355.475 -89.925 355.805 -89.595 ;
        RECT 355.475 -91.285 355.805 -90.955 ;
        RECT 355.475 -92.645 355.805 -92.315 ;
        RECT 355.475 -94.005 355.805 -93.675 ;
        RECT 355.475 -95.365 355.805 -95.035 ;
        RECT 355.475 -96.725 355.805 -96.395 ;
        RECT 355.475 -98.085 355.805 -97.755 ;
        RECT 355.475 -99.445 355.805 -99.115 ;
        RECT 355.475 -100.805 355.805 -100.475 ;
        RECT 355.475 -102.165 355.805 -101.835 ;
        RECT 355.475 -103.525 355.805 -103.195 ;
        RECT 355.475 -104.885 355.805 -104.555 ;
        RECT 355.475 -106.245 355.805 -105.915 ;
        RECT 355.475 -107.605 355.805 -107.275 ;
        RECT 355.475 -108.965 355.805 -108.635 ;
        RECT 355.475 -110.325 355.805 -109.995 ;
        RECT 355.475 -111.685 355.805 -111.355 ;
        RECT 355.475 -113.045 355.805 -112.715 ;
        RECT 355.475 -114.405 355.805 -114.075 ;
        RECT 355.475 -115.765 355.805 -115.435 ;
        RECT 355.475 -117.125 355.805 -116.795 ;
        RECT 355.475 -118.485 355.805 -118.155 ;
        RECT 355.475 -119.845 355.805 -119.515 ;
        RECT 355.475 -121.205 355.805 -120.875 ;
        RECT 355.475 -122.565 355.805 -122.235 ;
        RECT 355.475 -123.925 355.805 -123.595 ;
        RECT 355.475 -125.285 355.805 -124.955 ;
        RECT 355.475 -126.645 355.805 -126.315 ;
        RECT 355.475 -128.005 355.805 -127.675 ;
        RECT 355.475 -129.365 355.805 -129.035 ;
        RECT 355.475 -130.725 355.805 -130.395 ;
        RECT 355.475 -132.085 355.805 -131.755 ;
        RECT 355.475 -133.445 355.805 -133.115 ;
        RECT 355.475 -134.805 355.805 -134.475 ;
        RECT 355.475 -136.165 355.805 -135.835 ;
        RECT 355.475 -137.525 355.805 -137.195 ;
        RECT 355.475 -138.885 355.805 -138.555 ;
        RECT 355.475 -140.245 355.805 -139.915 ;
        RECT 355.475 -141.605 355.805 -141.275 ;
        RECT 355.475 -142.965 355.805 -142.635 ;
        RECT 355.475 -144.325 355.805 -143.995 ;
        RECT 355.475 -145.685 355.805 -145.355 ;
        RECT 355.475 -147.045 355.805 -146.715 ;
        RECT 355.475 -148.405 355.805 -148.075 ;
        RECT 355.475 -149.765 355.805 -149.435 ;
        RECT 355.475 -151.125 355.805 -150.795 ;
        RECT 355.475 -152.485 355.805 -152.155 ;
        RECT 355.475 -153.845 355.805 -153.515 ;
        RECT 355.475 -155.205 355.805 -154.875 ;
        RECT 355.475 -156.565 355.805 -156.235 ;
        RECT 355.475 -157.925 355.805 -157.595 ;
        RECT 355.475 -159.285 355.805 -158.955 ;
        RECT 355.475 -160.645 355.805 -160.315 ;
        RECT 355.475 -162.005 355.805 -161.675 ;
        RECT 355.475 -163.365 355.805 -163.035 ;
        RECT 355.475 -164.725 355.805 -164.395 ;
        RECT 355.475 -166.085 355.805 -165.755 ;
        RECT 355.475 -167.445 355.805 -167.115 ;
        RECT 355.475 -168.805 355.805 -168.475 ;
        RECT 355.475 -170.165 355.805 -169.835 ;
        RECT 355.475 -171.525 355.805 -171.195 ;
        RECT 355.475 -172.885 355.805 -172.555 ;
        RECT 355.475 -174.245 355.805 -173.915 ;
        RECT 355.475 -175.605 355.805 -175.275 ;
        RECT 355.475 -176.965 355.805 -176.635 ;
        RECT 355.475 -178.325 355.805 -177.995 ;
        RECT 355.475 -179.685 355.805 -179.355 ;
        RECT 355.475 -181.93 355.805 -180.8 ;
        RECT 355.48 -182.045 355.8 242.565 ;
        RECT 355.475 241.32 355.805 242.45 ;
        RECT 355.475 239.195 355.805 239.525 ;
        RECT 355.475 237.835 355.805 238.165 ;
        RECT 355.475 235.975 355.805 236.305 ;
        RECT 355.475 233.925 355.805 234.255 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.035 241.32 316.365 242.45 ;
        RECT 316.035 239.195 316.365 239.525 ;
        RECT 316.035 237.835 316.365 238.165 ;
        RECT 316.04 237.16 316.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.035 -1.525 316.365 -1.195 ;
        RECT 316.035 -2.885 316.365 -2.555 ;
        RECT 316.04 -3.56 316.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 316.035 -95.365 316.365 -95.035 ;
        RECT 316.035 -96.725 316.365 -96.395 ;
        RECT 316.035 -98.085 316.365 -97.755 ;
        RECT 316.035 -99.445 316.365 -99.115 ;
        RECT 316.035 -100.805 316.365 -100.475 ;
        RECT 316.035 -102.165 316.365 -101.835 ;
        RECT 316.035 -103.525 316.365 -103.195 ;
        RECT 316.035 -104.885 316.365 -104.555 ;
        RECT 316.035 -106.245 316.365 -105.915 ;
        RECT 316.035 -107.605 316.365 -107.275 ;
        RECT 316.035 -108.965 316.365 -108.635 ;
        RECT 316.035 -110.325 316.365 -109.995 ;
        RECT 316.035 -111.685 316.365 -111.355 ;
        RECT 316.035 -113.045 316.365 -112.715 ;
        RECT 316.035 -114.405 316.365 -114.075 ;
        RECT 316.035 -115.765 316.365 -115.435 ;
        RECT 316.035 -117.125 316.365 -116.795 ;
        RECT 316.035 -118.485 316.365 -118.155 ;
        RECT 316.035 -119.845 316.365 -119.515 ;
        RECT 316.035 -121.205 316.365 -120.875 ;
        RECT 316.035 -122.565 316.365 -122.235 ;
        RECT 316.035 -123.925 316.365 -123.595 ;
        RECT 316.035 -125.285 316.365 -124.955 ;
        RECT 316.035 -126.645 316.365 -126.315 ;
        RECT 316.035 -128.005 316.365 -127.675 ;
        RECT 316.035 -129.365 316.365 -129.035 ;
        RECT 316.035 -130.725 316.365 -130.395 ;
        RECT 316.035 -132.085 316.365 -131.755 ;
        RECT 316.035 -133.445 316.365 -133.115 ;
        RECT 316.035 -134.805 316.365 -134.475 ;
        RECT 316.035 -136.165 316.365 -135.835 ;
        RECT 316.035 -137.525 316.365 -137.195 ;
        RECT 316.035 -138.885 316.365 -138.555 ;
        RECT 316.035 -140.245 316.365 -139.915 ;
        RECT 316.035 -141.605 316.365 -141.275 ;
        RECT 316.035 -142.965 316.365 -142.635 ;
        RECT 316.035 -144.325 316.365 -143.995 ;
        RECT 316.035 -145.685 316.365 -145.355 ;
        RECT 316.035 -147.045 316.365 -146.715 ;
        RECT 316.035 -148.405 316.365 -148.075 ;
        RECT 316.035 -149.765 316.365 -149.435 ;
        RECT 316.035 -151.125 316.365 -150.795 ;
        RECT 316.035 -152.485 316.365 -152.155 ;
        RECT 316.035 -153.845 316.365 -153.515 ;
        RECT 316.035 -155.205 316.365 -154.875 ;
        RECT 316.035 -156.565 316.365 -156.235 ;
        RECT 316.035 -157.925 316.365 -157.595 ;
        RECT 316.035 -159.285 316.365 -158.955 ;
        RECT 316.035 -160.645 316.365 -160.315 ;
        RECT 316.035 -162.005 316.365 -161.675 ;
        RECT 316.035 -163.365 316.365 -163.035 ;
        RECT 316.035 -164.725 316.365 -164.395 ;
        RECT 316.035 -166.085 316.365 -165.755 ;
        RECT 316.035 -167.445 316.365 -167.115 ;
        RECT 316.035 -168.805 316.365 -168.475 ;
        RECT 316.035 -170.165 316.365 -169.835 ;
        RECT 316.035 -171.525 316.365 -171.195 ;
        RECT 316.035 -172.885 316.365 -172.555 ;
        RECT 316.035 -174.245 316.365 -173.915 ;
        RECT 316.035 -175.605 316.365 -175.275 ;
        RECT 316.035 -176.965 316.365 -176.635 ;
        RECT 316.035 -178.325 316.365 -177.995 ;
        RECT 316.035 -179.685 316.365 -179.355 ;
        RECT 316.035 -181.93 316.365 -180.8 ;
        RECT 316.04 -182.045 316.36 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.395 241.32 317.725 242.45 ;
        RECT 317.395 239.195 317.725 239.525 ;
        RECT 317.395 237.835 317.725 238.165 ;
        RECT 317.4 237.16 317.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.395 -1.525 317.725 -1.195 ;
        RECT 317.395 -2.885 317.725 -2.555 ;
        RECT 317.4 -3.56 317.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 317.395 -95.365 317.725 -95.035 ;
        RECT 317.395 -96.725 317.725 -96.395 ;
        RECT 317.395 -98.085 317.725 -97.755 ;
        RECT 317.395 -99.445 317.725 -99.115 ;
        RECT 317.395 -100.805 317.725 -100.475 ;
        RECT 317.395 -102.165 317.725 -101.835 ;
        RECT 317.395 -103.525 317.725 -103.195 ;
        RECT 317.395 -104.885 317.725 -104.555 ;
        RECT 317.395 -106.245 317.725 -105.915 ;
        RECT 317.395 -107.605 317.725 -107.275 ;
        RECT 317.395 -108.965 317.725 -108.635 ;
        RECT 317.395 -110.325 317.725 -109.995 ;
        RECT 317.395 -111.685 317.725 -111.355 ;
        RECT 317.395 -113.045 317.725 -112.715 ;
        RECT 317.395 -114.405 317.725 -114.075 ;
        RECT 317.395 -115.765 317.725 -115.435 ;
        RECT 317.395 -117.125 317.725 -116.795 ;
        RECT 317.395 -118.485 317.725 -118.155 ;
        RECT 317.395 -119.845 317.725 -119.515 ;
        RECT 317.395 -121.205 317.725 -120.875 ;
        RECT 317.395 -122.565 317.725 -122.235 ;
        RECT 317.395 -123.925 317.725 -123.595 ;
        RECT 317.395 -125.285 317.725 -124.955 ;
        RECT 317.395 -126.645 317.725 -126.315 ;
        RECT 317.395 -128.005 317.725 -127.675 ;
        RECT 317.395 -129.365 317.725 -129.035 ;
        RECT 317.395 -130.725 317.725 -130.395 ;
        RECT 317.395 -132.085 317.725 -131.755 ;
        RECT 317.395 -133.445 317.725 -133.115 ;
        RECT 317.395 -134.805 317.725 -134.475 ;
        RECT 317.395 -136.165 317.725 -135.835 ;
        RECT 317.395 -137.525 317.725 -137.195 ;
        RECT 317.395 -138.885 317.725 -138.555 ;
        RECT 317.395 -140.245 317.725 -139.915 ;
        RECT 317.395 -141.605 317.725 -141.275 ;
        RECT 317.395 -142.965 317.725 -142.635 ;
        RECT 317.395 -144.325 317.725 -143.995 ;
        RECT 317.395 -145.685 317.725 -145.355 ;
        RECT 317.395 -147.045 317.725 -146.715 ;
        RECT 317.395 -148.405 317.725 -148.075 ;
        RECT 317.395 -149.765 317.725 -149.435 ;
        RECT 317.395 -151.125 317.725 -150.795 ;
        RECT 317.395 -152.485 317.725 -152.155 ;
        RECT 317.395 -153.845 317.725 -153.515 ;
        RECT 317.395 -155.205 317.725 -154.875 ;
        RECT 317.395 -156.565 317.725 -156.235 ;
        RECT 317.395 -157.925 317.725 -157.595 ;
        RECT 317.395 -159.285 317.725 -158.955 ;
        RECT 317.395 -160.645 317.725 -160.315 ;
        RECT 317.395 -162.005 317.725 -161.675 ;
        RECT 317.395 -163.365 317.725 -163.035 ;
        RECT 317.395 -164.725 317.725 -164.395 ;
        RECT 317.395 -166.085 317.725 -165.755 ;
        RECT 317.395 -167.445 317.725 -167.115 ;
        RECT 317.395 -168.805 317.725 -168.475 ;
        RECT 317.395 -170.165 317.725 -169.835 ;
        RECT 317.395 -171.525 317.725 -171.195 ;
        RECT 317.395 -172.885 317.725 -172.555 ;
        RECT 317.395 -174.245 317.725 -173.915 ;
        RECT 317.395 -175.605 317.725 -175.275 ;
        RECT 317.395 -176.965 317.725 -176.635 ;
        RECT 317.395 -178.325 317.725 -177.995 ;
        RECT 317.395 -179.685 317.725 -179.355 ;
        RECT 317.395 -181.93 317.725 -180.8 ;
        RECT 317.4 -182.045 317.72 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.755 241.32 319.085 242.45 ;
        RECT 318.755 239.195 319.085 239.525 ;
        RECT 318.755 237.835 319.085 238.165 ;
        RECT 318.76 237.16 319.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 318.755 -99.445 319.085 -99.115 ;
        RECT 318.755 -100.805 319.085 -100.475 ;
        RECT 318.755 -102.165 319.085 -101.835 ;
        RECT 318.755 -103.525 319.085 -103.195 ;
        RECT 318.755 -104.885 319.085 -104.555 ;
        RECT 318.755 -106.245 319.085 -105.915 ;
        RECT 318.755 -107.605 319.085 -107.275 ;
        RECT 318.755 -108.965 319.085 -108.635 ;
        RECT 318.755 -110.325 319.085 -109.995 ;
        RECT 318.755 -111.685 319.085 -111.355 ;
        RECT 318.755 -113.045 319.085 -112.715 ;
        RECT 318.755 -114.405 319.085 -114.075 ;
        RECT 318.755 -115.765 319.085 -115.435 ;
        RECT 318.755 -117.125 319.085 -116.795 ;
        RECT 318.755 -118.485 319.085 -118.155 ;
        RECT 318.755 -119.845 319.085 -119.515 ;
        RECT 318.755 -121.205 319.085 -120.875 ;
        RECT 318.755 -122.565 319.085 -122.235 ;
        RECT 318.755 -123.925 319.085 -123.595 ;
        RECT 318.755 -125.285 319.085 -124.955 ;
        RECT 318.755 -126.645 319.085 -126.315 ;
        RECT 318.755 -128.005 319.085 -127.675 ;
        RECT 318.755 -129.365 319.085 -129.035 ;
        RECT 318.755 -130.725 319.085 -130.395 ;
        RECT 318.755 -132.085 319.085 -131.755 ;
        RECT 318.755 -133.445 319.085 -133.115 ;
        RECT 318.755 -134.805 319.085 -134.475 ;
        RECT 318.755 -136.165 319.085 -135.835 ;
        RECT 318.755 -137.525 319.085 -137.195 ;
        RECT 318.755 -138.885 319.085 -138.555 ;
        RECT 318.755 -140.245 319.085 -139.915 ;
        RECT 318.755 -141.605 319.085 -141.275 ;
        RECT 318.755 -142.965 319.085 -142.635 ;
        RECT 318.755 -144.325 319.085 -143.995 ;
        RECT 318.755 -145.685 319.085 -145.355 ;
        RECT 318.755 -147.045 319.085 -146.715 ;
        RECT 318.755 -148.405 319.085 -148.075 ;
        RECT 318.755 -149.765 319.085 -149.435 ;
        RECT 318.755 -151.125 319.085 -150.795 ;
        RECT 318.755 -152.485 319.085 -152.155 ;
        RECT 318.755 -153.845 319.085 -153.515 ;
        RECT 318.755 -155.205 319.085 -154.875 ;
        RECT 318.755 -156.565 319.085 -156.235 ;
        RECT 318.755 -157.925 319.085 -157.595 ;
        RECT 318.755 -159.285 319.085 -158.955 ;
        RECT 318.755 -160.645 319.085 -160.315 ;
        RECT 318.755 -162.005 319.085 -161.675 ;
        RECT 318.755 -163.365 319.085 -163.035 ;
        RECT 318.755 -164.725 319.085 -164.395 ;
        RECT 318.755 -166.085 319.085 -165.755 ;
        RECT 318.755 -167.445 319.085 -167.115 ;
        RECT 318.755 -168.805 319.085 -168.475 ;
        RECT 318.755 -170.165 319.085 -169.835 ;
        RECT 318.755 -171.525 319.085 -171.195 ;
        RECT 318.755 -172.885 319.085 -172.555 ;
        RECT 318.755 -174.245 319.085 -173.915 ;
        RECT 318.755 -175.605 319.085 -175.275 ;
        RECT 318.755 -176.965 319.085 -176.635 ;
        RECT 318.755 -178.325 319.085 -177.995 ;
        RECT 318.755 -179.685 319.085 -179.355 ;
        RECT 318.755 -181.93 319.085 -180.8 ;
        RECT 318.76 -182.045 319.08 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 319.41 -98.075 319.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.115 241.32 320.445 242.45 ;
        RECT 320.115 239.195 320.445 239.525 ;
        RECT 320.115 237.835 320.445 238.165 ;
        RECT 320.12 237.16 320.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 320.115 -1.525 320.445 -1.195 ;
        RECT 320.115 -2.885 320.445 -2.555 ;
        RECT 320.12 -3.56 320.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.475 241.32 321.805 242.45 ;
        RECT 321.475 239.195 321.805 239.525 ;
        RECT 321.475 237.835 321.805 238.165 ;
        RECT 321.48 237.16 321.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 321.475 -1.525 321.805 -1.195 ;
        RECT 321.475 -2.885 321.805 -2.555 ;
        RECT 321.48 -3.56 321.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.835 241.32 323.165 242.45 ;
        RECT 322.835 239.195 323.165 239.525 ;
        RECT 322.835 237.835 323.165 238.165 ;
        RECT 322.84 237.16 323.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.835 -1.525 323.165 -1.195 ;
        RECT 322.835 -2.885 323.165 -2.555 ;
        RECT 322.84 -3.56 323.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 322.835 -95.365 323.165 -95.035 ;
        RECT 322.835 -96.725 323.165 -96.395 ;
        RECT 322.835 -98.085 323.165 -97.755 ;
        RECT 322.835 -99.445 323.165 -99.115 ;
        RECT 322.835 -100.805 323.165 -100.475 ;
        RECT 322.835 -102.165 323.165 -101.835 ;
        RECT 322.835 -103.525 323.165 -103.195 ;
        RECT 322.835 -104.885 323.165 -104.555 ;
        RECT 322.835 -106.245 323.165 -105.915 ;
        RECT 322.835 -107.605 323.165 -107.275 ;
        RECT 322.835 -108.965 323.165 -108.635 ;
        RECT 322.835 -110.325 323.165 -109.995 ;
        RECT 322.835 -111.685 323.165 -111.355 ;
        RECT 322.835 -113.045 323.165 -112.715 ;
        RECT 322.835 -114.405 323.165 -114.075 ;
        RECT 322.835 -115.765 323.165 -115.435 ;
        RECT 322.835 -117.125 323.165 -116.795 ;
        RECT 322.835 -118.485 323.165 -118.155 ;
        RECT 322.835 -119.845 323.165 -119.515 ;
        RECT 322.835 -121.205 323.165 -120.875 ;
        RECT 322.835 -122.565 323.165 -122.235 ;
        RECT 322.835 -123.925 323.165 -123.595 ;
        RECT 322.835 -125.285 323.165 -124.955 ;
        RECT 322.835 -126.645 323.165 -126.315 ;
        RECT 322.835 -128.005 323.165 -127.675 ;
        RECT 322.835 -129.365 323.165 -129.035 ;
        RECT 322.835 -130.725 323.165 -130.395 ;
        RECT 322.835 -132.085 323.165 -131.755 ;
        RECT 322.835 -133.445 323.165 -133.115 ;
        RECT 322.835 -134.805 323.165 -134.475 ;
        RECT 322.835 -136.165 323.165 -135.835 ;
        RECT 322.835 -137.525 323.165 -137.195 ;
        RECT 322.835 -138.885 323.165 -138.555 ;
        RECT 322.835 -140.245 323.165 -139.915 ;
        RECT 322.835 -141.605 323.165 -141.275 ;
        RECT 322.835 -142.965 323.165 -142.635 ;
        RECT 322.835 -144.325 323.165 -143.995 ;
        RECT 322.835 -145.685 323.165 -145.355 ;
        RECT 322.835 -147.045 323.165 -146.715 ;
        RECT 322.835 -148.405 323.165 -148.075 ;
        RECT 322.835 -149.765 323.165 -149.435 ;
        RECT 322.835 -151.125 323.165 -150.795 ;
        RECT 322.835 -152.485 323.165 -152.155 ;
        RECT 322.835 -153.845 323.165 -153.515 ;
        RECT 322.835 -155.205 323.165 -154.875 ;
        RECT 322.835 -156.565 323.165 -156.235 ;
        RECT 322.835 -157.925 323.165 -157.595 ;
        RECT 322.835 -159.285 323.165 -158.955 ;
        RECT 322.835 -160.645 323.165 -160.315 ;
        RECT 322.835 -162.005 323.165 -161.675 ;
        RECT 322.835 -163.365 323.165 -163.035 ;
        RECT 322.835 -164.725 323.165 -164.395 ;
        RECT 322.835 -166.085 323.165 -165.755 ;
        RECT 322.835 -167.445 323.165 -167.115 ;
        RECT 322.835 -168.805 323.165 -168.475 ;
        RECT 322.835 -170.165 323.165 -169.835 ;
        RECT 322.835 -171.525 323.165 -171.195 ;
        RECT 322.835 -172.885 323.165 -172.555 ;
        RECT 322.835 -174.245 323.165 -173.915 ;
        RECT 322.835 -175.605 323.165 -175.275 ;
        RECT 322.835 -176.965 323.165 -176.635 ;
        RECT 322.835 -178.325 323.165 -177.995 ;
        RECT 322.835 -179.685 323.165 -179.355 ;
        RECT 322.835 -181.93 323.165 -180.8 ;
        RECT 322.84 -182.045 323.16 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.195 241.32 324.525 242.45 ;
        RECT 324.195 239.195 324.525 239.525 ;
        RECT 324.195 237.835 324.525 238.165 ;
        RECT 324.2 237.16 324.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.195 -1.525 324.525 -1.195 ;
        RECT 324.195 -2.885 324.525 -2.555 ;
        RECT 324.2 -3.56 324.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 324.195 -95.365 324.525 -95.035 ;
        RECT 324.195 -96.725 324.525 -96.395 ;
        RECT 324.195 -98.085 324.525 -97.755 ;
        RECT 324.195 -99.445 324.525 -99.115 ;
        RECT 324.195 -100.805 324.525 -100.475 ;
        RECT 324.195 -102.165 324.525 -101.835 ;
        RECT 324.195 -103.525 324.525 -103.195 ;
        RECT 324.195 -104.885 324.525 -104.555 ;
        RECT 324.195 -106.245 324.525 -105.915 ;
        RECT 324.195 -107.605 324.525 -107.275 ;
        RECT 324.195 -108.965 324.525 -108.635 ;
        RECT 324.195 -110.325 324.525 -109.995 ;
        RECT 324.195 -111.685 324.525 -111.355 ;
        RECT 324.195 -113.045 324.525 -112.715 ;
        RECT 324.195 -114.405 324.525 -114.075 ;
        RECT 324.195 -115.765 324.525 -115.435 ;
        RECT 324.195 -117.125 324.525 -116.795 ;
        RECT 324.195 -118.485 324.525 -118.155 ;
        RECT 324.195 -119.845 324.525 -119.515 ;
        RECT 324.195 -121.205 324.525 -120.875 ;
        RECT 324.195 -122.565 324.525 -122.235 ;
        RECT 324.195 -123.925 324.525 -123.595 ;
        RECT 324.195 -125.285 324.525 -124.955 ;
        RECT 324.195 -126.645 324.525 -126.315 ;
        RECT 324.195 -128.005 324.525 -127.675 ;
        RECT 324.195 -129.365 324.525 -129.035 ;
        RECT 324.195 -130.725 324.525 -130.395 ;
        RECT 324.195 -132.085 324.525 -131.755 ;
        RECT 324.195 -133.445 324.525 -133.115 ;
        RECT 324.195 -134.805 324.525 -134.475 ;
        RECT 324.195 -136.165 324.525 -135.835 ;
        RECT 324.195 -137.525 324.525 -137.195 ;
        RECT 324.195 -138.885 324.525 -138.555 ;
        RECT 324.195 -140.245 324.525 -139.915 ;
        RECT 324.195 -141.605 324.525 -141.275 ;
        RECT 324.195 -142.965 324.525 -142.635 ;
        RECT 324.195 -144.325 324.525 -143.995 ;
        RECT 324.195 -145.685 324.525 -145.355 ;
        RECT 324.195 -147.045 324.525 -146.715 ;
        RECT 324.195 -148.405 324.525 -148.075 ;
        RECT 324.195 -149.765 324.525 -149.435 ;
        RECT 324.195 -151.125 324.525 -150.795 ;
        RECT 324.195 -152.485 324.525 -152.155 ;
        RECT 324.195 -153.845 324.525 -153.515 ;
        RECT 324.195 -155.205 324.525 -154.875 ;
        RECT 324.195 -156.565 324.525 -156.235 ;
        RECT 324.195 -157.925 324.525 -157.595 ;
        RECT 324.195 -159.285 324.525 -158.955 ;
        RECT 324.195 -160.645 324.525 -160.315 ;
        RECT 324.195 -162.005 324.525 -161.675 ;
        RECT 324.195 -163.365 324.525 -163.035 ;
        RECT 324.195 -164.725 324.525 -164.395 ;
        RECT 324.195 -166.085 324.525 -165.755 ;
        RECT 324.195 -167.445 324.525 -167.115 ;
        RECT 324.195 -168.805 324.525 -168.475 ;
        RECT 324.195 -170.165 324.525 -169.835 ;
        RECT 324.195 -171.525 324.525 -171.195 ;
        RECT 324.195 -172.885 324.525 -172.555 ;
        RECT 324.195 -174.245 324.525 -173.915 ;
        RECT 324.195 -175.605 324.525 -175.275 ;
        RECT 324.195 -176.965 324.525 -176.635 ;
        RECT 324.195 -178.325 324.525 -177.995 ;
        RECT 324.195 -179.685 324.525 -179.355 ;
        RECT 324.195 -181.93 324.525 -180.8 ;
        RECT 324.2 -182.045 324.52 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.555 241.32 325.885 242.45 ;
        RECT 325.555 239.195 325.885 239.525 ;
        RECT 325.555 237.835 325.885 238.165 ;
        RECT 325.56 237.16 325.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.555 -1.525 325.885 -1.195 ;
        RECT 325.555 -2.885 325.885 -2.555 ;
        RECT 325.56 -3.56 325.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 325.555 -95.365 325.885 -95.035 ;
        RECT 325.555 -96.725 325.885 -96.395 ;
        RECT 325.555 -98.085 325.885 -97.755 ;
        RECT 325.555 -99.445 325.885 -99.115 ;
        RECT 325.555 -100.805 325.885 -100.475 ;
        RECT 325.555 -102.165 325.885 -101.835 ;
        RECT 325.555 -103.525 325.885 -103.195 ;
        RECT 325.555 -104.885 325.885 -104.555 ;
        RECT 325.555 -106.245 325.885 -105.915 ;
        RECT 325.555 -107.605 325.885 -107.275 ;
        RECT 325.555 -108.965 325.885 -108.635 ;
        RECT 325.555 -110.325 325.885 -109.995 ;
        RECT 325.555 -111.685 325.885 -111.355 ;
        RECT 325.555 -113.045 325.885 -112.715 ;
        RECT 325.555 -114.405 325.885 -114.075 ;
        RECT 325.555 -115.765 325.885 -115.435 ;
        RECT 325.555 -117.125 325.885 -116.795 ;
        RECT 325.555 -118.485 325.885 -118.155 ;
        RECT 325.555 -119.845 325.885 -119.515 ;
        RECT 325.555 -121.205 325.885 -120.875 ;
        RECT 325.555 -122.565 325.885 -122.235 ;
        RECT 325.555 -123.925 325.885 -123.595 ;
        RECT 325.555 -125.285 325.885 -124.955 ;
        RECT 325.555 -126.645 325.885 -126.315 ;
        RECT 325.555 -128.005 325.885 -127.675 ;
        RECT 325.555 -129.365 325.885 -129.035 ;
        RECT 325.555 -130.725 325.885 -130.395 ;
        RECT 325.555 -132.085 325.885 -131.755 ;
        RECT 325.555 -133.445 325.885 -133.115 ;
        RECT 325.555 -134.805 325.885 -134.475 ;
        RECT 325.555 -136.165 325.885 -135.835 ;
        RECT 325.555 -137.525 325.885 -137.195 ;
        RECT 325.555 -138.885 325.885 -138.555 ;
        RECT 325.555 -140.245 325.885 -139.915 ;
        RECT 325.555 -141.605 325.885 -141.275 ;
        RECT 325.555 -142.965 325.885 -142.635 ;
        RECT 325.555 -144.325 325.885 -143.995 ;
        RECT 325.555 -145.685 325.885 -145.355 ;
        RECT 325.555 -147.045 325.885 -146.715 ;
        RECT 325.555 -148.405 325.885 -148.075 ;
        RECT 325.555 -149.765 325.885 -149.435 ;
        RECT 325.555 -151.125 325.885 -150.795 ;
        RECT 325.555 -152.485 325.885 -152.155 ;
        RECT 325.555 -153.845 325.885 -153.515 ;
        RECT 325.555 -155.205 325.885 -154.875 ;
        RECT 325.555 -156.565 325.885 -156.235 ;
        RECT 325.555 -157.925 325.885 -157.595 ;
        RECT 325.555 -159.285 325.885 -158.955 ;
        RECT 325.555 -160.645 325.885 -160.315 ;
        RECT 325.555 -162.005 325.885 -161.675 ;
        RECT 325.555 -163.365 325.885 -163.035 ;
        RECT 325.555 -164.725 325.885 -164.395 ;
        RECT 325.555 -166.085 325.885 -165.755 ;
        RECT 325.555 -167.445 325.885 -167.115 ;
        RECT 325.555 -168.805 325.885 -168.475 ;
        RECT 325.555 -170.165 325.885 -169.835 ;
        RECT 325.555 -171.525 325.885 -171.195 ;
        RECT 325.555 -172.885 325.885 -172.555 ;
        RECT 325.555 -174.245 325.885 -173.915 ;
        RECT 325.555 -175.605 325.885 -175.275 ;
        RECT 325.555 -176.965 325.885 -176.635 ;
        RECT 325.555 -178.325 325.885 -177.995 ;
        RECT 325.555 -179.685 325.885 -179.355 ;
        RECT 325.555 -181.93 325.885 -180.8 ;
        RECT 325.56 -182.045 325.88 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.915 241.32 327.245 242.45 ;
        RECT 326.915 239.195 327.245 239.525 ;
        RECT 326.915 237.835 327.245 238.165 ;
        RECT 326.92 237.16 327.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.915 -1.525 327.245 -1.195 ;
        RECT 326.915 -2.885 327.245 -2.555 ;
        RECT 326.92 -3.56 327.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 326.915 -95.365 327.245 -95.035 ;
        RECT 326.915 -96.725 327.245 -96.395 ;
        RECT 326.915 -98.085 327.245 -97.755 ;
        RECT 326.915 -99.445 327.245 -99.115 ;
        RECT 326.915 -100.805 327.245 -100.475 ;
        RECT 326.915 -102.165 327.245 -101.835 ;
        RECT 326.915 -103.525 327.245 -103.195 ;
        RECT 326.915 -104.885 327.245 -104.555 ;
        RECT 326.915 -106.245 327.245 -105.915 ;
        RECT 326.915 -107.605 327.245 -107.275 ;
        RECT 326.915 -108.965 327.245 -108.635 ;
        RECT 326.915 -110.325 327.245 -109.995 ;
        RECT 326.915 -111.685 327.245 -111.355 ;
        RECT 326.915 -113.045 327.245 -112.715 ;
        RECT 326.915 -114.405 327.245 -114.075 ;
        RECT 326.915 -115.765 327.245 -115.435 ;
        RECT 326.915 -117.125 327.245 -116.795 ;
        RECT 326.915 -118.485 327.245 -118.155 ;
        RECT 326.915 -119.845 327.245 -119.515 ;
        RECT 326.915 -121.205 327.245 -120.875 ;
        RECT 326.915 -122.565 327.245 -122.235 ;
        RECT 326.915 -123.925 327.245 -123.595 ;
        RECT 326.915 -125.285 327.245 -124.955 ;
        RECT 326.915 -126.645 327.245 -126.315 ;
        RECT 326.915 -128.005 327.245 -127.675 ;
        RECT 326.915 -129.365 327.245 -129.035 ;
        RECT 326.915 -130.725 327.245 -130.395 ;
        RECT 326.915 -132.085 327.245 -131.755 ;
        RECT 326.915 -133.445 327.245 -133.115 ;
        RECT 326.915 -134.805 327.245 -134.475 ;
        RECT 326.915 -136.165 327.245 -135.835 ;
        RECT 326.915 -137.525 327.245 -137.195 ;
        RECT 326.915 -138.885 327.245 -138.555 ;
        RECT 326.915 -140.245 327.245 -139.915 ;
        RECT 326.915 -141.605 327.245 -141.275 ;
        RECT 326.915 -142.965 327.245 -142.635 ;
        RECT 326.915 -144.325 327.245 -143.995 ;
        RECT 326.915 -145.685 327.245 -145.355 ;
        RECT 326.915 -147.045 327.245 -146.715 ;
        RECT 326.915 -148.405 327.245 -148.075 ;
        RECT 326.915 -149.765 327.245 -149.435 ;
        RECT 326.915 -151.125 327.245 -150.795 ;
        RECT 326.915 -152.485 327.245 -152.155 ;
        RECT 326.915 -153.845 327.245 -153.515 ;
        RECT 326.915 -155.205 327.245 -154.875 ;
        RECT 326.915 -156.565 327.245 -156.235 ;
        RECT 326.915 -157.925 327.245 -157.595 ;
        RECT 326.915 -159.285 327.245 -158.955 ;
        RECT 326.915 -160.645 327.245 -160.315 ;
        RECT 326.915 -162.005 327.245 -161.675 ;
        RECT 326.915 -163.365 327.245 -163.035 ;
        RECT 326.915 -164.725 327.245 -164.395 ;
        RECT 326.915 -166.085 327.245 -165.755 ;
        RECT 326.915 -167.445 327.245 -167.115 ;
        RECT 326.915 -168.805 327.245 -168.475 ;
        RECT 326.915 -170.165 327.245 -169.835 ;
        RECT 326.915 -171.525 327.245 -171.195 ;
        RECT 326.915 -172.885 327.245 -172.555 ;
        RECT 326.915 -174.245 327.245 -173.915 ;
        RECT 326.915 -175.605 327.245 -175.275 ;
        RECT 326.915 -176.965 327.245 -176.635 ;
        RECT 326.915 -178.325 327.245 -177.995 ;
        RECT 326.915 -179.685 327.245 -179.355 ;
        RECT 326.915 -181.93 327.245 -180.8 ;
        RECT 326.92 -182.045 327.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.275 241.32 328.605 242.45 ;
        RECT 328.275 239.195 328.605 239.525 ;
        RECT 328.275 237.835 328.605 238.165 ;
        RECT 328.28 237.16 328.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.275 -1.525 328.605 -1.195 ;
        RECT 328.275 -2.885 328.605 -2.555 ;
        RECT 328.28 -3.56 328.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 328.275 -95.365 328.605 -95.035 ;
        RECT 328.275 -96.725 328.605 -96.395 ;
        RECT 328.275 -98.085 328.605 -97.755 ;
        RECT 328.275 -99.445 328.605 -99.115 ;
        RECT 328.275 -100.805 328.605 -100.475 ;
        RECT 328.275 -102.165 328.605 -101.835 ;
        RECT 328.275 -103.525 328.605 -103.195 ;
        RECT 328.275 -104.885 328.605 -104.555 ;
        RECT 328.275 -106.245 328.605 -105.915 ;
        RECT 328.275 -107.605 328.605 -107.275 ;
        RECT 328.275 -108.965 328.605 -108.635 ;
        RECT 328.275 -110.325 328.605 -109.995 ;
        RECT 328.275 -111.685 328.605 -111.355 ;
        RECT 328.275 -113.045 328.605 -112.715 ;
        RECT 328.275 -114.405 328.605 -114.075 ;
        RECT 328.275 -115.765 328.605 -115.435 ;
        RECT 328.275 -117.125 328.605 -116.795 ;
        RECT 328.275 -118.485 328.605 -118.155 ;
        RECT 328.275 -119.845 328.605 -119.515 ;
        RECT 328.275 -121.205 328.605 -120.875 ;
        RECT 328.275 -122.565 328.605 -122.235 ;
        RECT 328.275 -123.925 328.605 -123.595 ;
        RECT 328.275 -125.285 328.605 -124.955 ;
        RECT 328.275 -126.645 328.605 -126.315 ;
        RECT 328.275 -128.005 328.605 -127.675 ;
        RECT 328.275 -129.365 328.605 -129.035 ;
        RECT 328.275 -130.725 328.605 -130.395 ;
        RECT 328.275 -132.085 328.605 -131.755 ;
        RECT 328.275 -133.445 328.605 -133.115 ;
        RECT 328.275 -134.805 328.605 -134.475 ;
        RECT 328.275 -136.165 328.605 -135.835 ;
        RECT 328.275 -137.525 328.605 -137.195 ;
        RECT 328.275 -138.885 328.605 -138.555 ;
        RECT 328.275 -140.245 328.605 -139.915 ;
        RECT 328.275 -141.605 328.605 -141.275 ;
        RECT 328.275 -142.965 328.605 -142.635 ;
        RECT 328.275 -144.325 328.605 -143.995 ;
        RECT 328.275 -145.685 328.605 -145.355 ;
        RECT 328.275 -147.045 328.605 -146.715 ;
        RECT 328.275 -148.405 328.605 -148.075 ;
        RECT 328.275 -149.765 328.605 -149.435 ;
        RECT 328.275 -151.125 328.605 -150.795 ;
        RECT 328.275 -152.485 328.605 -152.155 ;
        RECT 328.275 -153.845 328.605 -153.515 ;
        RECT 328.275 -155.205 328.605 -154.875 ;
        RECT 328.275 -156.565 328.605 -156.235 ;
        RECT 328.275 -157.925 328.605 -157.595 ;
        RECT 328.275 -159.285 328.605 -158.955 ;
        RECT 328.275 -160.645 328.605 -160.315 ;
        RECT 328.275 -162.005 328.605 -161.675 ;
        RECT 328.275 -163.365 328.605 -163.035 ;
        RECT 328.275 -164.725 328.605 -164.395 ;
        RECT 328.275 -166.085 328.605 -165.755 ;
        RECT 328.275 -167.445 328.605 -167.115 ;
        RECT 328.275 -168.805 328.605 -168.475 ;
        RECT 328.275 -170.165 328.605 -169.835 ;
        RECT 328.275 -171.525 328.605 -171.195 ;
        RECT 328.275 -172.885 328.605 -172.555 ;
        RECT 328.275 -174.245 328.605 -173.915 ;
        RECT 328.275 -175.605 328.605 -175.275 ;
        RECT 328.275 -176.965 328.605 -176.635 ;
        RECT 328.275 -178.325 328.605 -177.995 ;
        RECT 328.275 -179.685 328.605 -179.355 ;
        RECT 328.275 -181.93 328.605 -180.8 ;
        RECT 328.28 -182.045 328.6 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.635 241.32 329.965 242.45 ;
        RECT 329.635 239.195 329.965 239.525 ;
        RECT 329.635 237.835 329.965 238.165 ;
        RECT 329.64 237.16 329.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 329.635 -99.445 329.965 -99.115 ;
        RECT 329.635 -100.805 329.965 -100.475 ;
        RECT 329.635 -102.165 329.965 -101.835 ;
        RECT 329.635 -103.525 329.965 -103.195 ;
        RECT 329.635 -104.885 329.965 -104.555 ;
        RECT 329.635 -106.245 329.965 -105.915 ;
        RECT 329.635 -107.605 329.965 -107.275 ;
        RECT 329.635 -108.965 329.965 -108.635 ;
        RECT 329.635 -110.325 329.965 -109.995 ;
        RECT 329.635 -111.685 329.965 -111.355 ;
        RECT 329.635 -113.045 329.965 -112.715 ;
        RECT 329.635 -114.405 329.965 -114.075 ;
        RECT 329.635 -115.765 329.965 -115.435 ;
        RECT 329.635 -117.125 329.965 -116.795 ;
        RECT 329.635 -118.485 329.965 -118.155 ;
        RECT 329.635 -119.845 329.965 -119.515 ;
        RECT 329.635 -121.205 329.965 -120.875 ;
        RECT 329.635 -122.565 329.965 -122.235 ;
        RECT 329.635 -123.925 329.965 -123.595 ;
        RECT 329.635 -125.285 329.965 -124.955 ;
        RECT 329.635 -126.645 329.965 -126.315 ;
        RECT 329.635 -128.005 329.965 -127.675 ;
        RECT 329.635 -129.365 329.965 -129.035 ;
        RECT 329.635 -130.725 329.965 -130.395 ;
        RECT 329.635 -132.085 329.965 -131.755 ;
        RECT 329.635 -133.445 329.965 -133.115 ;
        RECT 329.635 -134.805 329.965 -134.475 ;
        RECT 329.635 -136.165 329.965 -135.835 ;
        RECT 329.635 -137.525 329.965 -137.195 ;
        RECT 329.635 -138.885 329.965 -138.555 ;
        RECT 329.635 -140.245 329.965 -139.915 ;
        RECT 329.635 -141.605 329.965 -141.275 ;
        RECT 329.635 -142.965 329.965 -142.635 ;
        RECT 329.635 -144.325 329.965 -143.995 ;
        RECT 329.635 -145.685 329.965 -145.355 ;
        RECT 329.635 -147.045 329.965 -146.715 ;
        RECT 329.635 -148.405 329.965 -148.075 ;
        RECT 329.635 -149.765 329.965 -149.435 ;
        RECT 329.635 -151.125 329.965 -150.795 ;
        RECT 329.635 -152.485 329.965 -152.155 ;
        RECT 329.635 -153.845 329.965 -153.515 ;
        RECT 329.635 -155.205 329.965 -154.875 ;
        RECT 329.635 -156.565 329.965 -156.235 ;
        RECT 329.635 -157.925 329.965 -157.595 ;
        RECT 329.635 -159.285 329.965 -158.955 ;
        RECT 329.635 -160.645 329.965 -160.315 ;
        RECT 329.635 -162.005 329.965 -161.675 ;
        RECT 329.635 -163.365 329.965 -163.035 ;
        RECT 329.635 -164.725 329.965 -164.395 ;
        RECT 329.635 -166.085 329.965 -165.755 ;
        RECT 329.635 -167.445 329.965 -167.115 ;
        RECT 329.635 -168.805 329.965 -168.475 ;
        RECT 329.635 -170.165 329.965 -169.835 ;
        RECT 329.635 -171.525 329.965 -171.195 ;
        RECT 329.635 -172.885 329.965 -172.555 ;
        RECT 329.635 -174.245 329.965 -173.915 ;
        RECT 329.635 -175.605 329.965 -175.275 ;
        RECT 329.635 -176.965 329.965 -176.635 ;
        RECT 329.635 -178.325 329.965 -177.995 ;
        RECT 329.635 -179.685 329.965 -179.355 ;
        RECT 329.635 -181.93 329.965 -180.8 ;
        RECT 329.64 -182.045 329.96 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.31 -98.075 330.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.995 241.32 331.325 242.45 ;
        RECT 330.995 239.195 331.325 239.525 ;
        RECT 330.995 237.835 331.325 238.165 ;
        RECT 331 237.16 331.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 330.995 -1.525 331.325 -1.195 ;
        RECT 330.995 -2.885 331.325 -2.555 ;
        RECT 331 -3.56 331.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.355 241.32 332.685 242.45 ;
        RECT 332.355 239.195 332.685 239.525 ;
        RECT 332.355 237.835 332.685 238.165 ;
        RECT 332.36 237.16 332.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 332.355 -1.525 332.685 -1.195 ;
        RECT 332.355 -2.885 332.685 -2.555 ;
        RECT 332.36 -3.56 332.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.715 241.32 334.045 242.45 ;
        RECT 333.715 239.195 334.045 239.525 ;
        RECT 333.715 237.835 334.045 238.165 ;
        RECT 333.72 237.16 334.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.715 -1.525 334.045 -1.195 ;
        RECT 333.715 -2.885 334.045 -2.555 ;
        RECT 333.72 -3.56 334.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 333.715 -95.365 334.045 -95.035 ;
        RECT 333.715 -96.725 334.045 -96.395 ;
        RECT 333.715 -98.085 334.045 -97.755 ;
        RECT 333.715 -99.445 334.045 -99.115 ;
        RECT 333.715 -100.805 334.045 -100.475 ;
        RECT 333.715 -102.165 334.045 -101.835 ;
        RECT 333.715 -103.525 334.045 -103.195 ;
        RECT 333.715 -104.885 334.045 -104.555 ;
        RECT 333.715 -106.245 334.045 -105.915 ;
        RECT 333.715 -107.605 334.045 -107.275 ;
        RECT 333.715 -108.965 334.045 -108.635 ;
        RECT 333.715 -110.325 334.045 -109.995 ;
        RECT 333.715 -111.685 334.045 -111.355 ;
        RECT 333.715 -113.045 334.045 -112.715 ;
        RECT 333.715 -114.405 334.045 -114.075 ;
        RECT 333.715 -115.765 334.045 -115.435 ;
        RECT 333.715 -117.125 334.045 -116.795 ;
        RECT 333.715 -118.485 334.045 -118.155 ;
        RECT 333.715 -119.845 334.045 -119.515 ;
        RECT 333.715 -121.205 334.045 -120.875 ;
        RECT 333.715 -122.565 334.045 -122.235 ;
        RECT 333.715 -123.925 334.045 -123.595 ;
        RECT 333.715 -125.285 334.045 -124.955 ;
        RECT 333.715 -126.645 334.045 -126.315 ;
        RECT 333.715 -128.005 334.045 -127.675 ;
        RECT 333.715 -129.365 334.045 -129.035 ;
        RECT 333.715 -130.725 334.045 -130.395 ;
        RECT 333.715 -132.085 334.045 -131.755 ;
        RECT 333.715 -133.445 334.045 -133.115 ;
        RECT 333.715 -134.805 334.045 -134.475 ;
        RECT 333.715 -136.165 334.045 -135.835 ;
        RECT 333.715 -137.525 334.045 -137.195 ;
        RECT 333.715 -138.885 334.045 -138.555 ;
        RECT 333.715 -140.245 334.045 -139.915 ;
        RECT 333.715 -141.605 334.045 -141.275 ;
        RECT 333.715 -142.965 334.045 -142.635 ;
        RECT 333.715 -144.325 334.045 -143.995 ;
        RECT 333.715 -145.685 334.045 -145.355 ;
        RECT 333.715 -147.045 334.045 -146.715 ;
        RECT 333.715 -148.405 334.045 -148.075 ;
        RECT 333.715 -149.765 334.045 -149.435 ;
        RECT 333.715 -151.125 334.045 -150.795 ;
        RECT 333.715 -152.485 334.045 -152.155 ;
        RECT 333.715 -153.845 334.045 -153.515 ;
        RECT 333.715 -155.205 334.045 -154.875 ;
        RECT 333.715 -156.565 334.045 -156.235 ;
        RECT 333.715 -157.925 334.045 -157.595 ;
        RECT 333.715 -159.285 334.045 -158.955 ;
        RECT 333.715 -160.645 334.045 -160.315 ;
        RECT 333.715 -162.005 334.045 -161.675 ;
        RECT 333.715 -163.365 334.045 -163.035 ;
        RECT 333.715 -164.725 334.045 -164.395 ;
        RECT 333.715 -166.085 334.045 -165.755 ;
        RECT 333.715 -167.445 334.045 -167.115 ;
        RECT 333.715 -168.805 334.045 -168.475 ;
        RECT 333.715 -170.165 334.045 -169.835 ;
        RECT 333.715 -171.525 334.045 -171.195 ;
        RECT 333.715 -172.885 334.045 -172.555 ;
        RECT 333.715 -174.245 334.045 -173.915 ;
        RECT 333.715 -175.605 334.045 -175.275 ;
        RECT 333.715 -176.965 334.045 -176.635 ;
        RECT 333.715 -178.325 334.045 -177.995 ;
        RECT 333.715 -179.685 334.045 -179.355 ;
        RECT 333.715 -181.93 334.045 -180.8 ;
        RECT 333.72 -182.045 334.04 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.075 241.32 335.405 242.45 ;
        RECT 335.075 239.195 335.405 239.525 ;
        RECT 335.075 237.835 335.405 238.165 ;
        RECT 335.08 237.16 335.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.075 -1.525 335.405 -1.195 ;
        RECT 335.075 -2.885 335.405 -2.555 ;
        RECT 335.08 -3.56 335.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 335.075 -95.365 335.405 -95.035 ;
        RECT 335.075 -96.725 335.405 -96.395 ;
        RECT 335.075 -98.085 335.405 -97.755 ;
        RECT 335.075 -99.445 335.405 -99.115 ;
        RECT 335.075 -100.805 335.405 -100.475 ;
        RECT 335.075 -102.165 335.405 -101.835 ;
        RECT 335.075 -103.525 335.405 -103.195 ;
        RECT 335.075 -104.885 335.405 -104.555 ;
        RECT 335.075 -106.245 335.405 -105.915 ;
        RECT 335.075 -107.605 335.405 -107.275 ;
        RECT 335.075 -108.965 335.405 -108.635 ;
        RECT 335.075 -110.325 335.405 -109.995 ;
        RECT 335.075 -111.685 335.405 -111.355 ;
        RECT 335.075 -113.045 335.405 -112.715 ;
        RECT 335.075 -114.405 335.405 -114.075 ;
        RECT 335.075 -115.765 335.405 -115.435 ;
        RECT 335.075 -117.125 335.405 -116.795 ;
        RECT 335.075 -118.485 335.405 -118.155 ;
        RECT 335.075 -119.845 335.405 -119.515 ;
        RECT 335.075 -121.205 335.405 -120.875 ;
        RECT 335.075 -122.565 335.405 -122.235 ;
        RECT 335.075 -123.925 335.405 -123.595 ;
        RECT 335.075 -125.285 335.405 -124.955 ;
        RECT 335.075 -126.645 335.405 -126.315 ;
        RECT 335.075 -128.005 335.405 -127.675 ;
        RECT 335.075 -129.365 335.405 -129.035 ;
        RECT 335.075 -130.725 335.405 -130.395 ;
        RECT 335.075 -132.085 335.405 -131.755 ;
        RECT 335.075 -133.445 335.405 -133.115 ;
        RECT 335.075 -134.805 335.405 -134.475 ;
        RECT 335.075 -136.165 335.405 -135.835 ;
        RECT 335.075 -137.525 335.405 -137.195 ;
        RECT 335.075 -138.885 335.405 -138.555 ;
        RECT 335.075 -140.245 335.405 -139.915 ;
        RECT 335.075 -141.605 335.405 -141.275 ;
        RECT 335.075 -142.965 335.405 -142.635 ;
        RECT 335.075 -144.325 335.405 -143.995 ;
        RECT 335.075 -145.685 335.405 -145.355 ;
        RECT 335.075 -147.045 335.405 -146.715 ;
        RECT 335.075 -148.405 335.405 -148.075 ;
        RECT 335.075 -149.765 335.405 -149.435 ;
        RECT 335.075 -151.125 335.405 -150.795 ;
        RECT 335.075 -152.485 335.405 -152.155 ;
        RECT 335.075 -153.845 335.405 -153.515 ;
        RECT 335.075 -155.205 335.405 -154.875 ;
        RECT 335.075 -156.565 335.405 -156.235 ;
        RECT 335.075 -157.925 335.405 -157.595 ;
        RECT 335.075 -159.285 335.405 -158.955 ;
        RECT 335.075 -160.645 335.405 -160.315 ;
        RECT 335.075 -162.005 335.405 -161.675 ;
        RECT 335.075 -163.365 335.405 -163.035 ;
        RECT 335.075 -164.725 335.405 -164.395 ;
        RECT 335.075 -166.085 335.405 -165.755 ;
        RECT 335.075 -167.445 335.405 -167.115 ;
        RECT 335.075 -168.805 335.405 -168.475 ;
        RECT 335.075 -170.165 335.405 -169.835 ;
        RECT 335.075 -171.525 335.405 -171.195 ;
        RECT 335.075 -172.885 335.405 -172.555 ;
        RECT 335.075 -174.245 335.405 -173.915 ;
        RECT 335.075 -175.605 335.405 -175.275 ;
        RECT 335.075 -176.965 335.405 -176.635 ;
        RECT 335.075 -178.325 335.405 -177.995 ;
        RECT 335.075 -179.685 335.405 -179.355 ;
        RECT 335.075 -181.93 335.405 -180.8 ;
        RECT 335.08 -182.045 335.4 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.435 241.32 336.765 242.45 ;
        RECT 336.435 239.195 336.765 239.525 ;
        RECT 336.435 237.835 336.765 238.165 ;
        RECT 336.44 237.16 336.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.435 -1.525 336.765 -1.195 ;
        RECT 336.435 -2.885 336.765 -2.555 ;
        RECT 336.44 -3.56 336.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 336.435 -95.365 336.765 -95.035 ;
        RECT 336.435 -96.725 336.765 -96.395 ;
        RECT 336.435 -98.085 336.765 -97.755 ;
        RECT 336.435 -99.445 336.765 -99.115 ;
        RECT 336.435 -100.805 336.765 -100.475 ;
        RECT 336.435 -102.165 336.765 -101.835 ;
        RECT 336.435 -103.525 336.765 -103.195 ;
        RECT 336.435 -104.885 336.765 -104.555 ;
        RECT 336.435 -106.245 336.765 -105.915 ;
        RECT 336.435 -107.605 336.765 -107.275 ;
        RECT 336.435 -108.965 336.765 -108.635 ;
        RECT 336.435 -110.325 336.765 -109.995 ;
        RECT 336.435 -111.685 336.765 -111.355 ;
        RECT 336.435 -113.045 336.765 -112.715 ;
        RECT 336.435 -114.405 336.765 -114.075 ;
        RECT 336.435 -115.765 336.765 -115.435 ;
        RECT 336.435 -117.125 336.765 -116.795 ;
        RECT 336.435 -118.485 336.765 -118.155 ;
        RECT 336.435 -119.845 336.765 -119.515 ;
        RECT 336.435 -121.205 336.765 -120.875 ;
        RECT 336.435 -122.565 336.765 -122.235 ;
        RECT 336.435 -123.925 336.765 -123.595 ;
        RECT 336.435 -125.285 336.765 -124.955 ;
        RECT 336.435 -126.645 336.765 -126.315 ;
        RECT 336.435 -128.005 336.765 -127.675 ;
        RECT 336.435 -129.365 336.765 -129.035 ;
        RECT 336.435 -130.725 336.765 -130.395 ;
        RECT 336.435 -132.085 336.765 -131.755 ;
        RECT 336.435 -133.445 336.765 -133.115 ;
        RECT 336.435 -134.805 336.765 -134.475 ;
        RECT 336.435 -136.165 336.765 -135.835 ;
        RECT 336.435 -137.525 336.765 -137.195 ;
        RECT 336.435 -138.885 336.765 -138.555 ;
        RECT 336.435 -140.245 336.765 -139.915 ;
        RECT 336.435 -141.605 336.765 -141.275 ;
        RECT 336.435 -142.965 336.765 -142.635 ;
        RECT 336.435 -144.325 336.765 -143.995 ;
        RECT 336.435 -145.685 336.765 -145.355 ;
        RECT 336.435 -147.045 336.765 -146.715 ;
        RECT 336.435 -148.405 336.765 -148.075 ;
        RECT 336.435 -149.765 336.765 -149.435 ;
        RECT 336.435 -151.125 336.765 -150.795 ;
        RECT 336.435 -152.485 336.765 -152.155 ;
        RECT 336.435 -153.845 336.765 -153.515 ;
        RECT 336.435 -155.205 336.765 -154.875 ;
        RECT 336.435 -156.565 336.765 -156.235 ;
        RECT 336.435 -157.925 336.765 -157.595 ;
        RECT 336.435 -159.285 336.765 -158.955 ;
        RECT 336.435 -160.645 336.765 -160.315 ;
        RECT 336.435 -162.005 336.765 -161.675 ;
        RECT 336.435 -163.365 336.765 -163.035 ;
        RECT 336.435 -164.725 336.765 -164.395 ;
        RECT 336.435 -166.085 336.765 -165.755 ;
        RECT 336.435 -167.445 336.765 -167.115 ;
        RECT 336.435 -168.805 336.765 -168.475 ;
        RECT 336.435 -170.165 336.765 -169.835 ;
        RECT 336.435 -171.525 336.765 -171.195 ;
        RECT 336.435 -172.885 336.765 -172.555 ;
        RECT 336.435 -174.245 336.765 -173.915 ;
        RECT 336.435 -175.605 336.765 -175.275 ;
        RECT 336.435 -176.965 336.765 -176.635 ;
        RECT 336.435 -178.325 336.765 -177.995 ;
        RECT 336.435 -179.685 336.765 -179.355 ;
        RECT 336.435 -181.93 336.765 -180.8 ;
        RECT 336.44 -182.045 336.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.795 241.32 338.125 242.45 ;
        RECT 337.795 239.195 338.125 239.525 ;
        RECT 337.795 237.835 338.125 238.165 ;
        RECT 337.8 237.16 338.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.795 -1.525 338.125 -1.195 ;
        RECT 337.795 -2.885 338.125 -2.555 ;
        RECT 337.8 -3.56 338.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 337.795 -100.805 338.125 -100.475 ;
        RECT 337.795 -102.165 338.125 -101.835 ;
        RECT 337.795 -103.525 338.125 -103.195 ;
        RECT 337.795 -104.885 338.125 -104.555 ;
        RECT 337.795 -106.245 338.125 -105.915 ;
        RECT 337.795 -107.605 338.125 -107.275 ;
        RECT 337.795 -108.965 338.125 -108.635 ;
        RECT 337.795 -110.325 338.125 -109.995 ;
        RECT 337.795 -111.685 338.125 -111.355 ;
        RECT 337.795 -113.045 338.125 -112.715 ;
        RECT 337.795 -114.405 338.125 -114.075 ;
        RECT 337.795 -115.765 338.125 -115.435 ;
        RECT 337.795 -117.125 338.125 -116.795 ;
        RECT 337.795 -118.485 338.125 -118.155 ;
        RECT 337.795 -119.845 338.125 -119.515 ;
        RECT 337.795 -121.205 338.125 -120.875 ;
        RECT 337.795 -122.565 338.125 -122.235 ;
        RECT 337.795 -123.925 338.125 -123.595 ;
        RECT 337.795 -125.285 338.125 -124.955 ;
        RECT 337.795 -126.645 338.125 -126.315 ;
        RECT 337.795 -128.005 338.125 -127.675 ;
        RECT 337.795 -129.365 338.125 -129.035 ;
        RECT 337.795 -130.725 338.125 -130.395 ;
        RECT 337.795 -132.085 338.125 -131.755 ;
        RECT 337.795 -133.445 338.125 -133.115 ;
        RECT 337.795 -134.805 338.125 -134.475 ;
        RECT 337.795 -136.165 338.125 -135.835 ;
        RECT 337.795 -137.525 338.125 -137.195 ;
        RECT 337.795 -138.885 338.125 -138.555 ;
        RECT 337.795 -140.245 338.125 -139.915 ;
        RECT 337.795 -141.605 338.125 -141.275 ;
        RECT 337.795 -142.965 338.125 -142.635 ;
        RECT 337.795 -144.325 338.125 -143.995 ;
        RECT 337.795 -145.685 338.125 -145.355 ;
        RECT 337.795 -147.045 338.125 -146.715 ;
        RECT 337.795 -148.405 338.125 -148.075 ;
        RECT 337.795 -149.765 338.125 -149.435 ;
        RECT 337.795 -151.125 338.125 -150.795 ;
        RECT 337.795 -152.485 338.125 -152.155 ;
        RECT 337.795 -153.845 338.125 -153.515 ;
        RECT 337.795 -155.205 338.125 -154.875 ;
        RECT 337.795 -156.565 338.125 -156.235 ;
        RECT 337.795 -157.925 338.125 -157.595 ;
        RECT 337.795 -159.285 338.125 -158.955 ;
        RECT 337.795 -160.645 338.125 -160.315 ;
        RECT 337.795 -162.005 338.125 -161.675 ;
        RECT 337.795 -163.365 338.125 -163.035 ;
        RECT 337.795 -164.725 338.125 -164.395 ;
        RECT 337.795 -166.085 338.125 -165.755 ;
        RECT 337.795 -167.445 338.125 -167.115 ;
        RECT 337.795 -168.805 338.125 -168.475 ;
        RECT 337.795 -170.165 338.125 -169.835 ;
        RECT 337.795 -171.525 338.125 -171.195 ;
        RECT 337.795 -172.885 338.125 -172.555 ;
        RECT 337.795 -174.245 338.125 -173.915 ;
        RECT 337.795 -175.605 338.125 -175.275 ;
        RECT 337.795 -176.965 338.125 -176.635 ;
        RECT 337.795 -178.325 338.125 -177.995 ;
        RECT 337.795 -179.685 338.125 -179.355 ;
        RECT 337.795 -181.93 338.125 -180.8 ;
        RECT 337.8 -182.045 338.12 -95.035 ;
        RECT 337.795 -95.365 338.125 -95.035 ;
        RECT 337.795 -96.725 338.125 -96.395 ;
        RECT 337.795 -98.085 338.125 -97.755 ;
        RECT 337.795 -99.445 338.125 -99.115 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.555 241.32 291.885 242.45 ;
        RECT 291.555 239.195 291.885 239.525 ;
        RECT 291.555 237.835 291.885 238.165 ;
        RECT 291.56 237.16 291.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.555 -1.525 291.885 -1.195 ;
        RECT 291.555 -2.885 291.885 -2.555 ;
        RECT 291.56 -3.56 291.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 291.555 -95.365 291.885 -95.035 ;
        RECT 291.555 -96.725 291.885 -96.395 ;
        RECT 291.555 -98.085 291.885 -97.755 ;
        RECT 291.555 -99.445 291.885 -99.115 ;
        RECT 291.555 -100.805 291.885 -100.475 ;
        RECT 291.555 -102.165 291.885 -101.835 ;
        RECT 291.555 -103.525 291.885 -103.195 ;
        RECT 291.555 -104.885 291.885 -104.555 ;
        RECT 291.555 -106.245 291.885 -105.915 ;
        RECT 291.555 -107.605 291.885 -107.275 ;
        RECT 291.555 -108.965 291.885 -108.635 ;
        RECT 291.555 -110.325 291.885 -109.995 ;
        RECT 291.555 -111.685 291.885 -111.355 ;
        RECT 291.555 -113.045 291.885 -112.715 ;
        RECT 291.555 -114.405 291.885 -114.075 ;
        RECT 291.555 -115.765 291.885 -115.435 ;
        RECT 291.555 -117.125 291.885 -116.795 ;
        RECT 291.555 -118.485 291.885 -118.155 ;
        RECT 291.555 -119.845 291.885 -119.515 ;
        RECT 291.555 -121.205 291.885 -120.875 ;
        RECT 291.555 -122.565 291.885 -122.235 ;
        RECT 291.555 -123.925 291.885 -123.595 ;
        RECT 291.555 -125.285 291.885 -124.955 ;
        RECT 291.555 -126.645 291.885 -126.315 ;
        RECT 291.555 -128.005 291.885 -127.675 ;
        RECT 291.555 -129.365 291.885 -129.035 ;
        RECT 291.555 -130.725 291.885 -130.395 ;
        RECT 291.555 -132.085 291.885 -131.755 ;
        RECT 291.555 -133.445 291.885 -133.115 ;
        RECT 291.555 -134.805 291.885 -134.475 ;
        RECT 291.555 -136.165 291.885 -135.835 ;
        RECT 291.555 -137.525 291.885 -137.195 ;
        RECT 291.555 -138.885 291.885 -138.555 ;
        RECT 291.555 -140.245 291.885 -139.915 ;
        RECT 291.555 -141.605 291.885 -141.275 ;
        RECT 291.555 -142.965 291.885 -142.635 ;
        RECT 291.555 -144.325 291.885 -143.995 ;
        RECT 291.555 -145.685 291.885 -145.355 ;
        RECT 291.555 -147.045 291.885 -146.715 ;
        RECT 291.555 -148.405 291.885 -148.075 ;
        RECT 291.555 -149.765 291.885 -149.435 ;
        RECT 291.555 -151.125 291.885 -150.795 ;
        RECT 291.555 -152.485 291.885 -152.155 ;
        RECT 291.555 -153.845 291.885 -153.515 ;
        RECT 291.555 -155.205 291.885 -154.875 ;
        RECT 291.555 -156.565 291.885 -156.235 ;
        RECT 291.555 -157.925 291.885 -157.595 ;
        RECT 291.555 -159.285 291.885 -158.955 ;
        RECT 291.555 -160.645 291.885 -160.315 ;
        RECT 291.555 -162.005 291.885 -161.675 ;
        RECT 291.555 -163.365 291.885 -163.035 ;
        RECT 291.555 -164.725 291.885 -164.395 ;
        RECT 291.555 -166.085 291.885 -165.755 ;
        RECT 291.555 -167.445 291.885 -167.115 ;
        RECT 291.555 -168.805 291.885 -168.475 ;
        RECT 291.555 -170.165 291.885 -169.835 ;
        RECT 291.555 -171.525 291.885 -171.195 ;
        RECT 291.555 -172.885 291.885 -172.555 ;
        RECT 291.555 -174.245 291.885 -173.915 ;
        RECT 291.555 -175.605 291.885 -175.275 ;
        RECT 291.555 -176.965 291.885 -176.635 ;
        RECT 291.555 -178.325 291.885 -177.995 ;
        RECT 291.555 -179.685 291.885 -179.355 ;
        RECT 291.555 -181.93 291.885 -180.8 ;
        RECT 291.56 -182.045 291.88 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.915 241.32 293.245 242.45 ;
        RECT 292.915 239.195 293.245 239.525 ;
        RECT 292.915 237.835 293.245 238.165 ;
        RECT 292.92 237.16 293.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.915 -1.525 293.245 -1.195 ;
        RECT 292.915 -2.885 293.245 -2.555 ;
        RECT 292.92 -3.56 293.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 292.915 -95.365 293.245 -95.035 ;
        RECT 292.915 -96.725 293.245 -96.395 ;
        RECT 292.915 -98.085 293.245 -97.755 ;
        RECT 292.915 -99.445 293.245 -99.115 ;
        RECT 292.915 -100.805 293.245 -100.475 ;
        RECT 292.915 -102.165 293.245 -101.835 ;
        RECT 292.915 -103.525 293.245 -103.195 ;
        RECT 292.915 -104.885 293.245 -104.555 ;
        RECT 292.915 -106.245 293.245 -105.915 ;
        RECT 292.915 -107.605 293.245 -107.275 ;
        RECT 292.915 -108.965 293.245 -108.635 ;
        RECT 292.915 -110.325 293.245 -109.995 ;
        RECT 292.915 -111.685 293.245 -111.355 ;
        RECT 292.915 -113.045 293.245 -112.715 ;
        RECT 292.915 -114.405 293.245 -114.075 ;
        RECT 292.915 -115.765 293.245 -115.435 ;
        RECT 292.915 -117.125 293.245 -116.795 ;
        RECT 292.915 -118.485 293.245 -118.155 ;
        RECT 292.915 -119.845 293.245 -119.515 ;
        RECT 292.915 -121.205 293.245 -120.875 ;
        RECT 292.915 -122.565 293.245 -122.235 ;
        RECT 292.915 -123.925 293.245 -123.595 ;
        RECT 292.915 -125.285 293.245 -124.955 ;
        RECT 292.915 -126.645 293.245 -126.315 ;
        RECT 292.915 -128.005 293.245 -127.675 ;
        RECT 292.915 -129.365 293.245 -129.035 ;
        RECT 292.915 -130.725 293.245 -130.395 ;
        RECT 292.915 -132.085 293.245 -131.755 ;
        RECT 292.915 -133.445 293.245 -133.115 ;
        RECT 292.915 -134.805 293.245 -134.475 ;
        RECT 292.915 -136.165 293.245 -135.835 ;
        RECT 292.915 -137.525 293.245 -137.195 ;
        RECT 292.915 -138.885 293.245 -138.555 ;
        RECT 292.915 -140.245 293.245 -139.915 ;
        RECT 292.915 -141.605 293.245 -141.275 ;
        RECT 292.915 -142.965 293.245 -142.635 ;
        RECT 292.915 -144.325 293.245 -143.995 ;
        RECT 292.915 -145.685 293.245 -145.355 ;
        RECT 292.915 -147.045 293.245 -146.715 ;
        RECT 292.915 -148.405 293.245 -148.075 ;
        RECT 292.915 -149.765 293.245 -149.435 ;
        RECT 292.915 -151.125 293.245 -150.795 ;
        RECT 292.915 -152.485 293.245 -152.155 ;
        RECT 292.915 -153.845 293.245 -153.515 ;
        RECT 292.915 -155.205 293.245 -154.875 ;
        RECT 292.915 -156.565 293.245 -156.235 ;
        RECT 292.915 -157.925 293.245 -157.595 ;
        RECT 292.915 -159.285 293.245 -158.955 ;
        RECT 292.915 -160.645 293.245 -160.315 ;
        RECT 292.915 -162.005 293.245 -161.675 ;
        RECT 292.915 -163.365 293.245 -163.035 ;
        RECT 292.915 -164.725 293.245 -164.395 ;
        RECT 292.915 -166.085 293.245 -165.755 ;
        RECT 292.915 -167.445 293.245 -167.115 ;
        RECT 292.915 -168.805 293.245 -168.475 ;
        RECT 292.915 -170.165 293.245 -169.835 ;
        RECT 292.915 -171.525 293.245 -171.195 ;
        RECT 292.915 -172.885 293.245 -172.555 ;
        RECT 292.915 -174.245 293.245 -173.915 ;
        RECT 292.915 -175.605 293.245 -175.275 ;
        RECT 292.915 -176.965 293.245 -176.635 ;
        RECT 292.915 -178.325 293.245 -177.995 ;
        RECT 292.915 -179.685 293.245 -179.355 ;
        RECT 292.915 -181.93 293.245 -180.8 ;
        RECT 292.92 -182.045 293.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.275 241.32 294.605 242.45 ;
        RECT 294.275 239.195 294.605 239.525 ;
        RECT 294.275 237.835 294.605 238.165 ;
        RECT 294.28 237.16 294.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.275 -1.525 294.605 -1.195 ;
        RECT 294.275 -2.885 294.605 -2.555 ;
        RECT 294.28 -3.56 294.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 294.275 -95.365 294.605 -95.035 ;
        RECT 294.275 -96.725 294.605 -96.395 ;
        RECT 294.275 -98.085 294.605 -97.755 ;
        RECT 294.275 -99.445 294.605 -99.115 ;
        RECT 294.275 -100.805 294.605 -100.475 ;
        RECT 294.275 -102.165 294.605 -101.835 ;
        RECT 294.275 -103.525 294.605 -103.195 ;
        RECT 294.275 -104.885 294.605 -104.555 ;
        RECT 294.275 -106.245 294.605 -105.915 ;
        RECT 294.275 -107.605 294.605 -107.275 ;
        RECT 294.275 -108.965 294.605 -108.635 ;
        RECT 294.275 -110.325 294.605 -109.995 ;
        RECT 294.275 -111.685 294.605 -111.355 ;
        RECT 294.275 -113.045 294.605 -112.715 ;
        RECT 294.275 -114.405 294.605 -114.075 ;
        RECT 294.275 -115.765 294.605 -115.435 ;
        RECT 294.275 -117.125 294.605 -116.795 ;
        RECT 294.275 -118.485 294.605 -118.155 ;
        RECT 294.275 -119.845 294.605 -119.515 ;
        RECT 294.275 -121.205 294.605 -120.875 ;
        RECT 294.275 -122.565 294.605 -122.235 ;
        RECT 294.275 -123.925 294.605 -123.595 ;
        RECT 294.275 -125.285 294.605 -124.955 ;
        RECT 294.275 -126.645 294.605 -126.315 ;
        RECT 294.275 -128.005 294.605 -127.675 ;
        RECT 294.275 -129.365 294.605 -129.035 ;
        RECT 294.275 -130.725 294.605 -130.395 ;
        RECT 294.275 -132.085 294.605 -131.755 ;
        RECT 294.275 -133.445 294.605 -133.115 ;
        RECT 294.275 -134.805 294.605 -134.475 ;
        RECT 294.275 -136.165 294.605 -135.835 ;
        RECT 294.275 -137.525 294.605 -137.195 ;
        RECT 294.275 -138.885 294.605 -138.555 ;
        RECT 294.275 -140.245 294.605 -139.915 ;
        RECT 294.275 -141.605 294.605 -141.275 ;
        RECT 294.275 -142.965 294.605 -142.635 ;
        RECT 294.275 -144.325 294.605 -143.995 ;
        RECT 294.275 -145.685 294.605 -145.355 ;
        RECT 294.275 -147.045 294.605 -146.715 ;
        RECT 294.275 -148.405 294.605 -148.075 ;
        RECT 294.275 -149.765 294.605 -149.435 ;
        RECT 294.275 -151.125 294.605 -150.795 ;
        RECT 294.275 -152.485 294.605 -152.155 ;
        RECT 294.275 -153.845 294.605 -153.515 ;
        RECT 294.275 -155.205 294.605 -154.875 ;
        RECT 294.275 -156.565 294.605 -156.235 ;
        RECT 294.275 -157.925 294.605 -157.595 ;
        RECT 294.275 -159.285 294.605 -158.955 ;
        RECT 294.275 -160.645 294.605 -160.315 ;
        RECT 294.275 -162.005 294.605 -161.675 ;
        RECT 294.275 -163.365 294.605 -163.035 ;
        RECT 294.275 -164.725 294.605 -164.395 ;
        RECT 294.275 -166.085 294.605 -165.755 ;
        RECT 294.275 -167.445 294.605 -167.115 ;
        RECT 294.275 -168.805 294.605 -168.475 ;
        RECT 294.275 -170.165 294.605 -169.835 ;
        RECT 294.275 -171.525 294.605 -171.195 ;
        RECT 294.275 -172.885 294.605 -172.555 ;
        RECT 294.275 -174.245 294.605 -173.915 ;
        RECT 294.275 -175.605 294.605 -175.275 ;
        RECT 294.275 -176.965 294.605 -176.635 ;
        RECT 294.275 -178.325 294.605 -177.995 ;
        RECT 294.275 -179.685 294.605 -179.355 ;
        RECT 294.275 -181.93 294.605 -180.8 ;
        RECT 294.28 -182.045 294.6 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.635 241.32 295.965 242.45 ;
        RECT 295.635 239.195 295.965 239.525 ;
        RECT 295.635 237.835 295.965 238.165 ;
        RECT 295.64 237.16 295.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.635 -1.525 295.965 -1.195 ;
        RECT 295.635 -2.885 295.965 -2.555 ;
        RECT 295.64 -3.56 295.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 295.635 -95.365 295.965 -95.035 ;
        RECT 295.635 -96.725 295.965 -96.395 ;
        RECT 295.635 -98.085 295.965 -97.755 ;
        RECT 295.635 -99.445 295.965 -99.115 ;
        RECT 295.635 -100.805 295.965 -100.475 ;
        RECT 295.635 -102.165 295.965 -101.835 ;
        RECT 295.635 -103.525 295.965 -103.195 ;
        RECT 295.635 -104.885 295.965 -104.555 ;
        RECT 295.635 -106.245 295.965 -105.915 ;
        RECT 295.635 -107.605 295.965 -107.275 ;
        RECT 295.635 -108.965 295.965 -108.635 ;
        RECT 295.635 -110.325 295.965 -109.995 ;
        RECT 295.635 -111.685 295.965 -111.355 ;
        RECT 295.635 -113.045 295.965 -112.715 ;
        RECT 295.635 -114.405 295.965 -114.075 ;
        RECT 295.635 -115.765 295.965 -115.435 ;
        RECT 295.635 -117.125 295.965 -116.795 ;
        RECT 295.635 -118.485 295.965 -118.155 ;
        RECT 295.635 -119.845 295.965 -119.515 ;
        RECT 295.635 -121.205 295.965 -120.875 ;
        RECT 295.635 -122.565 295.965 -122.235 ;
        RECT 295.635 -123.925 295.965 -123.595 ;
        RECT 295.635 -125.285 295.965 -124.955 ;
        RECT 295.635 -126.645 295.965 -126.315 ;
        RECT 295.635 -128.005 295.965 -127.675 ;
        RECT 295.635 -129.365 295.965 -129.035 ;
        RECT 295.635 -130.725 295.965 -130.395 ;
        RECT 295.635 -132.085 295.965 -131.755 ;
        RECT 295.635 -133.445 295.965 -133.115 ;
        RECT 295.635 -134.805 295.965 -134.475 ;
        RECT 295.635 -136.165 295.965 -135.835 ;
        RECT 295.635 -137.525 295.965 -137.195 ;
        RECT 295.635 -138.885 295.965 -138.555 ;
        RECT 295.635 -140.245 295.965 -139.915 ;
        RECT 295.635 -141.605 295.965 -141.275 ;
        RECT 295.635 -142.965 295.965 -142.635 ;
        RECT 295.635 -144.325 295.965 -143.995 ;
        RECT 295.635 -145.685 295.965 -145.355 ;
        RECT 295.635 -147.045 295.965 -146.715 ;
        RECT 295.635 -148.405 295.965 -148.075 ;
        RECT 295.635 -149.765 295.965 -149.435 ;
        RECT 295.635 -151.125 295.965 -150.795 ;
        RECT 295.635 -152.485 295.965 -152.155 ;
        RECT 295.635 -153.845 295.965 -153.515 ;
        RECT 295.635 -155.205 295.965 -154.875 ;
        RECT 295.635 -156.565 295.965 -156.235 ;
        RECT 295.635 -157.925 295.965 -157.595 ;
        RECT 295.635 -159.285 295.965 -158.955 ;
        RECT 295.635 -160.645 295.965 -160.315 ;
        RECT 295.635 -162.005 295.965 -161.675 ;
        RECT 295.635 -163.365 295.965 -163.035 ;
        RECT 295.635 -164.725 295.965 -164.395 ;
        RECT 295.635 -166.085 295.965 -165.755 ;
        RECT 295.635 -167.445 295.965 -167.115 ;
        RECT 295.635 -168.805 295.965 -168.475 ;
        RECT 295.635 -170.165 295.965 -169.835 ;
        RECT 295.635 -171.525 295.965 -171.195 ;
        RECT 295.635 -172.885 295.965 -172.555 ;
        RECT 295.635 -174.245 295.965 -173.915 ;
        RECT 295.635 -175.605 295.965 -175.275 ;
        RECT 295.635 -176.965 295.965 -176.635 ;
        RECT 295.635 -178.325 295.965 -177.995 ;
        RECT 295.635 -179.685 295.965 -179.355 ;
        RECT 295.635 -181.93 295.965 -180.8 ;
        RECT 295.64 -182.045 295.96 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.995 241.32 297.325 242.45 ;
        RECT 296.995 239.195 297.325 239.525 ;
        RECT 296.995 237.835 297.325 238.165 ;
        RECT 297 237.16 297.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 296.995 -99.445 297.325 -99.115 ;
        RECT 296.995 -100.805 297.325 -100.475 ;
        RECT 296.995 -102.165 297.325 -101.835 ;
        RECT 296.995 -103.525 297.325 -103.195 ;
        RECT 296.995 -104.885 297.325 -104.555 ;
        RECT 296.995 -106.245 297.325 -105.915 ;
        RECT 296.995 -107.605 297.325 -107.275 ;
        RECT 296.995 -108.965 297.325 -108.635 ;
        RECT 296.995 -110.325 297.325 -109.995 ;
        RECT 296.995 -111.685 297.325 -111.355 ;
        RECT 296.995 -113.045 297.325 -112.715 ;
        RECT 296.995 -114.405 297.325 -114.075 ;
        RECT 296.995 -115.765 297.325 -115.435 ;
        RECT 296.995 -117.125 297.325 -116.795 ;
        RECT 296.995 -118.485 297.325 -118.155 ;
        RECT 296.995 -119.845 297.325 -119.515 ;
        RECT 296.995 -121.205 297.325 -120.875 ;
        RECT 296.995 -122.565 297.325 -122.235 ;
        RECT 296.995 -123.925 297.325 -123.595 ;
        RECT 296.995 -125.285 297.325 -124.955 ;
        RECT 296.995 -126.645 297.325 -126.315 ;
        RECT 296.995 -128.005 297.325 -127.675 ;
        RECT 296.995 -129.365 297.325 -129.035 ;
        RECT 296.995 -130.725 297.325 -130.395 ;
        RECT 296.995 -132.085 297.325 -131.755 ;
        RECT 296.995 -133.445 297.325 -133.115 ;
        RECT 296.995 -134.805 297.325 -134.475 ;
        RECT 296.995 -136.165 297.325 -135.835 ;
        RECT 296.995 -137.525 297.325 -137.195 ;
        RECT 296.995 -138.885 297.325 -138.555 ;
        RECT 296.995 -140.245 297.325 -139.915 ;
        RECT 296.995 -141.605 297.325 -141.275 ;
        RECT 296.995 -142.965 297.325 -142.635 ;
        RECT 296.995 -144.325 297.325 -143.995 ;
        RECT 296.995 -145.685 297.325 -145.355 ;
        RECT 296.995 -147.045 297.325 -146.715 ;
        RECT 296.995 -148.405 297.325 -148.075 ;
        RECT 296.995 -149.765 297.325 -149.435 ;
        RECT 296.995 -151.125 297.325 -150.795 ;
        RECT 296.995 -152.485 297.325 -152.155 ;
        RECT 296.995 -153.845 297.325 -153.515 ;
        RECT 296.995 -155.205 297.325 -154.875 ;
        RECT 296.995 -156.565 297.325 -156.235 ;
        RECT 296.995 -157.925 297.325 -157.595 ;
        RECT 296.995 -159.285 297.325 -158.955 ;
        RECT 296.995 -160.645 297.325 -160.315 ;
        RECT 296.995 -162.005 297.325 -161.675 ;
        RECT 296.995 -163.365 297.325 -163.035 ;
        RECT 296.995 -164.725 297.325 -164.395 ;
        RECT 296.995 -166.085 297.325 -165.755 ;
        RECT 296.995 -167.445 297.325 -167.115 ;
        RECT 296.995 -168.805 297.325 -168.475 ;
        RECT 296.995 -170.165 297.325 -169.835 ;
        RECT 296.995 -171.525 297.325 -171.195 ;
        RECT 296.995 -172.885 297.325 -172.555 ;
        RECT 296.995 -174.245 297.325 -173.915 ;
        RECT 296.995 -175.605 297.325 -175.275 ;
        RECT 296.995 -176.965 297.325 -176.635 ;
        RECT 296.995 -178.325 297.325 -177.995 ;
        RECT 296.995 -179.685 297.325 -179.355 ;
        RECT 296.995 -181.93 297.325 -180.8 ;
        RECT 297 -182.045 297.32 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 297.61 -98.075 297.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.355 241.32 298.685 242.45 ;
        RECT 298.355 239.195 298.685 239.525 ;
        RECT 298.355 237.835 298.685 238.165 ;
        RECT 298.36 237.16 298.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 298.355 -1.525 298.685 -1.195 ;
        RECT 298.355 -2.885 298.685 -2.555 ;
        RECT 298.36 -3.56 298.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.715 241.32 300.045 242.45 ;
        RECT 299.715 239.195 300.045 239.525 ;
        RECT 299.715 237.835 300.045 238.165 ;
        RECT 299.72 237.16 300.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 299.715 -1.525 300.045 -1.195 ;
        RECT 299.715 -2.885 300.045 -2.555 ;
        RECT 299.72 -3.56 300.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.075 241.32 301.405 242.45 ;
        RECT 301.075 239.195 301.405 239.525 ;
        RECT 301.075 237.835 301.405 238.165 ;
        RECT 301.08 237.16 301.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.075 -1.525 301.405 -1.195 ;
        RECT 301.075 -2.885 301.405 -2.555 ;
        RECT 301.08 -3.56 301.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 301.075 -95.365 301.405 -95.035 ;
        RECT 301.075 -96.725 301.405 -96.395 ;
        RECT 301.075 -98.085 301.405 -97.755 ;
        RECT 301.075 -99.445 301.405 -99.115 ;
        RECT 301.075 -100.805 301.405 -100.475 ;
        RECT 301.075 -102.165 301.405 -101.835 ;
        RECT 301.075 -103.525 301.405 -103.195 ;
        RECT 301.075 -104.885 301.405 -104.555 ;
        RECT 301.075 -106.245 301.405 -105.915 ;
        RECT 301.075 -107.605 301.405 -107.275 ;
        RECT 301.075 -108.965 301.405 -108.635 ;
        RECT 301.075 -110.325 301.405 -109.995 ;
        RECT 301.075 -111.685 301.405 -111.355 ;
        RECT 301.075 -113.045 301.405 -112.715 ;
        RECT 301.075 -114.405 301.405 -114.075 ;
        RECT 301.075 -115.765 301.405 -115.435 ;
        RECT 301.075 -117.125 301.405 -116.795 ;
        RECT 301.075 -118.485 301.405 -118.155 ;
        RECT 301.075 -119.845 301.405 -119.515 ;
        RECT 301.075 -121.205 301.405 -120.875 ;
        RECT 301.075 -122.565 301.405 -122.235 ;
        RECT 301.075 -123.925 301.405 -123.595 ;
        RECT 301.075 -125.285 301.405 -124.955 ;
        RECT 301.075 -126.645 301.405 -126.315 ;
        RECT 301.075 -128.005 301.405 -127.675 ;
        RECT 301.075 -129.365 301.405 -129.035 ;
        RECT 301.075 -130.725 301.405 -130.395 ;
        RECT 301.075 -132.085 301.405 -131.755 ;
        RECT 301.075 -133.445 301.405 -133.115 ;
        RECT 301.075 -134.805 301.405 -134.475 ;
        RECT 301.075 -136.165 301.405 -135.835 ;
        RECT 301.075 -137.525 301.405 -137.195 ;
        RECT 301.075 -138.885 301.405 -138.555 ;
        RECT 301.075 -140.245 301.405 -139.915 ;
        RECT 301.075 -141.605 301.405 -141.275 ;
        RECT 301.075 -142.965 301.405 -142.635 ;
        RECT 301.075 -144.325 301.405 -143.995 ;
        RECT 301.075 -145.685 301.405 -145.355 ;
        RECT 301.075 -147.045 301.405 -146.715 ;
        RECT 301.075 -148.405 301.405 -148.075 ;
        RECT 301.075 -149.765 301.405 -149.435 ;
        RECT 301.075 -151.125 301.405 -150.795 ;
        RECT 301.075 -152.485 301.405 -152.155 ;
        RECT 301.075 -153.845 301.405 -153.515 ;
        RECT 301.075 -155.205 301.405 -154.875 ;
        RECT 301.075 -156.565 301.405 -156.235 ;
        RECT 301.075 -157.925 301.405 -157.595 ;
        RECT 301.075 -159.285 301.405 -158.955 ;
        RECT 301.075 -160.645 301.405 -160.315 ;
        RECT 301.075 -162.005 301.405 -161.675 ;
        RECT 301.075 -163.365 301.405 -163.035 ;
        RECT 301.075 -164.725 301.405 -164.395 ;
        RECT 301.075 -166.085 301.405 -165.755 ;
        RECT 301.075 -167.445 301.405 -167.115 ;
        RECT 301.075 -168.805 301.405 -168.475 ;
        RECT 301.075 -170.165 301.405 -169.835 ;
        RECT 301.075 -171.525 301.405 -171.195 ;
        RECT 301.075 -172.885 301.405 -172.555 ;
        RECT 301.075 -174.245 301.405 -173.915 ;
        RECT 301.075 -175.605 301.405 -175.275 ;
        RECT 301.075 -176.965 301.405 -176.635 ;
        RECT 301.075 -178.325 301.405 -177.995 ;
        RECT 301.075 -179.685 301.405 -179.355 ;
        RECT 301.075 -181.93 301.405 -180.8 ;
        RECT 301.08 -182.045 301.4 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.435 241.32 302.765 242.45 ;
        RECT 302.435 239.195 302.765 239.525 ;
        RECT 302.435 237.835 302.765 238.165 ;
        RECT 302.44 237.16 302.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.435 -1.525 302.765 -1.195 ;
        RECT 302.435 -2.885 302.765 -2.555 ;
        RECT 302.44 -3.56 302.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 302.435 -95.365 302.765 -95.035 ;
        RECT 302.435 -96.725 302.765 -96.395 ;
        RECT 302.435 -98.085 302.765 -97.755 ;
        RECT 302.435 -99.445 302.765 -99.115 ;
        RECT 302.435 -100.805 302.765 -100.475 ;
        RECT 302.435 -102.165 302.765 -101.835 ;
        RECT 302.435 -103.525 302.765 -103.195 ;
        RECT 302.435 -104.885 302.765 -104.555 ;
        RECT 302.435 -106.245 302.765 -105.915 ;
        RECT 302.435 -107.605 302.765 -107.275 ;
        RECT 302.435 -108.965 302.765 -108.635 ;
        RECT 302.435 -110.325 302.765 -109.995 ;
        RECT 302.435 -111.685 302.765 -111.355 ;
        RECT 302.435 -113.045 302.765 -112.715 ;
        RECT 302.435 -114.405 302.765 -114.075 ;
        RECT 302.435 -115.765 302.765 -115.435 ;
        RECT 302.435 -117.125 302.765 -116.795 ;
        RECT 302.435 -118.485 302.765 -118.155 ;
        RECT 302.435 -119.845 302.765 -119.515 ;
        RECT 302.435 -121.205 302.765 -120.875 ;
        RECT 302.435 -122.565 302.765 -122.235 ;
        RECT 302.435 -123.925 302.765 -123.595 ;
        RECT 302.435 -125.285 302.765 -124.955 ;
        RECT 302.435 -126.645 302.765 -126.315 ;
        RECT 302.435 -128.005 302.765 -127.675 ;
        RECT 302.435 -129.365 302.765 -129.035 ;
        RECT 302.435 -130.725 302.765 -130.395 ;
        RECT 302.435 -132.085 302.765 -131.755 ;
        RECT 302.435 -133.445 302.765 -133.115 ;
        RECT 302.435 -134.805 302.765 -134.475 ;
        RECT 302.435 -136.165 302.765 -135.835 ;
        RECT 302.435 -137.525 302.765 -137.195 ;
        RECT 302.435 -138.885 302.765 -138.555 ;
        RECT 302.435 -140.245 302.765 -139.915 ;
        RECT 302.435 -141.605 302.765 -141.275 ;
        RECT 302.435 -142.965 302.765 -142.635 ;
        RECT 302.435 -144.325 302.765 -143.995 ;
        RECT 302.435 -145.685 302.765 -145.355 ;
        RECT 302.435 -147.045 302.765 -146.715 ;
        RECT 302.435 -148.405 302.765 -148.075 ;
        RECT 302.435 -149.765 302.765 -149.435 ;
        RECT 302.435 -151.125 302.765 -150.795 ;
        RECT 302.435 -152.485 302.765 -152.155 ;
        RECT 302.435 -153.845 302.765 -153.515 ;
        RECT 302.435 -155.205 302.765 -154.875 ;
        RECT 302.435 -156.565 302.765 -156.235 ;
        RECT 302.435 -157.925 302.765 -157.595 ;
        RECT 302.435 -159.285 302.765 -158.955 ;
        RECT 302.435 -160.645 302.765 -160.315 ;
        RECT 302.435 -162.005 302.765 -161.675 ;
        RECT 302.435 -163.365 302.765 -163.035 ;
        RECT 302.435 -164.725 302.765 -164.395 ;
        RECT 302.435 -166.085 302.765 -165.755 ;
        RECT 302.435 -167.445 302.765 -167.115 ;
        RECT 302.435 -168.805 302.765 -168.475 ;
        RECT 302.435 -170.165 302.765 -169.835 ;
        RECT 302.435 -171.525 302.765 -171.195 ;
        RECT 302.435 -172.885 302.765 -172.555 ;
        RECT 302.435 -174.245 302.765 -173.915 ;
        RECT 302.435 -175.605 302.765 -175.275 ;
        RECT 302.435 -176.965 302.765 -176.635 ;
        RECT 302.435 -178.325 302.765 -177.995 ;
        RECT 302.435 -179.685 302.765 -179.355 ;
        RECT 302.435 -181.93 302.765 -180.8 ;
        RECT 302.44 -182.045 302.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.795 241.32 304.125 242.45 ;
        RECT 303.795 239.195 304.125 239.525 ;
        RECT 303.795 237.835 304.125 238.165 ;
        RECT 303.8 237.16 304.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.795 -1.525 304.125 -1.195 ;
        RECT 303.795 -2.885 304.125 -2.555 ;
        RECT 303.8 -3.56 304.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 303.795 -95.365 304.125 -95.035 ;
        RECT 303.795 -96.725 304.125 -96.395 ;
        RECT 303.795 -98.085 304.125 -97.755 ;
        RECT 303.795 -99.445 304.125 -99.115 ;
        RECT 303.795 -100.805 304.125 -100.475 ;
        RECT 303.795 -102.165 304.125 -101.835 ;
        RECT 303.795 -103.525 304.125 -103.195 ;
        RECT 303.795 -104.885 304.125 -104.555 ;
        RECT 303.795 -106.245 304.125 -105.915 ;
        RECT 303.795 -107.605 304.125 -107.275 ;
        RECT 303.795 -108.965 304.125 -108.635 ;
        RECT 303.795 -110.325 304.125 -109.995 ;
        RECT 303.795 -111.685 304.125 -111.355 ;
        RECT 303.795 -113.045 304.125 -112.715 ;
        RECT 303.795 -114.405 304.125 -114.075 ;
        RECT 303.795 -115.765 304.125 -115.435 ;
        RECT 303.795 -117.125 304.125 -116.795 ;
        RECT 303.795 -118.485 304.125 -118.155 ;
        RECT 303.795 -119.845 304.125 -119.515 ;
        RECT 303.795 -121.205 304.125 -120.875 ;
        RECT 303.795 -122.565 304.125 -122.235 ;
        RECT 303.795 -123.925 304.125 -123.595 ;
        RECT 303.795 -125.285 304.125 -124.955 ;
        RECT 303.795 -126.645 304.125 -126.315 ;
        RECT 303.795 -128.005 304.125 -127.675 ;
        RECT 303.795 -129.365 304.125 -129.035 ;
        RECT 303.795 -130.725 304.125 -130.395 ;
        RECT 303.795 -132.085 304.125 -131.755 ;
        RECT 303.795 -133.445 304.125 -133.115 ;
        RECT 303.795 -134.805 304.125 -134.475 ;
        RECT 303.795 -136.165 304.125 -135.835 ;
        RECT 303.795 -137.525 304.125 -137.195 ;
        RECT 303.795 -138.885 304.125 -138.555 ;
        RECT 303.795 -140.245 304.125 -139.915 ;
        RECT 303.795 -141.605 304.125 -141.275 ;
        RECT 303.795 -142.965 304.125 -142.635 ;
        RECT 303.795 -144.325 304.125 -143.995 ;
        RECT 303.795 -145.685 304.125 -145.355 ;
        RECT 303.795 -147.045 304.125 -146.715 ;
        RECT 303.795 -148.405 304.125 -148.075 ;
        RECT 303.795 -149.765 304.125 -149.435 ;
        RECT 303.795 -151.125 304.125 -150.795 ;
        RECT 303.795 -152.485 304.125 -152.155 ;
        RECT 303.795 -153.845 304.125 -153.515 ;
        RECT 303.795 -155.205 304.125 -154.875 ;
        RECT 303.795 -156.565 304.125 -156.235 ;
        RECT 303.795 -157.925 304.125 -157.595 ;
        RECT 303.795 -159.285 304.125 -158.955 ;
        RECT 303.795 -160.645 304.125 -160.315 ;
        RECT 303.795 -162.005 304.125 -161.675 ;
        RECT 303.795 -163.365 304.125 -163.035 ;
        RECT 303.795 -164.725 304.125 -164.395 ;
        RECT 303.795 -166.085 304.125 -165.755 ;
        RECT 303.795 -167.445 304.125 -167.115 ;
        RECT 303.795 -168.805 304.125 -168.475 ;
        RECT 303.795 -170.165 304.125 -169.835 ;
        RECT 303.795 -171.525 304.125 -171.195 ;
        RECT 303.795 -172.885 304.125 -172.555 ;
        RECT 303.795 -174.245 304.125 -173.915 ;
        RECT 303.795 -175.605 304.125 -175.275 ;
        RECT 303.795 -176.965 304.125 -176.635 ;
        RECT 303.795 -178.325 304.125 -177.995 ;
        RECT 303.795 -179.685 304.125 -179.355 ;
        RECT 303.795 -181.93 304.125 -180.8 ;
        RECT 303.8 -182.045 304.12 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.155 241.32 305.485 242.45 ;
        RECT 305.155 239.195 305.485 239.525 ;
        RECT 305.155 237.835 305.485 238.165 ;
        RECT 305.16 237.16 305.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.155 -1.525 305.485 -1.195 ;
        RECT 305.155 -2.885 305.485 -2.555 ;
        RECT 305.16 -3.56 305.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 305.155 -95.365 305.485 -95.035 ;
        RECT 305.155 -96.725 305.485 -96.395 ;
        RECT 305.155 -98.085 305.485 -97.755 ;
        RECT 305.155 -99.445 305.485 -99.115 ;
        RECT 305.155 -100.805 305.485 -100.475 ;
        RECT 305.155 -102.165 305.485 -101.835 ;
        RECT 305.155 -103.525 305.485 -103.195 ;
        RECT 305.155 -104.885 305.485 -104.555 ;
        RECT 305.155 -106.245 305.485 -105.915 ;
        RECT 305.155 -107.605 305.485 -107.275 ;
        RECT 305.155 -108.965 305.485 -108.635 ;
        RECT 305.155 -110.325 305.485 -109.995 ;
        RECT 305.155 -111.685 305.485 -111.355 ;
        RECT 305.155 -113.045 305.485 -112.715 ;
        RECT 305.155 -114.405 305.485 -114.075 ;
        RECT 305.155 -115.765 305.485 -115.435 ;
        RECT 305.155 -117.125 305.485 -116.795 ;
        RECT 305.155 -118.485 305.485 -118.155 ;
        RECT 305.155 -119.845 305.485 -119.515 ;
        RECT 305.155 -121.205 305.485 -120.875 ;
        RECT 305.155 -122.565 305.485 -122.235 ;
        RECT 305.155 -123.925 305.485 -123.595 ;
        RECT 305.155 -125.285 305.485 -124.955 ;
        RECT 305.155 -126.645 305.485 -126.315 ;
        RECT 305.155 -128.005 305.485 -127.675 ;
        RECT 305.155 -129.365 305.485 -129.035 ;
        RECT 305.155 -130.725 305.485 -130.395 ;
        RECT 305.155 -132.085 305.485 -131.755 ;
        RECT 305.155 -133.445 305.485 -133.115 ;
        RECT 305.155 -134.805 305.485 -134.475 ;
        RECT 305.155 -136.165 305.485 -135.835 ;
        RECT 305.155 -137.525 305.485 -137.195 ;
        RECT 305.155 -138.885 305.485 -138.555 ;
        RECT 305.155 -140.245 305.485 -139.915 ;
        RECT 305.155 -141.605 305.485 -141.275 ;
        RECT 305.155 -142.965 305.485 -142.635 ;
        RECT 305.155 -144.325 305.485 -143.995 ;
        RECT 305.155 -145.685 305.485 -145.355 ;
        RECT 305.155 -147.045 305.485 -146.715 ;
        RECT 305.155 -148.405 305.485 -148.075 ;
        RECT 305.155 -149.765 305.485 -149.435 ;
        RECT 305.155 -151.125 305.485 -150.795 ;
        RECT 305.155 -152.485 305.485 -152.155 ;
        RECT 305.155 -153.845 305.485 -153.515 ;
        RECT 305.155 -155.205 305.485 -154.875 ;
        RECT 305.155 -156.565 305.485 -156.235 ;
        RECT 305.155 -157.925 305.485 -157.595 ;
        RECT 305.155 -159.285 305.485 -158.955 ;
        RECT 305.155 -160.645 305.485 -160.315 ;
        RECT 305.155 -162.005 305.485 -161.675 ;
        RECT 305.155 -163.365 305.485 -163.035 ;
        RECT 305.155 -164.725 305.485 -164.395 ;
        RECT 305.155 -166.085 305.485 -165.755 ;
        RECT 305.155 -167.445 305.485 -167.115 ;
        RECT 305.155 -168.805 305.485 -168.475 ;
        RECT 305.155 -170.165 305.485 -169.835 ;
        RECT 305.155 -171.525 305.485 -171.195 ;
        RECT 305.155 -172.885 305.485 -172.555 ;
        RECT 305.155 -174.245 305.485 -173.915 ;
        RECT 305.155 -175.605 305.485 -175.275 ;
        RECT 305.155 -176.965 305.485 -176.635 ;
        RECT 305.155 -178.325 305.485 -177.995 ;
        RECT 305.155 -179.685 305.485 -179.355 ;
        RECT 305.155 -181.93 305.485 -180.8 ;
        RECT 305.16 -182.045 305.48 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.515 241.32 306.845 242.45 ;
        RECT 306.515 239.195 306.845 239.525 ;
        RECT 306.515 237.835 306.845 238.165 ;
        RECT 306.52 237.16 306.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.515 -1.525 306.845 -1.195 ;
        RECT 306.515 -2.885 306.845 -2.555 ;
        RECT 306.52 -3.56 306.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 306.515 -95.365 306.845 -95.035 ;
        RECT 306.515 -96.725 306.845 -96.395 ;
        RECT 306.515 -98.085 306.845 -97.755 ;
        RECT 306.515 -99.445 306.845 -99.115 ;
        RECT 306.515 -100.805 306.845 -100.475 ;
        RECT 306.515 -102.165 306.845 -101.835 ;
        RECT 306.515 -103.525 306.845 -103.195 ;
        RECT 306.515 -104.885 306.845 -104.555 ;
        RECT 306.515 -106.245 306.845 -105.915 ;
        RECT 306.515 -107.605 306.845 -107.275 ;
        RECT 306.515 -108.965 306.845 -108.635 ;
        RECT 306.515 -110.325 306.845 -109.995 ;
        RECT 306.515 -111.685 306.845 -111.355 ;
        RECT 306.515 -113.045 306.845 -112.715 ;
        RECT 306.515 -114.405 306.845 -114.075 ;
        RECT 306.515 -115.765 306.845 -115.435 ;
        RECT 306.515 -117.125 306.845 -116.795 ;
        RECT 306.515 -118.485 306.845 -118.155 ;
        RECT 306.515 -119.845 306.845 -119.515 ;
        RECT 306.515 -121.205 306.845 -120.875 ;
        RECT 306.515 -122.565 306.845 -122.235 ;
        RECT 306.515 -123.925 306.845 -123.595 ;
        RECT 306.515 -125.285 306.845 -124.955 ;
        RECT 306.515 -126.645 306.845 -126.315 ;
        RECT 306.515 -128.005 306.845 -127.675 ;
        RECT 306.515 -129.365 306.845 -129.035 ;
        RECT 306.515 -130.725 306.845 -130.395 ;
        RECT 306.515 -132.085 306.845 -131.755 ;
        RECT 306.515 -133.445 306.845 -133.115 ;
        RECT 306.515 -134.805 306.845 -134.475 ;
        RECT 306.515 -136.165 306.845 -135.835 ;
        RECT 306.515 -137.525 306.845 -137.195 ;
        RECT 306.515 -138.885 306.845 -138.555 ;
        RECT 306.515 -140.245 306.845 -139.915 ;
        RECT 306.515 -141.605 306.845 -141.275 ;
        RECT 306.515 -142.965 306.845 -142.635 ;
        RECT 306.515 -144.325 306.845 -143.995 ;
        RECT 306.515 -145.685 306.845 -145.355 ;
        RECT 306.515 -147.045 306.845 -146.715 ;
        RECT 306.515 -148.405 306.845 -148.075 ;
        RECT 306.515 -149.765 306.845 -149.435 ;
        RECT 306.515 -151.125 306.845 -150.795 ;
        RECT 306.515 -152.485 306.845 -152.155 ;
        RECT 306.515 -153.845 306.845 -153.515 ;
        RECT 306.515 -155.205 306.845 -154.875 ;
        RECT 306.515 -156.565 306.845 -156.235 ;
        RECT 306.515 -157.925 306.845 -157.595 ;
        RECT 306.515 -159.285 306.845 -158.955 ;
        RECT 306.515 -160.645 306.845 -160.315 ;
        RECT 306.515 -162.005 306.845 -161.675 ;
        RECT 306.515 -163.365 306.845 -163.035 ;
        RECT 306.515 -164.725 306.845 -164.395 ;
        RECT 306.515 -166.085 306.845 -165.755 ;
        RECT 306.515 -167.445 306.845 -167.115 ;
        RECT 306.515 -168.805 306.845 -168.475 ;
        RECT 306.515 -170.165 306.845 -169.835 ;
        RECT 306.515 -171.525 306.845 -171.195 ;
        RECT 306.515 -172.885 306.845 -172.555 ;
        RECT 306.515 -174.245 306.845 -173.915 ;
        RECT 306.515 -175.605 306.845 -175.275 ;
        RECT 306.515 -176.965 306.845 -176.635 ;
        RECT 306.515 -178.325 306.845 -177.995 ;
        RECT 306.515 -179.685 306.845 -179.355 ;
        RECT 306.515 -181.93 306.845 -180.8 ;
        RECT 306.52 -182.045 306.84 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.875 241.32 308.205 242.45 ;
        RECT 307.875 239.195 308.205 239.525 ;
        RECT 307.875 237.835 308.205 238.165 ;
        RECT 307.88 237.16 308.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 307.875 -99.445 308.205 -99.115 ;
        RECT 307.875 -100.805 308.205 -100.475 ;
        RECT 307.875 -102.165 308.205 -101.835 ;
        RECT 307.875 -103.525 308.205 -103.195 ;
        RECT 307.875 -104.885 308.205 -104.555 ;
        RECT 307.875 -106.245 308.205 -105.915 ;
        RECT 307.875 -107.605 308.205 -107.275 ;
        RECT 307.875 -108.965 308.205 -108.635 ;
        RECT 307.875 -110.325 308.205 -109.995 ;
        RECT 307.875 -111.685 308.205 -111.355 ;
        RECT 307.875 -113.045 308.205 -112.715 ;
        RECT 307.875 -114.405 308.205 -114.075 ;
        RECT 307.875 -115.765 308.205 -115.435 ;
        RECT 307.875 -117.125 308.205 -116.795 ;
        RECT 307.875 -118.485 308.205 -118.155 ;
        RECT 307.875 -119.845 308.205 -119.515 ;
        RECT 307.875 -121.205 308.205 -120.875 ;
        RECT 307.875 -122.565 308.205 -122.235 ;
        RECT 307.875 -123.925 308.205 -123.595 ;
        RECT 307.875 -125.285 308.205 -124.955 ;
        RECT 307.875 -126.645 308.205 -126.315 ;
        RECT 307.875 -128.005 308.205 -127.675 ;
        RECT 307.875 -129.365 308.205 -129.035 ;
        RECT 307.875 -130.725 308.205 -130.395 ;
        RECT 307.875 -132.085 308.205 -131.755 ;
        RECT 307.875 -133.445 308.205 -133.115 ;
        RECT 307.875 -134.805 308.205 -134.475 ;
        RECT 307.875 -136.165 308.205 -135.835 ;
        RECT 307.875 -137.525 308.205 -137.195 ;
        RECT 307.875 -138.885 308.205 -138.555 ;
        RECT 307.875 -140.245 308.205 -139.915 ;
        RECT 307.875 -141.605 308.205 -141.275 ;
        RECT 307.875 -142.965 308.205 -142.635 ;
        RECT 307.875 -144.325 308.205 -143.995 ;
        RECT 307.875 -145.685 308.205 -145.355 ;
        RECT 307.875 -147.045 308.205 -146.715 ;
        RECT 307.875 -148.405 308.205 -148.075 ;
        RECT 307.875 -149.765 308.205 -149.435 ;
        RECT 307.875 -151.125 308.205 -150.795 ;
        RECT 307.875 -152.485 308.205 -152.155 ;
        RECT 307.875 -153.845 308.205 -153.515 ;
        RECT 307.875 -155.205 308.205 -154.875 ;
        RECT 307.875 -156.565 308.205 -156.235 ;
        RECT 307.875 -157.925 308.205 -157.595 ;
        RECT 307.875 -159.285 308.205 -158.955 ;
        RECT 307.875 -160.645 308.205 -160.315 ;
        RECT 307.875 -162.005 308.205 -161.675 ;
        RECT 307.875 -163.365 308.205 -163.035 ;
        RECT 307.875 -164.725 308.205 -164.395 ;
        RECT 307.875 -166.085 308.205 -165.755 ;
        RECT 307.875 -167.445 308.205 -167.115 ;
        RECT 307.875 -168.805 308.205 -168.475 ;
        RECT 307.875 -170.165 308.205 -169.835 ;
        RECT 307.875 -171.525 308.205 -171.195 ;
        RECT 307.875 -172.885 308.205 -172.555 ;
        RECT 307.875 -174.245 308.205 -173.915 ;
        RECT 307.875 -175.605 308.205 -175.275 ;
        RECT 307.875 -176.965 308.205 -176.635 ;
        RECT 307.875 -178.325 308.205 -177.995 ;
        RECT 307.875 -179.685 308.205 -179.355 ;
        RECT 307.875 -181.93 308.205 -180.8 ;
        RECT 307.88 -182.045 308.2 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 308.51 -98.075 308.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.235 241.32 309.565 242.45 ;
        RECT 309.235 239.195 309.565 239.525 ;
        RECT 309.235 237.835 309.565 238.165 ;
        RECT 309.24 237.16 309.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 309.235 -1.525 309.565 -1.195 ;
        RECT 309.235 -2.885 309.565 -2.555 ;
        RECT 309.24 -3.56 309.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.595 241.32 310.925 242.45 ;
        RECT 310.595 239.195 310.925 239.525 ;
        RECT 310.595 237.835 310.925 238.165 ;
        RECT 310.6 237.16 310.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 310.595 -1.525 310.925 -1.195 ;
        RECT 310.595 -2.885 310.925 -2.555 ;
        RECT 310.6 -3.56 310.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.955 241.32 312.285 242.45 ;
        RECT 311.955 239.195 312.285 239.525 ;
        RECT 311.955 237.835 312.285 238.165 ;
        RECT 311.96 237.16 312.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.955 -1.525 312.285 -1.195 ;
        RECT 311.955 -2.885 312.285 -2.555 ;
        RECT 311.96 -3.56 312.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 311.955 -95.365 312.285 -95.035 ;
        RECT 311.955 -96.725 312.285 -96.395 ;
        RECT 311.955 -98.085 312.285 -97.755 ;
        RECT 311.955 -99.445 312.285 -99.115 ;
        RECT 311.955 -100.805 312.285 -100.475 ;
        RECT 311.955 -102.165 312.285 -101.835 ;
        RECT 311.955 -103.525 312.285 -103.195 ;
        RECT 311.955 -104.885 312.285 -104.555 ;
        RECT 311.955 -106.245 312.285 -105.915 ;
        RECT 311.955 -107.605 312.285 -107.275 ;
        RECT 311.955 -108.965 312.285 -108.635 ;
        RECT 311.955 -110.325 312.285 -109.995 ;
        RECT 311.955 -111.685 312.285 -111.355 ;
        RECT 311.955 -113.045 312.285 -112.715 ;
        RECT 311.955 -114.405 312.285 -114.075 ;
        RECT 311.955 -115.765 312.285 -115.435 ;
        RECT 311.955 -117.125 312.285 -116.795 ;
        RECT 311.955 -118.485 312.285 -118.155 ;
        RECT 311.955 -119.845 312.285 -119.515 ;
        RECT 311.955 -121.205 312.285 -120.875 ;
        RECT 311.955 -122.565 312.285 -122.235 ;
        RECT 311.955 -123.925 312.285 -123.595 ;
        RECT 311.955 -125.285 312.285 -124.955 ;
        RECT 311.955 -126.645 312.285 -126.315 ;
        RECT 311.955 -128.005 312.285 -127.675 ;
        RECT 311.955 -129.365 312.285 -129.035 ;
        RECT 311.955 -130.725 312.285 -130.395 ;
        RECT 311.955 -132.085 312.285 -131.755 ;
        RECT 311.955 -133.445 312.285 -133.115 ;
        RECT 311.955 -134.805 312.285 -134.475 ;
        RECT 311.955 -136.165 312.285 -135.835 ;
        RECT 311.955 -137.525 312.285 -137.195 ;
        RECT 311.955 -138.885 312.285 -138.555 ;
        RECT 311.955 -140.245 312.285 -139.915 ;
        RECT 311.955 -141.605 312.285 -141.275 ;
        RECT 311.955 -142.965 312.285 -142.635 ;
        RECT 311.955 -144.325 312.285 -143.995 ;
        RECT 311.955 -145.685 312.285 -145.355 ;
        RECT 311.955 -147.045 312.285 -146.715 ;
        RECT 311.955 -148.405 312.285 -148.075 ;
        RECT 311.955 -149.765 312.285 -149.435 ;
        RECT 311.955 -151.125 312.285 -150.795 ;
        RECT 311.955 -152.485 312.285 -152.155 ;
        RECT 311.955 -153.845 312.285 -153.515 ;
        RECT 311.955 -155.205 312.285 -154.875 ;
        RECT 311.955 -156.565 312.285 -156.235 ;
        RECT 311.955 -157.925 312.285 -157.595 ;
        RECT 311.955 -159.285 312.285 -158.955 ;
        RECT 311.955 -160.645 312.285 -160.315 ;
        RECT 311.955 -162.005 312.285 -161.675 ;
        RECT 311.955 -163.365 312.285 -163.035 ;
        RECT 311.955 -164.725 312.285 -164.395 ;
        RECT 311.955 -166.085 312.285 -165.755 ;
        RECT 311.955 -167.445 312.285 -167.115 ;
        RECT 311.955 -168.805 312.285 -168.475 ;
        RECT 311.955 -170.165 312.285 -169.835 ;
        RECT 311.955 -171.525 312.285 -171.195 ;
        RECT 311.955 -172.885 312.285 -172.555 ;
        RECT 311.955 -174.245 312.285 -173.915 ;
        RECT 311.955 -175.605 312.285 -175.275 ;
        RECT 311.955 -176.965 312.285 -176.635 ;
        RECT 311.955 -178.325 312.285 -177.995 ;
        RECT 311.955 -179.685 312.285 -179.355 ;
        RECT 311.955 -181.93 312.285 -180.8 ;
        RECT 311.96 -182.045 312.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.315 241.32 313.645 242.45 ;
        RECT 313.315 239.195 313.645 239.525 ;
        RECT 313.315 237.835 313.645 238.165 ;
        RECT 313.32 237.16 313.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.315 -1.525 313.645 -1.195 ;
        RECT 313.315 -2.885 313.645 -2.555 ;
        RECT 313.32 -3.56 313.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 313.315 -95.365 313.645 -95.035 ;
        RECT 313.315 -96.725 313.645 -96.395 ;
        RECT 313.315 -98.085 313.645 -97.755 ;
        RECT 313.315 -99.445 313.645 -99.115 ;
        RECT 313.315 -100.805 313.645 -100.475 ;
        RECT 313.315 -102.165 313.645 -101.835 ;
        RECT 313.315 -103.525 313.645 -103.195 ;
        RECT 313.315 -104.885 313.645 -104.555 ;
        RECT 313.315 -106.245 313.645 -105.915 ;
        RECT 313.315 -107.605 313.645 -107.275 ;
        RECT 313.315 -108.965 313.645 -108.635 ;
        RECT 313.315 -110.325 313.645 -109.995 ;
        RECT 313.315 -111.685 313.645 -111.355 ;
        RECT 313.315 -113.045 313.645 -112.715 ;
        RECT 313.315 -114.405 313.645 -114.075 ;
        RECT 313.315 -115.765 313.645 -115.435 ;
        RECT 313.315 -117.125 313.645 -116.795 ;
        RECT 313.315 -118.485 313.645 -118.155 ;
        RECT 313.315 -119.845 313.645 -119.515 ;
        RECT 313.315 -121.205 313.645 -120.875 ;
        RECT 313.315 -122.565 313.645 -122.235 ;
        RECT 313.315 -123.925 313.645 -123.595 ;
        RECT 313.315 -125.285 313.645 -124.955 ;
        RECT 313.315 -126.645 313.645 -126.315 ;
        RECT 313.315 -128.005 313.645 -127.675 ;
        RECT 313.315 -129.365 313.645 -129.035 ;
        RECT 313.315 -130.725 313.645 -130.395 ;
        RECT 313.315 -132.085 313.645 -131.755 ;
        RECT 313.315 -133.445 313.645 -133.115 ;
        RECT 313.315 -134.805 313.645 -134.475 ;
        RECT 313.315 -136.165 313.645 -135.835 ;
        RECT 313.315 -137.525 313.645 -137.195 ;
        RECT 313.315 -138.885 313.645 -138.555 ;
        RECT 313.315 -140.245 313.645 -139.915 ;
        RECT 313.315 -141.605 313.645 -141.275 ;
        RECT 313.315 -142.965 313.645 -142.635 ;
        RECT 313.315 -144.325 313.645 -143.995 ;
        RECT 313.315 -145.685 313.645 -145.355 ;
        RECT 313.315 -147.045 313.645 -146.715 ;
        RECT 313.315 -148.405 313.645 -148.075 ;
        RECT 313.315 -149.765 313.645 -149.435 ;
        RECT 313.315 -151.125 313.645 -150.795 ;
        RECT 313.315 -152.485 313.645 -152.155 ;
        RECT 313.315 -153.845 313.645 -153.515 ;
        RECT 313.315 -155.205 313.645 -154.875 ;
        RECT 313.315 -156.565 313.645 -156.235 ;
        RECT 313.315 -157.925 313.645 -157.595 ;
        RECT 313.315 -159.285 313.645 -158.955 ;
        RECT 313.315 -160.645 313.645 -160.315 ;
        RECT 313.315 -162.005 313.645 -161.675 ;
        RECT 313.315 -163.365 313.645 -163.035 ;
        RECT 313.315 -164.725 313.645 -164.395 ;
        RECT 313.315 -166.085 313.645 -165.755 ;
        RECT 313.315 -167.445 313.645 -167.115 ;
        RECT 313.315 -168.805 313.645 -168.475 ;
        RECT 313.315 -170.165 313.645 -169.835 ;
        RECT 313.315 -171.525 313.645 -171.195 ;
        RECT 313.315 -172.885 313.645 -172.555 ;
        RECT 313.315 -174.245 313.645 -173.915 ;
        RECT 313.315 -175.605 313.645 -175.275 ;
        RECT 313.315 -176.965 313.645 -176.635 ;
        RECT 313.315 -178.325 313.645 -177.995 ;
        RECT 313.315 -179.685 313.645 -179.355 ;
        RECT 313.315 -181.93 313.645 -180.8 ;
        RECT 313.32 -182.045 313.64 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.675 241.32 315.005 242.45 ;
        RECT 314.675 239.195 315.005 239.525 ;
        RECT 314.675 237.835 315.005 238.165 ;
        RECT 314.68 237.16 315 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.675 -1.525 315.005 -1.195 ;
        RECT 314.675 -2.885 315.005 -2.555 ;
        RECT 314.68 -3.56 315 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 314.675 -163.365 315.005 -163.035 ;
        RECT 314.675 -164.725 315.005 -164.395 ;
        RECT 314.675 -166.085 315.005 -165.755 ;
        RECT 314.675 -167.445 315.005 -167.115 ;
        RECT 314.675 -168.805 315.005 -168.475 ;
        RECT 314.675 -170.165 315.005 -169.835 ;
        RECT 314.675 -171.525 315.005 -171.195 ;
        RECT 314.675 -172.885 315.005 -172.555 ;
        RECT 314.675 -174.245 315.005 -173.915 ;
        RECT 314.675 -175.605 315.005 -175.275 ;
        RECT 314.675 -176.965 315.005 -176.635 ;
        RECT 314.675 -178.325 315.005 -177.995 ;
        RECT 314.675 -179.685 315.005 -179.355 ;
        RECT 314.675 -181.93 315.005 -180.8 ;
        RECT 314.68 -182.045 315 -95.035 ;
        RECT 314.675 -95.365 315.005 -95.035 ;
        RECT 314.675 -96.725 315.005 -96.395 ;
        RECT 314.675 -98.085 315.005 -97.755 ;
        RECT 314.675 -99.445 315.005 -99.115 ;
        RECT 314.675 -100.805 315.005 -100.475 ;
        RECT 314.675 -102.165 315.005 -101.835 ;
        RECT 314.675 -103.525 315.005 -103.195 ;
        RECT 314.675 -104.885 315.005 -104.555 ;
        RECT 314.675 -106.245 315.005 -105.915 ;
        RECT 314.675 -107.605 315.005 -107.275 ;
        RECT 314.675 -108.965 315.005 -108.635 ;
        RECT 314.675 -110.325 315.005 -109.995 ;
        RECT 314.675 -111.685 315.005 -111.355 ;
        RECT 314.675 -113.045 315.005 -112.715 ;
        RECT 314.675 -114.405 315.005 -114.075 ;
        RECT 314.675 -115.765 315.005 -115.435 ;
        RECT 314.675 -117.125 315.005 -116.795 ;
        RECT 314.675 -118.485 315.005 -118.155 ;
        RECT 314.675 -119.845 315.005 -119.515 ;
        RECT 314.675 -121.205 315.005 -120.875 ;
        RECT 314.675 -122.565 315.005 -122.235 ;
        RECT 314.675 -123.925 315.005 -123.595 ;
        RECT 314.675 -125.285 315.005 -124.955 ;
        RECT 314.675 -126.645 315.005 -126.315 ;
        RECT 314.675 -128.005 315.005 -127.675 ;
        RECT 314.675 -129.365 315.005 -129.035 ;
        RECT 314.675 -130.725 315.005 -130.395 ;
        RECT 314.675 -132.085 315.005 -131.755 ;
        RECT 314.675 -133.445 315.005 -133.115 ;
        RECT 314.675 -134.805 315.005 -134.475 ;
        RECT 314.675 -136.165 315.005 -135.835 ;
        RECT 314.675 -137.525 315.005 -137.195 ;
        RECT 314.675 -138.885 315.005 -138.555 ;
        RECT 314.675 -140.245 315.005 -139.915 ;
        RECT 314.675 -141.605 315.005 -141.275 ;
        RECT 314.675 -142.965 315.005 -142.635 ;
        RECT 314.675 -144.325 315.005 -143.995 ;
        RECT 314.675 -145.685 315.005 -145.355 ;
        RECT 314.675 -147.045 315.005 -146.715 ;
        RECT 314.675 -148.405 315.005 -148.075 ;
        RECT 314.675 -149.765 315.005 -149.435 ;
        RECT 314.675 -151.125 315.005 -150.795 ;
        RECT 314.675 -152.485 315.005 -152.155 ;
        RECT 314.675 -153.845 315.005 -153.515 ;
        RECT 314.675 -155.205 315.005 -154.875 ;
        RECT 314.675 -156.565 315.005 -156.235 ;
        RECT 314.675 -157.925 315.005 -157.595 ;
        RECT 314.675 -159.285 315.005 -158.955 ;
        RECT 314.675 -160.645 315.005 -160.315 ;
        RECT 314.675 -162.005 315.005 -161.675 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.91 -98.075 265.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.715 241.32 266.045 242.45 ;
        RECT 265.715 239.195 266.045 239.525 ;
        RECT 265.715 237.835 266.045 238.165 ;
        RECT 265.72 237.16 266.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 265.715 -1.525 266.045 -1.195 ;
        RECT 265.715 -2.885 266.045 -2.555 ;
        RECT 265.72 -3.56 266.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.075 241.32 267.405 242.45 ;
        RECT 267.075 239.195 267.405 239.525 ;
        RECT 267.075 237.835 267.405 238.165 ;
        RECT 267.08 237.16 267.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 267.075 -1.525 267.405 -1.195 ;
        RECT 267.075 -2.885 267.405 -2.555 ;
        RECT 267.08 -3.56 267.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.435 241.32 268.765 242.45 ;
        RECT 268.435 239.195 268.765 239.525 ;
        RECT 268.435 237.835 268.765 238.165 ;
        RECT 268.44 237.16 268.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.435 -1.525 268.765 -1.195 ;
        RECT 268.435 -2.885 268.765 -2.555 ;
        RECT 268.44 -3.56 268.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 268.435 -95.365 268.765 -95.035 ;
        RECT 268.435 -96.725 268.765 -96.395 ;
        RECT 268.435 -98.085 268.765 -97.755 ;
        RECT 268.435 -99.445 268.765 -99.115 ;
        RECT 268.435 -100.805 268.765 -100.475 ;
        RECT 268.435 -102.165 268.765 -101.835 ;
        RECT 268.435 -103.525 268.765 -103.195 ;
        RECT 268.435 -104.885 268.765 -104.555 ;
        RECT 268.435 -106.245 268.765 -105.915 ;
        RECT 268.435 -107.605 268.765 -107.275 ;
        RECT 268.435 -108.965 268.765 -108.635 ;
        RECT 268.435 -110.325 268.765 -109.995 ;
        RECT 268.435 -111.685 268.765 -111.355 ;
        RECT 268.435 -113.045 268.765 -112.715 ;
        RECT 268.435 -114.405 268.765 -114.075 ;
        RECT 268.435 -115.765 268.765 -115.435 ;
        RECT 268.435 -117.125 268.765 -116.795 ;
        RECT 268.435 -118.485 268.765 -118.155 ;
        RECT 268.435 -119.845 268.765 -119.515 ;
        RECT 268.435 -121.205 268.765 -120.875 ;
        RECT 268.435 -122.565 268.765 -122.235 ;
        RECT 268.435 -123.925 268.765 -123.595 ;
        RECT 268.435 -125.285 268.765 -124.955 ;
        RECT 268.435 -126.645 268.765 -126.315 ;
        RECT 268.435 -128.005 268.765 -127.675 ;
        RECT 268.435 -129.365 268.765 -129.035 ;
        RECT 268.435 -130.725 268.765 -130.395 ;
        RECT 268.435 -132.085 268.765 -131.755 ;
        RECT 268.435 -133.445 268.765 -133.115 ;
        RECT 268.435 -134.805 268.765 -134.475 ;
        RECT 268.435 -136.165 268.765 -135.835 ;
        RECT 268.435 -137.525 268.765 -137.195 ;
        RECT 268.435 -138.885 268.765 -138.555 ;
        RECT 268.435 -140.245 268.765 -139.915 ;
        RECT 268.435 -141.605 268.765 -141.275 ;
        RECT 268.435 -142.965 268.765 -142.635 ;
        RECT 268.435 -144.325 268.765 -143.995 ;
        RECT 268.435 -145.685 268.765 -145.355 ;
        RECT 268.435 -147.045 268.765 -146.715 ;
        RECT 268.435 -148.405 268.765 -148.075 ;
        RECT 268.435 -149.765 268.765 -149.435 ;
        RECT 268.435 -151.125 268.765 -150.795 ;
        RECT 268.435 -152.485 268.765 -152.155 ;
        RECT 268.435 -153.845 268.765 -153.515 ;
        RECT 268.435 -155.205 268.765 -154.875 ;
        RECT 268.435 -156.565 268.765 -156.235 ;
        RECT 268.435 -157.925 268.765 -157.595 ;
        RECT 268.435 -159.285 268.765 -158.955 ;
        RECT 268.435 -160.645 268.765 -160.315 ;
        RECT 268.435 -162.005 268.765 -161.675 ;
        RECT 268.435 -163.365 268.765 -163.035 ;
        RECT 268.435 -164.725 268.765 -164.395 ;
        RECT 268.435 -166.085 268.765 -165.755 ;
        RECT 268.435 -167.445 268.765 -167.115 ;
        RECT 268.435 -168.805 268.765 -168.475 ;
        RECT 268.435 -170.165 268.765 -169.835 ;
        RECT 268.435 -171.525 268.765 -171.195 ;
        RECT 268.435 -172.885 268.765 -172.555 ;
        RECT 268.435 -174.245 268.765 -173.915 ;
        RECT 268.435 -175.605 268.765 -175.275 ;
        RECT 268.435 -176.965 268.765 -176.635 ;
        RECT 268.435 -178.325 268.765 -177.995 ;
        RECT 268.435 -179.685 268.765 -179.355 ;
        RECT 268.435 -181.93 268.765 -180.8 ;
        RECT 268.44 -182.045 268.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.795 241.32 270.125 242.45 ;
        RECT 269.795 239.195 270.125 239.525 ;
        RECT 269.795 237.835 270.125 238.165 ;
        RECT 269.8 237.16 270.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.795 -1.525 270.125 -1.195 ;
        RECT 269.795 -2.885 270.125 -2.555 ;
        RECT 269.8 -3.56 270.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 269.795 -95.365 270.125 -95.035 ;
        RECT 269.795 -96.725 270.125 -96.395 ;
        RECT 269.795 -98.085 270.125 -97.755 ;
        RECT 269.795 -99.445 270.125 -99.115 ;
        RECT 269.795 -100.805 270.125 -100.475 ;
        RECT 269.795 -102.165 270.125 -101.835 ;
        RECT 269.795 -103.525 270.125 -103.195 ;
        RECT 269.795 -104.885 270.125 -104.555 ;
        RECT 269.795 -106.245 270.125 -105.915 ;
        RECT 269.795 -107.605 270.125 -107.275 ;
        RECT 269.795 -108.965 270.125 -108.635 ;
        RECT 269.795 -110.325 270.125 -109.995 ;
        RECT 269.795 -111.685 270.125 -111.355 ;
        RECT 269.795 -113.045 270.125 -112.715 ;
        RECT 269.795 -114.405 270.125 -114.075 ;
        RECT 269.795 -115.765 270.125 -115.435 ;
        RECT 269.795 -117.125 270.125 -116.795 ;
        RECT 269.795 -118.485 270.125 -118.155 ;
        RECT 269.795 -119.845 270.125 -119.515 ;
        RECT 269.795 -121.205 270.125 -120.875 ;
        RECT 269.795 -122.565 270.125 -122.235 ;
        RECT 269.795 -123.925 270.125 -123.595 ;
        RECT 269.795 -125.285 270.125 -124.955 ;
        RECT 269.795 -126.645 270.125 -126.315 ;
        RECT 269.795 -128.005 270.125 -127.675 ;
        RECT 269.795 -129.365 270.125 -129.035 ;
        RECT 269.795 -130.725 270.125 -130.395 ;
        RECT 269.795 -132.085 270.125 -131.755 ;
        RECT 269.795 -133.445 270.125 -133.115 ;
        RECT 269.795 -134.805 270.125 -134.475 ;
        RECT 269.795 -136.165 270.125 -135.835 ;
        RECT 269.795 -137.525 270.125 -137.195 ;
        RECT 269.795 -138.885 270.125 -138.555 ;
        RECT 269.795 -140.245 270.125 -139.915 ;
        RECT 269.795 -141.605 270.125 -141.275 ;
        RECT 269.795 -142.965 270.125 -142.635 ;
        RECT 269.795 -144.325 270.125 -143.995 ;
        RECT 269.795 -145.685 270.125 -145.355 ;
        RECT 269.795 -147.045 270.125 -146.715 ;
        RECT 269.795 -148.405 270.125 -148.075 ;
        RECT 269.795 -149.765 270.125 -149.435 ;
        RECT 269.795 -151.125 270.125 -150.795 ;
        RECT 269.795 -152.485 270.125 -152.155 ;
        RECT 269.795 -153.845 270.125 -153.515 ;
        RECT 269.795 -155.205 270.125 -154.875 ;
        RECT 269.795 -156.565 270.125 -156.235 ;
        RECT 269.795 -157.925 270.125 -157.595 ;
        RECT 269.795 -159.285 270.125 -158.955 ;
        RECT 269.795 -160.645 270.125 -160.315 ;
        RECT 269.795 -162.005 270.125 -161.675 ;
        RECT 269.795 -163.365 270.125 -163.035 ;
        RECT 269.795 -164.725 270.125 -164.395 ;
        RECT 269.795 -166.085 270.125 -165.755 ;
        RECT 269.795 -167.445 270.125 -167.115 ;
        RECT 269.795 -168.805 270.125 -168.475 ;
        RECT 269.795 -170.165 270.125 -169.835 ;
        RECT 269.795 -171.525 270.125 -171.195 ;
        RECT 269.795 -172.885 270.125 -172.555 ;
        RECT 269.795 -174.245 270.125 -173.915 ;
        RECT 269.795 -175.605 270.125 -175.275 ;
        RECT 269.795 -176.965 270.125 -176.635 ;
        RECT 269.795 -178.325 270.125 -177.995 ;
        RECT 269.795 -179.685 270.125 -179.355 ;
        RECT 269.795 -181.93 270.125 -180.8 ;
        RECT 269.8 -182.045 270.12 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.155 241.32 271.485 242.45 ;
        RECT 271.155 239.195 271.485 239.525 ;
        RECT 271.155 237.835 271.485 238.165 ;
        RECT 271.16 237.16 271.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.155 -1.525 271.485 -1.195 ;
        RECT 271.155 -2.885 271.485 -2.555 ;
        RECT 271.16 -3.56 271.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 271.155 -95.365 271.485 -95.035 ;
        RECT 271.155 -96.725 271.485 -96.395 ;
        RECT 271.155 -98.085 271.485 -97.755 ;
        RECT 271.155 -99.445 271.485 -99.115 ;
        RECT 271.155 -100.805 271.485 -100.475 ;
        RECT 271.155 -102.165 271.485 -101.835 ;
        RECT 271.155 -103.525 271.485 -103.195 ;
        RECT 271.155 -104.885 271.485 -104.555 ;
        RECT 271.155 -106.245 271.485 -105.915 ;
        RECT 271.155 -107.605 271.485 -107.275 ;
        RECT 271.155 -108.965 271.485 -108.635 ;
        RECT 271.155 -110.325 271.485 -109.995 ;
        RECT 271.155 -111.685 271.485 -111.355 ;
        RECT 271.155 -113.045 271.485 -112.715 ;
        RECT 271.155 -114.405 271.485 -114.075 ;
        RECT 271.155 -115.765 271.485 -115.435 ;
        RECT 271.155 -117.125 271.485 -116.795 ;
        RECT 271.155 -118.485 271.485 -118.155 ;
        RECT 271.155 -119.845 271.485 -119.515 ;
        RECT 271.155 -121.205 271.485 -120.875 ;
        RECT 271.155 -122.565 271.485 -122.235 ;
        RECT 271.155 -123.925 271.485 -123.595 ;
        RECT 271.155 -125.285 271.485 -124.955 ;
        RECT 271.155 -126.645 271.485 -126.315 ;
        RECT 271.155 -128.005 271.485 -127.675 ;
        RECT 271.155 -129.365 271.485 -129.035 ;
        RECT 271.155 -130.725 271.485 -130.395 ;
        RECT 271.155 -132.085 271.485 -131.755 ;
        RECT 271.155 -133.445 271.485 -133.115 ;
        RECT 271.155 -134.805 271.485 -134.475 ;
        RECT 271.155 -136.165 271.485 -135.835 ;
        RECT 271.155 -137.525 271.485 -137.195 ;
        RECT 271.155 -138.885 271.485 -138.555 ;
        RECT 271.155 -140.245 271.485 -139.915 ;
        RECT 271.155 -141.605 271.485 -141.275 ;
        RECT 271.155 -142.965 271.485 -142.635 ;
        RECT 271.155 -144.325 271.485 -143.995 ;
        RECT 271.155 -145.685 271.485 -145.355 ;
        RECT 271.155 -147.045 271.485 -146.715 ;
        RECT 271.155 -148.405 271.485 -148.075 ;
        RECT 271.155 -149.765 271.485 -149.435 ;
        RECT 271.155 -151.125 271.485 -150.795 ;
        RECT 271.155 -152.485 271.485 -152.155 ;
        RECT 271.155 -153.845 271.485 -153.515 ;
        RECT 271.155 -155.205 271.485 -154.875 ;
        RECT 271.155 -156.565 271.485 -156.235 ;
        RECT 271.155 -157.925 271.485 -157.595 ;
        RECT 271.155 -159.285 271.485 -158.955 ;
        RECT 271.155 -160.645 271.485 -160.315 ;
        RECT 271.155 -162.005 271.485 -161.675 ;
        RECT 271.155 -163.365 271.485 -163.035 ;
        RECT 271.155 -164.725 271.485 -164.395 ;
        RECT 271.155 -166.085 271.485 -165.755 ;
        RECT 271.155 -167.445 271.485 -167.115 ;
        RECT 271.155 -168.805 271.485 -168.475 ;
        RECT 271.155 -170.165 271.485 -169.835 ;
        RECT 271.155 -171.525 271.485 -171.195 ;
        RECT 271.155 -172.885 271.485 -172.555 ;
        RECT 271.155 -174.245 271.485 -173.915 ;
        RECT 271.155 -175.605 271.485 -175.275 ;
        RECT 271.155 -176.965 271.485 -176.635 ;
        RECT 271.155 -178.325 271.485 -177.995 ;
        RECT 271.155 -179.685 271.485 -179.355 ;
        RECT 271.155 -181.93 271.485 -180.8 ;
        RECT 271.16 -182.045 271.48 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.515 241.32 272.845 242.45 ;
        RECT 272.515 239.195 272.845 239.525 ;
        RECT 272.515 237.835 272.845 238.165 ;
        RECT 272.52 237.16 272.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.515 -1.525 272.845 -1.195 ;
        RECT 272.515 -2.885 272.845 -2.555 ;
        RECT 272.52 -3.56 272.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 272.515 -95.365 272.845 -95.035 ;
        RECT 272.515 -96.725 272.845 -96.395 ;
        RECT 272.515 -98.085 272.845 -97.755 ;
        RECT 272.515 -99.445 272.845 -99.115 ;
        RECT 272.515 -100.805 272.845 -100.475 ;
        RECT 272.515 -102.165 272.845 -101.835 ;
        RECT 272.515 -103.525 272.845 -103.195 ;
        RECT 272.515 -104.885 272.845 -104.555 ;
        RECT 272.515 -106.245 272.845 -105.915 ;
        RECT 272.515 -107.605 272.845 -107.275 ;
        RECT 272.515 -108.965 272.845 -108.635 ;
        RECT 272.515 -110.325 272.845 -109.995 ;
        RECT 272.515 -111.685 272.845 -111.355 ;
        RECT 272.515 -113.045 272.845 -112.715 ;
        RECT 272.515 -114.405 272.845 -114.075 ;
        RECT 272.515 -115.765 272.845 -115.435 ;
        RECT 272.515 -117.125 272.845 -116.795 ;
        RECT 272.515 -118.485 272.845 -118.155 ;
        RECT 272.515 -119.845 272.845 -119.515 ;
        RECT 272.515 -121.205 272.845 -120.875 ;
        RECT 272.515 -122.565 272.845 -122.235 ;
        RECT 272.515 -123.925 272.845 -123.595 ;
        RECT 272.515 -125.285 272.845 -124.955 ;
        RECT 272.515 -126.645 272.845 -126.315 ;
        RECT 272.515 -128.005 272.845 -127.675 ;
        RECT 272.515 -129.365 272.845 -129.035 ;
        RECT 272.515 -130.725 272.845 -130.395 ;
        RECT 272.515 -132.085 272.845 -131.755 ;
        RECT 272.515 -133.445 272.845 -133.115 ;
        RECT 272.515 -134.805 272.845 -134.475 ;
        RECT 272.515 -136.165 272.845 -135.835 ;
        RECT 272.515 -137.525 272.845 -137.195 ;
        RECT 272.515 -138.885 272.845 -138.555 ;
        RECT 272.515 -140.245 272.845 -139.915 ;
        RECT 272.515 -141.605 272.845 -141.275 ;
        RECT 272.515 -142.965 272.845 -142.635 ;
        RECT 272.515 -144.325 272.845 -143.995 ;
        RECT 272.515 -145.685 272.845 -145.355 ;
        RECT 272.515 -147.045 272.845 -146.715 ;
        RECT 272.515 -148.405 272.845 -148.075 ;
        RECT 272.515 -149.765 272.845 -149.435 ;
        RECT 272.515 -151.125 272.845 -150.795 ;
        RECT 272.515 -152.485 272.845 -152.155 ;
        RECT 272.515 -153.845 272.845 -153.515 ;
        RECT 272.515 -155.205 272.845 -154.875 ;
        RECT 272.515 -156.565 272.845 -156.235 ;
        RECT 272.515 -157.925 272.845 -157.595 ;
        RECT 272.515 -159.285 272.845 -158.955 ;
        RECT 272.515 -160.645 272.845 -160.315 ;
        RECT 272.515 -162.005 272.845 -161.675 ;
        RECT 272.515 -163.365 272.845 -163.035 ;
        RECT 272.515 -164.725 272.845 -164.395 ;
        RECT 272.515 -166.085 272.845 -165.755 ;
        RECT 272.515 -167.445 272.845 -167.115 ;
        RECT 272.515 -168.805 272.845 -168.475 ;
        RECT 272.515 -170.165 272.845 -169.835 ;
        RECT 272.515 -171.525 272.845 -171.195 ;
        RECT 272.515 -172.885 272.845 -172.555 ;
        RECT 272.515 -174.245 272.845 -173.915 ;
        RECT 272.515 -175.605 272.845 -175.275 ;
        RECT 272.515 -176.965 272.845 -176.635 ;
        RECT 272.515 -178.325 272.845 -177.995 ;
        RECT 272.515 -179.685 272.845 -179.355 ;
        RECT 272.515 -181.93 272.845 -180.8 ;
        RECT 272.52 -182.045 272.84 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.875 241.32 274.205 242.45 ;
        RECT 273.875 239.195 274.205 239.525 ;
        RECT 273.875 237.835 274.205 238.165 ;
        RECT 273.88 237.16 274.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.875 -1.525 274.205 -1.195 ;
        RECT 273.875 -2.885 274.205 -2.555 ;
        RECT 273.88 -3.56 274.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 273.875 -95.365 274.205 -95.035 ;
        RECT 273.875 -96.725 274.205 -96.395 ;
        RECT 273.875 -98.085 274.205 -97.755 ;
        RECT 273.875 -99.445 274.205 -99.115 ;
        RECT 273.875 -100.805 274.205 -100.475 ;
        RECT 273.875 -102.165 274.205 -101.835 ;
        RECT 273.875 -103.525 274.205 -103.195 ;
        RECT 273.875 -104.885 274.205 -104.555 ;
        RECT 273.875 -106.245 274.205 -105.915 ;
        RECT 273.875 -107.605 274.205 -107.275 ;
        RECT 273.875 -108.965 274.205 -108.635 ;
        RECT 273.875 -110.325 274.205 -109.995 ;
        RECT 273.875 -111.685 274.205 -111.355 ;
        RECT 273.875 -113.045 274.205 -112.715 ;
        RECT 273.875 -114.405 274.205 -114.075 ;
        RECT 273.875 -115.765 274.205 -115.435 ;
        RECT 273.875 -117.125 274.205 -116.795 ;
        RECT 273.875 -118.485 274.205 -118.155 ;
        RECT 273.875 -119.845 274.205 -119.515 ;
        RECT 273.875 -121.205 274.205 -120.875 ;
        RECT 273.875 -122.565 274.205 -122.235 ;
        RECT 273.875 -123.925 274.205 -123.595 ;
        RECT 273.875 -125.285 274.205 -124.955 ;
        RECT 273.875 -126.645 274.205 -126.315 ;
        RECT 273.875 -128.005 274.205 -127.675 ;
        RECT 273.875 -129.365 274.205 -129.035 ;
        RECT 273.875 -130.725 274.205 -130.395 ;
        RECT 273.875 -132.085 274.205 -131.755 ;
        RECT 273.875 -133.445 274.205 -133.115 ;
        RECT 273.875 -134.805 274.205 -134.475 ;
        RECT 273.875 -136.165 274.205 -135.835 ;
        RECT 273.875 -137.525 274.205 -137.195 ;
        RECT 273.875 -138.885 274.205 -138.555 ;
        RECT 273.875 -140.245 274.205 -139.915 ;
        RECT 273.875 -141.605 274.205 -141.275 ;
        RECT 273.875 -142.965 274.205 -142.635 ;
        RECT 273.875 -144.325 274.205 -143.995 ;
        RECT 273.875 -145.685 274.205 -145.355 ;
        RECT 273.875 -147.045 274.205 -146.715 ;
        RECT 273.875 -148.405 274.205 -148.075 ;
        RECT 273.875 -149.765 274.205 -149.435 ;
        RECT 273.875 -151.125 274.205 -150.795 ;
        RECT 273.875 -152.485 274.205 -152.155 ;
        RECT 273.875 -153.845 274.205 -153.515 ;
        RECT 273.875 -155.205 274.205 -154.875 ;
        RECT 273.875 -156.565 274.205 -156.235 ;
        RECT 273.875 -157.925 274.205 -157.595 ;
        RECT 273.875 -159.285 274.205 -158.955 ;
        RECT 273.875 -160.645 274.205 -160.315 ;
        RECT 273.875 -162.005 274.205 -161.675 ;
        RECT 273.875 -163.365 274.205 -163.035 ;
        RECT 273.875 -164.725 274.205 -164.395 ;
        RECT 273.875 -166.085 274.205 -165.755 ;
        RECT 273.875 -167.445 274.205 -167.115 ;
        RECT 273.875 -168.805 274.205 -168.475 ;
        RECT 273.875 -170.165 274.205 -169.835 ;
        RECT 273.875 -171.525 274.205 -171.195 ;
        RECT 273.875 -172.885 274.205 -172.555 ;
        RECT 273.875 -174.245 274.205 -173.915 ;
        RECT 273.875 -175.605 274.205 -175.275 ;
        RECT 273.875 -176.965 274.205 -176.635 ;
        RECT 273.875 -178.325 274.205 -177.995 ;
        RECT 273.875 -179.685 274.205 -179.355 ;
        RECT 273.875 -181.93 274.205 -180.8 ;
        RECT 273.88 -182.045 274.2 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.235 241.32 275.565 242.45 ;
        RECT 275.235 239.195 275.565 239.525 ;
        RECT 275.235 237.835 275.565 238.165 ;
        RECT 275.24 237.16 275.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.235 -99.445 275.565 -99.115 ;
        RECT 275.235 -100.805 275.565 -100.475 ;
        RECT 275.235 -102.165 275.565 -101.835 ;
        RECT 275.235 -103.525 275.565 -103.195 ;
        RECT 275.235 -104.885 275.565 -104.555 ;
        RECT 275.235 -106.245 275.565 -105.915 ;
        RECT 275.235 -107.605 275.565 -107.275 ;
        RECT 275.235 -108.965 275.565 -108.635 ;
        RECT 275.235 -110.325 275.565 -109.995 ;
        RECT 275.235 -111.685 275.565 -111.355 ;
        RECT 275.235 -113.045 275.565 -112.715 ;
        RECT 275.235 -114.405 275.565 -114.075 ;
        RECT 275.235 -115.765 275.565 -115.435 ;
        RECT 275.235 -117.125 275.565 -116.795 ;
        RECT 275.235 -118.485 275.565 -118.155 ;
        RECT 275.235 -119.845 275.565 -119.515 ;
        RECT 275.235 -121.205 275.565 -120.875 ;
        RECT 275.235 -122.565 275.565 -122.235 ;
        RECT 275.235 -123.925 275.565 -123.595 ;
        RECT 275.235 -125.285 275.565 -124.955 ;
        RECT 275.235 -126.645 275.565 -126.315 ;
        RECT 275.235 -128.005 275.565 -127.675 ;
        RECT 275.235 -129.365 275.565 -129.035 ;
        RECT 275.235 -130.725 275.565 -130.395 ;
        RECT 275.235 -132.085 275.565 -131.755 ;
        RECT 275.235 -133.445 275.565 -133.115 ;
        RECT 275.235 -134.805 275.565 -134.475 ;
        RECT 275.235 -136.165 275.565 -135.835 ;
        RECT 275.235 -137.525 275.565 -137.195 ;
        RECT 275.235 -138.885 275.565 -138.555 ;
        RECT 275.235 -140.245 275.565 -139.915 ;
        RECT 275.235 -141.605 275.565 -141.275 ;
        RECT 275.235 -142.965 275.565 -142.635 ;
        RECT 275.235 -144.325 275.565 -143.995 ;
        RECT 275.235 -145.685 275.565 -145.355 ;
        RECT 275.235 -147.045 275.565 -146.715 ;
        RECT 275.235 -148.405 275.565 -148.075 ;
        RECT 275.235 -149.765 275.565 -149.435 ;
        RECT 275.235 -151.125 275.565 -150.795 ;
        RECT 275.235 -152.485 275.565 -152.155 ;
        RECT 275.235 -153.845 275.565 -153.515 ;
        RECT 275.235 -155.205 275.565 -154.875 ;
        RECT 275.235 -156.565 275.565 -156.235 ;
        RECT 275.235 -157.925 275.565 -157.595 ;
        RECT 275.235 -159.285 275.565 -158.955 ;
        RECT 275.235 -160.645 275.565 -160.315 ;
        RECT 275.235 -162.005 275.565 -161.675 ;
        RECT 275.235 -163.365 275.565 -163.035 ;
        RECT 275.235 -164.725 275.565 -164.395 ;
        RECT 275.235 -166.085 275.565 -165.755 ;
        RECT 275.235 -167.445 275.565 -167.115 ;
        RECT 275.235 -168.805 275.565 -168.475 ;
        RECT 275.235 -170.165 275.565 -169.835 ;
        RECT 275.235 -171.525 275.565 -171.195 ;
        RECT 275.235 -172.885 275.565 -172.555 ;
        RECT 275.235 -174.245 275.565 -173.915 ;
        RECT 275.235 -175.605 275.565 -175.275 ;
        RECT 275.235 -176.965 275.565 -176.635 ;
        RECT 275.235 -178.325 275.565 -177.995 ;
        RECT 275.235 -179.685 275.565 -179.355 ;
        RECT 275.235 -181.93 275.565 -180.8 ;
        RECT 275.24 -182.045 275.56 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 275.81 -98.075 276.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.595 241.32 276.925 242.45 ;
        RECT 276.595 239.195 276.925 239.525 ;
        RECT 276.595 237.835 276.925 238.165 ;
        RECT 276.6 237.16 276.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 276.595 -1.525 276.925 -1.195 ;
        RECT 276.595 -2.885 276.925 -2.555 ;
        RECT 276.6 -3.56 276.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.955 241.32 278.285 242.45 ;
        RECT 277.955 239.195 278.285 239.525 ;
        RECT 277.955 237.835 278.285 238.165 ;
        RECT 277.96 237.16 278.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 277.955 -1.525 278.285 -1.195 ;
        RECT 277.955 -2.885 278.285 -2.555 ;
        RECT 277.96 -3.56 278.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.315 241.32 279.645 242.45 ;
        RECT 279.315 239.195 279.645 239.525 ;
        RECT 279.315 237.835 279.645 238.165 ;
        RECT 279.32 237.16 279.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.315 -1.525 279.645 -1.195 ;
        RECT 279.315 -2.885 279.645 -2.555 ;
        RECT 279.32 -3.56 279.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 279.315 -95.365 279.645 -95.035 ;
        RECT 279.315 -96.725 279.645 -96.395 ;
        RECT 279.315 -98.085 279.645 -97.755 ;
        RECT 279.315 -99.445 279.645 -99.115 ;
        RECT 279.315 -100.805 279.645 -100.475 ;
        RECT 279.315 -102.165 279.645 -101.835 ;
        RECT 279.315 -103.525 279.645 -103.195 ;
        RECT 279.315 -104.885 279.645 -104.555 ;
        RECT 279.315 -106.245 279.645 -105.915 ;
        RECT 279.315 -107.605 279.645 -107.275 ;
        RECT 279.315 -108.965 279.645 -108.635 ;
        RECT 279.315 -110.325 279.645 -109.995 ;
        RECT 279.315 -111.685 279.645 -111.355 ;
        RECT 279.315 -113.045 279.645 -112.715 ;
        RECT 279.315 -114.405 279.645 -114.075 ;
        RECT 279.315 -115.765 279.645 -115.435 ;
        RECT 279.315 -117.125 279.645 -116.795 ;
        RECT 279.315 -118.485 279.645 -118.155 ;
        RECT 279.315 -119.845 279.645 -119.515 ;
        RECT 279.315 -121.205 279.645 -120.875 ;
        RECT 279.315 -122.565 279.645 -122.235 ;
        RECT 279.315 -123.925 279.645 -123.595 ;
        RECT 279.315 -125.285 279.645 -124.955 ;
        RECT 279.315 -126.645 279.645 -126.315 ;
        RECT 279.315 -128.005 279.645 -127.675 ;
        RECT 279.315 -129.365 279.645 -129.035 ;
        RECT 279.315 -130.725 279.645 -130.395 ;
        RECT 279.315 -132.085 279.645 -131.755 ;
        RECT 279.315 -133.445 279.645 -133.115 ;
        RECT 279.315 -134.805 279.645 -134.475 ;
        RECT 279.315 -136.165 279.645 -135.835 ;
        RECT 279.315 -137.525 279.645 -137.195 ;
        RECT 279.315 -138.885 279.645 -138.555 ;
        RECT 279.315 -140.245 279.645 -139.915 ;
        RECT 279.315 -141.605 279.645 -141.275 ;
        RECT 279.315 -142.965 279.645 -142.635 ;
        RECT 279.315 -144.325 279.645 -143.995 ;
        RECT 279.315 -145.685 279.645 -145.355 ;
        RECT 279.315 -147.045 279.645 -146.715 ;
        RECT 279.315 -148.405 279.645 -148.075 ;
        RECT 279.315 -149.765 279.645 -149.435 ;
        RECT 279.315 -151.125 279.645 -150.795 ;
        RECT 279.315 -152.485 279.645 -152.155 ;
        RECT 279.315 -153.845 279.645 -153.515 ;
        RECT 279.315 -155.205 279.645 -154.875 ;
        RECT 279.315 -156.565 279.645 -156.235 ;
        RECT 279.315 -157.925 279.645 -157.595 ;
        RECT 279.315 -159.285 279.645 -158.955 ;
        RECT 279.315 -160.645 279.645 -160.315 ;
        RECT 279.315 -162.005 279.645 -161.675 ;
        RECT 279.315 -163.365 279.645 -163.035 ;
        RECT 279.315 -164.725 279.645 -164.395 ;
        RECT 279.315 -166.085 279.645 -165.755 ;
        RECT 279.315 -167.445 279.645 -167.115 ;
        RECT 279.315 -168.805 279.645 -168.475 ;
        RECT 279.315 -170.165 279.645 -169.835 ;
        RECT 279.315 -171.525 279.645 -171.195 ;
        RECT 279.315 -172.885 279.645 -172.555 ;
        RECT 279.315 -174.245 279.645 -173.915 ;
        RECT 279.315 -175.605 279.645 -175.275 ;
        RECT 279.315 -176.965 279.645 -176.635 ;
        RECT 279.315 -178.325 279.645 -177.995 ;
        RECT 279.315 -179.685 279.645 -179.355 ;
        RECT 279.315 -181.93 279.645 -180.8 ;
        RECT 279.32 -182.045 279.64 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.675 241.32 281.005 242.45 ;
        RECT 280.675 239.195 281.005 239.525 ;
        RECT 280.675 237.835 281.005 238.165 ;
        RECT 280.68 237.16 281 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.675 -1.525 281.005 -1.195 ;
        RECT 280.675 -2.885 281.005 -2.555 ;
        RECT 280.68 -3.56 281 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 280.675 -95.365 281.005 -95.035 ;
        RECT 280.675 -96.725 281.005 -96.395 ;
        RECT 280.675 -98.085 281.005 -97.755 ;
        RECT 280.675 -99.445 281.005 -99.115 ;
        RECT 280.675 -100.805 281.005 -100.475 ;
        RECT 280.675 -102.165 281.005 -101.835 ;
        RECT 280.675 -103.525 281.005 -103.195 ;
        RECT 280.675 -104.885 281.005 -104.555 ;
        RECT 280.675 -106.245 281.005 -105.915 ;
        RECT 280.675 -107.605 281.005 -107.275 ;
        RECT 280.675 -108.965 281.005 -108.635 ;
        RECT 280.675 -110.325 281.005 -109.995 ;
        RECT 280.675 -111.685 281.005 -111.355 ;
        RECT 280.675 -113.045 281.005 -112.715 ;
        RECT 280.675 -114.405 281.005 -114.075 ;
        RECT 280.675 -115.765 281.005 -115.435 ;
        RECT 280.675 -117.125 281.005 -116.795 ;
        RECT 280.675 -118.485 281.005 -118.155 ;
        RECT 280.675 -119.845 281.005 -119.515 ;
        RECT 280.675 -121.205 281.005 -120.875 ;
        RECT 280.675 -122.565 281.005 -122.235 ;
        RECT 280.675 -123.925 281.005 -123.595 ;
        RECT 280.675 -125.285 281.005 -124.955 ;
        RECT 280.675 -126.645 281.005 -126.315 ;
        RECT 280.675 -128.005 281.005 -127.675 ;
        RECT 280.675 -129.365 281.005 -129.035 ;
        RECT 280.675 -130.725 281.005 -130.395 ;
        RECT 280.675 -132.085 281.005 -131.755 ;
        RECT 280.675 -133.445 281.005 -133.115 ;
        RECT 280.675 -134.805 281.005 -134.475 ;
        RECT 280.675 -136.165 281.005 -135.835 ;
        RECT 280.675 -137.525 281.005 -137.195 ;
        RECT 280.675 -138.885 281.005 -138.555 ;
        RECT 280.675 -140.245 281.005 -139.915 ;
        RECT 280.675 -141.605 281.005 -141.275 ;
        RECT 280.675 -142.965 281.005 -142.635 ;
        RECT 280.675 -144.325 281.005 -143.995 ;
        RECT 280.675 -145.685 281.005 -145.355 ;
        RECT 280.675 -147.045 281.005 -146.715 ;
        RECT 280.675 -148.405 281.005 -148.075 ;
        RECT 280.675 -149.765 281.005 -149.435 ;
        RECT 280.675 -151.125 281.005 -150.795 ;
        RECT 280.675 -152.485 281.005 -152.155 ;
        RECT 280.675 -153.845 281.005 -153.515 ;
        RECT 280.675 -155.205 281.005 -154.875 ;
        RECT 280.675 -156.565 281.005 -156.235 ;
        RECT 280.675 -157.925 281.005 -157.595 ;
        RECT 280.675 -159.285 281.005 -158.955 ;
        RECT 280.675 -160.645 281.005 -160.315 ;
        RECT 280.675 -162.005 281.005 -161.675 ;
        RECT 280.675 -163.365 281.005 -163.035 ;
        RECT 280.675 -164.725 281.005 -164.395 ;
        RECT 280.675 -166.085 281.005 -165.755 ;
        RECT 280.675 -167.445 281.005 -167.115 ;
        RECT 280.675 -168.805 281.005 -168.475 ;
        RECT 280.675 -170.165 281.005 -169.835 ;
        RECT 280.675 -171.525 281.005 -171.195 ;
        RECT 280.675 -172.885 281.005 -172.555 ;
        RECT 280.675 -174.245 281.005 -173.915 ;
        RECT 280.675 -175.605 281.005 -175.275 ;
        RECT 280.675 -176.965 281.005 -176.635 ;
        RECT 280.675 -178.325 281.005 -177.995 ;
        RECT 280.675 -179.685 281.005 -179.355 ;
        RECT 280.675 -181.93 281.005 -180.8 ;
        RECT 280.68 -182.045 281 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.035 241.32 282.365 242.45 ;
        RECT 282.035 239.195 282.365 239.525 ;
        RECT 282.035 237.835 282.365 238.165 ;
        RECT 282.04 237.16 282.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.035 -1.525 282.365 -1.195 ;
        RECT 282.035 -2.885 282.365 -2.555 ;
        RECT 282.04 -3.56 282.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 282.035 -95.365 282.365 -95.035 ;
        RECT 282.035 -96.725 282.365 -96.395 ;
        RECT 282.035 -98.085 282.365 -97.755 ;
        RECT 282.035 -99.445 282.365 -99.115 ;
        RECT 282.035 -100.805 282.365 -100.475 ;
        RECT 282.035 -102.165 282.365 -101.835 ;
        RECT 282.035 -103.525 282.365 -103.195 ;
        RECT 282.035 -104.885 282.365 -104.555 ;
        RECT 282.035 -106.245 282.365 -105.915 ;
        RECT 282.035 -107.605 282.365 -107.275 ;
        RECT 282.035 -108.965 282.365 -108.635 ;
        RECT 282.035 -110.325 282.365 -109.995 ;
        RECT 282.035 -111.685 282.365 -111.355 ;
        RECT 282.035 -113.045 282.365 -112.715 ;
        RECT 282.035 -114.405 282.365 -114.075 ;
        RECT 282.035 -115.765 282.365 -115.435 ;
        RECT 282.035 -117.125 282.365 -116.795 ;
        RECT 282.035 -118.485 282.365 -118.155 ;
        RECT 282.035 -119.845 282.365 -119.515 ;
        RECT 282.035 -121.205 282.365 -120.875 ;
        RECT 282.035 -122.565 282.365 -122.235 ;
        RECT 282.035 -123.925 282.365 -123.595 ;
        RECT 282.035 -125.285 282.365 -124.955 ;
        RECT 282.035 -126.645 282.365 -126.315 ;
        RECT 282.035 -128.005 282.365 -127.675 ;
        RECT 282.035 -129.365 282.365 -129.035 ;
        RECT 282.035 -130.725 282.365 -130.395 ;
        RECT 282.035 -132.085 282.365 -131.755 ;
        RECT 282.035 -133.445 282.365 -133.115 ;
        RECT 282.035 -134.805 282.365 -134.475 ;
        RECT 282.035 -136.165 282.365 -135.835 ;
        RECT 282.035 -137.525 282.365 -137.195 ;
        RECT 282.035 -138.885 282.365 -138.555 ;
        RECT 282.035 -140.245 282.365 -139.915 ;
        RECT 282.035 -141.605 282.365 -141.275 ;
        RECT 282.035 -142.965 282.365 -142.635 ;
        RECT 282.035 -144.325 282.365 -143.995 ;
        RECT 282.035 -145.685 282.365 -145.355 ;
        RECT 282.035 -147.045 282.365 -146.715 ;
        RECT 282.035 -148.405 282.365 -148.075 ;
        RECT 282.035 -149.765 282.365 -149.435 ;
        RECT 282.035 -151.125 282.365 -150.795 ;
        RECT 282.035 -152.485 282.365 -152.155 ;
        RECT 282.035 -153.845 282.365 -153.515 ;
        RECT 282.035 -155.205 282.365 -154.875 ;
        RECT 282.035 -156.565 282.365 -156.235 ;
        RECT 282.035 -157.925 282.365 -157.595 ;
        RECT 282.035 -159.285 282.365 -158.955 ;
        RECT 282.035 -160.645 282.365 -160.315 ;
        RECT 282.035 -162.005 282.365 -161.675 ;
        RECT 282.035 -163.365 282.365 -163.035 ;
        RECT 282.035 -164.725 282.365 -164.395 ;
        RECT 282.035 -166.085 282.365 -165.755 ;
        RECT 282.035 -167.445 282.365 -167.115 ;
        RECT 282.035 -168.805 282.365 -168.475 ;
        RECT 282.035 -170.165 282.365 -169.835 ;
        RECT 282.035 -171.525 282.365 -171.195 ;
        RECT 282.035 -172.885 282.365 -172.555 ;
        RECT 282.035 -174.245 282.365 -173.915 ;
        RECT 282.035 -175.605 282.365 -175.275 ;
        RECT 282.035 -176.965 282.365 -176.635 ;
        RECT 282.035 -178.325 282.365 -177.995 ;
        RECT 282.035 -179.685 282.365 -179.355 ;
        RECT 282.035 -181.93 282.365 -180.8 ;
        RECT 282.04 -182.045 282.36 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.395 241.32 283.725 242.45 ;
        RECT 283.395 239.195 283.725 239.525 ;
        RECT 283.395 237.835 283.725 238.165 ;
        RECT 283.4 237.16 283.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.395 -1.525 283.725 -1.195 ;
        RECT 283.395 -2.885 283.725 -2.555 ;
        RECT 283.4 -3.56 283.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 283.395 -95.365 283.725 -95.035 ;
        RECT 283.395 -96.725 283.725 -96.395 ;
        RECT 283.395 -98.085 283.725 -97.755 ;
        RECT 283.395 -99.445 283.725 -99.115 ;
        RECT 283.395 -100.805 283.725 -100.475 ;
        RECT 283.395 -102.165 283.725 -101.835 ;
        RECT 283.395 -103.525 283.725 -103.195 ;
        RECT 283.395 -104.885 283.725 -104.555 ;
        RECT 283.395 -106.245 283.725 -105.915 ;
        RECT 283.395 -107.605 283.725 -107.275 ;
        RECT 283.395 -108.965 283.725 -108.635 ;
        RECT 283.395 -110.325 283.725 -109.995 ;
        RECT 283.395 -111.685 283.725 -111.355 ;
        RECT 283.395 -113.045 283.725 -112.715 ;
        RECT 283.395 -114.405 283.725 -114.075 ;
        RECT 283.395 -115.765 283.725 -115.435 ;
        RECT 283.395 -117.125 283.725 -116.795 ;
        RECT 283.395 -118.485 283.725 -118.155 ;
        RECT 283.395 -119.845 283.725 -119.515 ;
        RECT 283.395 -121.205 283.725 -120.875 ;
        RECT 283.395 -122.565 283.725 -122.235 ;
        RECT 283.395 -123.925 283.725 -123.595 ;
        RECT 283.395 -125.285 283.725 -124.955 ;
        RECT 283.395 -126.645 283.725 -126.315 ;
        RECT 283.395 -128.005 283.725 -127.675 ;
        RECT 283.395 -129.365 283.725 -129.035 ;
        RECT 283.395 -130.725 283.725 -130.395 ;
        RECT 283.395 -132.085 283.725 -131.755 ;
        RECT 283.395 -133.445 283.725 -133.115 ;
        RECT 283.395 -134.805 283.725 -134.475 ;
        RECT 283.395 -136.165 283.725 -135.835 ;
        RECT 283.395 -137.525 283.725 -137.195 ;
        RECT 283.395 -138.885 283.725 -138.555 ;
        RECT 283.395 -140.245 283.725 -139.915 ;
        RECT 283.395 -141.605 283.725 -141.275 ;
        RECT 283.395 -142.965 283.725 -142.635 ;
        RECT 283.395 -144.325 283.725 -143.995 ;
        RECT 283.395 -145.685 283.725 -145.355 ;
        RECT 283.395 -147.045 283.725 -146.715 ;
        RECT 283.395 -148.405 283.725 -148.075 ;
        RECT 283.395 -149.765 283.725 -149.435 ;
        RECT 283.395 -151.125 283.725 -150.795 ;
        RECT 283.395 -152.485 283.725 -152.155 ;
        RECT 283.395 -153.845 283.725 -153.515 ;
        RECT 283.395 -155.205 283.725 -154.875 ;
        RECT 283.395 -156.565 283.725 -156.235 ;
        RECT 283.395 -157.925 283.725 -157.595 ;
        RECT 283.395 -159.285 283.725 -158.955 ;
        RECT 283.395 -160.645 283.725 -160.315 ;
        RECT 283.395 -162.005 283.725 -161.675 ;
        RECT 283.395 -163.365 283.725 -163.035 ;
        RECT 283.395 -164.725 283.725 -164.395 ;
        RECT 283.395 -166.085 283.725 -165.755 ;
        RECT 283.395 -167.445 283.725 -167.115 ;
        RECT 283.395 -168.805 283.725 -168.475 ;
        RECT 283.395 -170.165 283.725 -169.835 ;
        RECT 283.395 -171.525 283.725 -171.195 ;
        RECT 283.395 -172.885 283.725 -172.555 ;
        RECT 283.395 -174.245 283.725 -173.915 ;
        RECT 283.395 -175.605 283.725 -175.275 ;
        RECT 283.395 -176.965 283.725 -176.635 ;
        RECT 283.395 -178.325 283.725 -177.995 ;
        RECT 283.395 -179.685 283.725 -179.355 ;
        RECT 283.395 -181.93 283.725 -180.8 ;
        RECT 283.4 -182.045 283.72 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.755 241.32 285.085 242.45 ;
        RECT 284.755 239.195 285.085 239.525 ;
        RECT 284.755 237.835 285.085 238.165 ;
        RECT 284.76 237.16 285.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.755 -1.525 285.085 -1.195 ;
        RECT 284.755 -2.885 285.085 -2.555 ;
        RECT 284.76 -3.56 285.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 284.755 -95.365 285.085 -95.035 ;
        RECT 284.755 -96.725 285.085 -96.395 ;
        RECT 284.755 -98.085 285.085 -97.755 ;
        RECT 284.755 -99.445 285.085 -99.115 ;
        RECT 284.755 -100.805 285.085 -100.475 ;
        RECT 284.755 -102.165 285.085 -101.835 ;
        RECT 284.755 -103.525 285.085 -103.195 ;
        RECT 284.755 -104.885 285.085 -104.555 ;
        RECT 284.755 -106.245 285.085 -105.915 ;
        RECT 284.755 -107.605 285.085 -107.275 ;
        RECT 284.755 -108.965 285.085 -108.635 ;
        RECT 284.755 -110.325 285.085 -109.995 ;
        RECT 284.755 -111.685 285.085 -111.355 ;
        RECT 284.755 -113.045 285.085 -112.715 ;
        RECT 284.755 -114.405 285.085 -114.075 ;
        RECT 284.755 -115.765 285.085 -115.435 ;
        RECT 284.755 -117.125 285.085 -116.795 ;
        RECT 284.755 -118.485 285.085 -118.155 ;
        RECT 284.755 -119.845 285.085 -119.515 ;
        RECT 284.755 -121.205 285.085 -120.875 ;
        RECT 284.755 -122.565 285.085 -122.235 ;
        RECT 284.755 -123.925 285.085 -123.595 ;
        RECT 284.755 -125.285 285.085 -124.955 ;
        RECT 284.755 -126.645 285.085 -126.315 ;
        RECT 284.755 -128.005 285.085 -127.675 ;
        RECT 284.755 -129.365 285.085 -129.035 ;
        RECT 284.755 -130.725 285.085 -130.395 ;
        RECT 284.755 -132.085 285.085 -131.755 ;
        RECT 284.755 -133.445 285.085 -133.115 ;
        RECT 284.755 -134.805 285.085 -134.475 ;
        RECT 284.755 -136.165 285.085 -135.835 ;
        RECT 284.755 -137.525 285.085 -137.195 ;
        RECT 284.755 -138.885 285.085 -138.555 ;
        RECT 284.755 -140.245 285.085 -139.915 ;
        RECT 284.755 -141.605 285.085 -141.275 ;
        RECT 284.755 -142.965 285.085 -142.635 ;
        RECT 284.755 -144.325 285.085 -143.995 ;
        RECT 284.755 -145.685 285.085 -145.355 ;
        RECT 284.755 -147.045 285.085 -146.715 ;
        RECT 284.755 -148.405 285.085 -148.075 ;
        RECT 284.755 -149.765 285.085 -149.435 ;
        RECT 284.755 -151.125 285.085 -150.795 ;
        RECT 284.755 -152.485 285.085 -152.155 ;
        RECT 284.755 -153.845 285.085 -153.515 ;
        RECT 284.755 -155.205 285.085 -154.875 ;
        RECT 284.755 -156.565 285.085 -156.235 ;
        RECT 284.755 -157.925 285.085 -157.595 ;
        RECT 284.755 -159.285 285.085 -158.955 ;
        RECT 284.755 -160.645 285.085 -160.315 ;
        RECT 284.755 -162.005 285.085 -161.675 ;
        RECT 284.755 -163.365 285.085 -163.035 ;
        RECT 284.755 -164.725 285.085 -164.395 ;
        RECT 284.755 -166.085 285.085 -165.755 ;
        RECT 284.755 -167.445 285.085 -167.115 ;
        RECT 284.755 -168.805 285.085 -168.475 ;
        RECT 284.755 -170.165 285.085 -169.835 ;
        RECT 284.755 -171.525 285.085 -171.195 ;
        RECT 284.755 -172.885 285.085 -172.555 ;
        RECT 284.755 -174.245 285.085 -173.915 ;
        RECT 284.755 -175.605 285.085 -175.275 ;
        RECT 284.755 -176.965 285.085 -176.635 ;
        RECT 284.755 -178.325 285.085 -177.995 ;
        RECT 284.755 -179.685 285.085 -179.355 ;
        RECT 284.755 -181.93 285.085 -180.8 ;
        RECT 284.76 -182.045 285.08 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.115 241.32 286.445 242.45 ;
        RECT 286.115 239.195 286.445 239.525 ;
        RECT 286.115 237.835 286.445 238.165 ;
        RECT 286.12 237.16 286.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.115 -99.445 286.445 -99.115 ;
        RECT 286.115 -100.805 286.445 -100.475 ;
        RECT 286.115 -102.165 286.445 -101.835 ;
        RECT 286.115 -103.525 286.445 -103.195 ;
        RECT 286.115 -104.885 286.445 -104.555 ;
        RECT 286.115 -106.245 286.445 -105.915 ;
        RECT 286.115 -107.605 286.445 -107.275 ;
        RECT 286.115 -108.965 286.445 -108.635 ;
        RECT 286.115 -110.325 286.445 -109.995 ;
        RECT 286.115 -111.685 286.445 -111.355 ;
        RECT 286.115 -113.045 286.445 -112.715 ;
        RECT 286.115 -114.405 286.445 -114.075 ;
        RECT 286.115 -115.765 286.445 -115.435 ;
        RECT 286.115 -117.125 286.445 -116.795 ;
        RECT 286.115 -118.485 286.445 -118.155 ;
        RECT 286.115 -119.845 286.445 -119.515 ;
        RECT 286.115 -121.205 286.445 -120.875 ;
        RECT 286.115 -122.565 286.445 -122.235 ;
        RECT 286.115 -123.925 286.445 -123.595 ;
        RECT 286.115 -125.285 286.445 -124.955 ;
        RECT 286.115 -126.645 286.445 -126.315 ;
        RECT 286.115 -128.005 286.445 -127.675 ;
        RECT 286.115 -129.365 286.445 -129.035 ;
        RECT 286.115 -130.725 286.445 -130.395 ;
        RECT 286.115 -132.085 286.445 -131.755 ;
        RECT 286.115 -133.445 286.445 -133.115 ;
        RECT 286.115 -134.805 286.445 -134.475 ;
        RECT 286.115 -136.165 286.445 -135.835 ;
        RECT 286.115 -137.525 286.445 -137.195 ;
        RECT 286.115 -138.885 286.445 -138.555 ;
        RECT 286.115 -140.245 286.445 -139.915 ;
        RECT 286.115 -141.605 286.445 -141.275 ;
        RECT 286.115 -142.965 286.445 -142.635 ;
        RECT 286.115 -144.325 286.445 -143.995 ;
        RECT 286.115 -145.685 286.445 -145.355 ;
        RECT 286.115 -147.045 286.445 -146.715 ;
        RECT 286.115 -148.405 286.445 -148.075 ;
        RECT 286.115 -149.765 286.445 -149.435 ;
        RECT 286.115 -151.125 286.445 -150.795 ;
        RECT 286.115 -152.485 286.445 -152.155 ;
        RECT 286.115 -153.845 286.445 -153.515 ;
        RECT 286.115 -155.205 286.445 -154.875 ;
        RECT 286.115 -156.565 286.445 -156.235 ;
        RECT 286.115 -157.925 286.445 -157.595 ;
        RECT 286.115 -159.285 286.445 -158.955 ;
        RECT 286.115 -160.645 286.445 -160.315 ;
        RECT 286.115 -162.005 286.445 -161.675 ;
        RECT 286.115 -163.365 286.445 -163.035 ;
        RECT 286.115 -164.725 286.445 -164.395 ;
        RECT 286.115 -166.085 286.445 -165.755 ;
        RECT 286.115 -167.445 286.445 -167.115 ;
        RECT 286.115 -168.805 286.445 -168.475 ;
        RECT 286.115 -170.165 286.445 -169.835 ;
        RECT 286.115 -171.525 286.445 -171.195 ;
        RECT 286.115 -172.885 286.445 -172.555 ;
        RECT 286.115 -174.245 286.445 -173.915 ;
        RECT 286.115 -175.605 286.445 -175.275 ;
        RECT 286.115 -176.965 286.445 -176.635 ;
        RECT 286.115 -178.325 286.445 -177.995 ;
        RECT 286.115 -179.685 286.445 -179.355 ;
        RECT 286.115 -181.93 286.445 -180.8 ;
        RECT 286.12 -182.045 286.44 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 286.71 -98.075 287.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.475 241.32 287.805 242.45 ;
        RECT 287.475 239.195 287.805 239.525 ;
        RECT 287.475 237.835 287.805 238.165 ;
        RECT 287.48 237.16 287.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 287.475 -1.525 287.805 -1.195 ;
        RECT 287.475 -2.885 287.805 -2.555 ;
        RECT 287.48 -3.56 287.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.835 241.32 289.165 242.45 ;
        RECT 288.835 239.195 289.165 239.525 ;
        RECT 288.835 237.835 289.165 238.165 ;
        RECT 288.84 237.16 289.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 288.835 -1.525 289.165 -1.195 ;
        RECT 288.835 -2.885 289.165 -2.555 ;
        RECT 288.84 -3.56 289.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.195 241.32 290.525 242.45 ;
        RECT 290.195 239.195 290.525 239.525 ;
        RECT 290.195 237.835 290.525 238.165 ;
        RECT 290.2 237.16 290.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.195 -1.525 290.525 -1.195 ;
        RECT 290.195 -2.885 290.525 -2.555 ;
        RECT 290.2 -3.56 290.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 290.195 -128.005 290.525 -127.675 ;
        RECT 290.195 -129.365 290.525 -129.035 ;
        RECT 290.195 -130.725 290.525 -130.395 ;
        RECT 290.195 -132.085 290.525 -131.755 ;
        RECT 290.195 -133.445 290.525 -133.115 ;
        RECT 290.195 -134.805 290.525 -134.475 ;
        RECT 290.195 -136.165 290.525 -135.835 ;
        RECT 290.195 -137.525 290.525 -137.195 ;
        RECT 290.195 -138.885 290.525 -138.555 ;
        RECT 290.195 -140.245 290.525 -139.915 ;
        RECT 290.195 -141.605 290.525 -141.275 ;
        RECT 290.195 -142.965 290.525 -142.635 ;
        RECT 290.195 -144.325 290.525 -143.995 ;
        RECT 290.195 -145.685 290.525 -145.355 ;
        RECT 290.195 -147.045 290.525 -146.715 ;
        RECT 290.195 -148.405 290.525 -148.075 ;
        RECT 290.195 -149.765 290.525 -149.435 ;
        RECT 290.195 -151.125 290.525 -150.795 ;
        RECT 290.195 -152.485 290.525 -152.155 ;
        RECT 290.195 -153.845 290.525 -153.515 ;
        RECT 290.195 -155.205 290.525 -154.875 ;
        RECT 290.195 -156.565 290.525 -156.235 ;
        RECT 290.195 -157.925 290.525 -157.595 ;
        RECT 290.195 -159.285 290.525 -158.955 ;
        RECT 290.195 -160.645 290.525 -160.315 ;
        RECT 290.195 -162.005 290.525 -161.675 ;
        RECT 290.195 -163.365 290.525 -163.035 ;
        RECT 290.195 -164.725 290.525 -164.395 ;
        RECT 290.195 -166.085 290.525 -165.755 ;
        RECT 290.195 -167.445 290.525 -167.115 ;
        RECT 290.195 -168.805 290.525 -168.475 ;
        RECT 290.195 -170.165 290.525 -169.835 ;
        RECT 290.195 -171.525 290.525 -171.195 ;
        RECT 290.195 -172.885 290.525 -172.555 ;
        RECT 290.195 -174.245 290.525 -173.915 ;
        RECT 290.195 -175.605 290.525 -175.275 ;
        RECT 290.195 -176.965 290.525 -176.635 ;
        RECT 290.195 -178.325 290.525 -177.995 ;
        RECT 290.195 -179.685 290.525 -179.355 ;
        RECT 290.195 -181.93 290.525 -180.8 ;
        RECT 290.2 -182.045 290.52 -95.035 ;
        RECT 290.195 -95.365 290.525 -95.035 ;
        RECT 290.195 -96.725 290.525 -96.395 ;
        RECT 290.195 -98.085 290.525 -97.755 ;
        RECT 290.195 -99.445 290.525 -99.115 ;
        RECT 290.195 -100.805 290.525 -100.475 ;
        RECT 290.195 -102.165 290.525 -101.835 ;
        RECT 290.195 -103.525 290.525 -103.195 ;
        RECT 290.195 -104.885 290.525 -104.555 ;
        RECT 290.195 -106.245 290.525 -105.915 ;
        RECT 290.195 -107.605 290.525 -107.275 ;
        RECT 290.195 -108.965 290.525 -108.635 ;
        RECT 290.195 -110.325 290.525 -109.995 ;
        RECT 290.195 -111.685 290.525 -111.355 ;
        RECT 290.195 -113.045 290.525 -112.715 ;
        RECT 290.195 -114.405 290.525 -114.075 ;
        RECT 290.195 -115.765 290.525 -115.435 ;
        RECT 290.195 -117.125 290.525 -116.795 ;
        RECT 290.195 -118.485 290.525 -118.155 ;
        RECT 290.195 -119.845 290.525 -119.515 ;
        RECT 290.195 -121.205 290.525 -120.875 ;
        RECT 290.195 -122.565 290.525 -122.235 ;
        RECT 290.195 -123.925 290.525 -123.595 ;
        RECT 290.195 -125.285 290.525 -124.955 ;
        RECT 290.195 -126.645 290.525 -126.315 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.235 241.32 241.565 242.45 ;
        RECT 241.235 239.195 241.565 239.525 ;
        RECT 241.235 237.835 241.565 238.165 ;
        RECT 241.24 237.16 241.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.235 -1.525 241.565 -1.195 ;
        RECT 241.235 -2.885 241.565 -2.555 ;
        RECT 241.24 -3.56 241.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 241.235 -95.365 241.565 -95.035 ;
        RECT 241.235 -96.725 241.565 -96.395 ;
        RECT 241.235 -98.085 241.565 -97.755 ;
        RECT 241.235 -99.445 241.565 -99.115 ;
        RECT 241.235 -100.805 241.565 -100.475 ;
        RECT 241.235 -102.165 241.565 -101.835 ;
        RECT 241.235 -103.525 241.565 -103.195 ;
        RECT 241.235 -104.885 241.565 -104.555 ;
        RECT 241.235 -106.245 241.565 -105.915 ;
        RECT 241.235 -107.605 241.565 -107.275 ;
        RECT 241.235 -108.965 241.565 -108.635 ;
        RECT 241.235 -110.325 241.565 -109.995 ;
        RECT 241.235 -111.685 241.565 -111.355 ;
        RECT 241.235 -113.045 241.565 -112.715 ;
        RECT 241.235 -114.405 241.565 -114.075 ;
        RECT 241.235 -115.765 241.565 -115.435 ;
        RECT 241.235 -117.125 241.565 -116.795 ;
        RECT 241.235 -118.485 241.565 -118.155 ;
        RECT 241.235 -119.845 241.565 -119.515 ;
        RECT 241.235 -121.205 241.565 -120.875 ;
        RECT 241.235 -122.565 241.565 -122.235 ;
        RECT 241.235 -123.925 241.565 -123.595 ;
        RECT 241.235 -125.285 241.565 -124.955 ;
        RECT 241.235 -126.645 241.565 -126.315 ;
        RECT 241.235 -128.005 241.565 -127.675 ;
        RECT 241.235 -129.365 241.565 -129.035 ;
        RECT 241.235 -130.725 241.565 -130.395 ;
        RECT 241.235 -132.085 241.565 -131.755 ;
        RECT 241.235 -133.445 241.565 -133.115 ;
        RECT 241.235 -134.805 241.565 -134.475 ;
        RECT 241.235 -136.165 241.565 -135.835 ;
        RECT 241.235 -137.525 241.565 -137.195 ;
        RECT 241.235 -138.885 241.565 -138.555 ;
        RECT 241.235 -140.245 241.565 -139.915 ;
        RECT 241.235 -141.605 241.565 -141.275 ;
        RECT 241.235 -142.965 241.565 -142.635 ;
        RECT 241.235 -144.325 241.565 -143.995 ;
        RECT 241.235 -145.685 241.565 -145.355 ;
        RECT 241.235 -147.045 241.565 -146.715 ;
        RECT 241.235 -148.405 241.565 -148.075 ;
        RECT 241.235 -149.765 241.565 -149.435 ;
        RECT 241.235 -151.125 241.565 -150.795 ;
        RECT 241.235 -152.485 241.565 -152.155 ;
        RECT 241.235 -153.845 241.565 -153.515 ;
        RECT 241.235 -155.205 241.565 -154.875 ;
        RECT 241.235 -156.565 241.565 -156.235 ;
        RECT 241.235 -157.925 241.565 -157.595 ;
        RECT 241.235 -159.285 241.565 -158.955 ;
        RECT 241.235 -160.645 241.565 -160.315 ;
        RECT 241.235 -162.005 241.565 -161.675 ;
        RECT 241.235 -163.365 241.565 -163.035 ;
        RECT 241.235 -164.725 241.565 -164.395 ;
        RECT 241.235 -166.085 241.565 -165.755 ;
        RECT 241.235 -167.445 241.565 -167.115 ;
        RECT 241.235 -168.805 241.565 -168.475 ;
        RECT 241.235 -170.165 241.565 -169.835 ;
        RECT 241.235 -171.525 241.565 -171.195 ;
        RECT 241.235 -172.885 241.565 -172.555 ;
        RECT 241.235 -174.245 241.565 -173.915 ;
        RECT 241.235 -175.605 241.565 -175.275 ;
        RECT 241.235 -176.965 241.565 -176.635 ;
        RECT 241.235 -178.325 241.565 -177.995 ;
        RECT 241.235 -179.685 241.565 -179.355 ;
        RECT 241.235 -181.93 241.565 -180.8 ;
        RECT 241.24 -182.045 241.56 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.595 241.32 242.925 242.45 ;
        RECT 242.595 239.195 242.925 239.525 ;
        RECT 242.595 237.835 242.925 238.165 ;
        RECT 242.6 237.16 242.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 242.595 -99.445 242.925 -99.115 ;
        RECT 242.595 -100.805 242.925 -100.475 ;
        RECT 242.595 -102.165 242.925 -101.835 ;
        RECT 242.595 -103.525 242.925 -103.195 ;
        RECT 242.595 -104.885 242.925 -104.555 ;
        RECT 242.595 -106.245 242.925 -105.915 ;
        RECT 242.595 -107.605 242.925 -107.275 ;
        RECT 242.595 -108.965 242.925 -108.635 ;
        RECT 242.595 -110.325 242.925 -109.995 ;
        RECT 242.595 -111.685 242.925 -111.355 ;
        RECT 242.595 -113.045 242.925 -112.715 ;
        RECT 242.595 -114.405 242.925 -114.075 ;
        RECT 242.595 -115.765 242.925 -115.435 ;
        RECT 242.595 -117.125 242.925 -116.795 ;
        RECT 242.595 -118.485 242.925 -118.155 ;
        RECT 242.595 -119.845 242.925 -119.515 ;
        RECT 242.595 -121.205 242.925 -120.875 ;
        RECT 242.595 -122.565 242.925 -122.235 ;
        RECT 242.595 -123.925 242.925 -123.595 ;
        RECT 242.595 -125.285 242.925 -124.955 ;
        RECT 242.595 -126.645 242.925 -126.315 ;
        RECT 242.595 -128.005 242.925 -127.675 ;
        RECT 242.595 -129.365 242.925 -129.035 ;
        RECT 242.595 -130.725 242.925 -130.395 ;
        RECT 242.595 -132.085 242.925 -131.755 ;
        RECT 242.595 -133.445 242.925 -133.115 ;
        RECT 242.595 -134.805 242.925 -134.475 ;
        RECT 242.595 -136.165 242.925 -135.835 ;
        RECT 242.595 -137.525 242.925 -137.195 ;
        RECT 242.595 -138.885 242.925 -138.555 ;
        RECT 242.595 -140.245 242.925 -139.915 ;
        RECT 242.595 -141.605 242.925 -141.275 ;
        RECT 242.595 -142.965 242.925 -142.635 ;
        RECT 242.595 -144.325 242.925 -143.995 ;
        RECT 242.595 -145.685 242.925 -145.355 ;
        RECT 242.595 -147.045 242.925 -146.715 ;
        RECT 242.595 -148.405 242.925 -148.075 ;
        RECT 242.595 -149.765 242.925 -149.435 ;
        RECT 242.595 -151.125 242.925 -150.795 ;
        RECT 242.595 -152.485 242.925 -152.155 ;
        RECT 242.595 -153.845 242.925 -153.515 ;
        RECT 242.595 -155.205 242.925 -154.875 ;
        RECT 242.595 -156.565 242.925 -156.235 ;
        RECT 242.595 -157.925 242.925 -157.595 ;
        RECT 242.595 -159.285 242.925 -158.955 ;
        RECT 242.595 -160.645 242.925 -160.315 ;
        RECT 242.595 -162.005 242.925 -161.675 ;
        RECT 242.595 -163.365 242.925 -163.035 ;
        RECT 242.595 -164.725 242.925 -164.395 ;
        RECT 242.595 -166.085 242.925 -165.755 ;
        RECT 242.595 -167.445 242.925 -167.115 ;
        RECT 242.595 -168.805 242.925 -168.475 ;
        RECT 242.595 -170.165 242.925 -169.835 ;
        RECT 242.595 -171.525 242.925 -171.195 ;
        RECT 242.595 -172.885 242.925 -172.555 ;
        RECT 242.595 -174.245 242.925 -173.915 ;
        RECT 242.595 -175.605 242.925 -175.275 ;
        RECT 242.595 -176.965 242.925 -176.635 ;
        RECT 242.595 -178.325 242.925 -177.995 ;
        RECT 242.595 -179.685 242.925 -179.355 ;
        RECT 242.595 -181.93 242.925 -180.8 ;
        RECT 242.6 -182.045 242.92 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.11 -98.075 243.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.955 241.32 244.285 242.45 ;
        RECT 243.955 239.195 244.285 239.525 ;
        RECT 243.955 237.835 244.285 238.165 ;
        RECT 243.96 237.16 244.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 243.955 -1.525 244.285 -1.195 ;
        RECT 243.955 -2.885 244.285 -2.555 ;
        RECT 243.96 -3.56 244.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.315 241.32 245.645 242.45 ;
        RECT 245.315 239.195 245.645 239.525 ;
        RECT 245.315 237.835 245.645 238.165 ;
        RECT 245.32 237.16 245.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 245.315 -1.525 245.645 -1.195 ;
        RECT 245.315 -2.885 245.645 -2.555 ;
        RECT 245.32 -3.56 245.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.675 241.32 247.005 242.45 ;
        RECT 246.675 239.195 247.005 239.525 ;
        RECT 246.675 237.835 247.005 238.165 ;
        RECT 246.68 237.16 247 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.675 -1.525 247.005 -1.195 ;
        RECT 246.675 -2.885 247.005 -2.555 ;
        RECT 246.68 -3.56 247 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 246.675 -95.365 247.005 -95.035 ;
        RECT 246.675 -96.725 247.005 -96.395 ;
        RECT 246.675 -98.085 247.005 -97.755 ;
        RECT 246.675 -99.445 247.005 -99.115 ;
        RECT 246.675 -100.805 247.005 -100.475 ;
        RECT 246.675 -102.165 247.005 -101.835 ;
        RECT 246.675 -103.525 247.005 -103.195 ;
        RECT 246.675 -104.885 247.005 -104.555 ;
        RECT 246.675 -106.245 247.005 -105.915 ;
        RECT 246.675 -107.605 247.005 -107.275 ;
        RECT 246.675 -108.965 247.005 -108.635 ;
        RECT 246.675 -110.325 247.005 -109.995 ;
        RECT 246.675 -111.685 247.005 -111.355 ;
        RECT 246.675 -113.045 247.005 -112.715 ;
        RECT 246.675 -114.405 247.005 -114.075 ;
        RECT 246.675 -115.765 247.005 -115.435 ;
        RECT 246.675 -117.125 247.005 -116.795 ;
        RECT 246.675 -118.485 247.005 -118.155 ;
        RECT 246.675 -119.845 247.005 -119.515 ;
        RECT 246.675 -121.205 247.005 -120.875 ;
        RECT 246.675 -122.565 247.005 -122.235 ;
        RECT 246.675 -123.925 247.005 -123.595 ;
        RECT 246.675 -125.285 247.005 -124.955 ;
        RECT 246.675 -126.645 247.005 -126.315 ;
        RECT 246.675 -128.005 247.005 -127.675 ;
        RECT 246.675 -129.365 247.005 -129.035 ;
        RECT 246.675 -130.725 247.005 -130.395 ;
        RECT 246.675 -132.085 247.005 -131.755 ;
        RECT 246.675 -133.445 247.005 -133.115 ;
        RECT 246.675 -134.805 247.005 -134.475 ;
        RECT 246.675 -136.165 247.005 -135.835 ;
        RECT 246.675 -137.525 247.005 -137.195 ;
        RECT 246.675 -138.885 247.005 -138.555 ;
        RECT 246.675 -140.245 247.005 -139.915 ;
        RECT 246.675 -141.605 247.005 -141.275 ;
        RECT 246.675 -142.965 247.005 -142.635 ;
        RECT 246.675 -144.325 247.005 -143.995 ;
        RECT 246.675 -145.685 247.005 -145.355 ;
        RECT 246.675 -147.045 247.005 -146.715 ;
        RECT 246.675 -148.405 247.005 -148.075 ;
        RECT 246.675 -149.765 247.005 -149.435 ;
        RECT 246.675 -151.125 247.005 -150.795 ;
        RECT 246.675 -152.485 247.005 -152.155 ;
        RECT 246.675 -153.845 247.005 -153.515 ;
        RECT 246.675 -155.205 247.005 -154.875 ;
        RECT 246.675 -156.565 247.005 -156.235 ;
        RECT 246.675 -157.925 247.005 -157.595 ;
        RECT 246.675 -159.285 247.005 -158.955 ;
        RECT 246.675 -160.645 247.005 -160.315 ;
        RECT 246.675 -162.005 247.005 -161.675 ;
        RECT 246.675 -163.365 247.005 -163.035 ;
        RECT 246.675 -164.725 247.005 -164.395 ;
        RECT 246.675 -166.085 247.005 -165.755 ;
        RECT 246.675 -167.445 247.005 -167.115 ;
        RECT 246.675 -168.805 247.005 -168.475 ;
        RECT 246.675 -170.165 247.005 -169.835 ;
        RECT 246.675 -171.525 247.005 -171.195 ;
        RECT 246.675 -172.885 247.005 -172.555 ;
        RECT 246.675 -174.245 247.005 -173.915 ;
        RECT 246.675 -175.605 247.005 -175.275 ;
        RECT 246.675 -176.965 247.005 -176.635 ;
        RECT 246.675 -178.325 247.005 -177.995 ;
        RECT 246.675 -179.685 247.005 -179.355 ;
        RECT 246.675 -181.93 247.005 -180.8 ;
        RECT 246.68 -182.045 247 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.035 241.32 248.365 242.45 ;
        RECT 248.035 239.195 248.365 239.525 ;
        RECT 248.035 237.835 248.365 238.165 ;
        RECT 248.04 237.16 248.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.035 -1.525 248.365 -1.195 ;
        RECT 248.035 -2.885 248.365 -2.555 ;
        RECT 248.04 -3.56 248.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 248.035 -95.365 248.365 -95.035 ;
        RECT 248.035 -96.725 248.365 -96.395 ;
        RECT 248.035 -98.085 248.365 -97.755 ;
        RECT 248.035 -99.445 248.365 -99.115 ;
        RECT 248.035 -100.805 248.365 -100.475 ;
        RECT 248.035 -102.165 248.365 -101.835 ;
        RECT 248.035 -103.525 248.365 -103.195 ;
        RECT 248.035 -104.885 248.365 -104.555 ;
        RECT 248.035 -106.245 248.365 -105.915 ;
        RECT 248.035 -107.605 248.365 -107.275 ;
        RECT 248.035 -108.965 248.365 -108.635 ;
        RECT 248.035 -110.325 248.365 -109.995 ;
        RECT 248.035 -111.685 248.365 -111.355 ;
        RECT 248.035 -113.045 248.365 -112.715 ;
        RECT 248.035 -114.405 248.365 -114.075 ;
        RECT 248.035 -115.765 248.365 -115.435 ;
        RECT 248.035 -117.125 248.365 -116.795 ;
        RECT 248.035 -118.485 248.365 -118.155 ;
        RECT 248.035 -119.845 248.365 -119.515 ;
        RECT 248.035 -121.205 248.365 -120.875 ;
        RECT 248.035 -122.565 248.365 -122.235 ;
        RECT 248.035 -123.925 248.365 -123.595 ;
        RECT 248.035 -125.285 248.365 -124.955 ;
        RECT 248.035 -126.645 248.365 -126.315 ;
        RECT 248.035 -128.005 248.365 -127.675 ;
        RECT 248.035 -129.365 248.365 -129.035 ;
        RECT 248.035 -130.725 248.365 -130.395 ;
        RECT 248.035 -132.085 248.365 -131.755 ;
        RECT 248.035 -133.445 248.365 -133.115 ;
        RECT 248.035 -134.805 248.365 -134.475 ;
        RECT 248.035 -136.165 248.365 -135.835 ;
        RECT 248.035 -137.525 248.365 -137.195 ;
        RECT 248.035 -138.885 248.365 -138.555 ;
        RECT 248.035 -140.245 248.365 -139.915 ;
        RECT 248.035 -141.605 248.365 -141.275 ;
        RECT 248.035 -142.965 248.365 -142.635 ;
        RECT 248.035 -144.325 248.365 -143.995 ;
        RECT 248.035 -145.685 248.365 -145.355 ;
        RECT 248.035 -147.045 248.365 -146.715 ;
        RECT 248.035 -148.405 248.365 -148.075 ;
        RECT 248.035 -149.765 248.365 -149.435 ;
        RECT 248.035 -151.125 248.365 -150.795 ;
        RECT 248.035 -152.485 248.365 -152.155 ;
        RECT 248.035 -153.845 248.365 -153.515 ;
        RECT 248.035 -155.205 248.365 -154.875 ;
        RECT 248.035 -156.565 248.365 -156.235 ;
        RECT 248.035 -157.925 248.365 -157.595 ;
        RECT 248.035 -159.285 248.365 -158.955 ;
        RECT 248.035 -160.645 248.365 -160.315 ;
        RECT 248.035 -162.005 248.365 -161.675 ;
        RECT 248.035 -163.365 248.365 -163.035 ;
        RECT 248.035 -164.725 248.365 -164.395 ;
        RECT 248.035 -166.085 248.365 -165.755 ;
        RECT 248.035 -167.445 248.365 -167.115 ;
        RECT 248.035 -168.805 248.365 -168.475 ;
        RECT 248.035 -170.165 248.365 -169.835 ;
        RECT 248.035 -171.525 248.365 -171.195 ;
        RECT 248.035 -172.885 248.365 -172.555 ;
        RECT 248.035 -174.245 248.365 -173.915 ;
        RECT 248.035 -175.605 248.365 -175.275 ;
        RECT 248.035 -176.965 248.365 -176.635 ;
        RECT 248.035 -178.325 248.365 -177.995 ;
        RECT 248.035 -179.685 248.365 -179.355 ;
        RECT 248.035 -181.93 248.365 -180.8 ;
        RECT 248.04 -182.045 248.36 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.395 241.32 249.725 242.45 ;
        RECT 249.395 239.195 249.725 239.525 ;
        RECT 249.395 237.835 249.725 238.165 ;
        RECT 249.4 237.16 249.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.395 -1.525 249.725 -1.195 ;
        RECT 249.395 -2.885 249.725 -2.555 ;
        RECT 249.4 -3.56 249.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 249.395 -95.365 249.725 -95.035 ;
        RECT 249.395 -96.725 249.725 -96.395 ;
        RECT 249.395 -98.085 249.725 -97.755 ;
        RECT 249.395 -99.445 249.725 -99.115 ;
        RECT 249.395 -100.805 249.725 -100.475 ;
        RECT 249.395 -102.165 249.725 -101.835 ;
        RECT 249.395 -103.525 249.725 -103.195 ;
        RECT 249.395 -104.885 249.725 -104.555 ;
        RECT 249.395 -106.245 249.725 -105.915 ;
        RECT 249.395 -107.605 249.725 -107.275 ;
        RECT 249.395 -108.965 249.725 -108.635 ;
        RECT 249.395 -110.325 249.725 -109.995 ;
        RECT 249.395 -111.685 249.725 -111.355 ;
        RECT 249.395 -113.045 249.725 -112.715 ;
        RECT 249.395 -114.405 249.725 -114.075 ;
        RECT 249.395 -115.765 249.725 -115.435 ;
        RECT 249.395 -117.125 249.725 -116.795 ;
        RECT 249.395 -118.485 249.725 -118.155 ;
        RECT 249.395 -119.845 249.725 -119.515 ;
        RECT 249.395 -121.205 249.725 -120.875 ;
        RECT 249.395 -122.565 249.725 -122.235 ;
        RECT 249.395 -123.925 249.725 -123.595 ;
        RECT 249.395 -125.285 249.725 -124.955 ;
        RECT 249.395 -126.645 249.725 -126.315 ;
        RECT 249.395 -128.005 249.725 -127.675 ;
        RECT 249.395 -129.365 249.725 -129.035 ;
        RECT 249.395 -130.725 249.725 -130.395 ;
        RECT 249.395 -132.085 249.725 -131.755 ;
        RECT 249.395 -133.445 249.725 -133.115 ;
        RECT 249.395 -134.805 249.725 -134.475 ;
        RECT 249.395 -136.165 249.725 -135.835 ;
        RECT 249.395 -137.525 249.725 -137.195 ;
        RECT 249.395 -138.885 249.725 -138.555 ;
        RECT 249.395 -140.245 249.725 -139.915 ;
        RECT 249.395 -141.605 249.725 -141.275 ;
        RECT 249.395 -142.965 249.725 -142.635 ;
        RECT 249.395 -144.325 249.725 -143.995 ;
        RECT 249.395 -145.685 249.725 -145.355 ;
        RECT 249.395 -147.045 249.725 -146.715 ;
        RECT 249.395 -148.405 249.725 -148.075 ;
        RECT 249.395 -149.765 249.725 -149.435 ;
        RECT 249.395 -151.125 249.725 -150.795 ;
        RECT 249.395 -152.485 249.725 -152.155 ;
        RECT 249.395 -153.845 249.725 -153.515 ;
        RECT 249.395 -155.205 249.725 -154.875 ;
        RECT 249.395 -156.565 249.725 -156.235 ;
        RECT 249.395 -157.925 249.725 -157.595 ;
        RECT 249.395 -159.285 249.725 -158.955 ;
        RECT 249.395 -160.645 249.725 -160.315 ;
        RECT 249.395 -162.005 249.725 -161.675 ;
        RECT 249.395 -163.365 249.725 -163.035 ;
        RECT 249.395 -164.725 249.725 -164.395 ;
        RECT 249.395 -166.085 249.725 -165.755 ;
        RECT 249.395 -167.445 249.725 -167.115 ;
        RECT 249.395 -168.805 249.725 -168.475 ;
        RECT 249.395 -170.165 249.725 -169.835 ;
        RECT 249.395 -171.525 249.725 -171.195 ;
        RECT 249.395 -172.885 249.725 -172.555 ;
        RECT 249.395 -174.245 249.725 -173.915 ;
        RECT 249.395 -175.605 249.725 -175.275 ;
        RECT 249.395 -176.965 249.725 -176.635 ;
        RECT 249.395 -178.325 249.725 -177.995 ;
        RECT 249.395 -179.685 249.725 -179.355 ;
        RECT 249.395 -181.93 249.725 -180.8 ;
        RECT 249.4 -182.045 249.72 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.755 241.32 251.085 242.45 ;
        RECT 250.755 239.195 251.085 239.525 ;
        RECT 250.755 237.835 251.085 238.165 ;
        RECT 250.76 237.16 251.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.755 -1.525 251.085 -1.195 ;
        RECT 250.755 -2.885 251.085 -2.555 ;
        RECT 250.76 -3.56 251.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 250.755 -95.365 251.085 -95.035 ;
        RECT 250.755 -96.725 251.085 -96.395 ;
        RECT 250.755 -98.085 251.085 -97.755 ;
        RECT 250.755 -99.445 251.085 -99.115 ;
        RECT 250.755 -100.805 251.085 -100.475 ;
        RECT 250.755 -102.165 251.085 -101.835 ;
        RECT 250.755 -103.525 251.085 -103.195 ;
        RECT 250.755 -104.885 251.085 -104.555 ;
        RECT 250.755 -106.245 251.085 -105.915 ;
        RECT 250.755 -107.605 251.085 -107.275 ;
        RECT 250.755 -108.965 251.085 -108.635 ;
        RECT 250.755 -110.325 251.085 -109.995 ;
        RECT 250.755 -111.685 251.085 -111.355 ;
        RECT 250.755 -113.045 251.085 -112.715 ;
        RECT 250.755 -114.405 251.085 -114.075 ;
        RECT 250.755 -115.765 251.085 -115.435 ;
        RECT 250.755 -117.125 251.085 -116.795 ;
        RECT 250.755 -118.485 251.085 -118.155 ;
        RECT 250.755 -119.845 251.085 -119.515 ;
        RECT 250.755 -121.205 251.085 -120.875 ;
        RECT 250.755 -122.565 251.085 -122.235 ;
        RECT 250.755 -123.925 251.085 -123.595 ;
        RECT 250.755 -125.285 251.085 -124.955 ;
        RECT 250.755 -126.645 251.085 -126.315 ;
        RECT 250.755 -128.005 251.085 -127.675 ;
        RECT 250.755 -129.365 251.085 -129.035 ;
        RECT 250.755 -130.725 251.085 -130.395 ;
        RECT 250.755 -132.085 251.085 -131.755 ;
        RECT 250.755 -133.445 251.085 -133.115 ;
        RECT 250.755 -134.805 251.085 -134.475 ;
        RECT 250.755 -136.165 251.085 -135.835 ;
        RECT 250.755 -137.525 251.085 -137.195 ;
        RECT 250.755 -138.885 251.085 -138.555 ;
        RECT 250.755 -140.245 251.085 -139.915 ;
        RECT 250.755 -141.605 251.085 -141.275 ;
        RECT 250.755 -142.965 251.085 -142.635 ;
        RECT 250.755 -144.325 251.085 -143.995 ;
        RECT 250.755 -145.685 251.085 -145.355 ;
        RECT 250.755 -147.045 251.085 -146.715 ;
        RECT 250.755 -148.405 251.085 -148.075 ;
        RECT 250.755 -149.765 251.085 -149.435 ;
        RECT 250.755 -151.125 251.085 -150.795 ;
        RECT 250.755 -152.485 251.085 -152.155 ;
        RECT 250.755 -153.845 251.085 -153.515 ;
        RECT 250.755 -155.205 251.085 -154.875 ;
        RECT 250.755 -156.565 251.085 -156.235 ;
        RECT 250.755 -157.925 251.085 -157.595 ;
        RECT 250.755 -159.285 251.085 -158.955 ;
        RECT 250.755 -160.645 251.085 -160.315 ;
        RECT 250.755 -162.005 251.085 -161.675 ;
        RECT 250.755 -163.365 251.085 -163.035 ;
        RECT 250.755 -164.725 251.085 -164.395 ;
        RECT 250.755 -166.085 251.085 -165.755 ;
        RECT 250.755 -167.445 251.085 -167.115 ;
        RECT 250.755 -168.805 251.085 -168.475 ;
        RECT 250.755 -170.165 251.085 -169.835 ;
        RECT 250.755 -171.525 251.085 -171.195 ;
        RECT 250.755 -172.885 251.085 -172.555 ;
        RECT 250.755 -174.245 251.085 -173.915 ;
        RECT 250.755 -175.605 251.085 -175.275 ;
        RECT 250.755 -176.965 251.085 -176.635 ;
        RECT 250.755 -178.325 251.085 -177.995 ;
        RECT 250.755 -179.685 251.085 -179.355 ;
        RECT 250.755 -181.93 251.085 -180.8 ;
        RECT 250.76 -182.045 251.08 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.115 241.32 252.445 242.45 ;
        RECT 252.115 239.195 252.445 239.525 ;
        RECT 252.115 237.835 252.445 238.165 ;
        RECT 252.12 237.16 252.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.115 -1.525 252.445 -1.195 ;
        RECT 252.115 -2.885 252.445 -2.555 ;
        RECT 252.12 -3.56 252.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 252.115 -95.365 252.445 -95.035 ;
        RECT 252.115 -96.725 252.445 -96.395 ;
        RECT 252.115 -98.085 252.445 -97.755 ;
        RECT 252.115 -99.445 252.445 -99.115 ;
        RECT 252.115 -100.805 252.445 -100.475 ;
        RECT 252.115 -102.165 252.445 -101.835 ;
        RECT 252.115 -103.525 252.445 -103.195 ;
        RECT 252.115 -104.885 252.445 -104.555 ;
        RECT 252.115 -106.245 252.445 -105.915 ;
        RECT 252.115 -107.605 252.445 -107.275 ;
        RECT 252.115 -108.965 252.445 -108.635 ;
        RECT 252.115 -110.325 252.445 -109.995 ;
        RECT 252.115 -111.685 252.445 -111.355 ;
        RECT 252.115 -113.045 252.445 -112.715 ;
        RECT 252.115 -114.405 252.445 -114.075 ;
        RECT 252.115 -115.765 252.445 -115.435 ;
        RECT 252.115 -117.125 252.445 -116.795 ;
        RECT 252.115 -118.485 252.445 -118.155 ;
        RECT 252.115 -119.845 252.445 -119.515 ;
        RECT 252.115 -121.205 252.445 -120.875 ;
        RECT 252.115 -122.565 252.445 -122.235 ;
        RECT 252.115 -123.925 252.445 -123.595 ;
        RECT 252.115 -125.285 252.445 -124.955 ;
        RECT 252.115 -126.645 252.445 -126.315 ;
        RECT 252.115 -128.005 252.445 -127.675 ;
        RECT 252.115 -129.365 252.445 -129.035 ;
        RECT 252.115 -130.725 252.445 -130.395 ;
        RECT 252.115 -132.085 252.445 -131.755 ;
        RECT 252.115 -133.445 252.445 -133.115 ;
        RECT 252.115 -134.805 252.445 -134.475 ;
        RECT 252.115 -136.165 252.445 -135.835 ;
        RECT 252.115 -137.525 252.445 -137.195 ;
        RECT 252.115 -138.885 252.445 -138.555 ;
        RECT 252.115 -140.245 252.445 -139.915 ;
        RECT 252.115 -141.605 252.445 -141.275 ;
        RECT 252.115 -142.965 252.445 -142.635 ;
        RECT 252.115 -144.325 252.445 -143.995 ;
        RECT 252.115 -145.685 252.445 -145.355 ;
        RECT 252.115 -147.045 252.445 -146.715 ;
        RECT 252.115 -148.405 252.445 -148.075 ;
        RECT 252.115 -149.765 252.445 -149.435 ;
        RECT 252.115 -151.125 252.445 -150.795 ;
        RECT 252.115 -152.485 252.445 -152.155 ;
        RECT 252.115 -153.845 252.445 -153.515 ;
        RECT 252.115 -155.205 252.445 -154.875 ;
        RECT 252.115 -156.565 252.445 -156.235 ;
        RECT 252.115 -157.925 252.445 -157.595 ;
        RECT 252.115 -159.285 252.445 -158.955 ;
        RECT 252.115 -160.645 252.445 -160.315 ;
        RECT 252.115 -162.005 252.445 -161.675 ;
        RECT 252.115 -163.365 252.445 -163.035 ;
        RECT 252.115 -164.725 252.445 -164.395 ;
        RECT 252.115 -166.085 252.445 -165.755 ;
        RECT 252.115 -167.445 252.445 -167.115 ;
        RECT 252.115 -168.805 252.445 -168.475 ;
        RECT 252.115 -170.165 252.445 -169.835 ;
        RECT 252.115 -171.525 252.445 -171.195 ;
        RECT 252.115 -172.885 252.445 -172.555 ;
        RECT 252.115 -174.245 252.445 -173.915 ;
        RECT 252.115 -175.605 252.445 -175.275 ;
        RECT 252.115 -176.965 252.445 -176.635 ;
        RECT 252.115 -178.325 252.445 -177.995 ;
        RECT 252.115 -179.685 252.445 -179.355 ;
        RECT 252.115 -181.93 252.445 -180.8 ;
        RECT 252.12 -182.045 252.44 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.475 241.32 253.805 242.45 ;
        RECT 253.475 239.195 253.805 239.525 ;
        RECT 253.475 237.835 253.805 238.165 ;
        RECT 253.48 237.16 253.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 253.475 -99.445 253.805 -99.115 ;
        RECT 253.475 -100.805 253.805 -100.475 ;
        RECT 253.475 -102.165 253.805 -101.835 ;
        RECT 253.475 -103.525 253.805 -103.195 ;
        RECT 253.475 -104.885 253.805 -104.555 ;
        RECT 253.475 -106.245 253.805 -105.915 ;
        RECT 253.475 -107.605 253.805 -107.275 ;
        RECT 253.475 -108.965 253.805 -108.635 ;
        RECT 253.475 -110.325 253.805 -109.995 ;
        RECT 253.475 -111.685 253.805 -111.355 ;
        RECT 253.475 -113.045 253.805 -112.715 ;
        RECT 253.475 -114.405 253.805 -114.075 ;
        RECT 253.475 -115.765 253.805 -115.435 ;
        RECT 253.475 -117.125 253.805 -116.795 ;
        RECT 253.475 -118.485 253.805 -118.155 ;
        RECT 253.475 -119.845 253.805 -119.515 ;
        RECT 253.475 -121.205 253.805 -120.875 ;
        RECT 253.475 -122.565 253.805 -122.235 ;
        RECT 253.475 -123.925 253.805 -123.595 ;
        RECT 253.475 -125.285 253.805 -124.955 ;
        RECT 253.475 -126.645 253.805 -126.315 ;
        RECT 253.475 -128.005 253.805 -127.675 ;
        RECT 253.475 -129.365 253.805 -129.035 ;
        RECT 253.475 -130.725 253.805 -130.395 ;
        RECT 253.475 -132.085 253.805 -131.755 ;
        RECT 253.475 -133.445 253.805 -133.115 ;
        RECT 253.475 -134.805 253.805 -134.475 ;
        RECT 253.475 -136.165 253.805 -135.835 ;
        RECT 253.475 -137.525 253.805 -137.195 ;
        RECT 253.475 -138.885 253.805 -138.555 ;
        RECT 253.475 -140.245 253.805 -139.915 ;
        RECT 253.475 -141.605 253.805 -141.275 ;
        RECT 253.475 -142.965 253.805 -142.635 ;
        RECT 253.475 -144.325 253.805 -143.995 ;
        RECT 253.475 -145.685 253.805 -145.355 ;
        RECT 253.475 -147.045 253.805 -146.715 ;
        RECT 253.475 -148.405 253.805 -148.075 ;
        RECT 253.475 -149.765 253.805 -149.435 ;
        RECT 253.475 -151.125 253.805 -150.795 ;
        RECT 253.475 -152.485 253.805 -152.155 ;
        RECT 253.475 -153.845 253.805 -153.515 ;
        RECT 253.475 -155.205 253.805 -154.875 ;
        RECT 253.475 -156.565 253.805 -156.235 ;
        RECT 253.475 -157.925 253.805 -157.595 ;
        RECT 253.475 -159.285 253.805 -158.955 ;
        RECT 253.475 -160.645 253.805 -160.315 ;
        RECT 253.475 -162.005 253.805 -161.675 ;
        RECT 253.475 -163.365 253.805 -163.035 ;
        RECT 253.475 -164.725 253.805 -164.395 ;
        RECT 253.475 -166.085 253.805 -165.755 ;
        RECT 253.475 -167.445 253.805 -167.115 ;
        RECT 253.475 -168.805 253.805 -168.475 ;
        RECT 253.475 -170.165 253.805 -169.835 ;
        RECT 253.475 -171.525 253.805 -171.195 ;
        RECT 253.475 -172.885 253.805 -172.555 ;
        RECT 253.475 -174.245 253.805 -173.915 ;
        RECT 253.475 -175.605 253.805 -175.275 ;
        RECT 253.475 -176.965 253.805 -176.635 ;
        RECT 253.475 -178.325 253.805 -177.995 ;
        RECT 253.475 -179.685 253.805 -179.355 ;
        RECT 253.475 -181.93 253.805 -180.8 ;
        RECT 253.48 -182.045 253.8 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.01 -98.075 254.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.835 241.32 255.165 242.45 ;
        RECT 254.835 239.195 255.165 239.525 ;
        RECT 254.835 237.835 255.165 238.165 ;
        RECT 254.84 237.16 255.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 254.835 -1.525 255.165 -1.195 ;
        RECT 254.835 -2.885 255.165 -2.555 ;
        RECT 254.84 -3.56 255.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.195 241.32 256.525 242.45 ;
        RECT 256.195 239.195 256.525 239.525 ;
        RECT 256.195 237.835 256.525 238.165 ;
        RECT 256.2 237.16 256.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 256.195 -1.525 256.525 -1.195 ;
        RECT 256.195 -2.885 256.525 -2.555 ;
        RECT 256.2 -3.56 256.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.555 241.32 257.885 242.45 ;
        RECT 257.555 239.195 257.885 239.525 ;
        RECT 257.555 237.835 257.885 238.165 ;
        RECT 257.56 237.16 257.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.555 -1.525 257.885 -1.195 ;
        RECT 257.555 -2.885 257.885 -2.555 ;
        RECT 257.56 -3.56 257.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 257.555 -95.365 257.885 -95.035 ;
        RECT 257.555 -96.725 257.885 -96.395 ;
        RECT 257.555 -98.085 257.885 -97.755 ;
        RECT 257.555 -99.445 257.885 -99.115 ;
        RECT 257.555 -100.805 257.885 -100.475 ;
        RECT 257.555 -102.165 257.885 -101.835 ;
        RECT 257.555 -103.525 257.885 -103.195 ;
        RECT 257.555 -104.885 257.885 -104.555 ;
        RECT 257.555 -106.245 257.885 -105.915 ;
        RECT 257.555 -107.605 257.885 -107.275 ;
        RECT 257.555 -108.965 257.885 -108.635 ;
        RECT 257.555 -110.325 257.885 -109.995 ;
        RECT 257.555 -111.685 257.885 -111.355 ;
        RECT 257.555 -113.045 257.885 -112.715 ;
        RECT 257.555 -114.405 257.885 -114.075 ;
        RECT 257.555 -115.765 257.885 -115.435 ;
        RECT 257.555 -117.125 257.885 -116.795 ;
        RECT 257.555 -118.485 257.885 -118.155 ;
        RECT 257.555 -119.845 257.885 -119.515 ;
        RECT 257.555 -121.205 257.885 -120.875 ;
        RECT 257.555 -122.565 257.885 -122.235 ;
        RECT 257.555 -123.925 257.885 -123.595 ;
        RECT 257.555 -125.285 257.885 -124.955 ;
        RECT 257.555 -126.645 257.885 -126.315 ;
        RECT 257.555 -128.005 257.885 -127.675 ;
        RECT 257.555 -129.365 257.885 -129.035 ;
        RECT 257.555 -130.725 257.885 -130.395 ;
        RECT 257.555 -132.085 257.885 -131.755 ;
        RECT 257.555 -133.445 257.885 -133.115 ;
        RECT 257.555 -134.805 257.885 -134.475 ;
        RECT 257.555 -136.165 257.885 -135.835 ;
        RECT 257.555 -137.525 257.885 -137.195 ;
        RECT 257.555 -138.885 257.885 -138.555 ;
        RECT 257.555 -140.245 257.885 -139.915 ;
        RECT 257.555 -141.605 257.885 -141.275 ;
        RECT 257.555 -142.965 257.885 -142.635 ;
        RECT 257.555 -144.325 257.885 -143.995 ;
        RECT 257.555 -145.685 257.885 -145.355 ;
        RECT 257.555 -147.045 257.885 -146.715 ;
        RECT 257.555 -148.405 257.885 -148.075 ;
        RECT 257.555 -149.765 257.885 -149.435 ;
        RECT 257.555 -151.125 257.885 -150.795 ;
        RECT 257.555 -152.485 257.885 -152.155 ;
        RECT 257.555 -153.845 257.885 -153.515 ;
        RECT 257.555 -155.205 257.885 -154.875 ;
        RECT 257.555 -156.565 257.885 -156.235 ;
        RECT 257.555 -157.925 257.885 -157.595 ;
        RECT 257.555 -159.285 257.885 -158.955 ;
        RECT 257.555 -160.645 257.885 -160.315 ;
        RECT 257.555 -162.005 257.885 -161.675 ;
        RECT 257.555 -163.365 257.885 -163.035 ;
        RECT 257.555 -164.725 257.885 -164.395 ;
        RECT 257.555 -166.085 257.885 -165.755 ;
        RECT 257.555 -167.445 257.885 -167.115 ;
        RECT 257.555 -168.805 257.885 -168.475 ;
        RECT 257.555 -170.165 257.885 -169.835 ;
        RECT 257.555 -171.525 257.885 -171.195 ;
        RECT 257.555 -172.885 257.885 -172.555 ;
        RECT 257.555 -174.245 257.885 -173.915 ;
        RECT 257.555 -175.605 257.885 -175.275 ;
        RECT 257.555 -176.965 257.885 -176.635 ;
        RECT 257.555 -178.325 257.885 -177.995 ;
        RECT 257.555 -179.685 257.885 -179.355 ;
        RECT 257.555 -181.93 257.885 -180.8 ;
        RECT 257.56 -182.045 257.88 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.915 241.32 259.245 242.45 ;
        RECT 258.915 239.195 259.245 239.525 ;
        RECT 258.915 237.835 259.245 238.165 ;
        RECT 258.92 237.16 259.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.915 -1.525 259.245 -1.195 ;
        RECT 258.915 -2.885 259.245 -2.555 ;
        RECT 258.92 -3.56 259.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 258.915 -95.365 259.245 -95.035 ;
        RECT 258.915 -96.725 259.245 -96.395 ;
        RECT 258.915 -98.085 259.245 -97.755 ;
        RECT 258.915 -99.445 259.245 -99.115 ;
        RECT 258.915 -100.805 259.245 -100.475 ;
        RECT 258.915 -102.165 259.245 -101.835 ;
        RECT 258.915 -103.525 259.245 -103.195 ;
        RECT 258.915 -104.885 259.245 -104.555 ;
        RECT 258.915 -106.245 259.245 -105.915 ;
        RECT 258.915 -107.605 259.245 -107.275 ;
        RECT 258.915 -108.965 259.245 -108.635 ;
        RECT 258.915 -110.325 259.245 -109.995 ;
        RECT 258.915 -111.685 259.245 -111.355 ;
        RECT 258.915 -113.045 259.245 -112.715 ;
        RECT 258.915 -114.405 259.245 -114.075 ;
        RECT 258.915 -115.765 259.245 -115.435 ;
        RECT 258.915 -117.125 259.245 -116.795 ;
        RECT 258.915 -118.485 259.245 -118.155 ;
        RECT 258.915 -119.845 259.245 -119.515 ;
        RECT 258.915 -121.205 259.245 -120.875 ;
        RECT 258.915 -122.565 259.245 -122.235 ;
        RECT 258.915 -123.925 259.245 -123.595 ;
        RECT 258.915 -125.285 259.245 -124.955 ;
        RECT 258.915 -126.645 259.245 -126.315 ;
        RECT 258.915 -128.005 259.245 -127.675 ;
        RECT 258.915 -129.365 259.245 -129.035 ;
        RECT 258.915 -130.725 259.245 -130.395 ;
        RECT 258.915 -132.085 259.245 -131.755 ;
        RECT 258.915 -133.445 259.245 -133.115 ;
        RECT 258.915 -134.805 259.245 -134.475 ;
        RECT 258.915 -136.165 259.245 -135.835 ;
        RECT 258.915 -137.525 259.245 -137.195 ;
        RECT 258.915 -138.885 259.245 -138.555 ;
        RECT 258.915 -140.245 259.245 -139.915 ;
        RECT 258.915 -141.605 259.245 -141.275 ;
        RECT 258.915 -142.965 259.245 -142.635 ;
        RECT 258.915 -144.325 259.245 -143.995 ;
        RECT 258.915 -145.685 259.245 -145.355 ;
        RECT 258.915 -147.045 259.245 -146.715 ;
        RECT 258.915 -148.405 259.245 -148.075 ;
        RECT 258.915 -149.765 259.245 -149.435 ;
        RECT 258.915 -151.125 259.245 -150.795 ;
        RECT 258.915 -152.485 259.245 -152.155 ;
        RECT 258.915 -153.845 259.245 -153.515 ;
        RECT 258.915 -155.205 259.245 -154.875 ;
        RECT 258.915 -156.565 259.245 -156.235 ;
        RECT 258.915 -157.925 259.245 -157.595 ;
        RECT 258.915 -159.285 259.245 -158.955 ;
        RECT 258.915 -160.645 259.245 -160.315 ;
        RECT 258.915 -162.005 259.245 -161.675 ;
        RECT 258.915 -163.365 259.245 -163.035 ;
        RECT 258.915 -164.725 259.245 -164.395 ;
        RECT 258.915 -166.085 259.245 -165.755 ;
        RECT 258.915 -167.445 259.245 -167.115 ;
        RECT 258.915 -168.805 259.245 -168.475 ;
        RECT 258.915 -170.165 259.245 -169.835 ;
        RECT 258.915 -171.525 259.245 -171.195 ;
        RECT 258.915 -172.885 259.245 -172.555 ;
        RECT 258.915 -174.245 259.245 -173.915 ;
        RECT 258.915 -175.605 259.245 -175.275 ;
        RECT 258.915 -176.965 259.245 -176.635 ;
        RECT 258.915 -178.325 259.245 -177.995 ;
        RECT 258.915 -179.685 259.245 -179.355 ;
        RECT 258.915 -181.93 259.245 -180.8 ;
        RECT 258.92 -182.045 259.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.275 241.32 260.605 242.45 ;
        RECT 260.275 239.195 260.605 239.525 ;
        RECT 260.275 237.835 260.605 238.165 ;
        RECT 260.28 237.16 260.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.275 -1.525 260.605 -1.195 ;
        RECT 260.275 -2.885 260.605 -2.555 ;
        RECT 260.28 -3.56 260.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 260.275 -95.365 260.605 -95.035 ;
        RECT 260.275 -96.725 260.605 -96.395 ;
        RECT 260.275 -98.085 260.605 -97.755 ;
        RECT 260.275 -99.445 260.605 -99.115 ;
        RECT 260.275 -100.805 260.605 -100.475 ;
        RECT 260.275 -102.165 260.605 -101.835 ;
        RECT 260.275 -103.525 260.605 -103.195 ;
        RECT 260.275 -104.885 260.605 -104.555 ;
        RECT 260.275 -106.245 260.605 -105.915 ;
        RECT 260.275 -107.605 260.605 -107.275 ;
        RECT 260.275 -108.965 260.605 -108.635 ;
        RECT 260.275 -110.325 260.605 -109.995 ;
        RECT 260.275 -111.685 260.605 -111.355 ;
        RECT 260.275 -113.045 260.605 -112.715 ;
        RECT 260.275 -114.405 260.605 -114.075 ;
        RECT 260.275 -115.765 260.605 -115.435 ;
        RECT 260.275 -117.125 260.605 -116.795 ;
        RECT 260.275 -118.485 260.605 -118.155 ;
        RECT 260.275 -119.845 260.605 -119.515 ;
        RECT 260.275 -121.205 260.605 -120.875 ;
        RECT 260.275 -122.565 260.605 -122.235 ;
        RECT 260.275 -123.925 260.605 -123.595 ;
        RECT 260.275 -125.285 260.605 -124.955 ;
        RECT 260.275 -126.645 260.605 -126.315 ;
        RECT 260.275 -128.005 260.605 -127.675 ;
        RECT 260.275 -129.365 260.605 -129.035 ;
        RECT 260.275 -130.725 260.605 -130.395 ;
        RECT 260.275 -132.085 260.605 -131.755 ;
        RECT 260.275 -133.445 260.605 -133.115 ;
        RECT 260.275 -134.805 260.605 -134.475 ;
        RECT 260.275 -136.165 260.605 -135.835 ;
        RECT 260.275 -137.525 260.605 -137.195 ;
        RECT 260.275 -138.885 260.605 -138.555 ;
        RECT 260.275 -140.245 260.605 -139.915 ;
        RECT 260.275 -141.605 260.605 -141.275 ;
        RECT 260.275 -142.965 260.605 -142.635 ;
        RECT 260.275 -144.325 260.605 -143.995 ;
        RECT 260.275 -145.685 260.605 -145.355 ;
        RECT 260.275 -147.045 260.605 -146.715 ;
        RECT 260.275 -148.405 260.605 -148.075 ;
        RECT 260.275 -149.765 260.605 -149.435 ;
        RECT 260.275 -151.125 260.605 -150.795 ;
        RECT 260.275 -152.485 260.605 -152.155 ;
        RECT 260.275 -153.845 260.605 -153.515 ;
        RECT 260.275 -155.205 260.605 -154.875 ;
        RECT 260.275 -156.565 260.605 -156.235 ;
        RECT 260.275 -157.925 260.605 -157.595 ;
        RECT 260.275 -159.285 260.605 -158.955 ;
        RECT 260.275 -160.645 260.605 -160.315 ;
        RECT 260.275 -162.005 260.605 -161.675 ;
        RECT 260.275 -163.365 260.605 -163.035 ;
        RECT 260.275 -164.725 260.605 -164.395 ;
        RECT 260.275 -166.085 260.605 -165.755 ;
        RECT 260.275 -167.445 260.605 -167.115 ;
        RECT 260.275 -168.805 260.605 -168.475 ;
        RECT 260.275 -170.165 260.605 -169.835 ;
        RECT 260.275 -171.525 260.605 -171.195 ;
        RECT 260.275 -172.885 260.605 -172.555 ;
        RECT 260.275 -174.245 260.605 -173.915 ;
        RECT 260.275 -175.605 260.605 -175.275 ;
        RECT 260.275 -176.965 260.605 -176.635 ;
        RECT 260.275 -178.325 260.605 -177.995 ;
        RECT 260.275 -179.685 260.605 -179.355 ;
        RECT 260.275 -181.93 260.605 -180.8 ;
        RECT 260.28 -182.045 260.6 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.635 241.32 261.965 242.45 ;
        RECT 261.635 239.195 261.965 239.525 ;
        RECT 261.635 237.835 261.965 238.165 ;
        RECT 261.64 237.16 261.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.635 -1.525 261.965 -1.195 ;
        RECT 261.635 -2.885 261.965 -2.555 ;
        RECT 261.64 -3.56 261.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 261.635 -95.365 261.965 -95.035 ;
        RECT 261.635 -96.725 261.965 -96.395 ;
        RECT 261.635 -98.085 261.965 -97.755 ;
        RECT 261.635 -99.445 261.965 -99.115 ;
        RECT 261.635 -100.805 261.965 -100.475 ;
        RECT 261.635 -102.165 261.965 -101.835 ;
        RECT 261.635 -103.525 261.965 -103.195 ;
        RECT 261.635 -104.885 261.965 -104.555 ;
        RECT 261.635 -106.245 261.965 -105.915 ;
        RECT 261.635 -107.605 261.965 -107.275 ;
        RECT 261.635 -108.965 261.965 -108.635 ;
        RECT 261.635 -110.325 261.965 -109.995 ;
        RECT 261.635 -111.685 261.965 -111.355 ;
        RECT 261.635 -113.045 261.965 -112.715 ;
        RECT 261.635 -114.405 261.965 -114.075 ;
        RECT 261.635 -115.765 261.965 -115.435 ;
        RECT 261.635 -117.125 261.965 -116.795 ;
        RECT 261.635 -118.485 261.965 -118.155 ;
        RECT 261.635 -119.845 261.965 -119.515 ;
        RECT 261.635 -121.205 261.965 -120.875 ;
        RECT 261.635 -122.565 261.965 -122.235 ;
        RECT 261.635 -123.925 261.965 -123.595 ;
        RECT 261.635 -125.285 261.965 -124.955 ;
        RECT 261.635 -126.645 261.965 -126.315 ;
        RECT 261.635 -128.005 261.965 -127.675 ;
        RECT 261.635 -129.365 261.965 -129.035 ;
        RECT 261.635 -130.725 261.965 -130.395 ;
        RECT 261.635 -132.085 261.965 -131.755 ;
        RECT 261.635 -133.445 261.965 -133.115 ;
        RECT 261.635 -134.805 261.965 -134.475 ;
        RECT 261.635 -136.165 261.965 -135.835 ;
        RECT 261.635 -137.525 261.965 -137.195 ;
        RECT 261.635 -138.885 261.965 -138.555 ;
        RECT 261.635 -140.245 261.965 -139.915 ;
        RECT 261.635 -141.605 261.965 -141.275 ;
        RECT 261.635 -142.965 261.965 -142.635 ;
        RECT 261.635 -144.325 261.965 -143.995 ;
        RECT 261.635 -145.685 261.965 -145.355 ;
        RECT 261.635 -147.045 261.965 -146.715 ;
        RECT 261.635 -148.405 261.965 -148.075 ;
        RECT 261.635 -149.765 261.965 -149.435 ;
        RECT 261.635 -151.125 261.965 -150.795 ;
        RECT 261.635 -152.485 261.965 -152.155 ;
        RECT 261.635 -153.845 261.965 -153.515 ;
        RECT 261.635 -155.205 261.965 -154.875 ;
        RECT 261.635 -156.565 261.965 -156.235 ;
        RECT 261.635 -157.925 261.965 -157.595 ;
        RECT 261.635 -159.285 261.965 -158.955 ;
        RECT 261.635 -160.645 261.965 -160.315 ;
        RECT 261.635 -162.005 261.965 -161.675 ;
        RECT 261.635 -163.365 261.965 -163.035 ;
        RECT 261.635 -164.725 261.965 -164.395 ;
        RECT 261.635 -166.085 261.965 -165.755 ;
        RECT 261.635 -167.445 261.965 -167.115 ;
        RECT 261.635 -168.805 261.965 -168.475 ;
        RECT 261.635 -170.165 261.965 -169.835 ;
        RECT 261.635 -171.525 261.965 -171.195 ;
        RECT 261.635 -172.885 261.965 -172.555 ;
        RECT 261.635 -174.245 261.965 -173.915 ;
        RECT 261.635 -175.605 261.965 -175.275 ;
        RECT 261.635 -176.965 261.965 -176.635 ;
        RECT 261.635 -178.325 261.965 -177.995 ;
        RECT 261.635 -179.685 261.965 -179.355 ;
        RECT 261.635 -181.93 261.965 -180.8 ;
        RECT 261.64 -182.045 261.96 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.995 241.32 263.325 242.45 ;
        RECT 262.995 239.195 263.325 239.525 ;
        RECT 262.995 237.835 263.325 238.165 ;
        RECT 263 237.16 263.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.995 -1.525 263.325 -1.195 ;
        RECT 262.995 -2.885 263.325 -2.555 ;
        RECT 263 -3.56 263.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 262.995 -95.365 263.325 -95.035 ;
        RECT 262.995 -96.725 263.325 -96.395 ;
        RECT 262.995 -98.085 263.325 -97.755 ;
        RECT 262.995 -99.445 263.325 -99.115 ;
        RECT 262.995 -100.805 263.325 -100.475 ;
        RECT 262.995 -102.165 263.325 -101.835 ;
        RECT 262.995 -103.525 263.325 -103.195 ;
        RECT 262.995 -104.885 263.325 -104.555 ;
        RECT 262.995 -106.245 263.325 -105.915 ;
        RECT 262.995 -107.605 263.325 -107.275 ;
        RECT 262.995 -108.965 263.325 -108.635 ;
        RECT 262.995 -110.325 263.325 -109.995 ;
        RECT 262.995 -111.685 263.325 -111.355 ;
        RECT 262.995 -113.045 263.325 -112.715 ;
        RECT 262.995 -114.405 263.325 -114.075 ;
        RECT 262.995 -115.765 263.325 -115.435 ;
        RECT 262.995 -117.125 263.325 -116.795 ;
        RECT 262.995 -118.485 263.325 -118.155 ;
        RECT 262.995 -119.845 263.325 -119.515 ;
        RECT 262.995 -121.205 263.325 -120.875 ;
        RECT 262.995 -122.565 263.325 -122.235 ;
        RECT 262.995 -123.925 263.325 -123.595 ;
        RECT 262.995 -125.285 263.325 -124.955 ;
        RECT 262.995 -126.645 263.325 -126.315 ;
        RECT 262.995 -128.005 263.325 -127.675 ;
        RECT 262.995 -129.365 263.325 -129.035 ;
        RECT 262.995 -130.725 263.325 -130.395 ;
        RECT 262.995 -132.085 263.325 -131.755 ;
        RECT 262.995 -133.445 263.325 -133.115 ;
        RECT 262.995 -134.805 263.325 -134.475 ;
        RECT 262.995 -136.165 263.325 -135.835 ;
        RECT 262.995 -137.525 263.325 -137.195 ;
        RECT 262.995 -138.885 263.325 -138.555 ;
        RECT 262.995 -140.245 263.325 -139.915 ;
        RECT 262.995 -141.605 263.325 -141.275 ;
        RECT 262.995 -142.965 263.325 -142.635 ;
        RECT 262.995 -144.325 263.325 -143.995 ;
        RECT 262.995 -145.685 263.325 -145.355 ;
        RECT 262.995 -147.045 263.325 -146.715 ;
        RECT 262.995 -148.405 263.325 -148.075 ;
        RECT 262.995 -149.765 263.325 -149.435 ;
        RECT 262.995 -151.125 263.325 -150.795 ;
        RECT 262.995 -152.485 263.325 -152.155 ;
        RECT 262.995 -153.845 263.325 -153.515 ;
        RECT 262.995 -155.205 263.325 -154.875 ;
        RECT 262.995 -156.565 263.325 -156.235 ;
        RECT 262.995 -157.925 263.325 -157.595 ;
        RECT 262.995 -159.285 263.325 -158.955 ;
        RECT 262.995 -160.645 263.325 -160.315 ;
        RECT 262.995 -162.005 263.325 -161.675 ;
        RECT 262.995 -163.365 263.325 -163.035 ;
        RECT 262.995 -164.725 263.325 -164.395 ;
        RECT 262.995 -166.085 263.325 -165.755 ;
        RECT 262.995 -167.445 263.325 -167.115 ;
        RECT 262.995 -168.805 263.325 -168.475 ;
        RECT 262.995 -170.165 263.325 -169.835 ;
        RECT 262.995 -171.525 263.325 -171.195 ;
        RECT 262.995 -172.885 263.325 -172.555 ;
        RECT 262.995 -174.245 263.325 -173.915 ;
        RECT 262.995 -175.605 263.325 -175.275 ;
        RECT 262.995 -176.965 263.325 -176.635 ;
        RECT 262.995 -178.325 263.325 -177.995 ;
        RECT 262.995 -179.685 263.325 -179.355 ;
        RECT 262.995 -181.93 263.325 -180.8 ;
        RECT 263 -182.045 263.32 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.355 241.32 264.685 242.45 ;
        RECT 264.355 239.195 264.685 239.525 ;
        RECT 264.355 237.835 264.685 238.165 ;
        RECT 264.36 237.16 264.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 264.355 -174.245 264.685 -173.915 ;
        RECT 264.355 -175.605 264.685 -175.275 ;
        RECT 264.355 -176.965 264.685 -176.635 ;
        RECT 264.355 -178.325 264.685 -177.995 ;
        RECT 264.355 -179.685 264.685 -179.355 ;
        RECT 264.355 -181.93 264.685 -180.8 ;
        RECT 264.36 -182.045 264.68 -98.44 ;
        RECT 264.355 -99.445 264.685 -99.115 ;
        RECT 264.355 -100.805 264.685 -100.475 ;
        RECT 264.355 -102.165 264.685 -101.835 ;
        RECT 264.355 -103.525 264.685 -103.195 ;
        RECT 264.355 -104.885 264.685 -104.555 ;
        RECT 264.355 -106.245 264.685 -105.915 ;
        RECT 264.355 -107.605 264.685 -107.275 ;
        RECT 264.355 -108.965 264.685 -108.635 ;
        RECT 264.355 -110.325 264.685 -109.995 ;
        RECT 264.355 -111.685 264.685 -111.355 ;
        RECT 264.355 -113.045 264.685 -112.715 ;
        RECT 264.355 -114.405 264.685 -114.075 ;
        RECT 264.355 -115.765 264.685 -115.435 ;
        RECT 264.355 -117.125 264.685 -116.795 ;
        RECT 264.355 -118.485 264.685 -118.155 ;
        RECT 264.355 -119.845 264.685 -119.515 ;
        RECT 264.355 -121.205 264.685 -120.875 ;
        RECT 264.355 -122.565 264.685 -122.235 ;
        RECT 264.355 -123.925 264.685 -123.595 ;
        RECT 264.355 -125.285 264.685 -124.955 ;
        RECT 264.355 -126.645 264.685 -126.315 ;
        RECT 264.355 -128.005 264.685 -127.675 ;
        RECT 264.355 -129.365 264.685 -129.035 ;
        RECT 264.355 -130.725 264.685 -130.395 ;
        RECT 264.355 -132.085 264.685 -131.755 ;
        RECT 264.355 -133.445 264.685 -133.115 ;
        RECT 264.355 -134.805 264.685 -134.475 ;
        RECT 264.355 -136.165 264.685 -135.835 ;
        RECT 264.355 -137.525 264.685 -137.195 ;
        RECT 264.355 -138.885 264.685 -138.555 ;
        RECT 264.355 -140.245 264.685 -139.915 ;
        RECT 264.355 -141.605 264.685 -141.275 ;
        RECT 264.355 -142.965 264.685 -142.635 ;
        RECT 264.355 -144.325 264.685 -143.995 ;
        RECT 264.355 -145.685 264.685 -145.355 ;
        RECT 264.355 -147.045 264.685 -146.715 ;
        RECT 264.355 -148.405 264.685 -148.075 ;
        RECT 264.355 -149.765 264.685 -149.435 ;
        RECT 264.355 -151.125 264.685 -150.795 ;
        RECT 264.355 -152.485 264.685 -152.155 ;
        RECT 264.355 -153.845 264.685 -153.515 ;
        RECT 264.355 -155.205 264.685 -154.875 ;
        RECT 264.355 -156.565 264.685 -156.235 ;
        RECT 264.355 -157.925 264.685 -157.595 ;
        RECT 264.355 -159.285 264.685 -158.955 ;
        RECT 264.355 -160.645 264.685 -160.315 ;
        RECT 264.355 -162.005 264.685 -161.675 ;
        RECT 264.355 -163.365 264.685 -163.035 ;
        RECT 264.355 -164.725 264.685 -164.395 ;
        RECT 264.355 -166.085 264.685 -165.755 ;
        RECT 264.355 -167.445 264.685 -167.115 ;
        RECT 264.355 -168.805 264.685 -168.475 ;
        RECT 264.355 -170.165 264.685 -169.835 ;
        RECT 264.355 -171.525 264.685 -171.195 ;
        RECT 264.355 -172.885 264.685 -172.555 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.755 241.32 217.085 242.45 ;
        RECT 216.755 239.195 217.085 239.525 ;
        RECT 216.755 237.835 217.085 238.165 ;
        RECT 216.76 237.16 217.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.755 -1.525 217.085 -1.195 ;
        RECT 216.755 -2.885 217.085 -2.555 ;
        RECT 216.76 -3.56 217.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 216.755 -95.365 217.085 -95.035 ;
        RECT 216.755 -96.725 217.085 -96.395 ;
        RECT 216.755 -98.085 217.085 -97.755 ;
        RECT 216.755 -99.445 217.085 -99.115 ;
        RECT 216.755 -100.805 217.085 -100.475 ;
        RECT 216.755 -102.165 217.085 -101.835 ;
        RECT 216.755 -103.525 217.085 -103.195 ;
        RECT 216.755 -104.885 217.085 -104.555 ;
        RECT 216.755 -106.245 217.085 -105.915 ;
        RECT 216.755 -107.605 217.085 -107.275 ;
        RECT 216.755 -108.965 217.085 -108.635 ;
        RECT 216.755 -110.325 217.085 -109.995 ;
        RECT 216.755 -111.685 217.085 -111.355 ;
        RECT 216.755 -113.045 217.085 -112.715 ;
        RECT 216.755 -114.405 217.085 -114.075 ;
        RECT 216.755 -115.765 217.085 -115.435 ;
        RECT 216.755 -117.125 217.085 -116.795 ;
        RECT 216.755 -118.485 217.085 -118.155 ;
        RECT 216.755 -119.845 217.085 -119.515 ;
        RECT 216.755 -121.205 217.085 -120.875 ;
        RECT 216.755 -122.565 217.085 -122.235 ;
        RECT 216.755 -123.925 217.085 -123.595 ;
        RECT 216.755 -125.285 217.085 -124.955 ;
        RECT 216.755 -126.645 217.085 -126.315 ;
        RECT 216.755 -128.005 217.085 -127.675 ;
        RECT 216.755 -129.365 217.085 -129.035 ;
        RECT 216.755 -130.725 217.085 -130.395 ;
        RECT 216.755 -132.085 217.085 -131.755 ;
        RECT 216.755 -133.445 217.085 -133.115 ;
        RECT 216.755 -134.805 217.085 -134.475 ;
        RECT 216.755 -136.165 217.085 -135.835 ;
        RECT 216.755 -137.525 217.085 -137.195 ;
        RECT 216.755 -138.885 217.085 -138.555 ;
        RECT 216.755 -140.245 217.085 -139.915 ;
        RECT 216.755 -141.605 217.085 -141.275 ;
        RECT 216.755 -142.965 217.085 -142.635 ;
        RECT 216.755 -144.325 217.085 -143.995 ;
        RECT 216.755 -145.685 217.085 -145.355 ;
        RECT 216.755 -147.045 217.085 -146.715 ;
        RECT 216.755 -148.405 217.085 -148.075 ;
        RECT 216.755 -149.765 217.085 -149.435 ;
        RECT 216.755 -151.125 217.085 -150.795 ;
        RECT 216.755 -152.485 217.085 -152.155 ;
        RECT 216.755 -153.845 217.085 -153.515 ;
        RECT 216.755 -155.205 217.085 -154.875 ;
        RECT 216.755 -156.565 217.085 -156.235 ;
        RECT 216.755 -157.925 217.085 -157.595 ;
        RECT 216.755 -159.285 217.085 -158.955 ;
        RECT 216.755 -160.645 217.085 -160.315 ;
        RECT 216.755 -162.005 217.085 -161.675 ;
        RECT 216.755 -163.365 217.085 -163.035 ;
        RECT 216.755 -164.725 217.085 -164.395 ;
        RECT 216.755 -166.085 217.085 -165.755 ;
        RECT 216.755 -167.445 217.085 -167.115 ;
        RECT 216.755 -168.805 217.085 -168.475 ;
        RECT 216.755 -170.165 217.085 -169.835 ;
        RECT 216.755 -171.525 217.085 -171.195 ;
        RECT 216.755 -172.885 217.085 -172.555 ;
        RECT 216.755 -174.245 217.085 -173.915 ;
        RECT 216.755 -175.605 217.085 -175.275 ;
        RECT 216.755 -176.965 217.085 -176.635 ;
        RECT 216.755 -178.325 217.085 -177.995 ;
        RECT 216.755 -179.685 217.085 -179.355 ;
        RECT 216.755 -181.93 217.085 -180.8 ;
        RECT 216.76 -182.045 217.08 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.115 241.32 218.445 242.45 ;
        RECT 218.115 239.195 218.445 239.525 ;
        RECT 218.115 237.835 218.445 238.165 ;
        RECT 218.12 237.16 218.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.115 -1.525 218.445 -1.195 ;
        RECT 218.115 -2.885 218.445 -2.555 ;
        RECT 218.12 -3.56 218.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 218.115 -95.365 218.445 -95.035 ;
        RECT 218.115 -96.725 218.445 -96.395 ;
        RECT 218.115 -98.085 218.445 -97.755 ;
        RECT 218.115 -99.445 218.445 -99.115 ;
        RECT 218.115 -100.805 218.445 -100.475 ;
        RECT 218.115 -102.165 218.445 -101.835 ;
        RECT 218.115 -103.525 218.445 -103.195 ;
        RECT 218.115 -104.885 218.445 -104.555 ;
        RECT 218.115 -106.245 218.445 -105.915 ;
        RECT 218.115 -107.605 218.445 -107.275 ;
        RECT 218.115 -108.965 218.445 -108.635 ;
        RECT 218.115 -110.325 218.445 -109.995 ;
        RECT 218.115 -111.685 218.445 -111.355 ;
        RECT 218.115 -113.045 218.445 -112.715 ;
        RECT 218.115 -114.405 218.445 -114.075 ;
        RECT 218.115 -115.765 218.445 -115.435 ;
        RECT 218.115 -117.125 218.445 -116.795 ;
        RECT 218.115 -118.485 218.445 -118.155 ;
        RECT 218.115 -119.845 218.445 -119.515 ;
        RECT 218.115 -121.205 218.445 -120.875 ;
        RECT 218.115 -122.565 218.445 -122.235 ;
        RECT 218.115 -123.925 218.445 -123.595 ;
        RECT 218.115 -125.285 218.445 -124.955 ;
        RECT 218.115 -126.645 218.445 -126.315 ;
        RECT 218.115 -128.005 218.445 -127.675 ;
        RECT 218.115 -129.365 218.445 -129.035 ;
        RECT 218.115 -130.725 218.445 -130.395 ;
        RECT 218.115 -132.085 218.445 -131.755 ;
        RECT 218.115 -133.445 218.445 -133.115 ;
        RECT 218.115 -134.805 218.445 -134.475 ;
        RECT 218.115 -136.165 218.445 -135.835 ;
        RECT 218.115 -137.525 218.445 -137.195 ;
        RECT 218.115 -138.885 218.445 -138.555 ;
        RECT 218.115 -140.245 218.445 -139.915 ;
        RECT 218.115 -141.605 218.445 -141.275 ;
        RECT 218.115 -142.965 218.445 -142.635 ;
        RECT 218.115 -144.325 218.445 -143.995 ;
        RECT 218.115 -145.685 218.445 -145.355 ;
        RECT 218.115 -147.045 218.445 -146.715 ;
        RECT 218.115 -148.405 218.445 -148.075 ;
        RECT 218.115 -149.765 218.445 -149.435 ;
        RECT 218.115 -151.125 218.445 -150.795 ;
        RECT 218.115 -152.485 218.445 -152.155 ;
        RECT 218.115 -153.845 218.445 -153.515 ;
        RECT 218.115 -155.205 218.445 -154.875 ;
        RECT 218.115 -156.565 218.445 -156.235 ;
        RECT 218.115 -157.925 218.445 -157.595 ;
        RECT 218.115 -159.285 218.445 -158.955 ;
        RECT 218.115 -160.645 218.445 -160.315 ;
        RECT 218.115 -162.005 218.445 -161.675 ;
        RECT 218.115 -163.365 218.445 -163.035 ;
        RECT 218.115 -164.725 218.445 -164.395 ;
        RECT 218.115 -166.085 218.445 -165.755 ;
        RECT 218.115 -167.445 218.445 -167.115 ;
        RECT 218.115 -168.805 218.445 -168.475 ;
        RECT 218.115 -170.165 218.445 -169.835 ;
        RECT 218.115 -171.525 218.445 -171.195 ;
        RECT 218.115 -172.885 218.445 -172.555 ;
        RECT 218.115 -174.245 218.445 -173.915 ;
        RECT 218.115 -175.605 218.445 -175.275 ;
        RECT 218.115 -176.965 218.445 -176.635 ;
        RECT 218.115 -178.325 218.445 -177.995 ;
        RECT 218.115 -179.685 218.445 -179.355 ;
        RECT 218.115 -181.93 218.445 -180.8 ;
        RECT 218.12 -182.045 218.44 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.475 241.32 219.805 242.45 ;
        RECT 219.475 239.195 219.805 239.525 ;
        RECT 219.475 237.835 219.805 238.165 ;
        RECT 219.48 237.16 219.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.475 -1.525 219.805 -1.195 ;
        RECT 219.475 -2.885 219.805 -2.555 ;
        RECT 219.48 -3.56 219.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 219.475 -95.365 219.805 -95.035 ;
        RECT 219.475 -96.725 219.805 -96.395 ;
        RECT 219.475 -98.085 219.805 -97.755 ;
        RECT 219.475 -99.445 219.805 -99.115 ;
        RECT 219.475 -100.805 219.805 -100.475 ;
        RECT 219.475 -102.165 219.805 -101.835 ;
        RECT 219.475 -103.525 219.805 -103.195 ;
        RECT 219.475 -104.885 219.805 -104.555 ;
        RECT 219.475 -106.245 219.805 -105.915 ;
        RECT 219.475 -107.605 219.805 -107.275 ;
        RECT 219.475 -108.965 219.805 -108.635 ;
        RECT 219.475 -110.325 219.805 -109.995 ;
        RECT 219.475 -111.685 219.805 -111.355 ;
        RECT 219.475 -113.045 219.805 -112.715 ;
        RECT 219.475 -114.405 219.805 -114.075 ;
        RECT 219.475 -115.765 219.805 -115.435 ;
        RECT 219.475 -117.125 219.805 -116.795 ;
        RECT 219.475 -118.485 219.805 -118.155 ;
        RECT 219.475 -119.845 219.805 -119.515 ;
        RECT 219.475 -121.205 219.805 -120.875 ;
        RECT 219.475 -122.565 219.805 -122.235 ;
        RECT 219.475 -123.925 219.805 -123.595 ;
        RECT 219.475 -125.285 219.805 -124.955 ;
        RECT 219.475 -126.645 219.805 -126.315 ;
        RECT 219.475 -128.005 219.805 -127.675 ;
        RECT 219.475 -129.365 219.805 -129.035 ;
        RECT 219.475 -130.725 219.805 -130.395 ;
        RECT 219.475 -132.085 219.805 -131.755 ;
        RECT 219.475 -133.445 219.805 -133.115 ;
        RECT 219.475 -134.805 219.805 -134.475 ;
        RECT 219.475 -136.165 219.805 -135.835 ;
        RECT 219.475 -137.525 219.805 -137.195 ;
        RECT 219.475 -138.885 219.805 -138.555 ;
        RECT 219.475 -140.245 219.805 -139.915 ;
        RECT 219.475 -141.605 219.805 -141.275 ;
        RECT 219.475 -142.965 219.805 -142.635 ;
        RECT 219.475 -144.325 219.805 -143.995 ;
        RECT 219.475 -145.685 219.805 -145.355 ;
        RECT 219.475 -147.045 219.805 -146.715 ;
        RECT 219.475 -148.405 219.805 -148.075 ;
        RECT 219.475 -149.765 219.805 -149.435 ;
        RECT 219.475 -151.125 219.805 -150.795 ;
        RECT 219.475 -152.485 219.805 -152.155 ;
        RECT 219.475 -153.845 219.805 -153.515 ;
        RECT 219.475 -155.205 219.805 -154.875 ;
        RECT 219.475 -156.565 219.805 -156.235 ;
        RECT 219.475 -157.925 219.805 -157.595 ;
        RECT 219.475 -159.285 219.805 -158.955 ;
        RECT 219.475 -160.645 219.805 -160.315 ;
        RECT 219.475 -162.005 219.805 -161.675 ;
        RECT 219.475 -163.365 219.805 -163.035 ;
        RECT 219.475 -164.725 219.805 -164.395 ;
        RECT 219.475 -166.085 219.805 -165.755 ;
        RECT 219.475 -167.445 219.805 -167.115 ;
        RECT 219.475 -168.805 219.805 -168.475 ;
        RECT 219.475 -170.165 219.805 -169.835 ;
        RECT 219.475 -171.525 219.805 -171.195 ;
        RECT 219.475 -172.885 219.805 -172.555 ;
        RECT 219.475 -174.245 219.805 -173.915 ;
        RECT 219.475 -175.605 219.805 -175.275 ;
        RECT 219.475 -176.965 219.805 -176.635 ;
        RECT 219.475 -178.325 219.805 -177.995 ;
        RECT 219.475 -179.685 219.805 -179.355 ;
        RECT 219.475 -181.93 219.805 -180.8 ;
        RECT 219.48 -182.045 219.8 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.835 241.32 221.165 242.45 ;
        RECT 220.835 239.195 221.165 239.525 ;
        RECT 220.835 237.835 221.165 238.165 ;
        RECT 220.84 237.16 221.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 220.835 -99.445 221.165 -99.115 ;
        RECT 220.835 -100.805 221.165 -100.475 ;
        RECT 220.835 -102.165 221.165 -101.835 ;
        RECT 220.835 -103.525 221.165 -103.195 ;
        RECT 220.835 -104.885 221.165 -104.555 ;
        RECT 220.835 -106.245 221.165 -105.915 ;
        RECT 220.835 -107.605 221.165 -107.275 ;
        RECT 220.835 -108.965 221.165 -108.635 ;
        RECT 220.835 -110.325 221.165 -109.995 ;
        RECT 220.835 -111.685 221.165 -111.355 ;
        RECT 220.835 -113.045 221.165 -112.715 ;
        RECT 220.835 -114.405 221.165 -114.075 ;
        RECT 220.835 -115.765 221.165 -115.435 ;
        RECT 220.835 -117.125 221.165 -116.795 ;
        RECT 220.835 -118.485 221.165 -118.155 ;
        RECT 220.835 -119.845 221.165 -119.515 ;
        RECT 220.835 -121.205 221.165 -120.875 ;
        RECT 220.835 -122.565 221.165 -122.235 ;
        RECT 220.835 -123.925 221.165 -123.595 ;
        RECT 220.835 -125.285 221.165 -124.955 ;
        RECT 220.835 -126.645 221.165 -126.315 ;
        RECT 220.835 -128.005 221.165 -127.675 ;
        RECT 220.835 -129.365 221.165 -129.035 ;
        RECT 220.835 -130.725 221.165 -130.395 ;
        RECT 220.835 -132.085 221.165 -131.755 ;
        RECT 220.835 -133.445 221.165 -133.115 ;
        RECT 220.835 -134.805 221.165 -134.475 ;
        RECT 220.835 -136.165 221.165 -135.835 ;
        RECT 220.835 -137.525 221.165 -137.195 ;
        RECT 220.835 -138.885 221.165 -138.555 ;
        RECT 220.835 -140.245 221.165 -139.915 ;
        RECT 220.835 -141.605 221.165 -141.275 ;
        RECT 220.835 -142.965 221.165 -142.635 ;
        RECT 220.835 -144.325 221.165 -143.995 ;
        RECT 220.835 -145.685 221.165 -145.355 ;
        RECT 220.835 -147.045 221.165 -146.715 ;
        RECT 220.835 -148.405 221.165 -148.075 ;
        RECT 220.835 -149.765 221.165 -149.435 ;
        RECT 220.835 -151.125 221.165 -150.795 ;
        RECT 220.835 -152.485 221.165 -152.155 ;
        RECT 220.835 -153.845 221.165 -153.515 ;
        RECT 220.835 -155.205 221.165 -154.875 ;
        RECT 220.835 -156.565 221.165 -156.235 ;
        RECT 220.835 -157.925 221.165 -157.595 ;
        RECT 220.835 -159.285 221.165 -158.955 ;
        RECT 220.835 -160.645 221.165 -160.315 ;
        RECT 220.835 -162.005 221.165 -161.675 ;
        RECT 220.835 -163.365 221.165 -163.035 ;
        RECT 220.835 -164.725 221.165 -164.395 ;
        RECT 220.835 -166.085 221.165 -165.755 ;
        RECT 220.835 -167.445 221.165 -167.115 ;
        RECT 220.835 -168.805 221.165 -168.475 ;
        RECT 220.835 -170.165 221.165 -169.835 ;
        RECT 220.835 -171.525 221.165 -171.195 ;
        RECT 220.835 -172.885 221.165 -172.555 ;
        RECT 220.835 -174.245 221.165 -173.915 ;
        RECT 220.835 -175.605 221.165 -175.275 ;
        RECT 220.835 -176.965 221.165 -176.635 ;
        RECT 220.835 -178.325 221.165 -177.995 ;
        RECT 220.835 -179.685 221.165 -179.355 ;
        RECT 220.835 -181.93 221.165 -180.8 ;
        RECT 220.84 -182.045 221.16 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 221.31 -98.075 221.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.195 241.32 222.525 242.45 ;
        RECT 222.195 239.195 222.525 239.525 ;
        RECT 222.195 237.835 222.525 238.165 ;
        RECT 222.2 237.16 222.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 222.195 -1.525 222.525 -1.195 ;
        RECT 222.195 -2.885 222.525 -2.555 ;
        RECT 222.2 -3.56 222.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.555 241.32 223.885 242.45 ;
        RECT 223.555 239.195 223.885 239.525 ;
        RECT 223.555 237.835 223.885 238.165 ;
        RECT 223.56 237.16 223.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 223.555 -1.525 223.885 -1.195 ;
        RECT 223.555 -2.885 223.885 -2.555 ;
        RECT 223.56 -3.56 223.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.915 241.32 225.245 242.45 ;
        RECT 224.915 239.195 225.245 239.525 ;
        RECT 224.915 237.835 225.245 238.165 ;
        RECT 224.92 237.16 225.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.915 -1.525 225.245 -1.195 ;
        RECT 224.915 -2.885 225.245 -2.555 ;
        RECT 224.92 -3.56 225.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 224.915 -95.365 225.245 -95.035 ;
        RECT 224.915 -96.725 225.245 -96.395 ;
        RECT 224.915 -98.085 225.245 -97.755 ;
        RECT 224.915 -99.445 225.245 -99.115 ;
        RECT 224.915 -100.805 225.245 -100.475 ;
        RECT 224.915 -102.165 225.245 -101.835 ;
        RECT 224.915 -103.525 225.245 -103.195 ;
        RECT 224.915 -104.885 225.245 -104.555 ;
        RECT 224.915 -106.245 225.245 -105.915 ;
        RECT 224.915 -107.605 225.245 -107.275 ;
        RECT 224.915 -108.965 225.245 -108.635 ;
        RECT 224.915 -110.325 225.245 -109.995 ;
        RECT 224.915 -111.685 225.245 -111.355 ;
        RECT 224.915 -113.045 225.245 -112.715 ;
        RECT 224.915 -114.405 225.245 -114.075 ;
        RECT 224.915 -115.765 225.245 -115.435 ;
        RECT 224.915 -117.125 225.245 -116.795 ;
        RECT 224.915 -118.485 225.245 -118.155 ;
        RECT 224.915 -119.845 225.245 -119.515 ;
        RECT 224.915 -121.205 225.245 -120.875 ;
        RECT 224.915 -122.565 225.245 -122.235 ;
        RECT 224.915 -123.925 225.245 -123.595 ;
        RECT 224.915 -125.285 225.245 -124.955 ;
        RECT 224.915 -126.645 225.245 -126.315 ;
        RECT 224.915 -128.005 225.245 -127.675 ;
        RECT 224.915 -129.365 225.245 -129.035 ;
        RECT 224.915 -130.725 225.245 -130.395 ;
        RECT 224.915 -132.085 225.245 -131.755 ;
        RECT 224.915 -133.445 225.245 -133.115 ;
        RECT 224.915 -134.805 225.245 -134.475 ;
        RECT 224.915 -136.165 225.245 -135.835 ;
        RECT 224.915 -137.525 225.245 -137.195 ;
        RECT 224.915 -138.885 225.245 -138.555 ;
        RECT 224.915 -140.245 225.245 -139.915 ;
        RECT 224.915 -141.605 225.245 -141.275 ;
        RECT 224.915 -142.965 225.245 -142.635 ;
        RECT 224.915 -144.325 225.245 -143.995 ;
        RECT 224.915 -145.685 225.245 -145.355 ;
        RECT 224.915 -147.045 225.245 -146.715 ;
        RECT 224.915 -148.405 225.245 -148.075 ;
        RECT 224.915 -149.765 225.245 -149.435 ;
        RECT 224.915 -151.125 225.245 -150.795 ;
        RECT 224.915 -152.485 225.245 -152.155 ;
        RECT 224.915 -153.845 225.245 -153.515 ;
        RECT 224.915 -155.205 225.245 -154.875 ;
        RECT 224.915 -156.565 225.245 -156.235 ;
        RECT 224.915 -157.925 225.245 -157.595 ;
        RECT 224.915 -159.285 225.245 -158.955 ;
        RECT 224.915 -160.645 225.245 -160.315 ;
        RECT 224.915 -162.005 225.245 -161.675 ;
        RECT 224.915 -163.365 225.245 -163.035 ;
        RECT 224.915 -164.725 225.245 -164.395 ;
        RECT 224.915 -166.085 225.245 -165.755 ;
        RECT 224.915 -167.445 225.245 -167.115 ;
        RECT 224.915 -168.805 225.245 -168.475 ;
        RECT 224.915 -170.165 225.245 -169.835 ;
        RECT 224.915 -171.525 225.245 -171.195 ;
        RECT 224.915 -172.885 225.245 -172.555 ;
        RECT 224.915 -174.245 225.245 -173.915 ;
        RECT 224.915 -175.605 225.245 -175.275 ;
        RECT 224.915 -176.965 225.245 -176.635 ;
        RECT 224.915 -178.325 225.245 -177.995 ;
        RECT 224.915 -179.685 225.245 -179.355 ;
        RECT 224.915 -181.93 225.245 -180.8 ;
        RECT 224.92 -182.045 225.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 241.32 226.605 242.45 ;
        RECT 226.275 239.195 226.605 239.525 ;
        RECT 226.275 237.835 226.605 238.165 ;
        RECT 226.28 237.16 226.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 -1.525 226.605 -1.195 ;
        RECT 226.275 -2.885 226.605 -2.555 ;
        RECT 226.28 -3.56 226.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 226.275 -95.365 226.605 -95.035 ;
        RECT 226.275 -96.725 226.605 -96.395 ;
        RECT 226.275 -98.085 226.605 -97.755 ;
        RECT 226.275 -99.445 226.605 -99.115 ;
        RECT 226.275 -100.805 226.605 -100.475 ;
        RECT 226.275 -102.165 226.605 -101.835 ;
        RECT 226.275 -103.525 226.605 -103.195 ;
        RECT 226.275 -104.885 226.605 -104.555 ;
        RECT 226.275 -106.245 226.605 -105.915 ;
        RECT 226.275 -107.605 226.605 -107.275 ;
        RECT 226.275 -108.965 226.605 -108.635 ;
        RECT 226.275 -110.325 226.605 -109.995 ;
        RECT 226.275 -111.685 226.605 -111.355 ;
        RECT 226.275 -113.045 226.605 -112.715 ;
        RECT 226.275 -114.405 226.605 -114.075 ;
        RECT 226.275 -115.765 226.605 -115.435 ;
        RECT 226.275 -117.125 226.605 -116.795 ;
        RECT 226.275 -118.485 226.605 -118.155 ;
        RECT 226.275 -119.845 226.605 -119.515 ;
        RECT 226.275 -121.205 226.605 -120.875 ;
        RECT 226.275 -122.565 226.605 -122.235 ;
        RECT 226.275 -123.925 226.605 -123.595 ;
        RECT 226.275 -125.285 226.605 -124.955 ;
        RECT 226.275 -126.645 226.605 -126.315 ;
        RECT 226.275 -128.005 226.605 -127.675 ;
        RECT 226.275 -129.365 226.605 -129.035 ;
        RECT 226.275 -130.725 226.605 -130.395 ;
        RECT 226.275 -132.085 226.605 -131.755 ;
        RECT 226.275 -133.445 226.605 -133.115 ;
        RECT 226.275 -134.805 226.605 -134.475 ;
        RECT 226.275 -136.165 226.605 -135.835 ;
        RECT 226.275 -137.525 226.605 -137.195 ;
        RECT 226.275 -138.885 226.605 -138.555 ;
        RECT 226.275 -140.245 226.605 -139.915 ;
        RECT 226.275 -141.605 226.605 -141.275 ;
        RECT 226.275 -142.965 226.605 -142.635 ;
        RECT 226.275 -144.325 226.605 -143.995 ;
        RECT 226.275 -145.685 226.605 -145.355 ;
        RECT 226.275 -147.045 226.605 -146.715 ;
        RECT 226.275 -148.405 226.605 -148.075 ;
        RECT 226.275 -149.765 226.605 -149.435 ;
        RECT 226.275 -151.125 226.605 -150.795 ;
        RECT 226.275 -152.485 226.605 -152.155 ;
        RECT 226.275 -153.845 226.605 -153.515 ;
        RECT 226.275 -155.205 226.605 -154.875 ;
        RECT 226.275 -156.565 226.605 -156.235 ;
        RECT 226.275 -157.925 226.605 -157.595 ;
        RECT 226.275 -159.285 226.605 -158.955 ;
        RECT 226.275 -160.645 226.605 -160.315 ;
        RECT 226.275 -162.005 226.605 -161.675 ;
        RECT 226.275 -163.365 226.605 -163.035 ;
        RECT 226.275 -164.725 226.605 -164.395 ;
        RECT 226.275 -166.085 226.605 -165.755 ;
        RECT 226.275 -167.445 226.605 -167.115 ;
        RECT 226.275 -168.805 226.605 -168.475 ;
        RECT 226.275 -170.165 226.605 -169.835 ;
        RECT 226.275 -171.525 226.605 -171.195 ;
        RECT 226.275 -172.885 226.605 -172.555 ;
        RECT 226.275 -174.245 226.605 -173.915 ;
        RECT 226.275 -175.605 226.605 -175.275 ;
        RECT 226.275 -176.965 226.605 -176.635 ;
        RECT 226.275 -178.325 226.605 -177.995 ;
        RECT 226.275 -179.685 226.605 -179.355 ;
        RECT 226.275 -181.93 226.605 -180.8 ;
        RECT 226.28 -182.045 226.6 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.635 241.32 227.965 242.45 ;
        RECT 227.635 239.195 227.965 239.525 ;
        RECT 227.635 237.835 227.965 238.165 ;
        RECT 227.64 237.16 227.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.635 -1.525 227.965 -1.195 ;
        RECT 227.635 -2.885 227.965 -2.555 ;
        RECT 227.64 -3.56 227.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 227.635 -95.365 227.965 -95.035 ;
        RECT 227.635 -96.725 227.965 -96.395 ;
        RECT 227.635 -98.085 227.965 -97.755 ;
        RECT 227.635 -99.445 227.965 -99.115 ;
        RECT 227.635 -100.805 227.965 -100.475 ;
        RECT 227.635 -102.165 227.965 -101.835 ;
        RECT 227.635 -103.525 227.965 -103.195 ;
        RECT 227.635 -104.885 227.965 -104.555 ;
        RECT 227.635 -106.245 227.965 -105.915 ;
        RECT 227.635 -107.605 227.965 -107.275 ;
        RECT 227.635 -108.965 227.965 -108.635 ;
        RECT 227.635 -110.325 227.965 -109.995 ;
        RECT 227.635 -111.685 227.965 -111.355 ;
        RECT 227.635 -113.045 227.965 -112.715 ;
        RECT 227.635 -114.405 227.965 -114.075 ;
        RECT 227.635 -115.765 227.965 -115.435 ;
        RECT 227.635 -117.125 227.965 -116.795 ;
        RECT 227.635 -118.485 227.965 -118.155 ;
        RECT 227.635 -119.845 227.965 -119.515 ;
        RECT 227.635 -121.205 227.965 -120.875 ;
        RECT 227.635 -122.565 227.965 -122.235 ;
        RECT 227.635 -123.925 227.965 -123.595 ;
        RECT 227.635 -125.285 227.965 -124.955 ;
        RECT 227.635 -126.645 227.965 -126.315 ;
        RECT 227.635 -128.005 227.965 -127.675 ;
        RECT 227.635 -129.365 227.965 -129.035 ;
        RECT 227.635 -130.725 227.965 -130.395 ;
        RECT 227.635 -132.085 227.965 -131.755 ;
        RECT 227.635 -133.445 227.965 -133.115 ;
        RECT 227.635 -134.805 227.965 -134.475 ;
        RECT 227.635 -136.165 227.965 -135.835 ;
        RECT 227.635 -137.525 227.965 -137.195 ;
        RECT 227.635 -138.885 227.965 -138.555 ;
        RECT 227.635 -140.245 227.965 -139.915 ;
        RECT 227.635 -141.605 227.965 -141.275 ;
        RECT 227.635 -142.965 227.965 -142.635 ;
        RECT 227.635 -144.325 227.965 -143.995 ;
        RECT 227.635 -145.685 227.965 -145.355 ;
        RECT 227.635 -147.045 227.965 -146.715 ;
        RECT 227.635 -148.405 227.965 -148.075 ;
        RECT 227.635 -149.765 227.965 -149.435 ;
        RECT 227.635 -151.125 227.965 -150.795 ;
        RECT 227.635 -152.485 227.965 -152.155 ;
        RECT 227.635 -153.845 227.965 -153.515 ;
        RECT 227.635 -155.205 227.965 -154.875 ;
        RECT 227.635 -156.565 227.965 -156.235 ;
        RECT 227.635 -157.925 227.965 -157.595 ;
        RECT 227.635 -159.285 227.965 -158.955 ;
        RECT 227.635 -160.645 227.965 -160.315 ;
        RECT 227.635 -162.005 227.965 -161.675 ;
        RECT 227.635 -163.365 227.965 -163.035 ;
        RECT 227.635 -164.725 227.965 -164.395 ;
        RECT 227.635 -166.085 227.965 -165.755 ;
        RECT 227.635 -167.445 227.965 -167.115 ;
        RECT 227.635 -168.805 227.965 -168.475 ;
        RECT 227.635 -170.165 227.965 -169.835 ;
        RECT 227.635 -171.525 227.965 -171.195 ;
        RECT 227.635 -172.885 227.965 -172.555 ;
        RECT 227.635 -174.245 227.965 -173.915 ;
        RECT 227.635 -175.605 227.965 -175.275 ;
        RECT 227.635 -176.965 227.965 -176.635 ;
        RECT 227.635 -178.325 227.965 -177.995 ;
        RECT 227.635 -179.685 227.965 -179.355 ;
        RECT 227.635 -181.93 227.965 -180.8 ;
        RECT 227.64 -182.045 227.96 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.995 241.32 229.325 242.45 ;
        RECT 228.995 239.195 229.325 239.525 ;
        RECT 228.995 237.835 229.325 238.165 ;
        RECT 229 237.16 229.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.995 -1.525 229.325 -1.195 ;
        RECT 228.995 -2.885 229.325 -2.555 ;
        RECT 229 -3.56 229.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 228.995 -95.365 229.325 -95.035 ;
        RECT 228.995 -96.725 229.325 -96.395 ;
        RECT 228.995 -98.085 229.325 -97.755 ;
        RECT 228.995 -99.445 229.325 -99.115 ;
        RECT 228.995 -100.805 229.325 -100.475 ;
        RECT 228.995 -102.165 229.325 -101.835 ;
        RECT 228.995 -103.525 229.325 -103.195 ;
        RECT 228.995 -104.885 229.325 -104.555 ;
        RECT 228.995 -106.245 229.325 -105.915 ;
        RECT 228.995 -107.605 229.325 -107.275 ;
        RECT 228.995 -108.965 229.325 -108.635 ;
        RECT 228.995 -110.325 229.325 -109.995 ;
        RECT 228.995 -111.685 229.325 -111.355 ;
        RECT 228.995 -113.045 229.325 -112.715 ;
        RECT 228.995 -114.405 229.325 -114.075 ;
        RECT 228.995 -115.765 229.325 -115.435 ;
        RECT 228.995 -117.125 229.325 -116.795 ;
        RECT 228.995 -118.485 229.325 -118.155 ;
        RECT 228.995 -119.845 229.325 -119.515 ;
        RECT 228.995 -121.205 229.325 -120.875 ;
        RECT 228.995 -122.565 229.325 -122.235 ;
        RECT 228.995 -123.925 229.325 -123.595 ;
        RECT 228.995 -125.285 229.325 -124.955 ;
        RECT 228.995 -126.645 229.325 -126.315 ;
        RECT 228.995 -128.005 229.325 -127.675 ;
        RECT 228.995 -129.365 229.325 -129.035 ;
        RECT 228.995 -130.725 229.325 -130.395 ;
        RECT 228.995 -132.085 229.325 -131.755 ;
        RECT 228.995 -133.445 229.325 -133.115 ;
        RECT 228.995 -134.805 229.325 -134.475 ;
        RECT 228.995 -136.165 229.325 -135.835 ;
        RECT 228.995 -137.525 229.325 -137.195 ;
        RECT 228.995 -138.885 229.325 -138.555 ;
        RECT 228.995 -140.245 229.325 -139.915 ;
        RECT 228.995 -141.605 229.325 -141.275 ;
        RECT 228.995 -142.965 229.325 -142.635 ;
        RECT 228.995 -144.325 229.325 -143.995 ;
        RECT 228.995 -145.685 229.325 -145.355 ;
        RECT 228.995 -147.045 229.325 -146.715 ;
        RECT 228.995 -148.405 229.325 -148.075 ;
        RECT 228.995 -149.765 229.325 -149.435 ;
        RECT 228.995 -151.125 229.325 -150.795 ;
        RECT 228.995 -152.485 229.325 -152.155 ;
        RECT 228.995 -153.845 229.325 -153.515 ;
        RECT 228.995 -155.205 229.325 -154.875 ;
        RECT 228.995 -156.565 229.325 -156.235 ;
        RECT 228.995 -157.925 229.325 -157.595 ;
        RECT 228.995 -159.285 229.325 -158.955 ;
        RECT 228.995 -160.645 229.325 -160.315 ;
        RECT 228.995 -162.005 229.325 -161.675 ;
        RECT 228.995 -163.365 229.325 -163.035 ;
        RECT 228.995 -164.725 229.325 -164.395 ;
        RECT 228.995 -166.085 229.325 -165.755 ;
        RECT 228.995 -167.445 229.325 -167.115 ;
        RECT 228.995 -168.805 229.325 -168.475 ;
        RECT 228.995 -170.165 229.325 -169.835 ;
        RECT 228.995 -171.525 229.325 -171.195 ;
        RECT 228.995 -172.885 229.325 -172.555 ;
        RECT 228.995 -174.245 229.325 -173.915 ;
        RECT 228.995 -175.605 229.325 -175.275 ;
        RECT 228.995 -176.965 229.325 -176.635 ;
        RECT 228.995 -178.325 229.325 -177.995 ;
        RECT 228.995 -179.685 229.325 -179.355 ;
        RECT 228.995 -181.93 229.325 -180.8 ;
        RECT 229 -182.045 229.32 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.355 241.32 230.685 242.45 ;
        RECT 230.355 239.195 230.685 239.525 ;
        RECT 230.355 237.835 230.685 238.165 ;
        RECT 230.36 237.16 230.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.355 -1.525 230.685 -1.195 ;
        RECT 230.355 -2.885 230.685 -2.555 ;
        RECT 230.36 -3.56 230.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 230.355 -95.365 230.685 -95.035 ;
        RECT 230.355 -96.725 230.685 -96.395 ;
        RECT 230.355 -98.085 230.685 -97.755 ;
        RECT 230.355 -99.445 230.685 -99.115 ;
        RECT 230.355 -100.805 230.685 -100.475 ;
        RECT 230.355 -102.165 230.685 -101.835 ;
        RECT 230.355 -103.525 230.685 -103.195 ;
        RECT 230.355 -104.885 230.685 -104.555 ;
        RECT 230.355 -106.245 230.685 -105.915 ;
        RECT 230.355 -107.605 230.685 -107.275 ;
        RECT 230.355 -108.965 230.685 -108.635 ;
        RECT 230.355 -110.325 230.685 -109.995 ;
        RECT 230.355 -111.685 230.685 -111.355 ;
        RECT 230.355 -113.045 230.685 -112.715 ;
        RECT 230.355 -114.405 230.685 -114.075 ;
        RECT 230.355 -115.765 230.685 -115.435 ;
        RECT 230.355 -117.125 230.685 -116.795 ;
        RECT 230.355 -118.485 230.685 -118.155 ;
        RECT 230.355 -119.845 230.685 -119.515 ;
        RECT 230.355 -121.205 230.685 -120.875 ;
        RECT 230.355 -122.565 230.685 -122.235 ;
        RECT 230.355 -123.925 230.685 -123.595 ;
        RECT 230.355 -125.285 230.685 -124.955 ;
        RECT 230.355 -126.645 230.685 -126.315 ;
        RECT 230.355 -128.005 230.685 -127.675 ;
        RECT 230.355 -129.365 230.685 -129.035 ;
        RECT 230.355 -130.725 230.685 -130.395 ;
        RECT 230.355 -132.085 230.685 -131.755 ;
        RECT 230.355 -133.445 230.685 -133.115 ;
        RECT 230.355 -134.805 230.685 -134.475 ;
        RECT 230.355 -136.165 230.685 -135.835 ;
        RECT 230.355 -137.525 230.685 -137.195 ;
        RECT 230.355 -138.885 230.685 -138.555 ;
        RECT 230.355 -140.245 230.685 -139.915 ;
        RECT 230.355 -141.605 230.685 -141.275 ;
        RECT 230.355 -142.965 230.685 -142.635 ;
        RECT 230.355 -144.325 230.685 -143.995 ;
        RECT 230.355 -145.685 230.685 -145.355 ;
        RECT 230.355 -147.045 230.685 -146.715 ;
        RECT 230.355 -148.405 230.685 -148.075 ;
        RECT 230.355 -149.765 230.685 -149.435 ;
        RECT 230.355 -151.125 230.685 -150.795 ;
        RECT 230.355 -152.485 230.685 -152.155 ;
        RECT 230.355 -153.845 230.685 -153.515 ;
        RECT 230.355 -155.205 230.685 -154.875 ;
        RECT 230.355 -156.565 230.685 -156.235 ;
        RECT 230.355 -157.925 230.685 -157.595 ;
        RECT 230.355 -159.285 230.685 -158.955 ;
        RECT 230.355 -160.645 230.685 -160.315 ;
        RECT 230.355 -162.005 230.685 -161.675 ;
        RECT 230.355 -163.365 230.685 -163.035 ;
        RECT 230.355 -164.725 230.685 -164.395 ;
        RECT 230.355 -166.085 230.685 -165.755 ;
        RECT 230.355 -167.445 230.685 -167.115 ;
        RECT 230.355 -168.805 230.685 -168.475 ;
        RECT 230.355 -170.165 230.685 -169.835 ;
        RECT 230.355 -171.525 230.685 -171.195 ;
        RECT 230.355 -172.885 230.685 -172.555 ;
        RECT 230.355 -174.245 230.685 -173.915 ;
        RECT 230.355 -175.605 230.685 -175.275 ;
        RECT 230.355 -176.965 230.685 -176.635 ;
        RECT 230.355 -178.325 230.685 -177.995 ;
        RECT 230.355 -179.685 230.685 -179.355 ;
        RECT 230.355 -181.93 230.685 -180.8 ;
        RECT 230.36 -182.045 230.68 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.715 241.32 232.045 242.45 ;
        RECT 231.715 239.195 232.045 239.525 ;
        RECT 231.715 237.835 232.045 238.165 ;
        RECT 231.72 237.16 232.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 231.715 -99.445 232.045 -99.115 ;
        RECT 231.715 -100.805 232.045 -100.475 ;
        RECT 231.715 -102.165 232.045 -101.835 ;
        RECT 231.715 -103.525 232.045 -103.195 ;
        RECT 231.715 -104.885 232.045 -104.555 ;
        RECT 231.715 -106.245 232.045 -105.915 ;
        RECT 231.715 -107.605 232.045 -107.275 ;
        RECT 231.715 -108.965 232.045 -108.635 ;
        RECT 231.715 -110.325 232.045 -109.995 ;
        RECT 231.715 -111.685 232.045 -111.355 ;
        RECT 231.715 -113.045 232.045 -112.715 ;
        RECT 231.715 -114.405 232.045 -114.075 ;
        RECT 231.715 -115.765 232.045 -115.435 ;
        RECT 231.715 -117.125 232.045 -116.795 ;
        RECT 231.715 -118.485 232.045 -118.155 ;
        RECT 231.715 -119.845 232.045 -119.515 ;
        RECT 231.715 -121.205 232.045 -120.875 ;
        RECT 231.715 -122.565 232.045 -122.235 ;
        RECT 231.715 -123.925 232.045 -123.595 ;
        RECT 231.715 -125.285 232.045 -124.955 ;
        RECT 231.715 -126.645 232.045 -126.315 ;
        RECT 231.715 -128.005 232.045 -127.675 ;
        RECT 231.715 -129.365 232.045 -129.035 ;
        RECT 231.715 -130.725 232.045 -130.395 ;
        RECT 231.715 -132.085 232.045 -131.755 ;
        RECT 231.715 -133.445 232.045 -133.115 ;
        RECT 231.715 -134.805 232.045 -134.475 ;
        RECT 231.715 -136.165 232.045 -135.835 ;
        RECT 231.715 -137.525 232.045 -137.195 ;
        RECT 231.715 -138.885 232.045 -138.555 ;
        RECT 231.715 -140.245 232.045 -139.915 ;
        RECT 231.715 -141.605 232.045 -141.275 ;
        RECT 231.715 -142.965 232.045 -142.635 ;
        RECT 231.715 -144.325 232.045 -143.995 ;
        RECT 231.715 -145.685 232.045 -145.355 ;
        RECT 231.715 -147.045 232.045 -146.715 ;
        RECT 231.715 -148.405 232.045 -148.075 ;
        RECT 231.715 -149.765 232.045 -149.435 ;
        RECT 231.715 -151.125 232.045 -150.795 ;
        RECT 231.715 -152.485 232.045 -152.155 ;
        RECT 231.715 -153.845 232.045 -153.515 ;
        RECT 231.715 -155.205 232.045 -154.875 ;
        RECT 231.715 -156.565 232.045 -156.235 ;
        RECT 231.715 -157.925 232.045 -157.595 ;
        RECT 231.715 -159.285 232.045 -158.955 ;
        RECT 231.715 -160.645 232.045 -160.315 ;
        RECT 231.715 -162.005 232.045 -161.675 ;
        RECT 231.715 -163.365 232.045 -163.035 ;
        RECT 231.715 -164.725 232.045 -164.395 ;
        RECT 231.715 -166.085 232.045 -165.755 ;
        RECT 231.715 -167.445 232.045 -167.115 ;
        RECT 231.715 -168.805 232.045 -168.475 ;
        RECT 231.715 -170.165 232.045 -169.835 ;
        RECT 231.715 -171.525 232.045 -171.195 ;
        RECT 231.715 -172.885 232.045 -172.555 ;
        RECT 231.715 -174.245 232.045 -173.915 ;
        RECT 231.715 -175.605 232.045 -175.275 ;
        RECT 231.715 -176.965 232.045 -176.635 ;
        RECT 231.715 -178.325 232.045 -177.995 ;
        RECT 231.715 -179.685 232.045 -179.355 ;
        RECT 231.715 -181.93 232.045 -180.8 ;
        RECT 231.72 -182.045 232.04 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 232.21 -98.075 232.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.075 241.32 233.405 242.45 ;
        RECT 233.075 239.195 233.405 239.525 ;
        RECT 233.075 237.835 233.405 238.165 ;
        RECT 233.08 237.16 233.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 233.075 -1.525 233.405 -1.195 ;
        RECT 233.075 -2.885 233.405 -2.555 ;
        RECT 233.08 -3.56 233.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.435 241.32 234.765 242.45 ;
        RECT 234.435 239.195 234.765 239.525 ;
        RECT 234.435 237.835 234.765 238.165 ;
        RECT 234.44 237.16 234.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 234.435 -1.525 234.765 -1.195 ;
        RECT 234.435 -2.885 234.765 -2.555 ;
        RECT 234.44 -3.56 234.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.795 241.32 236.125 242.45 ;
        RECT 235.795 239.195 236.125 239.525 ;
        RECT 235.795 237.835 236.125 238.165 ;
        RECT 235.8 237.16 236.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.795 -1.525 236.125 -1.195 ;
        RECT 235.795 -2.885 236.125 -2.555 ;
        RECT 235.8 -3.56 236.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 235.795 -95.365 236.125 -95.035 ;
        RECT 235.795 -96.725 236.125 -96.395 ;
        RECT 235.795 -98.085 236.125 -97.755 ;
        RECT 235.795 -99.445 236.125 -99.115 ;
        RECT 235.795 -100.805 236.125 -100.475 ;
        RECT 235.795 -102.165 236.125 -101.835 ;
        RECT 235.795 -103.525 236.125 -103.195 ;
        RECT 235.795 -104.885 236.125 -104.555 ;
        RECT 235.795 -106.245 236.125 -105.915 ;
        RECT 235.795 -107.605 236.125 -107.275 ;
        RECT 235.795 -108.965 236.125 -108.635 ;
        RECT 235.795 -110.325 236.125 -109.995 ;
        RECT 235.795 -111.685 236.125 -111.355 ;
        RECT 235.795 -113.045 236.125 -112.715 ;
        RECT 235.795 -114.405 236.125 -114.075 ;
        RECT 235.795 -115.765 236.125 -115.435 ;
        RECT 235.795 -117.125 236.125 -116.795 ;
        RECT 235.795 -118.485 236.125 -118.155 ;
        RECT 235.795 -119.845 236.125 -119.515 ;
        RECT 235.795 -121.205 236.125 -120.875 ;
        RECT 235.795 -122.565 236.125 -122.235 ;
        RECT 235.795 -123.925 236.125 -123.595 ;
        RECT 235.795 -125.285 236.125 -124.955 ;
        RECT 235.795 -126.645 236.125 -126.315 ;
        RECT 235.795 -128.005 236.125 -127.675 ;
        RECT 235.795 -129.365 236.125 -129.035 ;
        RECT 235.795 -130.725 236.125 -130.395 ;
        RECT 235.795 -132.085 236.125 -131.755 ;
        RECT 235.795 -133.445 236.125 -133.115 ;
        RECT 235.795 -134.805 236.125 -134.475 ;
        RECT 235.795 -136.165 236.125 -135.835 ;
        RECT 235.795 -137.525 236.125 -137.195 ;
        RECT 235.795 -138.885 236.125 -138.555 ;
        RECT 235.795 -140.245 236.125 -139.915 ;
        RECT 235.795 -141.605 236.125 -141.275 ;
        RECT 235.795 -142.965 236.125 -142.635 ;
        RECT 235.795 -144.325 236.125 -143.995 ;
        RECT 235.795 -145.685 236.125 -145.355 ;
        RECT 235.795 -147.045 236.125 -146.715 ;
        RECT 235.795 -148.405 236.125 -148.075 ;
        RECT 235.795 -149.765 236.125 -149.435 ;
        RECT 235.795 -151.125 236.125 -150.795 ;
        RECT 235.795 -152.485 236.125 -152.155 ;
        RECT 235.795 -153.845 236.125 -153.515 ;
        RECT 235.795 -155.205 236.125 -154.875 ;
        RECT 235.795 -156.565 236.125 -156.235 ;
        RECT 235.795 -157.925 236.125 -157.595 ;
        RECT 235.795 -159.285 236.125 -158.955 ;
        RECT 235.795 -160.645 236.125 -160.315 ;
        RECT 235.795 -162.005 236.125 -161.675 ;
        RECT 235.795 -163.365 236.125 -163.035 ;
        RECT 235.795 -164.725 236.125 -164.395 ;
        RECT 235.795 -166.085 236.125 -165.755 ;
        RECT 235.795 -167.445 236.125 -167.115 ;
        RECT 235.795 -168.805 236.125 -168.475 ;
        RECT 235.795 -170.165 236.125 -169.835 ;
        RECT 235.795 -171.525 236.125 -171.195 ;
        RECT 235.795 -172.885 236.125 -172.555 ;
        RECT 235.795 -174.245 236.125 -173.915 ;
        RECT 235.795 -175.605 236.125 -175.275 ;
        RECT 235.795 -176.965 236.125 -176.635 ;
        RECT 235.795 -178.325 236.125 -177.995 ;
        RECT 235.795 -179.685 236.125 -179.355 ;
        RECT 235.795 -181.93 236.125 -180.8 ;
        RECT 235.8 -182.045 236.12 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.155 241.32 237.485 242.45 ;
        RECT 237.155 239.195 237.485 239.525 ;
        RECT 237.155 237.835 237.485 238.165 ;
        RECT 237.16 237.16 237.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.155 -1.525 237.485 -1.195 ;
        RECT 237.155 -2.885 237.485 -2.555 ;
        RECT 237.16 -3.56 237.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 237.155 -95.365 237.485 -95.035 ;
        RECT 237.155 -96.725 237.485 -96.395 ;
        RECT 237.155 -98.085 237.485 -97.755 ;
        RECT 237.155 -99.445 237.485 -99.115 ;
        RECT 237.155 -100.805 237.485 -100.475 ;
        RECT 237.155 -102.165 237.485 -101.835 ;
        RECT 237.155 -103.525 237.485 -103.195 ;
        RECT 237.155 -104.885 237.485 -104.555 ;
        RECT 237.155 -106.245 237.485 -105.915 ;
        RECT 237.155 -107.605 237.485 -107.275 ;
        RECT 237.155 -108.965 237.485 -108.635 ;
        RECT 237.155 -110.325 237.485 -109.995 ;
        RECT 237.155 -111.685 237.485 -111.355 ;
        RECT 237.155 -113.045 237.485 -112.715 ;
        RECT 237.155 -114.405 237.485 -114.075 ;
        RECT 237.155 -115.765 237.485 -115.435 ;
        RECT 237.155 -117.125 237.485 -116.795 ;
        RECT 237.155 -118.485 237.485 -118.155 ;
        RECT 237.155 -119.845 237.485 -119.515 ;
        RECT 237.155 -121.205 237.485 -120.875 ;
        RECT 237.155 -122.565 237.485 -122.235 ;
        RECT 237.155 -123.925 237.485 -123.595 ;
        RECT 237.155 -125.285 237.485 -124.955 ;
        RECT 237.155 -126.645 237.485 -126.315 ;
        RECT 237.155 -128.005 237.485 -127.675 ;
        RECT 237.155 -129.365 237.485 -129.035 ;
        RECT 237.155 -130.725 237.485 -130.395 ;
        RECT 237.155 -132.085 237.485 -131.755 ;
        RECT 237.155 -133.445 237.485 -133.115 ;
        RECT 237.155 -134.805 237.485 -134.475 ;
        RECT 237.155 -136.165 237.485 -135.835 ;
        RECT 237.155 -137.525 237.485 -137.195 ;
        RECT 237.155 -138.885 237.485 -138.555 ;
        RECT 237.155 -140.245 237.485 -139.915 ;
        RECT 237.155 -141.605 237.485 -141.275 ;
        RECT 237.155 -142.965 237.485 -142.635 ;
        RECT 237.155 -144.325 237.485 -143.995 ;
        RECT 237.155 -145.685 237.485 -145.355 ;
        RECT 237.155 -147.045 237.485 -146.715 ;
        RECT 237.155 -148.405 237.485 -148.075 ;
        RECT 237.155 -149.765 237.485 -149.435 ;
        RECT 237.155 -151.125 237.485 -150.795 ;
        RECT 237.155 -152.485 237.485 -152.155 ;
        RECT 237.155 -153.845 237.485 -153.515 ;
        RECT 237.155 -155.205 237.485 -154.875 ;
        RECT 237.155 -156.565 237.485 -156.235 ;
        RECT 237.155 -157.925 237.485 -157.595 ;
        RECT 237.155 -159.285 237.485 -158.955 ;
        RECT 237.155 -160.645 237.485 -160.315 ;
        RECT 237.155 -162.005 237.485 -161.675 ;
        RECT 237.155 -163.365 237.485 -163.035 ;
        RECT 237.155 -164.725 237.485 -164.395 ;
        RECT 237.155 -166.085 237.485 -165.755 ;
        RECT 237.155 -167.445 237.485 -167.115 ;
        RECT 237.155 -168.805 237.485 -168.475 ;
        RECT 237.155 -170.165 237.485 -169.835 ;
        RECT 237.155 -171.525 237.485 -171.195 ;
        RECT 237.155 -172.885 237.485 -172.555 ;
        RECT 237.155 -174.245 237.485 -173.915 ;
        RECT 237.155 -175.605 237.485 -175.275 ;
        RECT 237.155 -176.965 237.485 -176.635 ;
        RECT 237.155 -178.325 237.485 -177.995 ;
        RECT 237.155 -179.685 237.485 -179.355 ;
        RECT 237.155 -181.93 237.485 -180.8 ;
        RECT 237.16 -182.045 237.48 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.515 241.32 238.845 242.45 ;
        RECT 238.515 239.195 238.845 239.525 ;
        RECT 238.515 237.835 238.845 238.165 ;
        RECT 238.52 237.16 238.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.515 -1.525 238.845 -1.195 ;
        RECT 238.515 -2.885 238.845 -2.555 ;
        RECT 238.52 -3.56 238.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 238.515 -95.365 238.845 -95.035 ;
        RECT 238.515 -96.725 238.845 -96.395 ;
        RECT 238.515 -98.085 238.845 -97.755 ;
        RECT 238.515 -99.445 238.845 -99.115 ;
        RECT 238.515 -100.805 238.845 -100.475 ;
        RECT 238.515 -102.165 238.845 -101.835 ;
        RECT 238.515 -103.525 238.845 -103.195 ;
        RECT 238.515 -104.885 238.845 -104.555 ;
        RECT 238.515 -106.245 238.845 -105.915 ;
        RECT 238.515 -107.605 238.845 -107.275 ;
        RECT 238.515 -108.965 238.845 -108.635 ;
        RECT 238.515 -110.325 238.845 -109.995 ;
        RECT 238.515 -111.685 238.845 -111.355 ;
        RECT 238.515 -113.045 238.845 -112.715 ;
        RECT 238.515 -114.405 238.845 -114.075 ;
        RECT 238.515 -115.765 238.845 -115.435 ;
        RECT 238.515 -117.125 238.845 -116.795 ;
        RECT 238.515 -118.485 238.845 -118.155 ;
        RECT 238.515 -119.845 238.845 -119.515 ;
        RECT 238.515 -121.205 238.845 -120.875 ;
        RECT 238.515 -122.565 238.845 -122.235 ;
        RECT 238.515 -123.925 238.845 -123.595 ;
        RECT 238.515 -125.285 238.845 -124.955 ;
        RECT 238.515 -126.645 238.845 -126.315 ;
        RECT 238.515 -128.005 238.845 -127.675 ;
        RECT 238.515 -129.365 238.845 -129.035 ;
        RECT 238.515 -130.725 238.845 -130.395 ;
        RECT 238.515 -132.085 238.845 -131.755 ;
        RECT 238.515 -133.445 238.845 -133.115 ;
        RECT 238.515 -134.805 238.845 -134.475 ;
        RECT 238.515 -136.165 238.845 -135.835 ;
        RECT 238.515 -137.525 238.845 -137.195 ;
        RECT 238.515 -138.885 238.845 -138.555 ;
        RECT 238.515 -140.245 238.845 -139.915 ;
        RECT 238.515 -141.605 238.845 -141.275 ;
        RECT 238.515 -142.965 238.845 -142.635 ;
        RECT 238.515 -144.325 238.845 -143.995 ;
        RECT 238.515 -145.685 238.845 -145.355 ;
        RECT 238.515 -147.045 238.845 -146.715 ;
        RECT 238.515 -148.405 238.845 -148.075 ;
        RECT 238.515 -149.765 238.845 -149.435 ;
        RECT 238.515 -151.125 238.845 -150.795 ;
        RECT 238.515 -152.485 238.845 -152.155 ;
        RECT 238.515 -153.845 238.845 -153.515 ;
        RECT 238.515 -155.205 238.845 -154.875 ;
        RECT 238.515 -156.565 238.845 -156.235 ;
        RECT 238.515 -157.925 238.845 -157.595 ;
        RECT 238.515 -159.285 238.845 -158.955 ;
        RECT 238.515 -160.645 238.845 -160.315 ;
        RECT 238.515 -162.005 238.845 -161.675 ;
        RECT 238.515 -163.365 238.845 -163.035 ;
        RECT 238.515 -164.725 238.845 -164.395 ;
        RECT 238.515 -166.085 238.845 -165.755 ;
        RECT 238.515 -167.445 238.845 -167.115 ;
        RECT 238.515 -168.805 238.845 -168.475 ;
        RECT 238.515 -170.165 238.845 -169.835 ;
        RECT 238.515 -171.525 238.845 -171.195 ;
        RECT 238.515 -172.885 238.845 -172.555 ;
        RECT 238.515 -174.245 238.845 -173.915 ;
        RECT 238.515 -175.605 238.845 -175.275 ;
        RECT 238.515 -176.965 238.845 -176.635 ;
        RECT 238.515 -178.325 238.845 -177.995 ;
        RECT 238.515 -179.685 238.845 -179.355 ;
        RECT 238.515 -181.93 238.845 -180.8 ;
        RECT 238.52 -182.045 238.84 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.875 241.32 240.205 242.45 ;
        RECT 239.875 239.195 240.205 239.525 ;
        RECT 239.875 237.835 240.205 238.165 ;
        RECT 239.88 237.16 240.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.875 -1.525 240.205 -1.195 ;
        RECT 239.875 -2.885 240.205 -2.555 ;
        RECT 239.88 -3.56 240.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 239.875 -142.965 240.205 -142.635 ;
        RECT 239.875 -144.325 240.205 -143.995 ;
        RECT 239.875 -145.685 240.205 -145.355 ;
        RECT 239.875 -147.045 240.205 -146.715 ;
        RECT 239.875 -148.405 240.205 -148.075 ;
        RECT 239.875 -149.765 240.205 -149.435 ;
        RECT 239.875 -151.125 240.205 -150.795 ;
        RECT 239.875 -152.485 240.205 -152.155 ;
        RECT 239.875 -153.845 240.205 -153.515 ;
        RECT 239.875 -155.205 240.205 -154.875 ;
        RECT 239.875 -156.565 240.205 -156.235 ;
        RECT 239.875 -157.925 240.205 -157.595 ;
        RECT 239.875 -159.285 240.205 -158.955 ;
        RECT 239.875 -160.645 240.205 -160.315 ;
        RECT 239.875 -162.005 240.205 -161.675 ;
        RECT 239.875 -163.365 240.205 -163.035 ;
        RECT 239.875 -164.725 240.205 -164.395 ;
        RECT 239.875 -166.085 240.205 -165.755 ;
        RECT 239.875 -167.445 240.205 -167.115 ;
        RECT 239.875 -168.805 240.205 -168.475 ;
        RECT 239.875 -170.165 240.205 -169.835 ;
        RECT 239.875 -171.525 240.205 -171.195 ;
        RECT 239.875 -172.885 240.205 -172.555 ;
        RECT 239.875 -174.245 240.205 -173.915 ;
        RECT 239.875 -175.605 240.205 -175.275 ;
        RECT 239.875 -176.965 240.205 -176.635 ;
        RECT 239.875 -178.325 240.205 -177.995 ;
        RECT 239.875 -179.685 240.205 -179.355 ;
        RECT 239.875 -181.93 240.205 -180.8 ;
        RECT 239.88 -182.045 240.2 -95.035 ;
        RECT 239.875 -95.365 240.205 -95.035 ;
        RECT 239.875 -96.725 240.205 -96.395 ;
        RECT 239.875 -98.085 240.205 -97.755 ;
        RECT 239.875 -99.445 240.205 -99.115 ;
        RECT 239.875 -100.805 240.205 -100.475 ;
        RECT 239.875 -102.165 240.205 -101.835 ;
        RECT 239.875 -103.525 240.205 -103.195 ;
        RECT 239.875 -104.885 240.205 -104.555 ;
        RECT 239.875 -106.245 240.205 -105.915 ;
        RECT 239.875 -107.605 240.205 -107.275 ;
        RECT 239.875 -108.965 240.205 -108.635 ;
        RECT 239.875 -110.325 240.205 -109.995 ;
        RECT 239.875 -111.685 240.205 -111.355 ;
        RECT 239.875 -113.045 240.205 -112.715 ;
        RECT 239.875 -114.405 240.205 -114.075 ;
        RECT 239.875 -115.765 240.205 -115.435 ;
        RECT 239.875 -117.125 240.205 -116.795 ;
        RECT 239.875 -118.485 240.205 -118.155 ;
        RECT 239.875 -119.845 240.205 -119.515 ;
        RECT 239.875 -121.205 240.205 -120.875 ;
        RECT 239.875 -122.565 240.205 -122.235 ;
        RECT 239.875 -123.925 240.205 -123.595 ;
        RECT 239.875 -125.285 240.205 -124.955 ;
        RECT 239.875 -126.645 240.205 -126.315 ;
        RECT 239.875 -128.005 240.205 -127.675 ;
        RECT 239.875 -129.365 240.205 -129.035 ;
        RECT 239.875 -130.725 240.205 -130.395 ;
        RECT 239.875 -132.085 240.205 -131.755 ;
        RECT 239.875 -133.445 240.205 -133.115 ;
        RECT 239.875 -134.805 240.205 -134.475 ;
        RECT 239.875 -136.165 240.205 -135.835 ;
        RECT 239.875 -137.525 240.205 -137.195 ;
        RECT 239.875 -138.885 240.205 -138.555 ;
        RECT 239.875 -140.245 240.205 -139.915 ;
        RECT 239.875 -141.605 240.205 -141.275 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 241.32 193.965 242.45 ;
        RECT 193.635 239.195 193.965 239.525 ;
        RECT 193.635 237.835 193.965 238.165 ;
        RECT 193.64 237.16 193.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 -1.525 193.965 -1.195 ;
        RECT 193.635 -2.885 193.965 -2.555 ;
        RECT 193.64 -3.56 193.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 193.635 -95.365 193.965 -95.035 ;
        RECT 193.635 -96.725 193.965 -96.395 ;
        RECT 193.635 -98.085 193.965 -97.755 ;
        RECT 193.635 -99.445 193.965 -99.115 ;
        RECT 193.635 -100.805 193.965 -100.475 ;
        RECT 193.635 -102.165 193.965 -101.835 ;
        RECT 193.635 -103.525 193.965 -103.195 ;
        RECT 193.635 -104.885 193.965 -104.555 ;
        RECT 193.635 -106.245 193.965 -105.915 ;
        RECT 193.635 -107.605 193.965 -107.275 ;
        RECT 193.635 -108.965 193.965 -108.635 ;
        RECT 193.635 -110.325 193.965 -109.995 ;
        RECT 193.635 -111.685 193.965 -111.355 ;
        RECT 193.635 -113.045 193.965 -112.715 ;
        RECT 193.635 -114.405 193.965 -114.075 ;
        RECT 193.635 -115.765 193.965 -115.435 ;
        RECT 193.635 -117.125 193.965 -116.795 ;
        RECT 193.635 -118.485 193.965 -118.155 ;
        RECT 193.635 -119.845 193.965 -119.515 ;
        RECT 193.635 -121.205 193.965 -120.875 ;
        RECT 193.635 -122.565 193.965 -122.235 ;
        RECT 193.635 -123.925 193.965 -123.595 ;
        RECT 193.635 -125.285 193.965 -124.955 ;
        RECT 193.635 -126.645 193.965 -126.315 ;
        RECT 193.635 -128.005 193.965 -127.675 ;
        RECT 193.635 -129.365 193.965 -129.035 ;
        RECT 193.635 -130.725 193.965 -130.395 ;
        RECT 193.635 -132.085 193.965 -131.755 ;
        RECT 193.635 -133.445 193.965 -133.115 ;
        RECT 193.635 -134.805 193.965 -134.475 ;
        RECT 193.635 -136.165 193.965 -135.835 ;
        RECT 193.635 -137.525 193.965 -137.195 ;
        RECT 193.635 -138.885 193.965 -138.555 ;
        RECT 193.635 -140.245 193.965 -139.915 ;
        RECT 193.635 -141.605 193.965 -141.275 ;
        RECT 193.635 -142.965 193.965 -142.635 ;
        RECT 193.635 -144.325 193.965 -143.995 ;
        RECT 193.635 -145.685 193.965 -145.355 ;
        RECT 193.635 -147.045 193.965 -146.715 ;
        RECT 193.635 -148.405 193.965 -148.075 ;
        RECT 193.635 -149.765 193.965 -149.435 ;
        RECT 193.635 -151.125 193.965 -150.795 ;
        RECT 193.635 -152.485 193.965 -152.155 ;
        RECT 193.635 -153.845 193.965 -153.515 ;
        RECT 193.635 -155.205 193.965 -154.875 ;
        RECT 193.635 -156.565 193.965 -156.235 ;
        RECT 193.635 -157.925 193.965 -157.595 ;
        RECT 193.635 -159.285 193.965 -158.955 ;
        RECT 193.635 -160.645 193.965 -160.315 ;
        RECT 193.635 -162.005 193.965 -161.675 ;
        RECT 193.635 -163.365 193.965 -163.035 ;
        RECT 193.635 -164.725 193.965 -164.395 ;
        RECT 193.635 -166.085 193.965 -165.755 ;
        RECT 193.635 -167.445 193.965 -167.115 ;
        RECT 193.635 -168.805 193.965 -168.475 ;
        RECT 193.635 -170.165 193.965 -169.835 ;
        RECT 193.635 -171.525 193.965 -171.195 ;
        RECT 193.635 -172.885 193.965 -172.555 ;
        RECT 193.635 -174.245 193.965 -173.915 ;
        RECT 193.635 -175.605 193.965 -175.275 ;
        RECT 193.635 -176.965 193.965 -176.635 ;
        RECT 193.635 -178.325 193.965 -177.995 ;
        RECT 193.635 -179.685 193.965 -179.355 ;
        RECT 193.635 -181.93 193.965 -180.8 ;
        RECT 193.64 -182.045 193.96 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 241.32 195.325 242.45 ;
        RECT 194.995 239.195 195.325 239.525 ;
        RECT 194.995 237.835 195.325 238.165 ;
        RECT 195 237.16 195.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 -1.525 195.325 -1.195 ;
        RECT 194.995 -2.885 195.325 -2.555 ;
        RECT 195 -3.56 195.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 194.995 -95.365 195.325 -95.035 ;
        RECT 194.995 -96.725 195.325 -96.395 ;
        RECT 194.995 -98.085 195.325 -97.755 ;
        RECT 194.995 -99.445 195.325 -99.115 ;
        RECT 194.995 -100.805 195.325 -100.475 ;
        RECT 194.995 -102.165 195.325 -101.835 ;
        RECT 194.995 -103.525 195.325 -103.195 ;
        RECT 194.995 -104.885 195.325 -104.555 ;
        RECT 194.995 -106.245 195.325 -105.915 ;
        RECT 194.995 -107.605 195.325 -107.275 ;
        RECT 194.995 -108.965 195.325 -108.635 ;
        RECT 194.995 -110.325 195.325 -109.995 ;
        RECT 194.995 -111.685 195.325 -111.355 ;
        RECT 194.995 -113.045 195.325 -112.715 ;
        RECT 194.995 -114.405 195.325 -114.075 ;
        RECT 194.995 -115.765 195.325 -115.435 ;
        RECT 194.995 -117.125 195.325 -116.795 ;
        RECT 194.995 -118.485 195.325 -118.155 ;
        RECT 194.995 -119.845 195.325 -119.515 ;
        RECT 194.995 -121.205 195.325 -120.875 ;
        RECT 194.995 -122.565 195.325 -122.235 ;
        RECT 194.995 -123.925 195.325 -123.595 ;
        RECT 194.995 -125.285 195.325 -124.955 ;
        RECT 194.995 -126.645 195.325 -126.315 ;
        RECT 194.995 -128.005 195.325 -127.675 ;
        RECT 194.995 -129.365 195.325 -129.035 ;
        RECT 194.995 -130.725 195.325 -130.395 ;
        RECT 194.995 -132.085 195.325 -131.755 ;
        RECT 194.995 -133.445 195.325 -133.115 ;
        RECT 194.995 -134.805 195.325 -134.475 ;
        RECT 194.995 -136.165 195.325 -135.835 ;
        RECT 194.995 -137.525 195.325 -137.195 ;
        RECT 194.995 -138.885 195.325 -138.555 ;
        RECT 194.995 -140.245 195.325 -139.915 ;
        RECT 194.995 -141.605 195.325 -141.275 ;
        RECT 194.995 -142.965 195.325 -142.635 ;
        RECT 194.995 -144.325 195.325 -143.995 ;
        RECT 194.995 -145.685 195.325 -145.355 ;
        RECT 194.995 -147.045 195.325 -146.715 ;
        RECT 194.995 -148.405 195.325 -148.075 ;
        RECT 194.995 -149.765 195.325 -149.435 ;
        RECT 194.995 -151.125 195.325 -150.795 ;
        RECT 194.995 -152.485 195.325 -152.155 ;
        RECT 194.995 -153.845 195.325 -153.515 ;
        RECT 194.995 -155.205 195.325 -154.875 ;
        RECT 194.995 -156.565 195.325 -156.235 ;
        RECT 194.995 -157.925 195.325 -157.595 ;
        RECT 194.995 -159.285 195.325 -158.955 ;
        RECT 194.995 -160.645 195.325 -160.315 ;
        RECT 194.995 -162.005 195.325 -161.675 ;
        RECT 194.995 -163.365 195.325 -163.035 ;
        RECT 194.995 -164.725 195.325 -164.395 ;
        RECT 194.995 -166.085 195.325 -165.755 ;
        RECT 194.995 -167.445 195.325 -167.115 ;
        RECT 194.995 -168.805 195.325 -168.475 ;
        RECT 194.995 -170.165 195.325 -169.835 ;
        RECT 194.995 -171.525 195.325 -171.195 ;
        RECT 194.995 -172.885 195.325 -172.555 ;
        RECT 194.995 -174.245 195.325 -173.915 ;
        RECT 194.995 -175.605 195.325 -175.275 ;
        RECT 194.995 -176.965 195.325 -176.635 ;
        RECT 194.995 -178.325 195.325 -177.995 ;
        RECT 194.995 -179.685 195.325 -179.355 ;
        RECT 194.995 -181.93 195.325 -180.8 ;
        RECT 195 -182.045 195.32 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 241.32 196.685 242.45 ;
        RECT 196.355 239.195 196.685 239.525 ;
        RECT 196.355 237.835 196.685 238.165 ;
        RECT 196.36 237.16 196.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 -1.525 196.685 -1.195 ;
        RECT 196.355 -2.885 196.685 -2.555 ;
        RECT 196.36 -3.56 196.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 196.355 -95.365 196.685 -95.035 ;
        RECT 196.355 -96.725 196.685 -96.395 ;
        RECT 196.355 -98.085 196.685 -97.755 ;
        RECT 196.355 -99.445 196.685 -99.115 ;
        RECT 196.355 -100.805 196.685 -100.475 ;
        RECT 196.355 -102.165 196.685 -101.835 ;
        RECT 196.355 -103.525 196.685 -103.195 ;
        RECT 196.355 -104.885 196.685 -104.555 ;
        RECT 196.355 -106.245 196.685 -105.915 ;
        RECT 196.355 -107.605 196.685 -107.275 ;
        RECT 196.355 -108.965 196.685 -108.635 ;
        RECT 196.355 -110.325 196.685 -109.995 ;
        RECT 196.355 -111.685 196.685 -111.355 ;
        RECT 196.355 -113.045 196.685 -112.715 ;
        RECT 196.355 -114.405 196.685 -114.075 ;
        RECT 196.355 -115.765 196.685 -115.435 ;
        RECT 196.355 -117.125 196.685 -116.795 ;
        RECT 196.355 -118.485 196.685 -118.155 ;
        RECT 196.355 -119.845 196.685 -119.515 ;
        RECT 196.355 -121.205 196.685 -120.875 ;
        RECT 196.355 -122.565 196.685 -122.235 ;
        RECT 196.355 -123.925 196.685 -123.595 ;
        RECT 196.355 -125.285 196.685 -124.955 ;
        RECT 196.355 -126.645 196.685 -126.315 ;
        RECT 196.355 -128.005 196.685 -127.675 ;
        RECT 196.355 -129.365 196.685 -129.035 ;
        RECT 196.355 -130.725 196.685 -130.395 ;
        RECT 196.355 -132.085 196.685 -131.755 ;
        RECT 196.355 -133.445 196.685 -133.115 ;
        RECT 196.355 -134.805 196.685 -134.475 ;
        RECT 196.355 -136.165 196.685 -135.835 ;
        RECT 196.355 -137.525 196.685 -137.195 ;
        RECT 196.355 -138.885 196.685 -138.555 ;
        RECT 196.355 -140.245 196.685 -139.915 ;
        RECT 196.355 -141.605 196.685 -141.275 ;
        RECT 196.355 -142.965 196.685 -142.635 ;
        RECT 196.355 -144.325 196.685 -143.995 ;
        RECT 196.355 -145.685 196.685 -145.355 ;
        RECT 196.355 -147.045 196.685 -146.715 ;
        RECT 196.355 -148.405 196.685 -148.075 ;
        RECT 196.355 -149.765 196.685 -149.435 ;
        RECT 196.355 -151.125 196.685 -150.795 ;
        RECT 196.355 -152.485 196.685 -152.155 ;
        RECT 196.355 -153.845 196.685 -153.515 ;
        RECT 196.355 -155.205 196.685 -154.875 ;
        RECT 196.355 -156.565 196.685 -156.235 ;
        RECT 196.355 -157.925 196.685 -157.595 ;
        RECT 196.355 -159.285 196.685 -158.955 ;
        RECT 196.355 -160.645 196.685 -160.315 ;
        RECT 196.355 -162.005 196.685 -161.675 ;
        RECT 196.355 -163.365 196.685 -163.035 ;
        RECT 196.355 -164.725 196.685 -164.395 ;
        RECT 196.355 -166.085 196.685 -165.755 ;
        RECT 196.355 -167.445 196.685 -167.115 ;
        RECT 196.355 -168.805 196.685 -168.475 ;
        RECT 196.355 -170.165 196.685 -169.835 ;
        RECT 196.355 -171.525 196.685 -171.195 ;
        RECT 196.355 -172.885 196.685 -172.555 ;
        RECT 196.355 -174.245 196.685 -173.915 ;
        RECT 196.355 -175.605 196.685 -175.275 ;
        RECT 196.355 -176.965 196.685 -176.635 ;
        RECT 196.355 -178.325 196.685 -177.995 ;
        RECT 196.355 -179.685 196.685 -179.355 ;
        RECT 196.355 -181.93 196.685 -180.8 ;
        RECT 196.36 -182.045 196.68 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 241.32 198.045 242.45 ;
        RECT 197.715 239.195 198.045 239.525 ;
        RECT 197.715 237.835 198.045 238.165 ;
        RECT 197.72 237.16 198.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 -1.525 198.045 -1.195 ;
        RECT 197.715 -2.885 198.045 -2.555 ;
        RECT 197.72 -3.56 198.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 197.715 -95.365 198.045 -95.035 ;
        RECT 197.715 -96.725 198.045 -96.395 ;
        RECT 197.715 -98.085 198.045 -97.755 ;
        RECT 197.715 -99.445 198.045 -99.115 ;
        RECT 197.715 -100.805 198.045 -100.475 ;
        RECT 197.715 -102.165 198.045 -101.835 ;
        RECT 197.715 -103.525 198.045 -103.195 ;
        RECT 197.715 -104.885 198.045 -104.555 ;
        RECT 197.715 -106.245 198.045 -105.915 ;
        RECT 197.715 -107.605 198.045 -107.275 ;
        RECT 197.715 -108.965 198.045 -108.635 ;
        RECT 197.715 -110.325 198.045 -109.995 ;
        RECT 197.715 -111.685 198.045 -111.355 ;
        RECT 197.715 -113.045 198.045 -112.715 ;
        RECT 197.715 -114.405 198.045 -114.075 ;
        RECT 197.715 -115.765 198.045 -115.435 ;
        RECT 197.715 -117.125 198.045 -116.795 ;
        RECT 197.715 -118.485 198.045 -118.155 ;
        RECT 197.715 -119.845 198.045 -119.515 ;
        RECT 197.715 -121.205 198.045 -120.875 ;
        RECT 197.715 -122.565 198.045 -122.235 ;
        RECT 197.715 -123.925 198.045 -123.595 ;
        RECT 197.715 -125.285 198.045 -124.955 ;
        RECT 197.715 -126.645 198.045 -126.315 ;
        RECT 197.715 -128.005 198.045 -127.675 ;
        RECT 197.715 -129.365 198.045 -129.035 ;
        RECT 197.715 -130.725 198.045 -130.395 ;
        RECT 197.715 -132.085 198.045 -131.755 ;
        RECT 197.715 -133.445 198.045 -133.115 ;
        RECT 197.715 -134.805 198.045 -134.475 ;
        RECT 197.715 -136.165 198.045 -135.835 ;
        RECT 197.715 -137.525 198.045 -137.195 ;
        RECT 197.715 -138.885 198.045 -138.555 ;
        RECT 197.715 -140.245 198.045 -139.915 ;
        RECT 197.715 -141.605 198.045 -141.275 ;
        RECT 197.715 -142.965 198.045 -142.635 ;
        RECT 197.715 -144.325 198.045 -143.995 ;
        RECT 197.715 -145.685 198.045 -145.355 ;
        RECT 197.715 -147.045 198.045 -146.715 ;
        RECT 197.715 -148.405 198.045 -148.075 ;
        RECT 197.715 -149.765 198.045 -149.435 ;
        RECT 197.715 -151.125 198.045 -150.795 ;
        RECT 197.715 -152.485 198.045 -152.155 ;
        RECT 197.715 -153.845 198.045 -153.515 ;
        RECT 197.715 -155.205 198.045 -154.875 ;
        RECT 197.715 -156.565 198.045 -156.235 ;
        RECT 197.715 -157.925 198.045 -157.595 ;
        RECT 197.715 -159.285 198.045 -158.955 ;
        RECT 197.715 -160.645 198.045 -160.315 ;
        RECT 197.715 -162.005 198.045 -161.675 ;
        RECT 197.715 -163.365 198.045 -163.035 ;
        RECT 197.715 -164.725 198.045 -164.395 ;
        RECT 197.715 -166.085 198.045 -165.755 ;
        RECT 197.715 -167.445 198.045 -167.115 ;
        RECT 197.715 -168.805 198.045 -168.475 ;
        RECT 197.715 -170.165 198.045 -169.835 ;
        RECT 197.715 -171.525 198.045 -171.195 ;
        RECT 197.715 -172.885 198.045 -172.555 ;
        RECT 197.715 -174.245 198.045 -173.915 ;
        RECT 197.715 -175.605 198.045 -175.275 ;
        RECT 197.715 -176.965 198.045 -176.635 ;
        RECT 197.715 -178.325 198.045 -177.995 ;
        RECT 197.715 -179.685 198.045 -179.355 ;
        RECT 197.715 -181.93 198.045 -180.8 ;
        RECT 197.72 -182.045 198.04 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.075 241.32 199.405 242.45 ;
        RECT 199.075 239.195 199.405 239.525 ;
        RECT 199.075 237.835 199.405 238.165 ;
        RECT 199.08 237.16 199.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.075 -99.445 199.405 -99.115 ;
        RECT 199.075 -100.805 199.405 -100.475 ;
        RECT 199.075 -102.165 199.405 -101.835 ;
        RECT 199.075 -103.525 199.405 -103.195 ;
        RECT 199.075 -104.885 199.405 -104.555 ;
        RECT 199.075 -106.245 199.405 -105.915 ;
        RECT 199.075 -107.605 199.405 -107.275 ;
        RECT 199.075 -108.965 199.405 -108.635 ;
        RECT 199.075 -110.325 199.405 -109.995 ;
        RECT 199.075 -111.685 199.405 -111.355 ;
        RECT 199.075 -113.045 199.405 -112.715 ;
        RECT 199.075 -114.405 199.405 -114.075 ;
        RECT 199.075 -115.765 199.405 -115.435 ;
        RECT 199.075 -117.125 199.405 -116.795 ;
        RECT 199.075 -118.485 199.405 -118.155 ;
        RECT 199.075 -119.845 199.405 -119.515 ;
        RECT 199.075 -121.205 199.405 -120.875 ;
        RECT 199.075 -122.565 199.405 -122.235 ;
        RECT 199.075 -123.925 199.405 -123.595 ;
        RECT 199.075 -125.285 199.405 -124.955 ;
        RECT 199.075 -126.645 199.405 -126.315 ;
        RECT 199.075 -128.005 199.405 -127.675 ;
        RECT 199.075 -129.365 199.405 -129.035 ;
        RECT 199.075 -130.725 199.405 -130.395 ;
        RECT 199.075 -132.085 199.405 -131.755 ;
        RECT 199.075 -133.445 199.405 -133.115 ;
        RECT 199.075 -134.805 199.405 -134.475 ;
        RECT 199.075 -136.165 199.405 -135.835 ;
        RECT 199.075 -137.525 199.405 -137.195 ;
        RECT 199.075 -138.885 199.405 -138.555 ;
        RECT 199.075 -140.245 199.405 -139.915 ;
        RECT 199.075 -141.605 199.405 -141.275 ;
        RECT 199.075 -142.965 199.405 -142.635 ;
        RECT 199.075 -144.325 199.405 -143.995 ;
        RECT 199.075 -145.685 199.405 -145.355 ;
        RECT 199.075 -147.045 199.405 -146.715 ;
        RECT 199.075 -148.405 199.405 -148.075 ;
        RECT 199.075 -149.765 199.405 -149.435 ;
        RECT 199.075 -151.125 199.405 -150.795 ;
        RECT 199.075 -152.485 199.405 -152.155 ;
        RECT 199.075 -153.845 199.405 -153.515 ;
        RECT 199.075 -155.205 199.405 -154.875 ;
        RECT 199.075 -156.565 199.405 -156.235 ;
        RECT 199.075 -157.925 199.405 -157.595 ;
        RECT 199.075 -159.285 199.405 -158.955 ;
        RECT 199.075 -160.645 199.405 -160.315 ;
        RECT 199.075 -162.005 199.405 -161.675 ;
        RECT 199.075 -163.365 199.405 -163.035 ;
        RECT 199.075 -164.725 199.405 -164.395 ;
        RECT 199.075 -166.085 199.405 -165.755 ;
        RECT 199.075 -167.445 199.405 -167.115 ;
        RECT 199.075 -168.805 199.405 -168.475 ;
        RECT 199.075 -170.165 199.405 -169.835 ;
        RECT 199.075 -171.525 199.405 -171.195 ;
        RECT 199.075 -172.885 199.405 -172.555 ;
        RECT 199.075 -174.245 199.405 -173.915 ;
        RECT 199.075 -175.605 199.405 -175.275 ;
        RECT 199.075 -176.965 199.405 -176.635 ;
        RECT 199.075 -178.325 199.405 -177.995 ;
        RECT 199.075 -179.685 199.405 -179.355 ;
        RECT 199.075 -181.93 199.405 -180.8 ;
        RECT 199.08 -182.045 199.4 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 199.51 -98.075 199.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 241.32 200.765 242.45 ;
        RECT 200.435 239.195 200.765 239.525 ;
        RECT 200.435 237.835 200.765 238.165 ;
        RECT 200.44 237.16 200.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 200.435 -1.525 200.765 -1.195 ;
        RECT 200.435 -2.885 200.765 -2.555 ;
        RECT 200.44 -3.56 200.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 241.32 202.125 242.45 ;
        RECT 201.795 239.195 202.125 239.525 ;
        RECT 201.795 237.835 202.125 238.165 ;
        RECT 201.8 237.16 202.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 201.795 -1.525 202.125 -1.195 ;
        RECT 201.795 -2.885 202.125 -2.555 ;
        RECT 201.8 -3.56 202.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 241.32 203.485 242.45 ;
        RECT 203.155 239.195 203.485 239.525 ;
        RECT 203.155 237.835 203.485 238.165 ;
        RECT 203.16 237.16 203.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 -1.525 203.485 -1.195 ;
        RECT 203.155 -2.885 203.485 -2.555 ;
        RECT 203.16 -3.56 203.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 203.155 -95.365 203.485 -95.035 ;
        RECT 203.155 -96.725 203.485 -96.395 ;
        RECT 203.155 -98.085 203.485 -97.755 ;
        RECT 203.155 -99.445 203.485 -99.115 ;
        RECT 203.155 -100.805 203.485 -100.475 ;
        RECT 203.155 -102.165 203.485 -101.835 ;
        RECT 203.155 -103.525 203.485 -103.195 ;
        RECT 203.155 -104.885 203.485 -104.555 ;
        RECT 203.155 -106.245 203.485 -105.915 ;
        RECT 203.155 -107.605 203.485 -107.275 ;
        RECT 203.155 -108.965 203.485 -108.635 ;
        RECT 203.155 -110.325 203.485 -109.995 ;
        RECT 203.155 -111.685 203.485 -111.355 ;
        RECT 203.155 -113.045 203.485 -112.715 ;
        RECT 203.155 -114.405 203.485 -114.075 ;
        RECT 203.155 -115.765 203.485 -115.435 ;
        RECT 203.155 -117.125 203.485 -116.795 ;
        RECT 203.155 -118.485 203.485 -118.155 ;
        RECT 203.155 -119.845 203.485 -119.515 ;
        RECT 203.155 -121.205 203.485 -120.875 ;
        RECT 203.155 -122.565 203.485 -122.235 ;
        RECT 203.155 -123.925 203.485 -123.595 ;
        RECT 203.155 -125.285 203.485 -124.955 ;
        RECT 203.155 -126.645 203.485 -126.315 ;
        RECT 203.155 -128.005 203.485 -127.675 ;
        RECT 203.155 -129.365 203.485 -129.035 ;
        RECT 203.155 -130.725 203.485 -130.395 ;
        RECT 203.155 -132.085 203.485 -131.755 ;
        RECT 203.155 -133.445 203.485 -133.115 ;
        RECT 203.155 -134.805 203.485 -134.475 ;
        RECT 203.155 -136.165 203.485 -135.835 ;
        RECT 203.155 -137.525 203.485 -137.195 ;
        RECT 203.155 -138.885 203.485 -138.555 ;
        RECT 203.155 -140.245 203.485 -139.915 ;
        RECT 203.155 -141.605 203.485 -141.275 ;
        RECT 203.155 -142.965 203.485 -142.635 ;
        RECT 203.155 -144.325 203.485 -143.995 ;
        RECT 203.155 -145.685 203.485 -145.355 ;
        RECT 203.155 -147.045 203.485 -146.715 ;
        RECT 203.155 -148.405 203.485 -148.075 ;
        RECT 203.155 -149.765 203.485 -149.435 ;
        RECT 203.155 -151.125 203.485 -150.795 ;
        RECT 203.155 -152.485 203.485 -152.155 ;
        RECT 203.155 -153.845 203.485 -153.515 ;
        RECT 203.155 -155.205 203.485 -154.875 ;
        RECT 203.155 -156.565 203.485 -156.235 ;
        RECT 203.155 -157.925 203.485 -157.595 ;
        RECT 203.155 -159.285 203.485 -158.955 ;
        RECT 203.155 -160.645 203.485 -160.315 ;
        RECT 203.155 -162.005 203.485 -161.675 ;
        RECT 203.155 -163.365 203.485 -163.035 ;
        RECT 203.155 -164.725 203.485 -164.395 ;
        RECT 203.155 -166.085 203.485 -165.755 ;
        RECT 203.155 -167.445 203.485 -167.115 ;
        RECT 203.155 -168.805 203.485 -168.475 ;
        RECT 203.155 -170.165 203.485 -169.835 ;
        RECT 203.155 -171.525 203.485 -171.195 ;
        RECT 203.155 -172.885 203.485 -172.555 ;
        RECT 203.155 -174.245 203.485 -173.915 ;
        RECT 203.155 -175.605 203.485 -175.275 ;
        RECT 203.155 -176.965 203.485 -176.635 ;
        RECT 203.155 -178.325 203.485 -177.995 ;
        RECT 203.155 -179.685 203.485 -179.355 ;
        RECT 203.155 -181.93 203.485 -180.8 ;
        RECT 203.16 -182.045 203.48 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 241.32 204.845 242.45 ;
        RECT 204.515 239.195 204.845 239.525 ;
        RECT 204.515 237.835 204.845 238.165 ;
        RECT 204.52 237.16 204.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 -1.525 204.845 -1.195 ;
        RECT 204.515 -2.885 204.845 -2.555 ;
        RECT 204.52 -3.56 204.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 204.515 -95.365 204.845 -95.035 ;
        RECT 204.515 -96.725 204.845 -96.395 ;
        RECT 204.515 -98.085 204.845 -97.755 ;
        RECT 204.515 -99.445 204.845 -99.115 ;
        RECT 204.515 -100.805 204.845 -100.475 ;
        RECT 204.515 -102.165 204.845 -101.835 ;
        RECT 204.515 -103.525 204.845 -103.195 ;
        RECT 204.515 -104.885 204.845 -104.555 ;
        RECT 204.515 -106.245 204.845 -105.915 ;
        RECT 204.515 -107.605 204.845 -107.275 ;
        RECT 204.515 -108.965 204.845 -108.635 ;
        RECT 204.515 -110.325 204.845 -109.995 ;
        RECT 204.515 -111.685 204.845 -111.355 ;
        RECT 204.515 -113.045 204.845 -112.715 ;
        RECT 204.515 -114.405 204.845 -114.075 ;
        RECT 204.515 -115.765 204.845 -115.435 ;
        RECT 204.515 -117.125 204.845 -116.795 ;
        RECT 204.515 -118.485 204.845 -118.155 ;
        RECT 204.515 -119.845 204.845 -119.515 ;
        RECT 204.515 -121.205 204.845 -120.875 ;
        RECT 204.515 -122.565 204.845 -122.235 ;
        RECT 204.515 -123.925 204.845 -123.595 ;
        RECT 204.515 -125.285 204.845 -124.955 ;
        RECT 204.515 -126.645 204.845 -126.315 ;
        RECT 204.515 -128.005 204.845 -127.675 ;
        RECT 204.515 -129.365 204.845 -129.035 ;
        RECT 204.515 -130.725 204.845 -130.395 ;
        RECT 204.515 -132.085 204.845 -131.755 ;
        RECT 204.515 -133.445 204.845 -133.115 ;
        RECT 204.515 -134.805 204.845 -134.475 ;
        RECT 204.515 -136.165 204.845 -135.835 ;
        RECT 204.515 -137.525 204.845 -137.195 ;
        RECT 204.515 -138.885 204.845 -138.555 ;
        RECT 204.515 -140.245 204.845 -139.915 ;
        RECT 204.515 -141.605 204.845 -141.275 ;
        RECT 204.515 -142.965 204.845 -142.635 ;
        RECT 204.515 -144.325 204.845 -143.995 ;
        RECT 204.515 -145.685 204.845 -145.355 ;
        RECT 204.515 -147.045 204.845 -146.715 ;
        RECT 204.515 -148.405 204.845 -148.075 ;
        RECT 204.515 -149.765 204.845 -149.435 ;
        RECT 204.515 -151.125 204.845 -150.795 ;
        RECT 204.515 -152.485 204.845 -152.155 ;
        RECT 204.515 -153.845 204.845 -153.515 ;
        RECT 204.515 -155.205 204.845 -154.875 ;
        RECT 204.515 -156.565 204.845 -156.235 ;
        RECT 204.515 -157.925 204.845 -157.595 ;
        RECT 204.515 -159.285 204.845 -158.955 ;
        RECT 204.515 -160.645 204.845 -160.315 ;
        RECT 204.515 -162.005 204.845 -161.675 ;
        RECT 204.515 -163.365 204.845 -163.035 ;
        RECT 204.515 -164.725 204.845 -164.395 ;
        RECT 204.515 -166.085 204.845 -165.755 ;
        RECT 204.515 -167.445 204.845 -167.115 ;
        RECT 204.515 -168.805 204.845 -168.475 ;
        RECT 204.515 -170.165 204.845 -169.835 ;
        RECT 204.515 -171.525 204.845 -171.195 ;
        RECT 204.515 -172.885 204.845 -172.555 ;
        RECT 204.515 -174.245 204.845 -173.915 ;
        RECT 204.515 -175.605 204.845 -175.275 ;
        RECT 204.515 -176.965 204.845 -176.635 ;
        RECT 204.515 -178.325 204.845 -177.995 ;
        RECT 204.515 -179.685 204.845 -179.355 ;
        RECT 204.515 -181.93 204.845 -180.8 ;
        RECT 204.52 -182.045 204.84 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.875 241.32 206.205 242.45 ;
        RECT 205.875 239.195 206.205 239.525 ;
        RECT 205.875 237.835 206.205 238.165 ;
        RECT 205.88 237.16 206.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.875 -1.525 206.205 -1.195 ;
        RECT 205.875 -2.885 206.205 -2.555 ;
        RECT 205.88 -3.56 206.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 205.875 -95.365 206.205 -95.035 ;
        RECT 205.875 -96.725 206.205 -96.395 ;
        RECT 205.875 -98.085 206.205 -97.755 ;
        RECT 205.875 -99.445 206.205 -99.115 ;
        RECT 205.875 -100.805 206.205 -100.475 ;
        RECT 205.875 -102.165 206.205 -101.835 ;
        RECT 205.875 -103.525 206.205 -103.195 ;
        RECT 205.875 -104.885 206.205 -104.555 ;
        RECT 205.875 -106.245 206.205 -105.915 ;
        RECT 205.875 -107.605 206.205 -107.275 ;
        RECT 205.875 -108.965 206.205 -108.635 ;
        RECT 205.875 -110.325 206.205 -109.995 ;
        RECT 205.875 -111.685 206.205 -111.355 ;
        RECT 205.875 -113.045 206.205 -112.715 ;
        RECT 205.875 -114.405 206.205 -114.075 ;
        RECT 205.875 -115.765 206.205 -115.435 ;
        RECT 205.875 -117.125 206.205 -116.795 ;
        RECT 205.875 -118.485 206.205 -118.155 ;
        RECT 205.875 -119.845 206.205 -119.515 ;
        RECT 205.875 -121.205 206.205 -120.875 ;
        RECT 205.875 -122.565 206.205 -122.235 ;
        RECT 205.875 -123.925 206.205 -123.595 ;
        RECT 205.875 -125.285 206.205 -124.955 ;
        RECT 205.875 -126.645 206.205 -126.315 ;
        RECT 205.875 -128.005 206.205 -127.675 ;
        RECT 205.875 -129.365 206.205 -129.035 ;
        RECT 205.875 -130.725 206.205 -130.395 ;
        RECT 205.875 -132.085 206.205 -131.755 ;
        RECT 205.875 -133.445 206.205 -133.115 ;
        RECT 205.875 -134.805 206.205 -134.475 ;
        RECT 205.875 -136.165 206.205 -135.835 ;
        RECT 205.875 -137.525 206.205 -137.195 ;
        RECT 205.875 -138.885 206.205 -138.555 ;
        RECT 205.875 -140.245 206.205 -139.915 ;
        RECT 205.875 -141.605 206.205 -141.275 ;
        RECT 205.875 -142.965 206.205 -142.635 ;
        RECT 205.875 -144.325 206.205 -143.995 ;
        RECT 205.875 -145.685 206.205 -145.355 ;
        RECT 205.875 -147.045 206.205 -146.715 ;
        RECT 205.875 -148.405 206.205 -148.075 ;
        RECT 205.875 -149.765 206.205 -149.435 ;
        RECT 205.875 -151.125 206.205 -150.795 ;
        RECT 205.875 -152.485 206.205 -152.155 ;
        RECT 205.875 -153.845 206.205 -153.515 ;
        RECT 205.875 -155.205 206.205 -154.875 ;
        RECT 205.875 -156.565 206.205 -156.235 ;
        RECT 205.875 -157.925 206.205 -157.595 ;
        RECT 205.875 -159.285 206.205 -158.955 ;
        RECT 205.875 -160.645 206.205 -160.315 ;
        RECT 205.875 -162.005 206.205 -161.675 ;
        RECT 205.875 -163.365 206.205 -163.035 ;
        RECT 205.875 -164.725 206.205 -164.395 ;
        RECT 205.875 -166.085 206.205 -165.755 ;
        RECT 205.875 -167.445 206.205 -167.115 ;
        RECT 205.875 -168.805 206.205 -168.475 ;
        RECT 205.875 -170.165 206.205 -169.835 ;
        RECT 205.875 -171.525 206.205 -171.195 ;
        RECT 205.875 -172.885 206.205 -172.555 ;
        RECT 205.875 -174.245 206.205 -173.915 ;
        RECT 205.875 -175.605 206.205 -175.275 ;
        RECT 205.875 -176.965 206.205 -176.635 ;
        RECT 205.875 -178.325 206.205 -177.995 ;
        RECT 205.875 -179.685 206.205 -179.355 ;
        RECT 205.875 -181.93 206.205 -180.8 ;
        RECT 205.88 -182.045 206.2 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 241.32 207.565 242.45 ;
        RECT 207.235 239.195 207.565 239.525 ;
        RECT 207.235 237.835 207.565 238.165 ;
        RECT 207.24 237.16 207.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 -1.525 207.565 -1.195 ;
        RECT 207.235 -2.885 207.565 -2.555 ;
        RECT 207.24 -3.56 207.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 207.235 -95.365 207.565 -95.035 ;
        RECT 207.235 -96.725 207.565 -96.395 ;
        RECT 207.235 -98.085 207.565 -97.755 ;
        RECT 207.235 -99.445 207.565 -99.115 ;
        RECT 207.235 -100.805 207.565 -100.475 ;
        RECT 207.235 -102.165 207.565 -101.835 ;
        RECT 207.235 -103.525 207.565 -103.195 ;
        RECT 207.235 -104.885 207.565 -104.555 ;
        RECT 207.235 -106.245 207.565 -105.915 ;
        RECT 207.235 -107.605 207.565 -107.275 ;
        RECT 207.235 -108.965 207.565 -108.635 ;
        RECT 207.235 -110.325 207.565 -109.995 ;
        RECT 207.235 -111.685 207.565 -111.355 ;
        RECT 207.235 -113.045 207.565 -112.715 ;
        RECT 207.235 -114.405 207.565 -114.075 ;
        RECT 207.235 -115.765 207.565 -115.435 ;
        RECT 207.235 -117.125 207.565 -116.795 ;
        RECT 207.235 -118.485 207.565 -118.155 ;
        RECT 207.235 -119.845 207.565 -119.515 ;
        RECT 207.235 -121.205 207.565 -120.875 ;
        RECT 207.235 -122.565 207.565 -122.235 ;
        RECT 207.235 -123.925 207.565 -123.595 ;
        RECT 207.235 -125.285 207.565 -124.955 ;
        RECT 207.235 -126.645 207.565 -126.315 ;
        RECT 207.235 -128.005 207.565 -127.675 ;
        RECT 207.235 -129.365 207.565 -129.035 ;
        RECT 207.235 -130.725 207.565 -130.395 ;
        RECT 207.235 -132.085 207.565 -131.755 ;
        RECT 207.235 -133.445 207.565 -133.115 ;
        RECT 207.235 -134.805 207.565 -134.475 ;
        RECT 207.235 -136.165 207.565 -135.835 ;
        RECT 207.235 -137.525 207.565 -137.195 ;
        RECT 207.235 -138.885 207.565 -138.555 ;
        RECT 207.235 -140.245 207.565 -139.915 ;
        RECT 207.235 -141.605 207.565 -141.275 ;
        RECT 207.235 -142.965 207.565 -142.635 ;
        RECT 207.235 -144.325 207.565 -143.995 ;
        RECT 207.235 -145.685 207.565 -145.355 ;
        RECT 207.235 -147.045 207.565 -146.715 ;
        RECT 207.235 -148.405 207.565 -148.075 ;
        RECT 207.235 -149.765 207.565 -149.435 ;
        RECT 207.235 -151.125 207.565 -150.795 ;
        RECT 207.235 -152.485 207.565 -152.155 ;
        RECT 207.235 -153.845 207.565 -153.515 ;
        RECT 207.235 -155.205 207.565 -154.875 ;
        RECT 207.235 -156.565 207.565 -156.235 ;
        RECT 207.235 -157.925 207.565 -157.595 ;
        RECT 207.235 -159.285 207.565 -158.955 ;
        RECT 207.235 -160.645 207.565 -160.315 ;
        RECT 207.235 -162.005 207.565 -161.675 ;
        RECT 207.235 -163.365 207.565 -163.035 ;
        RECT 207.235 -164.725 207.565 -164.395 ;
        RECT 207.235 -166.085 207.565 -165.755 ;
        RECT 207.235 -167.445 207.565 -167.115 ;
        RECT 207.235 -168.805 207.565 -168.475 ;
        RECT 207.235 -170.165 207.565 -169.835 ;
        RECT 207.235 -171.525 207.565 -171.195 ;
        RECT 207.235 -172.885 207.565 -172.555 ;
        RECT 207.235 -174.245 207.565 -173.915 ;
        RECT 207.235 -175.605 207.565 -175.275 ;
        RECT 207.235 -176.965 207.565 -176.635 ;
        RECT 207.235 -178.325 207.565 -177.995 ;
        RECT 207.235 -179.685 207.565 -179.355 ;
        RECT 207.235 -181.93 207.565 -180.8 ;
        RECT 207.24 -182.045 207.56 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 241.32 208.925 242.45 ;
        RECT 208.595 239.195 208.925 239.525 ;
        RECT 208.595 237.835 208.925 238.165 ;
        RECT 208.6 237.16 208.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 -1.525 208.925 -1.195 ;
        RECT 208.595 -2.885 208.925 -2.555 ;
        RECT 208.6 -3.56 208.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 208.595 -95.365 208.925 -95.035 ;
        RECT 208.595 -96.725 208.925 -96.395 ;
        RECT 208.595 -98.085 208.925 -97.755 ;
        RECT 208.595 -99.445 208.925 -99.115 ;
        RECT 208.595 -100.805 208.925 -100.475 ;
        RECT 208.595 -102.165 208.925 -101.835 ;
        RECT 208.595 -103.525 208.925 -103.195 ;
        RECT 208.595 -104.885 208.925 -104.555 ;
        RECT 208.595 -106.245 208.925 -105.915 ;
        RECT 208.595 -107.605 208.925 -107.275 ;
        RECT 208.595 -108.965 208.925 -108.635 ;
        RECT 208.595 -110.325 208.925 -109.995 ;
        RECT 208.595 -111.685 208.925 -111.355 ;
        RECT 208.595 -113.045 208.925 -112.715 ;
        RECT 208.595 -114.405 208.925 -114.075 ;
        RECT 208.595 -115.765 208.925 -115.435 ;
        RECT 208.595 -117.125 208.925 -116.795 ;
        RECT 208.595 -118.485 208.925 -118.155 ;
        RECT 208.595 -119.845 208.925 -119.515 ;
        RECT 208.595 -121.205 208.925 -120.875 ;
        RECT 208.595 -122.565 208.925 -122.235 ;
        RECT 208.595 -123.925 208.925 -123.595 ;
        RECT 208.595 -125.285 208.925 -124.955 ;
        RECT 208.595 -126.645 208.925 -126.315 ;
        RECT 208.595 -128.005 208.925 -127.675 ;
        RECT 208.595 -129.365 208.925 -129.035 ;
        RECT 208.595 -130.725 208.925 -130.395 ;
        RECT 208.595 -132.085 208.925 -131.755 ;
        RECT 208.595 -133.445 208.925 -133.115 ;
        RECT 208.595 -134.805 208.925 -134.475 ;
        RECT 208.595 -136.165 208.925 -135.835 ;
        RECT 208.595 -137.525 208.925 -137.195 ;
        RECT 208.595 -138.885 208.925 -138.555 ;
        RECT 208.595 -140.245 208.925 -139.915 ;
        RECT 208.595 -141.605 208.925 -141.275 ;
        RECT 208.595 -142.965 208.925 -142.635 ;
        RECT 208.595 -144.325 208.925 -143.995 ;
        RECT 208.595 -145.685 208.925 -145.355 ;
        RECT 208.595 -147.045 208.925 -146.715 ;
        RECT 208.595 -148.405 208.925 -148.075 ;
        RECT 208.595 -149.765 208.925 -149.435 ;
        RECT 208.595 -151.125 208.925 -150.795 ;
        RECT 208.595 -152.485 208.925 -152.155 ;
        RECT 208.595 -153.845 208.925 -153.515 ;
        RECT 208.595 -155.205 208.925 -154.875 ;
        RECT 208.595 -156.565 208.925 -156.235 ;
        RECT 208.595 -157.925 208.925 -157.595 ;
        RECT 208.595 -159.285 208.925 -158.955 ;
        RECT 208.595 -160.645 208.925 -160.315 ;
        RECT 208.595 -162.005 208.925 -161.675 ;
        RECT 208.595 -163.365 208.925 -163.035 ;
        RECT 208.595 -164.725 208.925 -164.395 ;
        RECT 208.595 -166.085 208.925 -165.755 ;
        RECT 208.595 -167.445 208.925 -167.115 ;
        RECT 208.595 -168.805 208.925 -168.475 ;
        RECT 208.595 -170.165 208.925 -169.835 ;
        RECT 208.595 -171.525 208.925 -171.195 ;
        RECT 208.595 -172.885 208.925 -172.555 ;
        RECT 208.595 -174.245 208.925 -173.915 ;
        RECT 208.595 -175.605 208.925 -175.275 ;
        RECT 208.595 -176.965 208.925 -176.635 ;
        RECT 208.595 -178.325 208.925 -177.995 ;
        RECT 208.595 -179.685 208.925 -179.355 ;
        RECT 208.595 -181.93 208.925 -180.8 ;
        RECT 208.6 -182.045 208.92 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.955 241.32 210.285 242.45 ;
        RECT 209.955 239.195 210.285 239.525 ;
        RECT 209.955 237.835 210.285 238.165 ;
        RECT 209.96 237.16 210.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 209.955 -99.445 210.285 -99.115 ;
        RECT 209.955 -100.805 210.285 -100.475 ;
        RECT 209.955 -102.165 210.285 -101.835 ;
        RECT 209.955 -103.525 210.285 -103.195 ;
        RECT 209.955 -104.885 210.285 -104.555 ;
        RECT 209.955 -106.245 210.285 -105.915 ;
        RECT 209.955 -107.605 210.285 -107.275 ;
        RECT 209.955 -108.965 210.285 -108.635 ;
        RECT 209.955 -110.325 210.285 -109.995 ;
        RECT 209.955 -111.685 210.285 -111.355 ;
        RECT 209.955 -113.045 210.285 -112.715 ;
        RECT 209.955 -114.405 210.285 -114.075 ;
        RECT 209.955 -115.765 210.285 -115.435 ;
        RECT 209.955 -117.125 210.285 -116.795 ;
        RECT 209.955 -118.485 210.285 -118.155 ;
        RECT 209.955 -119.845 210.285 -119.515 ;
        RECT 209.955 -121.205 210.285 -120.875 ;
        RECT 209.955 -122.565 210.285 -122.235 ;
        RECT 209.955 -123.925 210.285 -123.595 ;
        RECT 209.955 -125.285 210.285 -124.955 ;
        RECT 209.955 -126.645 210.285 -126.315 ;
        RECT 209.955 -128.005 210.285 -127.675 ;
        RECT 209.955 -129.365 210.285 -129.035 ;
        RECT 209.955 -130.725 210.285 -130.395 ;
        RECT 209.955 -132.085 210.285 -131.755 ;
        RECT 209.955 -133.445 210.285 -133.115 ;
        RECT 209.955 -134.805 210.285 -134.475 ;
        RECT 209.955 -136.165 210.285 -135.835 ;
        RECT 209.955 -137.525 210.285 -137.195 ;
        RECT 209.955 -138.885 210.285 -138.555 ;
        RECT 209.955 -140.245 210.285 -139.915 ;
        RECT 209.955 -141.605 210.285 -141.275 ;
        RECT 209.955 -142.965 210.285 -142.635 ;
        RECT 209.955 -144.325 210.285 -143.995 ;
        RECT 209.955 -145.685 210.285 -145.355 ;
        RECT 209.955 -147.045 210.285 -146.715 ;
        RECT 209.955 -148.405 210.285 -148.075 ;
        RECT 209.955 -149.765 210.285 -149.435 ;
        RECT 209.955 -151.125 210.285 -150.795 ;
        RECT 209.955 -152.485 210.285 -152.155 ;
        RECT 209.955 -153.845 210.285 -153.515 ;
        RECT 209.955 -155.205 210.285 -154.875 ;
        RECT 209.955 -156.565 210.285 -156.235 ;
        RECT 209.955 -157.925 210.285 -157.595 ;
        RECT 209.955 -159.285 210.285 -158.955 ;
        RECT 209.955 -160.645 210.285 -160.315 ;
        RECT 209.955 -162.005 210.285 -161.675 ;
        RECT 209.955 -163.365 210.285 -163.035 ;
        RECT 209.955 -164.725 210.285 -164.395 ;
        RECT 209.955 -166.085 210.285 -165.755 ;
        RECT 209.955 -167.445 210.285 -167.115 ;
        RECT 209.955 -168.805 210.285 -168.475 ;
        RECT 209.955 -170.165 210.285 -169.835 ;
        RECT 209.955 -171.525 210.285 -171.195 ;
        RECT 209.955 -172.885 210.285 -172.555 ;
        RECT 209.955 -174.245 210.285 -173.915 ;
        RECT 209.955 -175.605 210.285 -175.275 ;
        RECT 209.955 -176.965 210.285 -176.635 ;
        RECT 209.955 -178.325 210.285 -177.995 ;
        RECT 209.955 -179.685 210.285 -179.355 ;
        RECT 209.955 -181.93 210.285 -180.8 ;
        RECT 209.96 -182.045 210.28 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 210.41 -98.075 210.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.315 241.32 211.645 242.45 ;
        RECT 211.315 239.195 211.645 239.525 ;
        RECT 211.315 237.835 211.645 238.165 ;
        RECT 211.32 237.16 211.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 211.315 -1.525 211.645 -1.195 ;
        RECT 211.315 -2.885 211.645 -2.555 ;
        RECT 211.32 -3.56 211.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.675 241.32 213.005 242.45 ;
        RECT 212.675 239.195 213.005 239.525 ;
        RECT 212.675 237.835 213.005 238.165 ;
        RECT 212.68 237.16 213 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 212.675 -1.525 213.005 -1.195 ;
        RECT 212.675 -2.885 213.005 -2.555 ;
        RECT 212.68 -3.56 213 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.035 241.32 214.365 242.45 ;
        RECT 214.035 239.195 214.365 239.525 ;
        RECT 214.035 237.835 214.365 238.165 ;
        RECT 214.04 237.16 214.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.035 -1.525 214.365 -1.195 ;
        RECT 214.035 -2.885 214.365 -2.555 ;
        RECT 214.04 -3.56 214.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 214.035 -95.365 214.365 -95.035 ;
        RECT 214.035 -96.725 214.365 -96.395 ;
        RECT 214.035 -98.085 214.365 -97.755 ;
        RECT 214.035 -99.445 214.365 -99.115 ;
        RECT 214.035 -100.805 214.365 -100.475 ;
        RECT 214.035 -102.165 214.365 -101.835 ;
        RECT 214.035 -103.525 214.365 -103.195 ;
        RECT 214.035 -104.885 214.365 -104.555 ;
        RECT 214.035 -106.245 214.365 -105.915 ;
        RECT 214.035 -107.605 214.365 -107.275 ;
        RECT 214.035 -108.965 214.365 -108.635 ;
        RECT 214.035 -110.325 214.365 -109.995 ;
        RECT 214.035 -111.685 214.365 -111.355 ;
        RECT 214.035 -113.045 214.365 -112.715 ;
        RECT 214.035 -114.405 214.365 -114.075 ;
        RECT 214.035 -115.765 214.365 -115.435 ;
        RECT 214.035 -117.125 214.365 -116.795 ;
        RECT 214.035 -118.485 214.365 -118.155 ;
        RECT 214.035 -119.845 214.365 -119.515 ;
        RECT 214.035 -121.205 214.365 -120.875 ;
        RECT 214.035 -122.565 214.365 -122.235 ;
        RECT 214.035 -123.925 214.365 -123.595 ;
        RECT 214.035 -125.285 214.365 -124.955 ;
        RECT 214.035 -126.645 214.365 -126.315 ;
        RECT 214.035 -128.005 214.365 -127.675 ;
        RECT 214.035 -129.365 214.365 -129.035 ;
        RECT 214.035 -130.725 214.365 -130.395 ;
        RECT 214.035 -132.085 214.365 -131.755 ;
        RECT 214.035 -133.445 214.365 -133.115 ;
        RECT 214.035 -134.805 214.365 -134.475 ;
        RECT 214.035 -136.165 214.365 -135.835 ;
        RECT 214.035 -137.525 214.365 -137.195 ;
        RECT 214.035 -138.885 214.365 -138.555 ;
        RECT 214.035 -140.245 214.365 -139.915 ;
        RECT 214.035 -141.605 214.365 -141.275 ;
        RECT 214.035 -142.965 214.365 -142.635 ;
        RECT 214.035 -144.325 214.365 -143.995 ;
        RECT 214.035 -145.685 214.365 -145.355 ;
        RECT 214.035 -147.045 214.365 -146.715 ;
        RECT 214.035 -148.405 214.365 -148.075 ;
        RECT 214.035 -149.765 214.365 -149.435 ;
        RECT 214.035 -151.125 214.365 -150.795 ;
        RECT 214.035 -152.485 214.365 -152.155 ;
        RECT 214.035 -153.845 214.365 -153.515 ;
        RECT 214.035 -155.205 214.365 -154.875 ;
        RECT 214.035 -156.565 214.365 -156.235 ;
        RECT 214.035 -157.925 214.365 -157.595 ;
        RECT 214.035 -159.285 214.365 -158.955 ;
        RECT 214.035 -160.645 214.365 -160.315 ;
        RECT 214.035 -162.005 214.365 -161.675 ;
        RECT 214.035 -163.365 214.365 -163.035 ;
        RECT 214.035 -164.725 214.365 -164.395 ;
        RECT 214.035 -166.085 214.365 -165.755 ;
        RECT 214.035 -167.445 214.365 -167.115 ;
        RECT 214.035 -168.805 214.365 -168.475 ;
        RECT 214.035 -170.165 214.365 -169.835 ;
        RECT 214.035 -171.525 214.365 -171.195 ;
        RECT 214.035 -172.885 214.365 -172.555 ;
        RECT 214.035 -174.245 214.365 -173.915 ;
        RECT 214.035 -175.605 214.365 -175.275 ;
        RECT 214.035 -176.965 214.365 -176.635 ;
        RECT 214.035 -178.325 214.365 -177.995 ;
        RECT 214.035 -179.685 214.365 -179.355 ;
        RECT 214.035 -181.93 214.365 -180.8 ;
        RECT 214.04 -182.045 214.36 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.395 241.32 215.725 242.45 ;
        RECT 215.395 239.195 215.725 239.525 ;
        RECT 215.395 237.835 215.725 238.165 ;
        RECT 215.4 237.16 215.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.395 -1.525 215.725 -1.195 ;
        RECT 215.395 -2.885 215.725 -2.555 ;
        RECT 215.4 -3.56 215.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 215.395 -107.605 215.725 -107.275 ;
        RECT 215.395 -108.965 215.725 -108.635 ;
        RECT 215.395 -110.325 215.725 -109.995 ;
        RECT 215.395 -111.685 215.725 -111.355 ;
        RECT 215.395 -113.045 215.725 -112.715 ;
        RECT 215.395 -114.405 215.725 -114.075 ;
        RECT 215.395 -115.765 215.725 -115.435 ;
        RECT 215.395 -117.125 215.725 -116.795 ;
        RECT 215.395 -118.485 215.725 -118.155 ;
        RECT 215.395 -119.845 215.725 -119.515 ;
        RECT 215.395 -121.205 215.725 -120.875 ;
        RECT 215.395 -122.565 215.725 -122.235 ;
        RECT 215.395 -123.925 215.725 -123.595 ;
        RECT 215.395 -125.285 215.725 -124.955 ;
        RECT 215.395 -126.645 215.725 -126.315 ;
        RECT 215.395 -128.005 215.725 -127.675 ;
        RECT 215.395 -129.365 215.725 -129.035 ;
        RECT 215.395 -130.725 215.725 -130.395 ;
        RECT 215.395 -132.085 215.725 -131.755 ;
        RECT 215.395 -133.445 215.725 -133.115 ;
        RECT 215.395 -134.805 215.725 -134.475 ;
        RECT 215.395 -136.165 215.725 -135.835 ;
        RECT 215.395 -137.525 215.725 -137.195 ;
        RECT 215.395 -138.885 215.725 -138.555 ;
        RECT 215.395 -140.245 215.725 -139.915 ;
        RECT 215.395 -141.605 215.725 -141.275 ;
        RECT 215.395 -142.965 215.725 -142.635 ;
        RECT 215.395 -144.325 215.725 -143.995 ;
        RECT 215.395 -145.685 215.725 -145.355 ;
        RECT 215.395 -147.045 215.725 -146.715 ;
        RECT 215.395 -148.405 215.725 -148.075 ;
        RECT 215.395 -149.765 215.725 -149.435 ;
        RECT 215.395 -151.125 215.725 -150.795 ;
        RECT 215.395 -152.485 215.725 -152.155 ;
        RECT 215.395 -153.845 215.725 -153.515 ;
        RECT 215.395 -155.205 215.725 -154.875 ;
        RECT 215.395 -156.565 215.725 -156.235 ;
        RECT 215.395 -157.925 215.725 -157.595 ;
        RECT 215.395 -159.285 215.725 -158.955 ;
        RECT 215.395 -160.645 215.725 -160.315 ;
        RECT 215.395 -162.005 215.725 -161.675 ;
        RECT 215.395 -163.365 215.725 -163.035 ;
        RECT 215.395 -164.725 215.725 -164.395 ;
        RECT 215.395 -166.085 215.725 -165.755 ;
        RECT 215.395 -167.445 215.725 -167.115 ;
        RECT 215.395 -168.805 215.725 -168.475 ;
        RECT 215.395 -170.165 215.725 -169.835 ;
        RECT 215.395 -171.525 215.725 -171.195 ;
        RECT 215.395 -172.885 215.725 -172.555 ;
        RECT 215.395 -174.245 215.725 -173.915 ;
        RECT 215.395 -175.605 215.725 -175.275 ;
        RECT 215.395 -176.965 215.725 -176.635 ;
        RECT 215.395 -178.325 215.725 -177.995 ;
        RECT 215.395 -179.685 215.725 -179.355 ;
        RECT 215.395 -181.93 215.725 -180.8 ;
        RECT 215.4 -182.045 215.72 -95.035 ;
        RECT 215.395 -95.365 215.725 -95.035 ;
        RECT 215.395 -96.725 215.725 -96.395 ;
        RECT 215.395 -98.085 215.725 -97.755 ;
        RECT 215.395 -99.445 215.725 -99.115 ;
        RECT 215.395 -100.805 215.725 -100.475 ;
        RECT 215.395 -102.165 215.725 -101.835 ;
        RECT 215.395 -103.525 215.725 -103.195 ;
        RECT 215.395 -104.885 215.725 -104.555 ;
        RECT 215.395 -106.245 215.725 -105.915 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 241.32 166.765 242.45 ;
        RECT 166.435 239.195 166.765 239.525 ;
        RECT 166.435 237.835 166.765 238.165 ;
        RECT 166.44 237.16 166.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.435 -99.445 166.765 -99.115 ;
        RECT 166.435 -100.805 166.765 -100.475 ;
        RECT 166.435 -102.165 166.765 -101.835 ;
        RECT 166.435 -103.525 166.765 -103.195 ;
        RECT 166.435 -104.885 166.765 -104.555 ;
        RECT 166.435 -106.245 166.765 -105.915 ;
        RECT 166.435 -107.605 166.765 -107.275 ;
        RECT 166.435 -108.965 166.765 -108.635 ;
        RECT 166.435 -110.325 166.765 -109.995 ;
        RECT 166.435 -111.685 166.765 -111.355 ;
        RECT 166.435 -113.045 166.765 -112.715 ;
        RECT 166.435 -114.405 166.765 -114.075 ;
        RECT 166.435 -115.765 166.765 -115.435 ;
        RECT 166.435 -117.125 166.765 -116.795 ;
        RECT 166.435 -118.485 166.765 -118.155 ;
        RECT 166.435 -119.845 166.765 -119.515 ;
        RECT 166.435 -121.205 166.765 -120.875 ;
        RECT 166.435 -122.565 166.765 -122.235 ;
        RECT 166.435 -123.925 166.765 -123.595 ;
        RECT 166.435 -125.285 166.765 -124.955 ;
        RECT 166.435 -126.645 166.765 -126.315 ;
        RECT 166.435 -128.005 166.765 -127.675 ;
        RECT 166.435 -129.365 166.765 -129.035 ;
        RECT 166.435 -130.725 166.765 -130.395 ;
        RECT 166.435 -132.085 166.765 -131.755 ;
        RECT 166.435 -133.445 166.765 -133.115 ;
        RECT 166.435 -134.805 166.765 -134.475 ;
        RECT 166.435 -136.165 166.765 -135.835 ;
        RECT 166.435 -137.525 166.765 -137.195 ;
        RECT 166.435 -138.885 166.765 -138.555 ;
        RECT 166.435 -140.245 166.765 -139.915 ;
        RECT 166.435 -141.605 166.765 -141.275 ;
        RECT 166.435 -142.965 166.765 -142.635 ;
        RECT 166.435 -144.325 166.765 -143.995 ;
        RECT 166.435 -145.685 166.765 -145.355 ;
        RECT 166.435 -147.045 166.765 -146.715 ;
        RECT 166.435 -148.405 166.765 -148.075 ;
        RECT 166.435 -149.765 166.765 -149.435 ;
        RECT 166.435 -151.125 166.765 -150.795 ;
        RECT 166.435 -152.485 166.765 -152.155 ;
        RECT 166.435 -153.845 166.765 -153.515 ;
        RECT 166.435 -155.205 166.765 -154.875 ;
        RECT 166.435 -156.565 166.765 -156.235 ;
        RECT 166.435 -157.925 166.765 -157.595 ;
        RECT 166.435 -159.285 166.765 -158.955 ;
        RECT 166.435 -160.645 166.765 -160.315 ;
        RECT 166.435 -162.005 166.765 -161.675 ;
        RECT 166.435 -163.365 166.765 -163.035 ;
        RECT 166.435 -164.725 166.765 -164.395 ;
        RECT 166.435 -166.085 166.765 -165.755 ;
        RECT 166.435 -167.445 166.765 -167.115 ;
        RECT 166.435 -168.805 166.765 -168.475 ;
        RECT 166.435 -170.165 166.765 -169.835 ;
        RECT 166.435 -171.525 166.765 -171.195 ;
        RECT 166.435 -172.885 166.765 -172.555 ;
        RECT 166.435 -174.245 166.765 -173.915 ;
        RECT 166.435 -175.605 166.765 -175.275 ;
        RECT 166.435 -176.965 166.765 -176.635 ;
        RECT 166.435 -178.325 166.765 -177.995 ;
        RECT 166.435 -179.685 166.765 -179.355 ;
        RECT 166.435 -181.93 166.765 -180.8 ;
        RECT 166.44 -182.045 166.76 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 166.81 -98.075 167.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 241.32 168.125 242.45 ;
        RECT 167.795 239.195 168.125 239.525 ;
        RECT 167.795 237.835 168.125 238.165 ;
        RECT 167.8 237.16 168.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 167.795 -1.525 168.125 -1.195 ;
        RECT 167.795 -2.885 168.125 -2.555 ;
        RECT 167.8 -3.56 168.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 241.32 169.485 242.45 ;
        RECT 169.155 239.195 169.485 239.525 ;
        RECT 169.155 237.835 169.485 238.165 ;
        RECT 169.16 237.16 169.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 169.155 -1.525 169.485 -1.195 ;
        RECT 169.155 -2.885 169.485 -2.555 ;
        RECT 169.16 -3.56 169.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 241.32 170.845 242.45 ;
        RECT 170.515 239.195 170.845 239.525 ;
        RECT 170.515 237.835 170.845 238.165 ;
        RECT 170.52 237.16 170.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 -1.525 170.845 -1.195 ;
        RECT 170.515 -2.885 170.845 -2.555 ;
        RECT 170.52 -3.56 170.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 170.515 -95.365 170.845 -95.035 ;
        RECT 170.515 -96.725 170.845 -96.395 ;
        RECT 170.515 -98.085 170.845 -97.755 ;
        RECT 170.515 -99.445 170.845 -99.115 ;
        RECT 170.515 -100.805 170.845 -100.475 ;
        RECT 170.515 -102.165 170.845 -101.835 ;
        RECT 170.515 -103.525 170.845 -103.195 ;
        RECT 170.515 -104.885 170.845 -104.555 ;
        RECT 170.515 -106.245 170.845 -105.915 ;
        RECT 170.515 -107.605 170.845 -107.275 ;
        RECT 170.515 -108.965 170.845 -108.635 ;
        RECT 170.515 -110.325 170.845 -109.995 ;
        RECT 170.515 -111.685 170.845 -111.355 ;
        RECT 170.515 -113.045 170.845 -112.715 ;
        RECT 170.515 -114.405 170.845 -114.075 ;
        RECT 170.515 -115.765 170.845 -115.435 ;
        RECT 170.515 -117.125 170.845 -116.795 ;
        RECT 170.515 -118.485 170.845 -118.155 ;
        RECT 170.515 -119.845 170.845 -119.515 ;
        RECT 170.515 -121.205 170.845 -120.875 ;
        RECT 170.515 -122.565 170.845 -122.235 ;
        RECT 170.515 -123.925 170.845 -123.595 ;
        RECT 170.515 -125.285 170.845 -124.955 ;
        RECT 170.515 -126.645 170.845 -126.315 ;
        RECT 170.515 -128.005 170.845 -127.675 ;
        RECT 170.515 -129.365 170.845 -129.035 ;
        RECT 170.515 -130.725 170.845 -130.395 ;
        RECT 170.515 -132.085 170.845 -131.755 ;
        RECT 170.515 -133.445 170.845 -133.115 ;
        RECT 170.515 -134.805 170.845 -134.475 ;
        RECT 170.515 -136.165 170.845 -135.835 ;
        RECT 170.515 -137.525 170.845 -137.195 ;
        RECT 170.515 -138.885 170.845 -138.555 ;
        RECT 170.515 -140.245 170.845 -139.915 ;
        RECT 170.515 -141.605 170.845 -141.275 ;
        RECT 170.515 -142.965 170.845 -142.635 ;
        RECT 170.515 -144.325 170.845 -143.995 ;
        RECT 170.515 -145.685 170.845 -145.355 ;
        RECT 170.515 -147.045 170.845 -146.715 ;
        RECT 170.515 -148.405 170.845 -148.075 ;
        RECT 170.515 -149.765 170.845 -149.435 ;
        RECT 170.515 -151.125 170.845 -150.795 ;
        RECT 170.515 -152.485 170.845 -152.155 ;
        RECT 170.515 -153.845 170.845 -153.515 ;
        RECT 170.515 -155.205 170.845 -154.875 ;
        RECT 170.515 -156.565 170.845 -156.235 ;
        RECT 170.515 -157.925 170.845 -157.595 ;
        RECT 170.515 -159.285 170.845 -158.955 ;
        RECT 170.515 -160.645 170.845 -160.315 ;
        RECT 170.515 -162.005 170.845 -161.675 ;
        RECT 170.515 -163.365 170.845 -163.035 ;
        RECT 170.515 -164.725 170.845 -164.395 ;
        RECT 170.515 -166.085 170.845 -165.755 ;
        RECT 170.515 -167.445 170.845 -167.115 ;
        RECT 170.515 -168.805 170.845 -168.475 ;
        RECT 170.515 -170.165 170.845 -169.835 ;
        RECT 170.515 -171.525 170.845 -171.195 ;
        RECT 170.515 -172.885 170.845 -172.555 ;
        RECT 170.515 -174.245 170.845 -173.915 ;
        RECT 170.515 -175.605 170.845 -175.275 ;
        RECT 170.515 -176.965 170.845 -176.635 ;
        RECT 170.515 -178.325 170.845 -177.995 ;
        RECT 170.515 -179.685 170.845 -179.355 ;
        RECT 170.515 -181.93 170.845 -180.8 ;
        RECT 170.52 -182.045 170.84 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 241.32 172.205 242.45 ;
        RECT 171.875 239.195 172.205 239.525 ;
        RECT 171.875 237.835 172.205 238.165 ;
        RECT 171.88 237.16 172.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 -1.525 172.205 -1.195 ;
        RECT 171.875 -2.885 172.205 -2.555 ;
        RECT 171.88 -3.56 172.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 171.875 -95.365 172.205 -95.035 ;
        RECT 171.875 -96.725 172.205 -96.395 ;
        RECT 171.875 -98.085 172.205 -97.755 ;
        RECT 171.875 -99.445 172.205 -99.115 ;
        RECT 171.875 -100.805 172.205 -100.475 ;
        RECT 171.875 -102.165 172.205 -101.835 ;
        RECT 171.875 -103.525 172.205 -103.195 ;
        RECT 171.875 -104.885 172.205 -104.555 ;
        RECT 171.875 -106.245 172.205 -105.915 ;
        RECT 171.875 -107.605 172.205 -107.275 ;
        RECT 171.875 -108.965 172.205 -108.635 ;
        RECT 171.875 -110.325 172.205 -109.995 ;
        RECT 171.875 -111.685 172.205 -111.355 ;
        RECT 171.875 -113.045 172.205 -112.715 ;
        RECT 171.875 -114.405 172.205 -114.075 ;
        RECT 171.875 -115.765 172.205 -115.435 ;
        RECT 171.875 -117.125 172.205 -116.795 ;
        RECT 171.875 -118.485 172.205 -118.155 ;
        RECT 171.875 -119.845 172.205 -119.515 ;
        RECT 171.875 -121.205 172.205 -120.875 ;
        RECT 171.875 -122.565 172.205 -122.235 ;
        RECT 171.875 -123.925 172.205 -123.595 ;
        RECT 171.875 -125.285 172.205 -124.955 ;
        RECT 171.875 -126.645 172.205 -126.315 ;
        RECT 171.875 -128.005 172.205 -127.675 ;
        RECT 171.875 -129.365 172.205 -129.035 ;
        RECT 171.875 -130.725 172.205 -130.395 ;
        RECT 171.875 -132.085 172.205 -131.755 ;
        RECT 171.875 -133.445 172.205 -133.115 ;
        RECT 171.875 -134.805 172.205 -134.475 ;
        RECT 171.875 -136.165 172.205 -135.835 ;
        RECT 171.875 -137.525 172.205 -137.195 ;
        RECT 171.875 -138.885 172.205 -138.555 ;
        RECT 171.875 -140.245 172.205 -139.915 ;
        RECT 171.875 -141.605 172.205 -141.275 ;
        RECT 171.875 -142.965 172.205 -142.635 ;
        RECT 171.875 -144.325 172.205 -143.995 ;
        RECT 171.875 -145.685 172.205 -145.355 ;
        RECT 171.875 -147.045 172.205 -146.715 ;
        RECT 171.875 -148.405 172.205 -148.075 ;
        RECT 171.875 -149.765 172.205 -149.435 ;
        RECT 171.875 -151.125 172.205 -150.795 ;
        RECT 171.875 -152.485 172.205 -152.155 ;
        RECT 171.875 -153.845 172.205 -153.515 ;
        RECT 171.875 -155.205 172.205 -154.875 ;
        RECT 171.875 -156.565 172.205 -156.235 ;
        RECT 171.875 -157.925 172.205 -157.595 ;
        RECT 171.875 -159.285 172.205 -158.955 ;
        RECT 171.875 -160.645 172.205 -160.315 ;
        RECT 171.875 -162.005 172.205 -161.675 ;
        RECT 171.875 -163.365 172.205 -163.035 ;
        RECT 171.875 -164.725 172.205 -164.395 ;
        RECT 171.875 -166.085 172.205 -165.755 ;
        RECT 171.875 -167.445 172.205 -167.115 ;
        RECT 171.875 -168.805 172.205 -168.475 ;
        RECT 171.875 -170.165 172.205 -169.835 ;
        RECT 171.875 -171.525 172.205 -171.195 ;
        RECT 171.875 -172.885 172.205 -172.555 ;
        RECT 171.875 -174.245 172.205 -173.915 ;
        RECT 171.875 -175.605 172.205 -175.275 ;
        RECT 171.875 -176.965 172.205 -176.635 ;
        RECT 171.875 -178.325 172.205 -177.995 ;
        RECT 171.875 -179.685 172.205 -179.355 ;
        RECT 171.875 -181.93 172.205 -180.8 ;
        RECT 171.88 -182.045 172.2 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 241.32 173.565 242.45 ;
        RECT 173.235 239.195 173.565 239.525 ;
        RECT 173.235 237.835 173.565 238.165 ;
        RECT 173.24 237.16 173.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 -1.525 173.565 -1.195 ;
        RECT 173.235 -2.885 173.565 -2.555 ;
        RECT 173.24 -3.56 173.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 173.235 -95.365 173.565 -95.035 ;
        RECT 173.235 -96.725 173.565 -96.395 ;
        RECT 173.235 -98.085 173.565 -97.755 ;
        RECT 173.235 -99.445 173.565 -99.115 ;
        RECT 173.235 -100.805 173.565 -100.475 ;
        RECT 173.235 -102.165 173.565 -101.835 ;
        RECT 173.235 -103.525 173.565 -103.195 ;
        RECT 173.235 -104.885 173.565 -104.555 ;
        RECT 173.235 -106.245 173.565 -105.915 ;
        RECT 173.235 -107.605 173.565 -107.275 ;
        RECT 173.235 -108.965 173.565 -108.635 ;
        RECT 173.235 -110.325 173.565 -109.995 ;
        RECT 173.235 -111.685 173.565 -111.355 ;
        RECT 173.235 -113.045 173.565 -112.715 ;
        RECT 173.235 -114.405 173.565 -114.075 ;
        RECT 173.235 -115.765 173.565 -115.435 ;
        RECT 173.235 -117.125 173.565 -116.795 ;
        RECT 173.235 -118.485 173.565 -118.155 ;
        RECT 173.235 -119.845 173.565 -119.515 ;
        RECT 173.235 -121.205 173.565 -120.875 ;
        RECT 173.235 -122.565 173.565 -122.235 ;
        RECT 173.235 -123.925 173.565 -123.595 ;
        RECT 173.235 -125.285 173.565 -124.955 ;
        RECT 173.235 -126.645 173.565 -126.315 ;
        RECT 173.235 -128.005 173.565 -127.675 ;
        RECT 173.235 -129.365 173.565 -129.035 ;
        RECT 173.235 -130.725 173.565 -130.395 ;
        RECT 173.235 -132.085 173.565 -131.755 ;
        RECT 173.235 -133.445 173.565 -133.115 ;
        RECT 173.235 -134.805 173.565 -134.475 ;
        RECT 173.235 -136.165 173.565 -135.835 ;
        RECT 173.235 -137.525 173.565 -137.195 ;
        RECT 173.235 -138.885 173.565 -138.555 ;
        RECT 173.235 -140.245 173.565 -139.915 ;
        RECT 173.235 -141.605 173.565 -141.275 ;
        RECT 173.235 -142.965 173.565 -142.635 ;
        RECT 173.235 -144.325 173.565 -143.995 ;
        RECT 173.235 -145.685 173.565 -145.355 ;
        RECT 173.235 -147.045 173.565 -146.715 ;
        RECT 173.235 -148.405 173.565 -148.075 ;
        RECT 173.235 -149.765 173.565 -149.435 ;
        RECT 173.235 -151.125 173.565 -150.795 ;
        RECT 173.235 -152.485 173.565 -152.155 ;
        RECT 173.235 -153.845 173.565 -153.515 ;
        RECT 173.235 -155.205 173.565 -154.875 ;
        RECT 173.235 -156.565 173.565 -156.235 ;
        RECT 173.235 -157.925 173.565 -157.595 ;
        RECT 173.235 -159.285 173.565 -158.955 ;
        RECT 173.235 -160.645 173.565 -160.315 ;
        RECT 173.235 -162.005 173.565 -161.675 ;
        RECT 173.235 -163.365 173.565 -163.035 ;
        RECT 173.235 -164.725 173.565 -164.395 ;
        RECT 173.235 -166.085 173.565 -165.755 ;
        RECT 173.235 -167.445 173.565 -167.115 ;
        RECT 173.235 -168.805 173.565 -168.475 ;
        RECT 173.235 -170.165 173.565 -169.835 ;
        RECT 173.235 -171.525 173.565 -171.195 ;
        RECT 173.235 -172.885 173.565 -172.555 ;
        RECT 173.235 -174.245 173.565 -173.915 ;
        RECT 173.235 -175.605 173.565 -175.275 ;
        RECT 173.235 -176.965 173.565 -176.635 ;
        RECT 173.235 -178.325 173.565 -177.995 ;
        RECT 173.235 -179.685 173.565 -179.355 ;
        RECT 173.235 -181.93 173.565 -180.8 ;
        RECT 173.24 -182.045 173.56 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.595 241.32 174.925 242.45 ;
        RECT 174.595 239.195 174.925 239.525 ;
        RECT 174.595 237.835 174.925 238.165 ;
        RECT 174.6 237.16 174.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.595 -1.525 174.925 -1.195 ;
        RECT 174.595 -2.885 174.925 -2.555 ;
        RECT 174.6 -3.56 174.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 174.595 -95.365 174.925 -95.035 ;
        RECT 174.595 -96.725 174.925 -96.395 ;
        RECT 174.595 -98.085 174.925 -97.755 ;
        RECT 174.595 -99.445 174.925 -99.115 ;
        RECT 174.595 -100.805 174.925 -100.475 ;
        RECT 174.595 -102.165 174.925 -101.835 ;
        RECT 174.595 -103.525 174.925 -103.195 ;
        RECT 174.595 -104.885 174.925 -104.555 ;
        RECT 174.595 -106.245 174.925 -105.915 ;
        RECT 174.595 -107.605 174.925 -107.275 ;
        RECT 174.595 -108.965 174.925 -108.635 ;
        RECT 174.595 -110.325 174.925 -109.995 ;
        RECT 174.595 -111.685 174.925 -111.355 ;
        RECT 174.595 -113.045 174.925 -112.715 ;
        RECT 174.595 -114.405 174.925 -114.075 ;
        RECT 174.595 -115.765 174.925 -115.435 ;
        RECT 174.595 -117.125 174.925 -116.795 ;
        RECT 174.595 -118.485 174.925 -118.155 ;
        RECT 174.595 -119.845 174.925 -119.515 ;
        RECT 174.595 -121.205 174.925 -120.875 ;
        RECT 174.595 -122.565 174.925 -122.235 ;
        RECT 174.595 -123.925 174.925 -123.595 ;
        RECT 174.595 -125.285 174.925 -124.955 ;
        RECT 174.595 -126.645 174.925 -126.315 ;
        RECT 174.595 -128.005 174.925 -127.675 ;
        RECT 174.595 -129.365 174.925 -129.035 ;
        RECT 174.595 -130.725 174.925 -130.395 ;
        RECT 174.595 -132.085 174.925 -131.755 ;
        RECT 174.595 -133.445 174.925 -133.115 ;
        RECT 174.595 -134.805 174.925 -134.475 ;
        RECT 174.595 -136.165 174.925 -135.835 ;
        RECT 174.595 -137.525 174.925 -137.195 ;
        RECT 174.595 -138.885 174.925 -138.555 ;
        RECT 174.595 -140.245 174.925 -139.915 ;
        RECT 174.595 -141.605 174.925 -141.275 ;
        RECT 174.595 -142.965 174.925 -142.635 ;
        RECT 174.595 -144.325 174.925 -143.995 ;
        RECT 174.595 -145.685 174.925 -145.355 ;
        RECT 174.595 -147.045 174.925 -146.715 ;
        RECT 174.595 -148.405 174.925 -148.075 ;
        RECT 174.595 -149.765 174.925 -149.435 ;
        RECT 174.595 -151.125 174.925 -150.795 ;
        RECT 174.595 -152.485 174.925 -152.155 ;
        RECT 174.595 -153.845 174.925 -153.515 ;
        RECT 174.595 -155.205 174.925 -154.875 ;
        RECT 174.595 -156.565 174.925 -156.235 ;
        RECT 174.595 -157.925 174.925 -157.595 ;
        RECT 174.595 -159.285 174.925 -158.955 ;
        RECT 174.595 -160.645 174.925 -160.315 ;
        RECT 174.595 -162.005 174.925 -161.675 ;
        RECT 174.595 -163.365 174.925 -163.035 ;
        RECT 174.595 -164.725 174.925 -164.395 ;
        RECT 174.595 -166.085 174.925 -165.755 ;
        RECT 174.595 -167.445 174.925 -167.115 ;
        RECT 174.595 -168.805 174.925 -168.475 ;
        RECT 174.595 -170.165 174.925 -169.835 ;
        RECT 174.595 -171.525 174.925 -171.195 ;
        RECT 174.595 -172.885 174.925 -172.555 ;
        RECT 174.595 -174.245 174.925 -173.915 ;
        RECT 174.595 -175.605 174.925 -175.275 ;
        RECT 174.595 -176.965 174.925 -176.635 ;
        RECT 174.595 -178.325 174.925 -177.995 ;
        RECT 174.595 -179.685 174.925 -179.355 ;
        RECT 174.595 -181.93 174.925 -180.8 ;
        RECT 174.6 -182.045 174.92 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 241.32 176.285 242.45 ;
        RECT 175.955 239.195 176.285 239.525 ;
        RECT 175.955 237.835 176.285 238.165 ;
        RECT 175.96 237.16 176.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 -1.525 176.285 -1.195 ;
        RECT 175.955 -2.885 176.285 -2.555 ;
        RECT 175.96 -3.56 176.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 175.955 -95.365 176.285 -95.035 ;
        RECT 175.955 -96.725 176.285 -96.395 ;
        RECT 175.955 -98.085 176.285 -97.755 ;
        RECT 175.955 -99.445 176.285 -99.115 ;
        RECT 175.955 -100.805 176.285 -100.475 ;
        RECT 175.955 -102.165 176.285 -101.835 ;
        RECT 175.955 -103.525 176.285 -103.195 ;
        RECT 175.955 -104.885 176.285 -104.555 ;
        RECT 175.955 -106.245 176.285 -105.915 ;
        RECT 175.955 -107.605 176.285 -107.275 ;
        RECT 175.955 -108.965 176.285 -108.635 ;
        RECT 175.955 -110.325 176.285 -109.995 ;
        RECT 175.955 -111.685 176.285 -111.355 ;
        RECT 175.955 -113.045 176.285 -112.715 ;
        RECT 175.955 -114.405 176.285 -114.075 ;
        RECT 175.955 -115.765 176.285 -115.435 ;
        RECT 175.955 -117.125 176.285 -116.795 ;
        RECT 175.955 -118.485 176.285 -118.155 ;
        RECT 175.955 -119.845 176.285 -119.515 ;
        RECT 175.955 -121.205 176.285 -120.875 ;
        RECT 175.955 -122.565 176.285 -122.235 ;
        RECT 175.955 -123.925 176.285 -123.595 ;
        RECT 175.955 -125.285 176.285 -124.955 ;
        RECT 175.955 -126.645 176.285 -126.315 ;
        RECT 175.955 -128.005 176.285 -127.675 ;
        RECT 175.955 -129.365 176.285 -129.035 ;
        RECT 175.955 -130.725 176.285 -130.395 ;
        RECT 175.955 -132.085 176.285 -131.755 ;
        RECT 175.955 -133.445 176.285 -133.115 ;
        RECT 175.955 -134.805 176.285 -134.475 ;
        RECT 175.955 -136.165 176.285 -135.835 ;
        RECT 175.955 -137.525 176.285 -137.195 ;
        RECT 175.955 -138.885 176.285 -138.555 ;
        RECT 175.955 -140.245 176.285 -139.915 ;
        RECT 175.955 -141.605 176.285 -141.275 ;
        RECT 175.955 -142.965 176.285 -142.635 ;
        RECT 175.955 -144.325 176.285 -143.995 ;
        RECT 175.955 -145.685 176.285 -145.355 ;
        RECT 175.955 -147.045 176.285 -146.715 ;
        RECT 175.955 -148.405 176.285 -148.075 ;
        RECT 175.955 -149.765 176.285 -149.435 ;
        RECT 175.955 -151.125 176.285 -150.795 ;
        RECT 175.955 -152.485 176.285 -152.155 ;
        RECT 175.955 -153.845 176.285 -153.515 ;
        RECT 175.955 -155.205 176.285 -154.875 ;
        RECT 175.955 -156.565 176.285 -156.235 ;
        RECT 175.955 -157.925 176.285 -157.595 ;
        RECT 175.955 -159.285 176.285 -158.955 ;
        RECT 175.955 -160.645 176.285 -160.315 ;
        RECT 175.955 -162.005 176.285 -161.675 ;
        RECT 175.955 -163.365 176.285 -163.035 ;
        RECT 175.955 -164.725 176.285 -164.395 ;
        RECT 175.955 -166.085 176.285 -165.755 ;
        RECT 175.955 -167.445 176.285 -167.115 ;
        RECT 175.955 -168.805 176.285 -168.475 ;
        RECT 175.955 -170.165 176.285 -169.835 ;
        RECT 175.955 -171.525 176.285 -171.195 ;
        RECT 175.955 -172.885 176.285 -172.555 ;
        RECT 175.955 -174.245 176.285 -173.915 ;
        RECT 175.955 -175.605 176.285 -175.275 ;
        RECT 175.955 -176.965 176.285 -176.635 ;
        RECT 175.955 -178.325 176.285 -177.995 ;
        RECT 175.955 -179.685 176.285 -179.355 ;
        RECT 175.955 -181.93 176.285 -180.8 ;
        RECT 175.96 -182.045 176.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 241.32 177.645 242.45 ;
        RECT 177.315 239.195 177.645 239.525 ;
        RECT 177.315 237.835 177.645 238.165 ;
        RECT 177.32 237.16 177.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.315 -99.445 177.645 -99.115 ;
        RECT 177.315 -100.805 177.645 -100.475 ;
        RECT 177.315 -102.165 177.645 -101.835 ;
        RECT 177.315 -103.525 177.645 -103.195 ;
        RECT 177.315 -104.885 177.645 -104.555 ;
        RECT 177.315 -106.245 177.645 -105.915 ;
        RECT 177.315 -107.605 177.645 -107.275 ;
        RECT 177.315 -108.965 177.645 -108.635 ;
        RECT 177.315 -110.325 177.645 -109.995 ;
        RECT 177.315 -111.685 177.645 -111.355 ;
        RECT 177.315 -113.045 177.645 -112.715 ;
        RECT 177.315 -114.405 177.645 -114.075 ;
        RECT 177.315 -115.765 177.645 -115.435 ;
        RECT 177.315 -117.125 177.645 -116.795 ;
        RECT 177.315 -118.485 177.645 -118.155 ;
        RECT 177.315 -119.845 177.645 -119.515 ;
        RECT 177.315 -121.205 177.645 -120.875 ;
        RECT 177.315 -122.565 177.645 -122.235 ;
        RECT 177.315 -123.925 177.645 -123.595 ;
        RECT 177.315 -125.285 177.645 -124.955 ;
        RECT 177.315 -126.645 177.645 -126.315 ;
        RECT 177.315 -128.005 177.645 -127.675 ;
        RECT 177.315 -129.365 177.645 -129.035 ;
        RECT 177.315 -130.725 177.645 -130.395 ;
        RECT 177.315 -132.085 177.645 -131.755 ;
        RECT 177.315 -133.445 177.645 -133.115 ;
        RECT 177.315 -134.805 177.645 -134.475 ;
        RECT 177.315 -136.165 177.645 -135.835 ;
        RECT 177.315 -137.525 177.645 -137.195 ;
        RECT 177.315 -138.885 177.645 -138.555 ;
        RECT 177.315 -140.245 177.645 -139.915 ;
        RECT 177.315 -141.605 177.645 -141.275 ;
        RECT 177.315 -142.965 177.645 -142.635 ;
        RECT 177.315 -144.325 177.645 -143.995 ;
        RECT 177.315 -145.685 177.645 -145.355 ;
        RECT 177.315 -147.045 177.645 -146.715 ;
        RECT 177.315 -148.405 177.645 -148.075 ;
        RECT 177.315 -149.765 177.645 -149.435 ;
        RECT 177.315 -151.125 177.645 -150.795 ;
        RECT 177.315 -152.485 177.645 -152.155 ;
        RECT 177.315 -153.845 177.645 -153.515 ;
        RECT 177.315 -155.205 177.645 -154.875 ;
        RECT 177.315 -156.565 177.645 -156.235 ;
        RECT 177.315 -157.925 177.645 -157.595 ;
        RECT 177.315 -159.285 177.645 -158.955 ;
        RECT 177.315 -160.645 177.645 -160.315 ;
        RECT 177.315 -162.005 177.645 -161.675 ;
        RECT 177.315 -163.365 177.645 -163.035 ;
        RECT 177.315 -164.725 177.645 -164.395 ;
        RECT 177.315 -166.085 177.645 -165.755 ;
        RECT 177.315 -167.445 177.645 -167.115 ;
        RECT 177.315 -168.805 177.645 -168.475 ;
        RECT 177.315 -170.165 177.645 -169.835 ;
        RECT 177.315 -171.525 177.645 -171.195 ;
        RECT 177.315 -172.885 177.645 -172.555 ;
        RECT 177.315 -174.245 177.645 -173.915 ;
        RECT 177.315 -175.605 177.645 -175.275 ;
        RECT 177.315 -176.965 177.645 -176.635 ;
        RECT 177.315 -178.325 177.645 -177.995 ;
        RECT 177.315 -179.685 177.645 -179.355 ;
        RECT 177.315 -181.93 177.645 -180.8 ;
        RECT 177.32 -182.045 177.64 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 177.71 -98.075 178.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 241.32 179.005 242.45 ;
        RECT 178.675 239.195 179.005 239.525 ;
        RECT 178.675 237.835 179.005 238.165 ;
        RECT 178.68 237.16 179 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 178.675 -1.525 179.005 -1.195 ;
        RECT 178.675 -2.885 179.005 -2.555 ;
        RECT 178.68 -3.56 179 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 241.32 180.365 242.45 ;
        RECT 180.035 239.195 180.365 239.525 ;
        RECT 180.035 237.835 180.365 238.165 ;
        RECT 180.04 237.16 180.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 180.035 -1.525 180.365 -1.195 ;
        RECT 180.035 -2.885 180.365 -2.555 ;
        RECT 180.04 -3.56 180.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 241.32 181.725 242.45 ;
        RECT 181.395 239.195 181.725 239.525 ;
        RECT 181.395 237.835 181.725 238.165 ;
        RECT 181.4 237.16 181.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 -1.525 181.725 -1.195 ;
        RECT 181.395 -2.885 181.725 -2.555 ;
        RECT 181.4 -3.56 181.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 181.395 -95.365 181.725 -95.035 ;
        RECT 181.395 -96.725 181.725 -96.395 ;
        RECT 181.395 -98.085 181.725 -97.755 ;
        RECT 181.395 -99.445 181.725 -99.115 ;
        RECT 181.395 -100.805 181.725 -100.475 ;
        RECT 181.395 -102.165 181.725 -101.835 ;
        RECT 181.395 -103.525 181.725 -103.195 ;
        RECT 181.395 -104.885 181.725 -104.555 ;
        RECT 181.395 -106.245 181.725 -105.915 ;
        RECT 181.395 -107.605 181.725 -107.275 ;
        RECT 181.395 -108.965 181.725 -108.635 ;
        RECT 181.395 -110.325 181.725 -109.995 ;
        RECT 181.395 -111.685 181.725 -111.355 ;
        RECT 181.395 -113.045 181.725 -112.715 ;
        RECT 181.395 -114.405 181.725 -114.075 ;
        RECT 181.395 -115.765 181.725 -115.435 ;
        RECT 181.395 -117.125 181.725 -116.795 ;
        RECT 181.395 -118.485 181.725 -118.155 ;
        RECT 181.395 -119.845 181.725 -119.515 ;
        RECT 181.395 -121.205 181.725 -120.875 ;
        RECT 181.395 -122.565 181.725 -122.235 ;
        RECT 181.395 -123.925 181.725 -123.595 ;
        RECT 181.395 -125.285 181.725 -124.955 ;
        RECT 181.395 -126.645 181.725 -126.315 ;
        RECT 181.395 -128.005 181.725 -127.675 ;
        RECT 181.395 -129.365 181.725 -129.035 ;
        RECT 181.395 -130.725 181.725 -130.395 ;
        RECT 181.395 -132.085 181.725 -131.755 ;
        RECT 181.395 -133.445 181.725 -133.115 ;
        RECT 181.395 -134.805 181.725 -134.475 ;
        RECT 181.395 -136.165 181.725 -135.835 ;
        RECT 181.395 -137.525 181.725 -137.195 ;
        RECT 181.395 -138.885 181.725 -138.555 ;
        RECT 181.395 -140.245 181.725 -139.915 ;
        RECT 181.395 -141.605 181.725 -141.275 ;
        RECT 181.395 -142.965 181.725 -142.635 ;
        RECT 181.395 -144.325 181.725 -143.995 ;
        RECT 181.395 -145.685 181.725 -145.355 ;
        RECT 181.395 -147.045 181.725 -146.715 ;
        RECT 181.395 -148.405 181.725 -148.075 ;
        RECT 181.395 -149.765 181.725 -149.435 ;
        RECT 181.395 -151.125 181.725 -150.795 ;
        RECT 181.395 -152.485 181.725 -152.155 ;
        RECT 181.395 -153.845 181.725 -153.515 ;
        RECT 181.395 -155.205 181.725 -154.875 ;
        RECT 181.395 -156.565 181.725 -156.235 ;
        RECT 181.395 -157.925 181.725 -157.595 ;
        RECT 181.395 -159.285 181.725 -158.955 ;
        RECT 181.395 -160.645 181.725 -160.315 ;
        RECT 181.395 -162.005 181.725 -161.675 ;
        RECT 181.395 -163.365 181.725 -163.035 ;
        RECT 181.395 -164.725 181.725 -164.395 ;
        RECT 181.395 -166.085 181.725 -165.755 ;
        RECT 181.395 -167.445 181.725 -167.115 ;
        RECT 181.395 -168.805 181.725 -168.475 ;
        RECT 181.395 -170.165 181.725 -169.835 ;
        RECT 181.395 -171.525 181.725 -171.195 ;
        RECT 181.395 -172.885 181.725 -172.555 ;
        RECT 181.395 -174.245 181.725 -173.915 ;
        RECT 181.395 -175.605 181.725 -175.275 ;
        RECT 181.395 -176.965 181.725 -176.635 ;
        RECT 181.395 -178.325 181.725 -177.995 ;
        RECT 181.395 -179.685 181.725 -179.355 ;
        RECT 181.395 -181.93 181.725 -180.8 ;
        RECT 181.4 -182.045 181.72 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 241.32 183.085 242.45 ;
        RECT 182.755 239.195 183.085 239.525 ;
        RECT 182.755 237.835 183.085 238.165 ;
        RECT 182.76 237.16 183.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 -1.525 183.085 -1.195 ;
        RECT 182.755 -2.885 183.085 -2.555 ;
        RECT 182.76 -3.56 183.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 182.755 -95.365 183.085 -95.035 ;
        RECT 182.755 -96.725 183.085 -96.395 ;
        RECT 182.755 -98.085 183.085 -97.755 ;
        RECT 182.755 -99.445 183.085 -99.115 ;
        RECT 182.755 -100.805 183.085 -100.475 ;
        RECT 182.755 -102.165 183.085 -101.835 ;
        RECT 182.755 -103.525 183.085 -103.195 ;
        RECT 182.755 -104.885 183.085 -104.555 ;
        RECT 182.755 -106.245 183.085 -105.915 ;
        RECT 182.755 -107.605 183.085 -107.275 ;
        RECT 182.755 -108.965 183.085 -108.635 ;
        RECT 182.755 -110.325 183.085 -109.995 ;
        RECT 182.755 -111.685 183.085 -111.355 ;
        RECT 182.755 -113.045 183.085 -112.715 ;
        RECT 182.755 -114.405 183.085 -114.075 ;
        RECT 182.755 -115.765 183.085 -115.435 ;
        RECT 182.755 -117.125 183.085 -116.795 ;
        RECT 182.755 -118.485 183.085 -118.155 ;
        RECT 182.755 -119.845 183.085 -119.515 ;
        RECT 182.755 -121.205 183.085 -120.875 ;
        RECT 182.755 -122.565 183.085 -122.235 ;
        RECT 182.755 -123.925 183.085 -123.595 ;
        RECT 182.755 -125.285 183.085 -124.955 ;
        RECT 182.755 -126.645 183.085 -126.315 ;
        RECT 182.755 -128.005 183.085 -127.675 ;
        RECT 182.755 -129.365 183.085 -129.035 ;
        RECT 182.755 -130.725 183.085 -130.395 ;
        RECT 182.755 -132.085 183.085 -131.755 ;
        RECT 182.755 -133.445 183.085 -133.115 ;
        RECT 182.755 -134.805 183.085 -134.475 ;
        RECT 182.755 -136.165 183.085 -135.835 ;
        RECT 182.755 -137.525 183.085 -137.195 ;
        RECT 182.755 -138.885 183.085 -138.555 ;
        RECT 182.755 -140.245 183.085 -139.915 ;
        RECT 182.755 -141.605 183.085 -141.275 ;
        RECT 182.755 -142.965 183.085 -142.635 ;
        RECT 182.755 -144.325 183.085 -143.995 ;
        RECT 182.755 -145.685 183.085 -145.355 ;
        RECT 182.755 -147.045 183.085 -146.715 ;
        RECT 182.755 -148.405 183.085 -148.075 ;
        RECT 182.755 -149.765 183.085 -149.435 ;
        RECT 182.755 -151.125 183.085 -150.795 ;
        RECT 182.755 -152.485 183.085 -152.155 ;
        RECT 182.755 -153.845 183.085 -153.515 ;
        RECT 182.755 -155.205 183.085 -154.875 ;
        RECT 182.755 -156.565 183.085 -156.235 ;
        RECT 182.755 -157.925 183.085 -157.595 ;
        RECT 182.755 -159.285 183.085 -158.955 ;
        RECT 182.755 -160.645 183.085 -160.315 ;
        RECT 182.755 -162.005 183.085 -161.675 ;
        RECT 182.755 -163.365 183.085 -163.035 ;
        RECT 182.755 -164.725 183.085 -164.395 ;
        RECT 182.755 -166.085 183.085 -165.755 ;
        RECT 182.755 -167.445 183.085 -167.115 ;
        RECT 182.755 -168.805 183.085 -168.475 ;
        RECT 182.755 -170.165 183.085 -169.835 ;
        RECT 182.755 -171.525 183.085 -171.195 ;
        RECT 182.755 -172.885 183.085 -172.555 ;
        RECT 182.755 -174.245 183.085 -173.915 ;
        RECT 182.755 -175.605 183.085 -175.275 ;
        RECT 182.755 -176.965 183.085 -176.635 ;
        RECT 182.755 -178.325 183.085 -177.995 ;
        RECT 182.755 -179.685 183.085 -179.355 ;
        RECT 182.755 -181.93 183.085 -180.8 ;
        RECT 182.76 -182.045 183.08 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 241.32 184.445 242.45 ;
        RECT 184.115 239.195 184.445 239.525 ;
        RECT 184.115 237.835 184.445 238.165 ;
        RECT 184.12 237.16 184.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 -1.525 184.445 -1.195 ;
        RECT 184.115 -2.885 184.445 -2.555 ;
        RECT 184.12 -3.56 184.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 184.115 -95.365 184.445 -95.035 ;
        RECT 184.115 -96.725 184.445 -96.395 ;
        RECT 184.115 -98.085 184.445 -97.755 ;
        RECT 184.115 -99.445 184.445 -99.115 ;
        RECT 184.115 -100.805 184.445 -100.475 ;
        RECT 184.115 -102.165 184.445 -101.835 ;
        RECT 184.115 -103.525 184.445 -103.195 ;
        RECT 184.115 -104.885 184.445 -104.555 ;
        RECT 184.115 -106.245 184.445 -105.915 ;
        RECT 184.115 -107.605 184.445 -107.275 ;
        RECT 184.115 -108.965 184.445 -108.635 ;
        RECT 184.115 -110.325 184.445 -109.995 ;
        RECT 184.115 -111.685 184.445 -111.355 ;
        RECT 184.115 -113.045 184.445 -112.715 ;
        RECT 184.115 -114.405 184.445 -114.075 ;
        RECT 184.115 -115.765 184.445 -115.435 ;
        RECT 184.115 -117.125 184.445 -116.795 ;
        RECT 184.115 -118.485 184.445 -118.155 ;
        RECT 184.115 -119.845 184.445 -119.515 ;
        RECT 184.115 -121.205 184.445 -120.875 ;
        RECT 184.115 -122.565 184.445 -122.235 ;
        RECT 184.115 -123.925 184.445 -123.595 ;
        RECT 184.115 -125.285 184.445 -124.955 ;
        RECT 184.115 -126.645 184.445 -126.315 ;
        RECT 184.115 -128.005 184.445 -127.675 ;
        RECT 184.115 -129.365 184.445 -129.035 ;
        RECT 184.115 -130.725 184.445 -130.395 ;
        RECT 184.115 -132.085 184.445 -131.755 ;
        RECT 184.115 -133.445 184.445 -133.115 ;
        RECT 184.115 -134.805 184.445 -134.475 ;
        RECT 184.115 -136.165 184.445 -135.835 ;
        RECT 184.115 -137.525 184.445 -137.195 ;
        RECT 184.115 -138.885 184.445 -138.555 ;
        RECT 184.115 -140.245 184.445 -139.915 ;
        RECT 184.115 -141.605 184.445 -141.275 ;
        RECT 184.115 -142.965 184.445 -142.635 ;
        RECT 184.115 -144.325 184.445 -143.995 ;
        RECT 184.115 -145.685 184.445 -145.355 ;
        RECT 184.115 -147.045 184.445 -146.715 ;
        RECT 184.115 -148.405 184.445 -148.075 ;
        RECT 184.115 -149.765 184.445 -149.435 ;
        RECT 184.115 -151.125 184.445 -150.795 ;
        RECT 184.115 -152.485 184.445 -152.155 ;
        RECT 184.115 -153.845 184.445 -153.515 ;
        RECT 184.115 -155.205 184.445 -154.875 ;
        RECT 184.115 -156.565 184.445 -156.235 ;
        RECT 184.115 -157.925 184.445 -157.595 ;
        RECT 184.115 -159.285 184.445 -158.955 ;
        RECT 184.115 -160.645 184.445 -160.315 ;
        RECT 184.115 -162.005 184.445 -161.675 ;
        RECT 184.115 -163.365 184.445 -163.035 ;
        RECT 184.115 -164.725 184.445 -164.395 ;
        RECT 184.115 -166.085 184.445 -165.755 ;
        RECT 184.115 -167.445 184.445 -167.115 ;
        RECT 184.115 -168.805 184.445 -168.475 ;
        RECT 184.115 -170.165 184.445 -169.835 ;
        RECT 184.115 -171.525 184.445 -171.195 ;
        RECT 184.115 -172.885 184.445 -172.555 ;
        RECT 184.115 -174.245 184.445 -173.915 ;
        RECT 184.115 -175.605 184.445 -175.275 ;
        RECT 184.115 -176.965 184.445 -176.635 ;
        RECT 184.115 -178.325 184.445 -177.995 ;
        RECT 184.115 -179.685 184.445 -179.355 ;
        RECT 184.115 -181.93 184.445 -180.8 ;
        RECT 184.12 -182.045 184.44 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 241.32 185.805 242.45 ;
        RECT 185.475 239.195 185.805 239.525 ;
        RECT 185.475 237.835 185.805 238.165 ;
        RECT 185.48 237.16 185.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 -1.525 185.805 -1.195 ;
        RECT 185.475 -2.885 185.805 -2.555 ;
        RECT 185.48 -3.56 185.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 185.475 -95.365 185.805 -95.035 ;
        RECT 185.475 -96.725 185.805 -96.395 ;
        RECT 185.475 -98.085 185.805 -97.755 ;
        RECT 185.475 -99.445 185.805 -99.115 ;
        RECT 185.475 -100.805 185.805 -100.475 ;
        RECT 185.475 -102.165 185.805 -101.835 ;
        RECT 185.475 -103.525 185.805 -103.195 ;
        RECT 185.475 -104.885 185.805 -104.555 ;
        RECT 185.475 -106.245 185.805 -105.915 ;
        RECT 185.475 -107.605 185.805 -107.275 ;
        RECT 185.475 -108.965 185.805 -108.635 ;
        RECT 185.475 -110.325 185.805 -109.995 ;
        RECT 185.475 -111.685 185.805 -111.355 ;
        RECT 185.475 -113.045 185.805 -112.715 ;
        RECT 185.475 -114.405 185.805 -114.075 ;
        RECT 185.475 -115.765 185.805 -115.435 ;
        RECT 185.475 -117.125 185.805 -116.795 ;
        RECT 185.475 -118.485 185.805 -118.155 ;
        RECT 185.475 -119.845 185.805 -119.515 ;
        RECT 185.475 -121.205 185.805 -120.875 ;
        RECT 185.475 -122.565 185.805 -122.235 ;
        RECT 185.475 -123.925 185.805 -123.595 ;
        RECT 185.475 -125.285 185.805 -124.955 ;
        RECT 185.475 -126.645 185.805 -126.315 ;
        RECT 185.475 -128.005 185.805 -127.675 ;
        RECT 185.475 -129.365 185.805 -129.035 ;
        RECT 185.475 -130.725 185.805 -130.395 ;
        RECT 185.475 -132.085 185.805 -131.755 ;
        RECT 185.475 -133.445 185.805 -133.115 ;
        RECT 185.475 -134.805 185.805 -134.475 ;
        RECT 185.475 -136.165 185.805 -135.835 ;
        RECT 185.475 -137.525 185.805 -137.195 ;
        RECT 185.475 -138.885 185.805 -138.555 ;
        RECT 185.475 -140.245 185.805 -139.915 ;
        RECT 185.475 -141.605 185.805 -141.275 ;
        RECT 185.475 -142.965 185.805 -142.635 ;
        RECT 185.475 -144.325 185.805 -143.995 ;
        RECT 185.475 -145.685 185.805 -145.355 ;
        RECT 185.475 -147.045 185.805 -146.715 ;
        RECT 185.475 -148.405 185.805 -148.075 ;
        RECT 185.475 -149.765 185.805 -149.435 ;
        RECT 185.475 -151.125 185.805 -150.795 ;
        RECT 185.475 -152.485 185.805 -152.155 ;
        RECT 185.475 -153.845 185.805 -153.515 ;
        RECT 185.475 -155.205 185.805 -154.875 ;
        RECT 185.475 -156.565 185.805 -156.235 ;
        RECT 185.475 -157.925 185.805 -157.595 ;
        RECT 185.475 -159.285 185.805 -158.955 ;
        RECT 185.475 -160.645 185.805 -160.315 ;
        RECT 185.475 -162.005 185.805 -161.675 ;
        RECT 185.475 -163.365 185.805 -163.035 ;
        RECT 185.475 -164.725 185.805 -164.395 ;
        RECT 185.475 -166.085 185.805 -165.755 ;
        RECT 185.475 -167.445 185.805 -167.115 ;
        RECT 185.475 -168.805 185.805 -168.475 ;
        RECT 185.475 -170.165 185.805 -169.835 ;
        RECT 185.475 -171.525 185.805 -171.195 ;
        RECT 185.475 -172.885 185.805 -172.555 ;
        RECT 185.475 -174.245 185.805 -173.915 ;
        RECT 185.475 -175.605 185.805 -175.275 ;
        RECT 185.475 -176.965 185.805 -176.635 ;
        RECT 185.475 -178.325 185.805 -177.995 ;
        RECT 185.475 -179.685 185.805 -179.355 ;
        RECT 185.475 -181.93 185.805 -180.8 ;
        RECT 185.48 -182.045 185.8 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.835 241.32 187.165 242.45 ;
        RECT 186.835 239.195 187.165 239.525 ;
        RECT 186.835 237.835 187.165 238.165 ;
        RECT 186.84 237.16 187.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.835 -1.525 187.165 -1.195 ;
        RECT 186.835 -2.885 187.165 -2.555 ;
        RECT 186.84 -3.56 187.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 186.835 -95.365 187.165 -95.035 ;
        RECT 186.835 -96.725 187.165 -96.395 ;
        RECT 186.835 -98.085 187.165 -97.755 ;
        RECT 186.835 -99.445 187.165 -99.115 ;
        RECT 186.835 -100.805 187.165 -100.475 ;
        RECT 186.835 -102.165 187.165 -101.835 ;
        RECT 186.835 -103.525 187.165 -103.195 ;
        RECT 186.835 -104.885 187.165 -104.555 ;
        RECT 186.835 -106.245 187.165 -105.915 ;
        RECT 186.835 -107.605 187.165 -107.275 ;
        RECT 186.835 -108.965 187.165 -108.635 ;
        RECT 186.835 -110.325 187.165 -109.995 ;
        RECT 186.835 -111.685 187.165 -111.355 ;
        RECT 186.835 -113.045 187.165 -112.715 ;
        RECT 186.835 -114.405 187.165 -114.075 ;
        RECT 186.835 -115.765 187.165 -115.435 ;
        RECT 186.835 -117.125 187.165 -116.795 ;
        RECT 186.835 -118.485 187.165 -118.155 ;
        RECT 186.835 -119.845 187.165 -119.515 ;
        RECT 186.835 -121.205 187.165 -120.875 ;
        RECT 186.835 -122.565 187.165 -122.235 ;
        RECT 186.835 -123.925 187.165 -123.595 ;
        RECT 186.835 -125.285 187.165 -124.955 ;
        RECT 186.835 -126.645 187.165 -126.315 ;
        RECT 186.835 -128.005 187.165 -127.675 ;
        RECT 186.835 -129.365 187.165 -129.035 ;
        RECT 186.835 -130.725 187.165 -130.395 ;
        RECT 186.835 -132.085 187.165 -131.755 ;
        RECT 186.835 -133.445 187.165 -133.115 ;
        RECT 186.835 -134.805 187.165 -134.475 ;
        RECT 186.835 -136.165 187.165 -135.835 ;
        RECT 186.835 -137.525 187.165 -137.195 ;
        RECT 186.835 -138.885 187.165 -138.555 ;
        RECT 186.835 -140.245 187.165 -139.915 ;
        RECT 186.835 -141.605 187.165 -141.275 ;
        RECT 186.835 -142.965 187.165 -142.635 ;
        RECT 186.835 -144.325 187.165 -143.995 ;
        RECT 186.835 -145.685 187.165 -145.355 ;
        RECT 186.835 -147.045 187.165 -146.715 ;
        RECT 186.835 -148.405 187.165 -148.075 ;
        RECT 186.835 -149.765 187.165 -149.435 ;
        RECT 186.835 -151.125 187.165 -150.795 ;
        RECT 186.835 -152.485 187.165 -152.155 ;
        RECT 186.835 -153.845 187.165 -153.515 ;
        RECT 186.835 -155.205 187.165 -154.875 ;
        RECT 186.835 -156.565 187.165 -156.235 ;
        RECT 186.835 -157.925 187.165 -157.595 ;
        RECT 186.835 -159.285 187.165 -158.955 ;
        RECT 186.835 -160.645 187.165 -160.315 ;
        RECT 186.835 -162.005 187.165 -161.675 ;
        RECT 186.835 -163.365 187.165 -163.035 ;
        RECT 186.835 -164.725 187.165 -164.395 ;
        RECT 186.835 -166.085 187.165 -165.755 ;
        RECT 186.835 -167.445 187.165 -167.115 ;
        RECT 186.835 -168.805 187.165 -168.475 ;
        RECT 186.835 -170.165 187.165 -169.835 ;
        RECT 186.835 -171.525 187.165 -171.195 ;
        RECT 186.835 -172.885 187.165 -172.555 ;
        RECT 186.835 -174.245 187.165 -173.915 ;
        RECT 186.835 -175.605 187.165 -175.275 ;
        RECT 186.835 -176.965 187.165 -176.635 ;
        RECT 186.835 -178.325 187.165 -177.995 ;
        RECT 186.835 -179.685 187.165 -179.355 ;
        RECT 186.835 -181.93 187.165 -180.8 ;
        RECT 186.84 -182.045 187.16 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 241.32 188.525 242.45 ;
        RECT 188.195 239.195 188.525 239.525 ;
        RECT 188.195 237.835 188.525 238.165 ;
        RECT 188.2 237.16 188.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.195 -99.445 188.525 -99.115 ;
        RECT 188.195 -100.805 188.525 -100.475 ;
        RECT 188.195 -102.165 188.525 -101.835 ;
        RECT 188.195 -103.525 188.525 -103.195 ;
        RECT 188.195 -104.885 188.525 -104.555 ;
        RECT 188.195 -106.245 188.525 -105.915 ;
        RECT 188.195 -107.605 188.525 -107.275 ;
        RECT 188.195 -108.965 188.525 -108.635 ;
        RECT 188.195 -110.325 188.525 -109.995 ;
        RECT 188.195 -111.685 188.525 -111.355 ;
        RECT 188.195 -113.045 188.525 -112.715 ;
        RECT 188.195 -114.405 188.525 -114.075 ;
        RECT 188.195 -115.765 188.525 -115.435 ;
        RECT 188.195 -117.125 188.525 -116.795 ;
        RECT 188.195 -118.485 188.525 -118.155 ;
        RECT 188.195 -119.845 188.525 -119.515 ;
        RECT 188.195 -121.205 188.525 -120.875 ;
        RECT 188.195 -122.565 188.525 -122.235 ;
        RECT 188.195 -123.925 188.525 -123.595 ;
        RECT 188.195 -125.285 188.525 -124.955 ;
        RECT 188.195 -126.645 188.525 -126.315 ;
        RECT 188.195 -128.005 188.525 -127.675 ;
        RECT 188.195 -129.365 188.525 -129.035 ;
        RECT 188.195 -130.725 188.525 -130.395 ;
        RECT 188.195 -132.085 188.525 -131.755 ;
        RECT 188.195 -133.445 188.525 -133.115 ;
        RECT 188.195 -134.805 188.525 -134.475 ;
        RECT 188.195 -136.165 188.525 -135.835 ;
        RECT 188.195 -137.525 188.525 -137.195 ;
        RECT 188.195 -138.885 188.525 -138.555 ;
        RECT 188.195 -140.245 188.525 -139.915 ;
        RECT 188.195 -141.605 188.525 -141.275 ;
        RECT 188.195 -142.965 188.525 -142.635 ;
        RECT 188.195 -144.325 188.525 -143.995 ;
        RECT 188.195 -145.685 188.525 -145.355 ;
        RECT 188.195 -147.045 188.525 -146.715 ;
        RECT 188.195 -148.405 188.525 -148.075 ;
        RECT 188.195 -149.765 188.525 -149.435 ;
        RECT 188.195 -151.125 188.525 -150.795 ;
        RECT 188.195 -152.485 188.525 -152.155 ;
        RECT 188.195 -153.845 188.525 -153.515 ;
        RECT 188.195 -155.205 188.525 -154.875 ;
        RECT 188.195 -156.565 188.525 -156.235 ;
        RECT 188.195 -157.925 188.525 -157.595 ;
        RECT 188.195 -159.285 188.525 -158.955 ;
        RECT 188.195 -160.645 188.525 -160.315 ;
        RECT 188.195 -162.005 188.525 -161.675 ;
        RECT 188.195 -163.365 188.525 -163.035 ;
        RECT 188.195 -164.725 188.525 -164.395 ;
        RECT 188.195 -166.085 188.525 -165.755 ;
        RECT 188.195 -167.445 188.525 -167.115 ;
        RECT 188.195 -168.805 188.525 -168.475 ;
        RECT 188.195 -170.165 188.525 -169.835 ;
        RECT 188.195 -171.525 188.525 -171.195 ;
        RECT 188.195 -172.885 188.525 -172.555 ;
        RECT 188.195 -174.245 188.525 -173.915 ;
        RECT 188.195 -175.605 188.525 -175.275 ;
        RECT 188.195 -176.965 188.525 -176.635 ;
        RECT 188.195 -178.325 188.525 -177.995 ;
        RECT 188.195 -179.685 188.525 -179.355 ;
        RECT 188.195 -181.93 188.525 -180.8 ;
        RECT 188.2 -182.045 188.52 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 188.61 -98.075 188.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 241.32 189.885 242.45 ;
        RECT 189.555 239.195 189.885 239.525 ;
        RECT 189.555 237.835 189.885 238.165 ;
        RECT 189.56 237.16 189.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 189.555 -1.525 189.885 -1.195 ;
        RECT 189.555 -2.885 189.885 -2.555 ;
        RECT 189.56 -3.56 189.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 241.32 191.245 242.45 ;
        RECT 190.915 239.195 191.245 239.525 ;
        RECT 190.915 237.835 191.245 238.165 ;
        RECT 190.92 237.16 191.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 190.915 -1.525 191.245 -1.195 ;
        RECT 190.915 -2.885 191.245 -2.555 ;
        RECT 190.92 -3.56 191.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 241.32 192.605 242.45 ;
        RECT 192.275 239.195 192.605 239.525 ;
        RECT 192.275 237.835 192.605 238.165 ;
        RECT 192.28 237.16 192.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 -1.525 192.605 -1.195 ;
        RECT 192.275 -2.885 192.605 -2.555 ;
        RECT 192.28 -3.56 192.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 192.275 -170.165 192.605 -169.835 ;
        RECT 192.275 -171.525 192.605 -171.195 ;
        RECT 192.275 -172.885 192.605 -172.555 ;
        RECT 192.275 -174.245 192.605 -173.915 ;
        RECT 192.275 -175.605 192.605 -175.275 ;
        RECT 192.275 -176.965 192.605 -176.635 ;
        RECT 192.275 -178.325 192.605 -177.995 ;
        RECT 192.275 -179.685 192.605 -179.355 ;
        RECT 192.275 -181.93 192.605 -180.8 ;
        RECT 192.28 -182.045 192.6 -95.035 ;
        RECT 192.275 -95.365 192.605 -95.035 ;
        RECT 192.275 -96.725 192.605 -96.395 ;
        RECT 192.275 -98.085 192.605 -97.755 ;
        RECT 192.275 -99.445 192.605 -99.115 ;
        RECT 192.275 -100.805 192.605 -100.475 ;
        RECT 192.275 -102.165 192.605 -101.835 ;
        RECT 192.275 -103.525 192.605 -103.195 ;
        RECT 192.275 -104.885 192.605 -104.555 ;
        RECT 192.275 -106.245 192.605 -105.915 ;
        RECT 192.275 -107.605 192.605 -107.275 ;
        RECT 192.275 -108.965 192.605 -108.635 ;
        RECT 192.275 -110.325 192.605 -109.995 ;
        RECT 192.275 -111.685 192.605 -111.355 ;
        RECT 192.275 -113.045 192.605 -112.715 ;
        RECT 192.275 -114.405 192.605 -114.075 ;
        RECT 192.275 -115.765 192.605 -115.435 ;
        RECT 192.275 -117.125 192.605 -116.795 ;
        RECT 192.275 -118.485 192.605 -118.155 ;
        RECT 192.275 -119.845 192.605 -119.515 ;
        RECT 192.275 -121.205 192.605 -120.875 ;
        RECT 192.275 -122.565 192.605 -122.235 ;
        RECT 192.275 -123.925 192.605 -123.595 ;
        RECT 192.275 -125.285 192.605 -124.955 ;
        RECT 192.275 -126.645 192.605 -126.315 ;
        RECT 192.275 -128.005 192.605 -127.675 ;
        RECT 192.275 -129.365 192.605 -129.035 ;
        RECT 192.275 -130.725 192.605 -130.395 ;
        RECT 192.275 -132.085 192.605 -131.755 ;
        RECT 192.275 -133.445 192.605 -133.115 ;
        RECT 192.275 -134.805 192.605 -134.475 ;
        RECT 192.275 -136.165 192.605 -135.835 ;
        RECT 192.275 -137.525 192.605 -137.195 ;
        RECT 192.275 -138.885 192.605 -138.555 ;
        RECT 192.275 -140.245 192.605 -139.915 ;
        RECT 192.275 -141.605 192.605 -141.275 ;
        RECT 192.275 -142.965 192.605 -142.635 ;
        RECT 192.275 -144.325 192.605 -143.995 ;
        RECT 192.275 -145.685 192.605 -145.355 ;
        RECT 192.275 -147.045 192.605 -146.715 ;
        RECT 192.275 -148.405 192.605 -148.075 ;
        RECT 192.275 -149.765 192.605 -149.435 ;
        RECT 192.275 -151.125 192.605 -150.795 ;
        RECT 192.275 -152.485 192.605 -152.155 ;
        RECT 192.275 -153.845 192.605 -153.515 ;
        RECT 192.275 -155.205 192.605 -154.875 ;
        RECT 192.275 -156.565 192.605 -156.235 ;
        RECT 192.275 -157.925 192.605 -157.595 ;
        RECT 192.275 -159.285 192.605 -158.955 ;
        RECT 192.275 -160.645 192.605 -160.315 ;
        RECT 192.275 -162.005 192.605 -161.675 ;
        RECT 192.275 -163.365 192.605 -163.035 ;
        RECT 192.275 -164.725 192.605 -164.395 ;
        RECT 192.275 -166.085 192.605 -165.755 ;
        RECT 192.275 -167.445 192.605 -167.115 ;
        RECT 192.275 -168.805 192.605 -168.475 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 -95.365 142.285 -95.035 ;
        RECT 141.955 -96.725 142.285 -96.395 ;
        RECT 141.955 -98.085 142.285 -97.755 ;
        RECT 141.955 -99.445 142.285 -99.115 ;
        RECT 141.955 -100.805 142.285 -100.475 ;
        RECT 141.955 -102.165 142.285 -101.835 ;
        RECT 141.955 -103.525 142.285 -103.195 ;
        RECT 141.955 -104.885 142.285 -104.555 ;
        RECT 141.955 -106.245 142.285 -105.915 ;
        RECT 141.955 -107.605 142.285 -107.275 ;
        RECT 141.955 -108.965 142.285 -108.635 ;
        RECT 141.955 -110.325 142.285 -109.995 ;
        RECT 141.955 -111.685 142.285 -111.355 ;
        RECT 141.955 -113.045 142.285 -112.715 ;
        RECT 141.955 -114.405 142.285 -114.075 ;
        RECT 141.955 -115.765 142.285 -115.435 ;
        RECT 141.955 -117.125 142.285 -116.795 ;
        RECT 141.955 -118.485 142.285 -118.155 ;
        RECT 141.955 -119.845 142.285 -119.515 ;
        RECT 141.955 -121.205 142.285 -120.875 ;
        RECT 141.955 -122.565 142.285 -122.235 ;
        RECT 141.955 -123.925 142.285 -123.595 ;
        RECT 141.955 -125.285 142.285 -124.955 ;
        RECT 141.955 -126.645 142.285 -126.315 ;
        RECT 141.955 -128.005 142.285 -127.675 ;
        RECT 141.955 -129.365 142.285 -129.035 ;
        RECT 141.955 -130.725 142.285 -130.395 ;
        RECT 141.955 -132.085 142.285 -131.755 ;
        RECT 141.955 -133.445 142.285 -133.115 ;
        RECT 141.955 -134.805 142.285 -134.475 ;
        RECT 141.955 -136.165 142.285 -135.835 ;
        RECT 141.955 -137.525 142.285 -137.195 ;
        RECT 141.955 -138.885 142.285 -138.555 ;
        RECT 141.955 -140.245 142.285 -139.915 ;
        RECT 141.955 -141.605 142.285 -141.275 ;
        RECT 141.955 -142.965 142.285 -142.635 ;
        RECT 141.955 -144.325 142.285 -143.995 ;
        RECT 141.955 -145.685 142.285 -145.355 ;
        RECT 141.955 -147.045 142.285 -146.715 ;
        RECT 141.955 -148.405 142.285 -148.075 ;
        RECT 141.955 -149.765 142.285 -149.435 ;
        RECT 141.955 -151.125 142.285 -150.795 ;
        RECT 141.955 -152.485 142.285 -152.155 ;
        RECT 141.955 -153.845 142.285 -153.515 ;
        RECT 141.955 -155.205 142.285 -154.875 ;
        RECT 141.955 -156.565 142.285 -156.235 ;
        RECT 141.955 -157.925 142.285 -157.595 ;
        RECT 141.955 -159.285 142.285 -158.955 ;
        RECT 141.955 -160.645 142.285 -160.315 ;
        RECT 141.955 -162.005 142.285 -161.675 ;
        RECT 141.955 -163.365 142.285 -163.035 ;
        RECT 141.955 -164.725 142.285 -164.395 ;
        RECT 141.955 -166.085 142.285 -165.755 ;
        RECT 141.955 -167.445 142.285 -167.115 ;
        RECT 141.955 -168.805 142.285 -168.475 ;
        RECT 141.955 -170.165 142.285 -169.835 ;
        RECT 141.955 -171.525 142.285 -171.195 ;
        RECT 141.955 -172.885 142.285 -172.555 ;
        RECT 141.955 -174.245 142.285 -173.915 ;
        RECT 141.955 -175.605 142.285 -175.275 ;
        RECT 141.955 -176.965 142.285 -176.635 ;
        RECT 141.955 -178.325 142.285 -177.995 ;
        RECT 141.955 -179.685 142.285 -179.355 ;
        RECT 141.955 -181.93 142.285 -180.8 ;
        RECT 141.96 -182.045 142.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 241.32 143.645 242.45 ;
        RECT 143.315 239.195 143.645 239.525 ;
        RECT 143.315 237.835 143.645 238.165 ;
        RECT 143.32 237.16 143.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 -1.525 143.645 -1.195 ;
        RECT 143.315 -2.885 143.645 -2.555 ;
        RECT 143.32 -3.56 143.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 143.315 -95.365 143.645 -95.035 ;
        RECT 143.315 -96.725 143.645 -96.395 ;
        RECT 143.315 -98.085 143.645 -97.755 ;
        RECT 143.315 -99.445 143.645 -99.115 ;
        RECT 143.315 -100.805 143.645 -100.475 ;
        RECT 143.315 -102.165 143.645 -101.835 ;
        RECT 143.315 -103.525 143.645 -103.195 ;
        RECT 143.315 -104.885 143.645 -104.555 ;
        RECT 143.315 -106.245 143.645 -105.915 ;
        RECT 143.315 -107.605 143.645 -107.275 ;
        RECT 143.315 -108.965 143.645 -108.635 ;
        RECT 143.315 -110.325 143.645 -109.995 ;
        RECT 143.315 -111.685 143.645 -111.355 ;
        RECT 143.315 -113.045 143.645 -112.715 ;
        RECT 143.315 -114.405 143.645 -114.075 ;
        RECT 143.315 -115.765 143.645 -115.435 ;
        RECT 143.315 -117.125 143.645 -116.795 ;
        RECT 143.315 -118.485 143.645 -118.155 ;
        RECT 143.315 -119.845 143.645 -119.515 ;
        RECT 143.315 -121.205 143.645 -120.875 ;
        RECT 143.315 -122.565 143.645 -122.235 ;
        RECT 143.315 -123.925 143.645 -123.595 ;
        RECT 143.315 -125.285 143.645 -124.955 ;
        RECT 143.315 -126.645 143.645 -126.315 ;
        RECT 143.315 -128.005 143.645 -127.675 ;
        RECT 143.315 -129.365 143.645 -129.035 ;
        RECT 143.315 -130.725 143.645 -130.395 ;
        RECT 143.315 -132.085 143.645 -131.755 ;
        RECT 143.315 -133.445 143.645 -133.115 ;
        RECT 143.315 -134.805 143.645 -134.475 ;
        RECT 143.315 -136.165 143.645 -135.835 ;
        RECT 143.315 -137.525 143.645 -137.195 ;
        RECT 143.315 -138.885 143.645 -138.555 ;
        RECT 143.315 -140.245 143.645 -139.915 ;
        RECT 143.315 -141.605 143.645 -141.275 ;
        RECT 143.315 -142.965 143.645 -142.635 ;
        RECT 143.315 -144.325 143.645 -143.995 ;
        RECT 143.315 -145.685 143.645 -145.355 ;
        RECT 143.315 -147.045 143.645 -146.715 ;
        RECT 143.315 -148.405 143.645 -148.075 ;
        RECT 143.315 -149.765 143.645 -149.435 ;
        RECT 143.315 -151.125 143.645 -150.795 ;
        RECT 143.315 -152.485 143.645 -152.155 ;
        RECT 143.315 -153.845 143.645 -153.515 ;
        RECT 143.315 -155.205 143.645 -154.875 ;
        RECT 143.315 -156.565 143.645 -156.235 ;
        RECT 143.315 -157.925 143.645 -157.595 ;
        RECT 143.315 -159.285 143.645 -158.955 ;
        RECT 143.315 -160.645 143.645 -160.315 ;
        RECT 143.315 -162.005 143.645 -161.675 ;
        RECT 143.315 -163.365 143.645 -163.035 ;
        RECT 143.315 -164.725 143.645 -164.395 ;
        RECT 143.315 -166.085 143.645 -165.755 ;
        RECT 143.315 -167.445 143.645 -167.115 ;
        RECT 143.315 -168.805 143.645 -168.475 ;
        RECT 143.315 -170.165 143.645 -169.835 ;
        RECT 143.315 -171.525 143.645 -171.195 ;
        RECT 143.315 -172.885 143.645 -172.555 ;
        RECT 143.315 -174.245 143.645 -173.915 ;
        RECT 143.315 -175.605 143.645 -175.275 ;
        RECT 143.315 -176.965 143.645 -176.635 ;
        RECT 143.315 -178.325 143.645 -177.995 ;
        RECT 143.315 -179.685 143.645 -179.355 ;
        RECT 143.315 -181.93 143.645 -180.8 ;
        RECT 143.32 -182.045 143.64 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 241.32 145.005 242.45 ;
        RECT 144.675 239.195 145.005 239.525 ;
        RECT 144.675 237.835 145.005 238.165 ;
        RECT 144.68 237.16 145 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 144.675 -99.445 145.005 -99.115 ;
        RECT 144.675 -100.805 145.005 -100.475 ;
        RECT 144.675 -102.165 145.005 -101.835 ;
        RECT 144.675 -103.525 145.005 -103.195 ;
        RECT 144.675 -104.885 145.005 -104.555 ;
        RECT 144.675 -106.245 145.005 -105.915 ;
        RECT 144.675 -107.605 145.005 -107.275 ;
        RECT 144.675 -108.965 145.005 -108.635 ;
        RECT 144.675 -110.325 145.005 -109.995 ;
        RECT 144.675 -111.685 145.005 -111.355 ;
        RECT 144.675 -113.045 145.005 -112.715 ;
        RECT 144.675 -114.405 145.005 -114.075 ;
        RECT 144.675 -115.765 145.005 -115.435 ;
        RECT 144.675 -117.125 145.005 -116.795 ;
        RECT 144.675 -118.485 145.005 -118.155 ;
        RECT 144.675 -119.845 145.005 -119.515 ;
        RECT 144.675 -121.205 145.005 -120.875 ;
        RECT 144.675 -122.565 145.005 -122.235 ;
        RECT 144.675 -123.925 145.005 -123.595 ;
        RECT 144.675 -125.285 145.005 -124.955 ;
        RECT 144.675 -126.645 145.005 -126.315 ;
        RECT 144.675 -128.005 145.005 -127.675 ;
        RECT 144.675 -129.365 145.005 -129.035 ;
        RECT 144.675 -130.725 145.005 -130.395 ;
        RECT 144.675 -132.085 145.005 -131.755 ;
        RECT 144.675 -133.445 145.005 -133.115 ;
        RECT 144.675 -134.805 145.005 -134.475 ;
        RECT 144.675 -136.165 145.005 -135.835 ;
        RECT 144.675 -137.525 145.005 -137.195 ;
        RECT 144.675 -138.885 145.005 -138.555 ;
        RECT 144.675 -140.245 145.005 -139.915 ;
        RECT 144.675 -141.605 145.005 -141.275 ;
        RECT 144.675 -142.965 145.005 -142.635 ;
        RECT 144.675 -144.325 145.005 -143.995 ;
        RECT 144.675 -145.685 145.005 -145.355 ;
        RECT 144.675 -147.045 145.005 -146.715 ;
        RECT 144.675 -148.405 145.005 -148.075 ;
        RECT 144.675 -149.765 145.005 -149.435 ;
        RECT 144.675 -151.125 145.005 -150.795 ;
        RECT 144.675 -152.485 145.005 -152.155 ;
        RECT 144.675 -153.845 145.005 -153.515 ;
        RECT 144.675 -155.205 145.005 -154.875 ;
        RECT 144.675 -156.565 145.005 -156.235 ;
        RECT 144.675 -157.925 145.005 -157.595 ;
        RECT 144.675 -159.285 145.005 -158.955 ;
        RECT 144.675 -160.645 145.005 -160.315 ;
        RECT 144.675 -162.005 145.005 -161.675 ;
        RECT 144.675 -163.365 145.005 -163.035 ;
        RECT 144.675 -164.725 145.005 -164.395 ;
        RECT 144.675 -166.085 145.005 -165.755 ;
        RECT 144.675 -167.445 145.005 -167.115 ;
        RECT 144.675 -168.805 145.005 -168.475 ;
        RECT 144.675 -170.165 145.005 -169.835 ;
        RECT 144.675 -171.525 145.005 -171.195 ;
        RECT 144.675 -172.885 145.005 -172.555 ;
        RECT 144.675 -174.245 145.005 -173.915 ;
        RECT 144.675 -175.605 145.005 -175.275 ;
        RECT 144.675 -176.965 145.005 -176.635 ;
        RECT 144.675 -178.325 145.005 -177.995 ;
        RECT 144.675 -179.685 145.005 -179.355 ;
        RECT 144.675 -181.93 145.005 -180.8 ;
        RECT 144.68 -182.045 145 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 145.01 -98.075 145.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 241.32 146.365 242.45 ;
        RECT 146.035 239.195 146.365 239.525 ;
        RECT 146.035 237.835 146.365 238.165 ;
        RECT 146.04 237.16 146.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 146.035 -1.525 146.365 -1.195 ;
        RECT 146.035 -2.885 146.365 -2.555 ;
        RECT 146.04 -3.56 146.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 241.32 147.725 242.45 ;
        RECT 147.395 239.195 147.725 239.525 ;
        RECT 147.395 237.835 147.725 238.165 ;
        RECT 147.4 237.16 147.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 147.395 -1.525 147.725 -1.195 ;
        RECT 147.395 -2.885 147.725 -2.555 ;
        RECT 147.4 -3.56 147.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 241.32 149.085 242.45 ;
        RECT 148.755 239.195 149.085 239.525 ;
        RECT 148.755 237.835 149.085 238.165 ;
        RECT 148.76 237.16 149.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 -1.525 149.085 -1.195 ;
        RECT 148.755 -2.885 149.085 -2.555 ;
        RECT 148.76 -3.56 149.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 148.755 -95.365 149.085 -95.035 ;
        RECT 148.755 -96.725 149.085 -96.395 ;
        RECT 148.755 -98.085 149.085 -97.755 ;
        RECT 148.755 -99.445 149.085 -99.115 ;
        RECT 148.755 -100.805 149.085 -100.475 ;
        RECT 148.755 -102.165 149.085 -101.835 ;
        RECT 148.755 -103.525 149.085 -103.195 ;
        RECT 148.755 -104.885 149.085 -104.555 ;
        RECT 148.755 -106.245 149.085 -105.915 ;
        RECT 148.755 -107.605 149.085 -107.275 ;
        RECT 148.755 -108.965 149.085 -108.635 ;
        RECT 148.755 -110.325 149.085 -109.995 ;
        RECT 148.755 -111.685 149.085 -111.355 ;
        RECT 148.755 -113.045 149.085 -112.715 ;
        RECT 148.755 -114.405 149.085 -114.075 ;
        RECT 148.755 -115.765 149.085 -115.435 ;
        RECT 148.755 -117.125 149.085 -116.795 ;
        RECT 148.755 -118.485 149.085 -118.155 ;
        RECT 148.755 -119.845 149.085 -119.515 ;
        RECT 148.755 -121.205 149.085 -120.875 ;
        RECT 148.755 -122.565 149.085 -122.235 ;
        RECT 148.755 -123.925 149.085 -123.595 ;
        RECT 148.755 -125.285 149.085 -124.955 ;
        RECT 148.755 -126.645 149.085 -126.315 ;
        RECT 148.755 -128.005 149.085 -127.675 ;
        RECT 148.755 -129.365 149.085 -129.035 ;
        RECT 148.755 -130.725 149.085 -130.395 ;
        RECT 148.755 -132.085 149.085 -131.755 ;
        RECT 148.755 -133.445 149.085 -133.115 ;
        RECT 148.755 -134.805 149.085 -134.475 ;
        RECT 148.755 -136.165 149.085 -135.835 ;
        RECT 148.755 -137.525 149.085 -137.195 ;
        RECT 148.755 -138.885 149.085 -138.555 ;
        RECT 148.755 -140.245 149.085 -139.915 ;
        RECT 148.755 -141.605 149.085 -141.275 ;
        RECT 148.755 -142.965 149.085 -142.635 ;
        RECT 148.755 -144.325 149.085 -143.995 ;
        RECT 148.755 -145.685 149.085 -145.355 ;
        RECT 148.755 -147.045 149.085 -146.715 ;
        RECT 148.755 -148.405 149.085 -148.075 ;
        RECT 148.755 -149.765 149.085 -149.435 ;
        RECT 148.755 -151.125 149.085 -150.795 ;
        RECT 148.755 -152.485 149.085 -152.155 ;
        RECT 148.755 -153.845 149.085 -153.515 ;
        RECT 148.755 -155.205 149.085 -154.875 ;
        RECT 148.755 -156.565 149.085 -156.235 ;
        RECT 148.755 -157.925 149.085 -157.595 ;
        RECT 148.755 -159.285 149.085 -158.955 ;
        RECT 148.755 -160.645 149.085 -160.315 ;
        RECT 148.755 -162.005 149.085 -161.675 ;
        RECT 148.755 -163.365 149.085 -163.035 ;
        RECT 148.755 -164.725 149.085 -164.395 ;
        RECT 148.755 -166.085 149.085 -165.755 ;
        RECT 148.755 -167.445 149.085 -167.115 ;
        RECT 148.755 -168.805 149.085 -168.475 ;
        RECT 148.755 -170.165 149.085 -169.835 ;
        RECT 148.755 -171.525 149.085 -171.195 ;
        RECT 148.755 -172.885 149.085 -172.555 ;
        RECT 148.755 -174.245 149.085 -173.915 ;
        RECT 148.755 -175.605 149.085 -175.275 ;
        RECT 148.755 -176.965 149.085 -176.635 ;
        RECT 148.755 -178.325 149.085 -177.995 ;
        RECT 148.755 -179.685 149.085 -179.355 ;
        RECT 148.755 -181.93 149.085 -180.8 ;
        RECT 148.76 -182.045 149.08 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.115 241.32 150.445 242.45 ;
        RECT 150.115 239.195 150.445 239.525 ;
        RECT 150.115 237.835 150.445 238.165 ;
        RECT 150.12 237.16 150.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.115 -1.525 150.445 -1.195 ;
        RECT 150.115 -2.885 150.445 -2.555 ;
        RECT 150.12 -3.56 150.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 150.115 -95.365 150.445 -95.035 ;
        RECT 150.115 -96.725 150.445 -96.395 ;
        RECT 150.115 -98.085 150.445 -97.755 ;
        RECT 150.115 -99.445 150.445 -99.115 ;
        RECT 150.115 -100.805 150.445 -100.475 ;
        RECT 150.115 -102.165 150.445 -101.835 ;
        RECT 150.115 -103.525 150.445 -103.195 ;
        RECT 150.115 -104.885 150.445 -104.555 ;
        RECT 150.115 -106.245 150.445 -105.915 ;
        RECT 150.115 -107.605 150.445 -107.275 ;
        RECT 150.115 -108.965 150.445 -108.635 ;
        RECT 150.115 -110.325 150.445 -109.995 ;
        RECT 150.115 -111.685 150.445 -111.355 ;
        RECT 150.115 -113.045 150.445 -112.715 ;
        RECT 150.115 -114.405 150.445 -114.075 ;
        RECT 150.115 -115.765 150.445 -115.435 ;
        RECT 150.115 -117.125 150.445 -116.795 ;
        RECT 150.115 -118.485 150.445 -118.155 ;
        RECT 150.115 -119.845 150.445 -119.515 ;
        RECT 150.115 -121.205 150.445 -120.875 ;
        RECT 150.115 -122.565 150.445 -122.235 ;
        RECT 150.115 -123.925 150.445 -123.595 ;
        RECT 150.115 -125.285 150.445 -124.955 ;
        RECT 150.115 -126.645 150.445 -126.315 ;
        RECT 150.115 -128.005 150.445 -127.675 ;
        RECT 150.115 -129.365 150.445 -129.035 ;
        RECT 150.115 -130.725 150.445 -130.395 ;
        RECT 150.115 -132.085 150.445 -131.755 ;
        RECT 150.115 -133.445 150.445 -133.115 ;
        RECT 150.115 -134.805 150.445 -134.475 ;
        RECT 150.115 -136.165 150.445 -135.835 ;
        RECT 150.115 -137.525 150.445 -137.195 ;
        RECT 150.115 -138.885 150.445 -138.555 ;
        RECT 150.115 -140.245 150.445 -139.915 ;
        RECT 150.115 -141.605 150.445 -141.275 ;
        RECT 150.115 -142.965 150.445 -142.635 ;
        RECT 150.115 -144.325 150.445 -143.995 ;
        RECT 150.115 -145.685 150.445 -145.355 ;
        RECT 150.115 -147.045 150.445 -146.715 ;
        RECT 150.115 -148.405 150.445 -148.075 ;
        RECT 150.115 -149.765 150.445 -149.435 ;
        RECT 150.115 -151.125 150.445 -150.795 ;
        RECT 150.115 -152.485 150.445 -152.155 ;
        RECT 150.115 -153.845 150.445 -153.515 ;
        RECT 150.115 -155.205 150.445 -154.875 ;
        RECT 150.115 -156.565 150.445 -156.235 ;
        RECT 150.115 -157.925 150.445 -157.595 ;
        RECT 150.115 -159.285 150.445 -158.955 ;
        RECT 150.115 -160.645 150.445 -160.315 ;
        RECT 150.115 -162.005 150.445 -161.675 ;
        RECT 150.115 -163.365 150.445 -163.035 ;
        RECT 150.115 -164.725 150.445 -164.395 ;
        RECT 150.115 -166.085 150.445 -165.755 ;
        RECT 150.115 -167.445 150.445 -167.115 ;
        RECT 150.115 -168.805 150.445 -168.475 ;
        RECT 150.115 -170.165 150.445 -169.835 ;
        RECT 150.115 -171.525 150.445 -171.195 ;
        RECT 150.115 -172.885 150.445 -172.555 ;
        RECT 150.115 -174.245 150.445 -173.915 ;
        RECT 150.115 -175.605 150.445 -175.275 ;
        RECT 150.115 -176.965 150.445 -176.635 ;
        RECT 150.115 -178.325 150.445 -177.995 ;
        RECT 150.115 -179.685 150.445 -179.355 ;
        RECT 150.115 -181.93 150.445 -180.8 ;
        RECT 150.12 -182.045 150.44 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 241.32 151.805 242.45 ;
        RECT 151.475 239.195 151.805 239.525 ;
        RECT 151.475 237.835 151.805 238.165 ;
        RECT 151.48 237.16 151.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 -1.525 151.805 -1.195 ;
        RECT 151.475 -2.885 151.805 -2.555 ;
        RECT 151.48 -3.56 151.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 151.475 -95.365 151.805 -95.035 ;
        RECT 151.475 -96.725 151.805 -96.395 ;
        RECT 151.475 -98.085 151.805 -97.755 ;
        RECT 151.475 -99.445 151.805 -99.115 ;
        RECT 151.475 -100.805 151.805 -100.475 ;
        RECT 151.475 -102.165 151.805 -101.835 ;
        RECT 151.475 -103.525 151.805 -103.195 ;
        RECT 151.475 -104.885 151.805 -104.555 ;
        RECT 151.475 -106.245 151.805 -105.915 ;
        RECT 151.475 -107.605 151.805 -107.275 ;
        RECT 151.475 -108.965 151.805 -108.635 ;
        RECT 151.475 -110.325 151.805 -109.995 ;
        RECT 151.475 -111.685 151.805 -111.355 ;
        RECT 151.475 -113.045 151.805 -112.715 ;
        RECT 151.475 -114.405 151.805 -114.075 ;
        RECT 151.475 -115.765 151.805 -115.435 ;
        RECT 151.475 -117.125 151.805 -116.795 ;
        RECT 151.475 -118.485 151.805 -118.155 ;
        RECT 151.475 -119.845 151.805 -119.515 ;
        RECT 151.475 -121.205 151.805 -120.875 ;
        RECT 151.475 -122.565 151.805 -122.235 ;
        RECT 151.475 -123.925 151.805 -123.595 ;
        RECT 151.475 -125.285 151.805 -124.955 ;
        RECT 151.475 -126.645 151.805 -126.315 ;
        RECT 151.475 -128.005 151.805 -127.675 ;
        RECT 151.475 -129.365 151.805 -129.035 ;
        RECT 151.475 -130.725 151.805 -130.395 ;
        RECT 151.475 -132.085 151.805 -131.755 ;
        RECT 151.475 -133.445 151.805 -133.115 ;
        RECT 151.475 -134.805 151.805 -134.475 ;
        RECT 151.475 -136.165 151.805 -135.835 ;
        RECT 151.475 -137.525 151.805 -137.195 ;
        RECT 151.475 -138.885 151.805 -138.555 ;
        RECT 151.475 -140.245 151.805 -139.915 ;
        RECT 151.475 -141.605 151.805 -141.275 ;
        RECT 151.475 -142.965 151.805 -142.635 ;
        RECT 151.475 -144.325 151.805 -143.995 ;
        RECT 151.475 -145.685 151.805 -145.355 ;
        RECT 151.475 -147.045 151.805 -146.715 ;
        RECT 151.475 -148.405 151.805 -148.075 ;
        RECT 151.475 -149.765 151.805 -149.435 ;
        RECT 151.475 -151.125 151.805 -150.795 ;
        RECT 151.475 -152.485 151.805 -152.155 ;
        RECT 151.475 -153.845 151.805 -153.515 ;
        RECT 151.475 -155.205 151.805 -154.875 ;
        RECT 151.475 -156.565 151.805 -156.235 ;
        RECT 151.475 -157.925 151.805 -157.595 ;
        RECT 151.475 -159.285 151.805 -158.955 ;
        RECT 151.475 -160.645 151.805 -160.315 ;
        RECT 151.475 -162.005 151.805 -161.675 ;
        RECT 151.475 -163.365 151.805 -163.035 ;
        RECT 151.475 -164.725 151.805 -164.395 ;
        RECT 151.475 -166.085 151.805 -165.755 ;
        RECT 151.475 -167.445 151.805 -167.115 ;
        RECT 151.475 -168.805 151.805 -168.475 ;
        RECT 151.475 -170.165 151.805 -169.835 ;
        RECT 151.475 -171.525 151.805 -171.195 ;
        RECT 151.475 -172.885 151.805 -172.555 ;
        RECT 151.475 -174.245 151.805 -173.915 ;
        RECT 151.475 -175.605 151.805 -175.275 ;
        RECT 151.475 -176.965 151.805 -176.635 ;
        RECT 151.475 -178.325 151.805 -177.995 ;
        RECT 151.475 -179.685 151.805 -179.355 ;
        RECT 151.475 -181.93 151.805 -180.8 ;
        RECT 151.48 -182.045 151.8 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 241.32 153.165 242.45 ;
        RECT 152.835 239.195 153.165 239.525 ;
        RECT 152.835 237.835 153.165 238.165 ;
        RECT 152.84 237.16 153.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 -1.525 153.165 -1.195 ;
        RECT 152.835 -2.885 153.165 -2.555 ;
        RECT 152.84 -3.56 153.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 152.835 -95.365 153.165 -95.035 ;
        RECT 152.835 -96.725 153.165 -96.395 ;
        RECT 152.835 -98.085 153.165 -97.755 ;
        RECT 152.835 -99.445 153.165 -99.115 ;
        RECT 152.835 -100.805 153.165 -100.475 ;
        RECT 152.835 -102.165 153.165 -101.835 ;
        RECT 152.835 -103.525 153.165 -103.195 ;
        RECT 152.835 -104.885 153.165 -104.555 ;
        RECT 152.835 -106.245 153.165 -105.915 ;
        RECT 152.835 -107.605 153.165 -107.275 ;
        RECT 152.835 -108.965 153.165 -108.635 ;
        RECT 152.835 -110.325 153.165 -109.995 ;
        RECT 152.835 -111.685 153.165 -111.355 ;
        RECT 152.835 -113.045 153.165 -112.715 ;
        RECT 152.835 -114.405 153.165 -114.075 ;
        RECT 152.835 -115.765 153.165 -115.435 ;
        RECT 152.835 -117.125 153.165 -116.795 ;
        RECT 152.835 -118.485 153.165 -118.155 ;
        RECT 152.835 -119.845 153.165 -119.515 ;
        RECT 152.835 -121.205 153.165 -120.875 ;
        RECT 152.835 -122.565 153.165 -122.235 ;
        RECT 152.835 -123.925 153.165 -123.595 ;
        RECT 152.835 -125.285 153.165 -124.955 ;
        RECT 152.835 -126.645 153.165 -126.315 ;
        RECT 152.835 -128.005 153.165 -127.675 ;
        RECT 152.835 -129.365 153.165 -129.035 ;
        RECT 152.835 -130.725 153.165 -130.395 ;
        RECT 152.835 -132.085 153.165 -131.755 ;
        RECT 152.835 -133.445 153.165 -133.115 ;
        RECT 152.835 -134.805 153.165 -134.475 ;
        RECT 152.835 -136.165 153.165 -135.835 ;
        RECT 152.835 -137.525 153.165 -137.195 ;
        RECT 152.835 -138.885 153.165 -138.555 ;
        RECT 152.835 -140.245 153.165 -139.915 ;
        RECT 152.835 -141.605 153.165 -141.275 ;
        RECT 152.835 -142.965 153.165 -142.635 ;
        RECT 152.835 -144.325 153.165 -143.995 ;
        RECT 152.835 -145.685 153.165 -145.355 ;
        RECT 152.835 -147.045 153.165 -146.715 ;
        RECT 152.835 -148.405 153.165 -148.075 ;
        RECT 152.835 -149.765 153.165 -149.435 ;
        RECT 152.835 -151.125 153.165 -150.795 ;
        RECT 152.835 -152.485 153.165 -152.155 ;
        RECT 152.835 -153.845 153.165 -153.515 ;
        RECT 152.835 -155.205 153.165 -154.875 ;
        RECT 152.835 -156.565 153.165 -156.235 ;
        RECT 152.835 -157.925 153.165 -157.595 ;
        RECT 152.835 -159.285 153.165 -158.955 ;
        RECT 152.835 -160.645 153.165 -160.315 ;
        RECT 152.835 -162.005 153.165 -161.675 ;
        RECT 152.835 -163.365 153.165 -163.035 ;
        RECT 152.835 -164.725 153.165 -164.395 ;
        RECT 152.835 -166.085 153.165 -165.755 ;
        RECT 152.835 -167.445 153.165 -167.115 ;
        RECT 152.835 -168.805 153.165 -168.475 ;
        RECT 152.835 -170.165 153.165 -169.835 ;
        RECT 152.835 -171.525 153.165 -171.195 ;
        RECT 152.835 -172.885 153.165 -172.555 ;
        RECT 152.835 -174.245 153.165 -173.915 ;
        RECT 152.835 -175.605 153.165 -175.275 ;
        RECT 152.835 -176.965 153.165 -176.635 ;
        RECT 152.835 -178.325 153.165 -177.995 ;
        RECT 152.835 -179.685 153.165 -179.355 ;
        RECT 152.835 -181.93 153.165 -180.8 ;
        RECT 152.84 -182.045 153.16 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 241.32 154.525 242.45 ;
        RECT 154.195 239.195 154.525 239.525 ;
        RECT 154.195 237.835 154.525 238.165 ;
        RECT 154.2 237.16 154.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 -1.525 154.525 -1.195 ;
        RECT 154.195 -2.885 154.525 -2.555 ;
        RECT 154.2 -3.56 154.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 154.195 -95.365 154.525 -95.035 ;
        RECT 154.195 -96.725 154.525 -96.395 ;
        RECT 154.195 -98.085 154.525 -97.755 ;
        RECT 154.195 -99.445 154.525 -99.115 ;
        RECT 154.195 -100.805 154.525 -100.475 ;
        RECT 154.195 -102.165 154.525 -101.835 ;
        RECT 154.195 -103.525 154.525 -103.195 ;
        RECT 154.195 -104.885 154.525 -104.555 ;
        RECT 154.195 -106.245 154.525 -105.915 ;
        RECT 154.195 -107.605 154.525 -107.275 ;
        RECT 154.195 -108.965 154.525 -108.635 ;
        RECT 154.195 -110.325 154.525 -109.995 ;
        RECT 154.195 -111.685 154.525 -111.355 ;
        RECT 154.195 -113.045 154.525 -112.715 ;
        RECT 154.195 -114.405 154.525 -114.075 ;
        RECT 154.195 -115.765 154.525 -115.435 ;
        RECT 154.195 -117.125 154.525 -116.795 ;
        RECT 154.195 -118.485 154.525 -118.155 ;
        RECT 154.195 -119.845 154.525 -119.515 ;
        RECT 154.195 -121.205 154.525 -120.875 ;
        RECT 154.195 -122.565 154.525 -122.235 ;
        RECT 154.195 -123.925 154.525 -123.595 ;
        RECT 154.195 -125.285 154.525 -124.955 ;
        RECT 154.195 -126.645 154.525 -126.315 ;
        RECT 154.195 -128.005 154.525 -127.675 ;
        RECT 154.195 -129.365 154.525 -129.035 ;
        RECT 154.195 -130.725 154.525 -130.395 ;
        RECT 154.195 -132.085 154.525 -131.755 ;
        RECT 154.195 -133.445 154.525 -133.115 ;
        RECT 154.195 -134.805 154.525 -134.475 ;
        RECT 154.195 -136.165 154.525 -135.835 ;
        RECT 154.195 -137.525 154.525 -137.195 ;
        RECT 154.195 -138.885 154.525 -138.555 ;
        RECT 154.195 -140.245 154.525 -139.915 ;
        RECT 154.195 -141.605 154.525 -141.275 ;
        RECT 154.195 -142.965 154.525 -142.635 ;
        RECT 154.195 -144.325 154.525 -143.995 ;
        RECT 154.195 -145.685 154.525 -145.355 ;
        RECT 154.195 -147.045 154.525 -146.715 ;
        RECT 154.195 -148.405 154.525 -148.075 ;
        RECT 154.195 -149.765 154.525 -149.435 ;
        RECT 154.195 -151.125 154.525 -150.795 ;
        RECT 154.195 -152.485 154.525 -152.155 ;
        RECT 154.195 -153.845 154.525 -153.515 ;
        RECT 154.195 -155.205 154.525 -154.875 ;
        RECT 154.195 -156.565 154.525 -156.235 ;
        RECT 154.195 -157.925 154.525 -157.595 ;
        RECT 154.195 -159.285 154.525 -158.955 ;
        RECT 154.195 -160.645 154.525 -160.315 ;
        RECT 154.195 -162.005 154.525 -161.675 ;
        RECT 154.195 -163.365 154.525 -163.035 ;
        RECT 154.195 -164.725 154.525 -164.395 ;
        RECT 154.195 -166.085 154.525 -165.755 ;
        RECT 154.195 -167.445 154.525 -167.115 ;
        RECT 154.195 -168.805 154.525 -168.475 ;
        RECT 154.195 -170.165 154.525 -169.835 ;
        RECT 154.195 -171.525 154.525 -171.195 ;
        RECT 154.195 -172.885 154.525 -172.555 ;
        RECT 154.195 -174.245 154.525 -173.915 ;
        RECT 154.195 -175.605 154.525 -175.275 ;
        RECT 154.195 -176.965 154.525 -176.635 ;
        RECT 154.195 -178.325 154.525 -177.995 ;
        RECT 154.195 -179.685 154.525 -179.355 ;
        RECT 154.195 -181.93 154.525 -180.8 ;
        RECT 154.2 -182.045 154.52 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 241.32 155.885 242.45 ;
        RECT 155.555 239.195 155.885 239.525 ;
        RECT 155.555 237.835 155.885 238.165 ;
        RECT 155.56 237.16 155.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.555 -99.445 155.885 -99.115 ;
        RECT 155.555 -100.805 155.885 -100.475 ;
        RECT 155.555 -102.165 155.885 -101.835 ;
        RECT 155.555 -103.525 155.885 -103.195 ;
        RECT 155.555 -104.885 155.885 -104.555 ;
        RECT 155.555 -106.245 155.885 -105.915 ;
        RECT 155.555 -107.605 155.885 -107.275 ;
        RECT 155.555 -108.965 155.885 -108.635 ;
        RECT 155.555 -110.325 155.885 -109.995 ;
        RECT 155.555 -111.685 155.885 -111.355 ;
        RECT 155.555 -113.045 155.885 -112.715 ;
        RECT 155.555 -114.405 155.885 -114.075 ;
        RECT 155.555 -115.765 155.885 -115.435 ;
        RECT 155.555 -117.125 155.885 -116.795 ;
        RECT 155.555 -118.485 155.885 -118.155 ;
        RECT 155.555 -119.845 155.885 -119.515 ;
        RECT 155.555 -121.205 155.885 -120.875 ;
        RECT 155.555 -122.565 155.885 -122.235 ;
        RECT 155.555 -123.925 155.885 -123.595 ;
        RECT 155.555 -125.285 155.885 -124.955 ;
        RECT 155.555 -126.645 155.885 -126.315 ;
        RECT 155.555 -128.005 155.885 -127.675 ;
        RECT 155.555 -129.365 155.885 -129.035 ;
        RECT 155.555 -130.725 155.885 -130.395 ;
        RECT 155.555 -132.085 155.885 -131.755 ;
        RECT 155.555 -133.445 155.885 -133.115 ;
        RECT 155.555 -134.805 155.885 -134.475 ;
        RECT 155.555 -136.165 155.885 -135.835 ;
        RECT 155.555 -137.525 155.885 -137.195 ;
        RECT 155.555 -138.885 155.885 -138.555 ;
        RECT 155.555 -140.245 155.885 -139.915 ;
        RECT 155.555 -141.605 155.885 -141.275 ;
        RECT 155.555 -142.965 155.885 -142.635 ;
        RECT 155.555 -144.325 155.885 -143.995 ;
        RECT 155.555 -145.685 155.885 -145.355 ;
        RECT 155.555 -147.045 155.885 -146.715 ;
        RECT 155.555 -148.405 155.885 -148.075 ;
        RECT 155.555 -149.765 155.885 -149.435 ;
        RECT 155.555 -151.125 155.885 -150.795 ;
        RECT 155.555 -152.485 155.885 -152.155 ;
        RECT 155.555 -153.845 155.885 -153.515 ;
        RECT 155.555 -155.205 155.885 -154.875 ;
        RECT 155.555 -156.565 155.885 -156.235 ;
        RECT 155.555 -157.925 155.885 -157.595 ;
        RECT 155.555 -159.285 155.885 -158.955 ;
        RECT 155.555 -160.645 155.885 -160.315 ;
        RECT 155.555 -162.005 155.885 -161.675 ;
        RECT 155.555 -163.365 155.885 -163.035 ;
        RECT 155.555 -164.725 155.885 -164.395 ;
        RECT 155.555 -166.085 155.885 -165.755 ;
        RECT 155.555 -167.445 155.885 -167.115 ;
        RECT 155.555 -168.805 155.885 -168.475 ;
        RECT 155.555 -170.165 155.885 -169.835 ;
        RECT 155.555 -171.525 155.885 -171.195 ;
        RECT 155.555 -172.885 155.885 -172.555 ;
        RECT 155.555 -174.245 155.885 -173.915 ;
        RECT 155.555 -175.605 155.885 -175.275 ;
        RECT 155.555 -176.965 155.885 -176.635 ;
        RECT 155.555 -178.325 155.885 -177.995 ;
        RECT 155.555 -179.685 155.885 -179.355 ;
        RECT 155.555 -181.93 155.885 -180.8 ;
        RECT 155.56 -182.045 155.88 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 155.91 -98.075 156.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 241.32 157.245 242.45 ;
        RECT 156.915 239.195 157.245 239.525 ;
        RECT 156.915 237.835 157.245 238.165 ;
        RECT 156.92 237.16 157.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 156.915 -1.525 157.245 -1.195 ;
        RECT 156.915 -2.885 157.245 -2.555 ;
        RECT 156.92 -3.56 157.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 241.32 158.605 242.45 ;
        RECT 158.275 239.195 158.605 239.525 ;
        RECT 158.275 237.835 158.605 238.165 ;
        RECT 158.28 237.16 158.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 158.275 -1.525 158.605 -1.195 ;
        RECT 158.275 -2.885 158.605 -2.555 ;
        RECT 158.28 -3.56 158.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 241.32 159.965 242.45 ;
        RECT 159.635 239.195 159.965 239.525 ;
        RECT 159.635 237.835 159.965 238.165 ;
        RECT 159.64 237.16 159.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 -1.525 159.965 -1.195 ;
        RECT 159.635 -2.885 159.965 -2.555 ;
        RECT 159.64 -3.56 159.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 159.635 -95.365 159.965 -95.035 ;
        RECT 159.635 -96.725 159.965 -96.395 ;
        RECT 159.635 -98.085 159.965 -97.755 ;
        RECT 159.635 -99.445 159.965 -99.115 ;
        RECT 159.635 -100.805 159.965 -100.475 ;
        RECT 159.635 -102.165 159.965 -101.835 ;
        RECT 159.635 -103.525 159.965 -103.195 ;
        RECT 159.635 -104.885 159.965 -104.555 ;
        RECT 159.635 -106.245 159.965 -105.915 ;
        RECT 159.635 -107.605 159.965 -107.275 ;
        RECT 159.635 -108.965 159.965 -108.635 ;
        RECT 159.635 -110.325 159.965 -109.995 ;
        RECT 159.635 -111.685 159.965 -111.355 ;
        RECT 159.635 -113.045 159.965 -112.715 ;
        RECT 159.635 -114.405 159.965 -114.075 ;
        RECT 159.635 -115.765 159.965 -115.435 ;
        RECT 159.635 -117.125 159.965 -116.795 ;
        RECT 159.635 -118.485 159.965 -118.155 ;
        RECT 159.635 -119.845 159.965 -119.515 ;
        RECT 159.635 -121.205 159.965 -120.875 ;
        RECT 159.635 -122.565 159.965 -122.235 ;
        RECT 159.635 -123.925 159.965 -123.595 ;
        RECT 159.635 -125.285 159.965 -124.955 ;
        RECT 159.635 -126.645 159.965 -126.315 ;
        RECT 159.635 -128.005 159.965 -127.675 ;
        RECT 159.635 -129.365 159.965 -129.035 ;
        RECT 159.635 -130.725 159.965 -130.395 ;
        RECT 159.635 -132.085 159.965 -131.755 ;
        RECT 159.635 -133.445 159.965 -133.115 ;
        RECT 159.635 -134.805 159.965 -134.475 ;
        RECT 159.635 -136.165 159.965 -135.835 ;
        RECT 159.635 -137.525 159.965 -137.195 ;
        RECT 159.635 -138.885 159.965 -138.555 ;
        RECT 159.635 -140.245 159.965 -139.915 ;
        RECT 159.635 -141.605 159.965 -141.275 ;
        RECT 159.635 -142.965 159.965 -142.635 ;
        RECT 159.635 -144.325 159.965 -143.995 ;
        RECT 159.635 -145.685 159.965 -145.355 ;
        RECT 159.635 -147.045 159.965 -146.715 ;
        RECT 159.635 -148.405 159.965 -148.075 ;
        RECT 159.635 -149.765 159.965 -149.435 ;
        RECT 159.635 -151.125 159.965 -150.795 ;
        RECT 159.635 -152.485 159.965 -152.155 ;
        RECT 159.635 -153.845 159.965 -153.515 ;
        RECT 159.635 -155.205 159.965 -154.875 ;
        RECT 159.635 -156.565 159.965 -156.235 ;
        RECT 159.635 -157.925 159.965 -157.595 ;
        RECT 159.635 -159.285 159.965 -158.955 ;
        RECT 159.635 -160.645 159.965 -160.315 ;
        RECT 159.635 -162.005 159.965 -161.675 ;
        RECT 159.635 -163.365 159.965 -163.035 ;
        RECT 159.635 -164.725 159.965 -164.395 ;
        RECT 159.635 -166.085 159.965 -165.755 ;
        RECT 159.635 -167.445 159.965 -167.115 ;
        RECT 159.635 -168.805 159.965 -168.475 ;
        RECT 159.635 -170.165 159.965 -169.835 ;
        RECT 159.635 -171.525 159.965 -171.195 ;
        RECT 159.635 -172.885 159.965 -172.555 ;
        RECT 159.635 -174.245 159.965 -173.915 ;
        RECT 159.635 -175.605 159.965 -175.275 ;
        RECT 159.635 -176.965 159.965 -176.635 ;
        RECT 159.635 -178.325 159.965 -177.995 ;
        RECT 159.635 -179.685 159.965 -179.355 ;
        RECT 159.635 -181.93 159.965 -180.8 ;
        RECT 159.64 -182.045 159.96 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 241.32 161.325 242.45 ;
        RECT 160.995 239.195 161.325 239.525 ;
        RECT 160.995 237.835 161.325 238.165 ;
        RECT 161 237.16 161.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 -1.525 161.325 -1.195 ;
        RECT 160.995 -2.885 161.325 -2.555 ;
        RECT 161 -3.56 161.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 160.995 -95.365 161.325 -95.035 ;
        RECT 160.995 -96.725 161.325 -96.395 ;
        RECT 160.995 -98.085 161.325 -97.755 ;
        RECT 160.995 -99.445 161.325 -99.115 ;
        RECT 160.995 -100.805 161.325 -100.475 ;
        RECT 160.995 -102.165 161.325 -101.835 ;
        RECT 160.995 -103.525 161.325 -103.195 ;
        RECT 160.995 -104.885 161.325 -104.555 ;
        RECT 160.995 -106.245 161.325 -105.915 ;
        RECT 160.995 -107.605 161.325 -107.275 ;
        RECT 160.995 -108.965 161.325 -108.635 ;
        RECT 160.995 -110.325 161.325 -109.995 ;
        RECT 160.995 -111.685 161.325 -111.355 ;
        RECT 160.995 -113.045 161.325 -112.715 ;
        RECT 160.995 -114.405 161.325 -114.075 ;
        RECT 160.995 -115.765 161.325 -115.435 ;
        RECT 160.995 -117.125 161.325 -116.795 ;
        RECT 160.995 -118.485 161.325 -118.155 ;
        RECT 160.995 -119.845 161.325 -119.515 ;
        RECT 160.995 -121.205 161.325 -120.875 ;
        RECT 160.995 -122.565 161.325 -122.235 ;
        RECT 160.995 -123.925 161.325 -123.595 ;
        RECT 160.995 -125.285 161.325 -124.955 ;
        RECT 160.995 -126.645 161.325 -126.315 ;
        RECT 160.995 -128.005 161.325 -127.675 ;
        RECT 160.995 -129.365 161.325 -129.035 ;
        RECT 160.995 -130.725 161.325 -130.395 ;
        RECT 160.995 -132.085 161.325 -131.755 ;
        RECT 160.995 -133.445 161.325 -133.115 ;
        RECT 160.995 -134.805 161.325 -134.475 ;
        RECT 160.995 -136.165 161.325 -135.835 ;
        RECT 160.995 -137.525 161.325 -137.195 ;
        RECT 160.995 -138.885 161.325 -138.555 ;
        RECT 160.995 -140.245 161.325 -139.915 ;
        RECT 160.995 -141.605 161.325 -141.275 ;
        RECT 160.995 -142.965 161.325 -142.635 ;
        RECT 160.995 -144.325 161.325 -143.995 ;
        RECT 160.995 -145.685 161.325 -145.355 ;
        RECT 160.995 -147.045 161.325 -146.715 ;
        RECT 160.995 -148.405 161.325 -148.075 ;
        RECT 160.995 -149.765 161.325 -149.435 ;
        RECT 160.995 -151.125 161.325 -150.795 ;
        RECT 160.995 -152.485 161.325 -152.155 ;
        RECT 160.995 -153.845 161.325 -153.515 ;
        RECT 160.995 -155.205 161.325 -154.875 ;
        RECT 160.995 -156.565 161.325 -156.235 ;
        RECT 160.995 -157.925 161.325 -157.595 ;
        RECT 160.995 -159.285 161.325 -158.955 ;
        RECT 160.995 -160.645 161.325 -160.315 ;
        RECT 160.995 -162.005 161.325 -161.675 ;
        RECT 160.995 -163.365 161.325 -163.035 ;
        RECT 160.995 -164.725 161.325 -164.395 ;
        RECT 160.995 -166.085 161.325 -165.755 ;
        RECT 160.995 -167.445 161.325 -167.115 ;
        RECT 160.995 -168.805 161.325 -168.475 ;
        RECT 160.995 -170.165 161.325 -169.835 ;
        RECT 160.995 -171.525 161.325 -171.195 ;
        RECT 160.995 -172.885 161.325 -172.555 ;
        RECT 160.995 -174.245 161.325 -173.915 ;
        RECT 160.995 -175.605 161.325 -175.275 ;
        RECT 160.995 -176.965 161.325 -176.635 ;
        RECT 160.995 -178.325 161.325 -177.995 ;
        RECT 160.995 -179.685 161.325 -179.355 ;
        RECT 160.995 -181.93 161.325 -180.8 ;
        RECT 161 -182.045 161.32 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.355 241.32 162.685 242.45 ;
        RECT 162.355 239.195 162.685 239.525 ;
        RECT 162.355 237.835 162.685 238.165 ;
        RECT 162.36 237.16 162.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.355 -1.525 162.685 -1.195 ;
        RECT 162.355 -2.885 162.685 -2.555 ;
        RECT 162.36 -3.56 162.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 162.355 -95.365 162.685 -95.035 ;
        RECT 162.355 -96.725 162.685 -96.395 ;
        RECT 162.355 -98.085 162.685 -97.755 ;
        RECT 162.355 -99.445 162.685 -99.115 ;
        RECT 162.355 -100.805 162.685 -100.475 ;
        RECT 162.355 -102.165 162.685 -101.835 ;
        RECT 162.355 -103.525 162.685 -103.195 ;
        RECT 162.355 -104.885 162.685 -104.555 ;
        RECT 162.355 -106.245 162.685 -105.915 ;
        RECT 162.355 -107.605 162.685 -107.275 ;
        RECT 162.355 -108.965 162.685 -108.635 ;
        RECT 162.355 -110.325 162.685 -109.995 ;
        RECT 162.355 -111.685 162.685 -111.355 ;
        RECT 162.355 -113.045 162.685 -112.715 ;
        RECT 162.355 -114.405 162.685 -114.075 ;
        RECT 162.355 -115.765 162.685 -115.435 ;
        RECT 162.355 -117.125 162.685 -116.795 ;
        RECT 162.355 -118.485 162.685 -118.155 ;
        RECT 162.355 -119.845 162.685 -119.515 ;
        RECT 162.355 -121.205 162.685 -120.875 ;
        RECT 162.355 -122.565 162.685 -122.235 ;
        RECT 162.355 -123.925 162.685 -123.595 ;
        RECT 162.355 -125.285 162.685 -124.955 ;
        RECT 162.355 -126.645 162.685 -126.315 ;
        RECT 162.355 -128.005 162.685 -127.675 ;
        RECT 162.355 -129.365 162.685 -129.035 ;
        RECT 162.355 -130.725 162.685 -130.395 ;
        RECT 162.355 -132.085 162.685 -131.755 ;
        RECT 162.355 -133.445 162.685 -133.115 ;
        RECT 162.355 -134.805 162.685 -134.475 ;
        RECT 162.355 -136.165 162.685 -135.835 ;
        RECT 162.355 -137.525 162.685 -137.195 ;
        RECT 162.355 -138.885 162.685 -138.555 ;
        RECT 162.355 -140.245 162.685 -139.915 ;
        RECT 162.355 -141.605 162.685 -141.275 ;
        RECT 162.355 -142.965 162.685 -142.635 ;
        RECT 162.355 -144.325 162.685 -143.995 ;
        RECT 162.355 -145.685 162.685 -145.355 ;
        RECT 162.355 -147.045 162.685 -146.715 ;
        RECT 162.355 -148.405 162.685 -148.075 ;
        RECT 162.355 -149.765 162.685 -149.435 ;
        RECT 162.355 -151.125 162.685 -150.795 ;
        RECT 162.355 -152.485 162.685 -152.155 ;
        RECT 162.355 -153.845 162.685 -153.515 ;
        RECT 162.355 -155.205 162.685 -154.875 ;
        RECT 162.355 -156.565 162.685 -156.235 ;
        RECT 162.355 -157.925 162.685 -157.595 ;
        RECT 162.355 -159.285 162.685 -158.955 ;
        RECT 162.355 -160.645 162.685 -160.315 ;
        RECT 162.355 -162.005 162.685 -161.675 ;
        RECT 162.355 -163.365 162.685 -163.035 ;
        RECT 162.355 -164.725 162.685 -164.395 ;
        RECT 162.355 -166.085 162.685 -165.755 ;
        RECT 162.355 -167.445 162.685 -167.115 ;
        RECT 162.355 -168.805 162.685 -168.475 ;
        RECT 162.355 -170.165 162.685 -169.835 ;
        RECT 162.355 -171.525 162.685 -171.195 ;
        RECT 162.355 -172.885 162.685 -172.555 ;
        RECT 162.355 -174.245 162.685 -173.915 ;
        RECT 162.355 -175.605 162.685 -175.275 ;
        RECT 162.355 -176.965 162.685 -176.635 ;
        RECT 162.355 -178.325 162.685 -177.995 ;
        RECT 162.355 -179.685 162.685 -179.355 ;
        RECT 162.355 -181.93 162.685 -180.8 ;
        RECT 162.36 -182.045 162.68 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 241.32 164.045 242.45 ;
        RECT 163.715 239.195 164.045 239.525 ;
        RECT 163.715 237.835 164.045 238.165 ;
        RECT 163.72 237.16 164.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 -1.525 164.045 -1.195 ;
        RECT 163.715 -2.885 164.045 -2.555 ;
        RECT 163.72 -3.56 164.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 163.715 -95.365 164.045 -95.035 ;
        RECT 163.715 -96.725 164.045 -96.395 ;
        RECT 163.715 -98.085 164.045 -97.755 ;
        RECT 163.715 -99.445 164.045 -99.115 ;
        RECT 163.715 -100.805 164.045 -100.475 ;
        RECT 163.715 -102.165 164.045 -101.835 ;
        RECT 163.715 -103.525 164.045 -103.195 ;
        RECT 163.715 -104.885 164.045 -104.555 ;
        RECT 163.715 -106.245 164.045 -105.915 ;
        RECT 163.715 -107.605 164.045 -107.275 ;
        RECT 163.715 -108.965 164.045 -108.635 ;
        RECT 163.715 -110.325 164.045 -109.995 ;
        RECT 163.715 -111.685 164.045 -111.355 ;
        RECT 163.715 -113.045 164.045 -112.715 ;
        RECT 163.715 -114.405 164.045 -114.075 ;
        RECT 163.715 -115.765 164.045 -115.435 ;
        RECT 163.715 -117.125 164.045 -116.795 ;
        RECT 163.715 -118.485 164.045 -118.155 ;
        RECT 163.715 -119.845 164.045 -119.515 ;
        RECT 163.715 -121.205 164.045 -120.875 ;
        RECT 163.715 -122.565 164.045 -122.235 ;
        RECT 163.715 -123.925 164.045 -123.595 ;
        RECT 163.715 -125.285 164.045 -124.955 ;
        RECT 163.715 -126.645 164.045 -126.315 ;
        RECT 163.715 -128.005 164.045 -127.675 ;
        RECT 163.715 -129.365 164.045 -129.035 ;
        RECT 163.715 -130.725 164.045 -130.395 ;
        RECT 163.715 -132.085 164.045 -131.755 ;
        RECT 163.715 -133.445 164.045 -133.115 ;
        RECT 163.715 -134.805 164.045 -134.475 ;
        RECT 163.715 -136.165 164.045 -135.835 ;
        RECT 163.715 -137.525 164.045 -137.195 ;
        RECT 163.715 -138.885 164.045 -138.555 ;
        RECT 163.715 -140.245 164.045 -139.915 ;
        RECT 163.715 -141.605 164.045 -141.275 ;
        RECT 163.715 -142.965 164.045 -142.635 ;
        RECT 163.715 -144.325 164.045 -143.995 ;
        RECT 163.715 -145.685 164.045 -145.355 ;
        RECT 163.715 -147.045 164.045 -146.715 ;
        RECT 163.715 -148.405 164.045 -148.075 ;
        RECT 163.715 -149.765 164.045 -149.435 ;
        RECT 163.715 -151.125 164.045 -150.795 ;
        RECT 163.715 -152.485 164.045 -152.155 ;
        RECT 163.715 -153.845 164.045 -153.515 ;
        RECT 163.715 -155.205 164.045 -154.875 ;
        RECT 163.715 -156.565 164.045 -156.235 ;
        RECT 163.715 -157.925 164.045 -157.595 ;
        RECT 163.715 -159.285 164.045 -158.955 ;
        RECT 163.715 -160.645 164.045 -160.315 ;
        RECT 163.715 -162.005 164.045 -161.675 ;
        RECT 163.715 -163.365 164.045 -163.035 ;
        RECT 163.715 -164.725 164.045 -164.395 ;
        RECT 163.715 -166.085 164.045 -165.755 ;
        RECT 163.715 -167.445 164.045 -167.115 ;
        RECT 163.715 -168.805 164.045 -168.475 ;
        RECT 163.715 -170.165 164.045 -169.835 ;
        RECT 163.715 -171.525 164.045 -171.195 ;
        RECT 163.715 -172.885 164.045 -172.555 ;
        RECT 163.715 -174.245 164.045 -173.915 ;
        RECT 163.715 -175.605 164.045 -175.275 ;
        RECT 163.715 -176.965 164.045 -176.635 ;
        RECT 163.715 -178.325 164.045 -177.995 ;
        RECT 163.715 -179.685 164.045 -179.355 ;
        RECT 163.715 -181.93 164.045 -180.8 ;
        RECT 163.72 -182.045 164.04 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 241.32 165.405 242.45 ;
        RECT 165.075 239.195 165.405 239.525 ;
        RECT 165.075 237.835 165.405 238.165 ;
        RECT 165.08 237.16 165.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 -1.525 165.405 -1.195 ;
        RECT 165.075 -2.885 165.405 -2.555 ;
        RECT 165.08 -3.56 165.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 165.075 -122.565 165.405 -122.235 ;
        RECT 165.075 -123.925 165.405 -123.595 ;
        RECT 165.075 -125.285 165.405 -124.955 ;
        RECT 165.075 -126.645 165.405 -126.315 ;
        RECT 165.075 -128.005 165.405 -127.675 ;
        RECT 165.075 -129.365 165.405 -129.035 ;
        RECT 165.075 -130.725 165.405 -130.395 ;
        RECT 165.075 -132.085 165.405 -131.755 ;
        RECT 165.075 -133.445 165.405 -133.115 ;
        RECT 165.075 -134.805 165.405 -134.475 ;
        RECT 165.075 -136.165 165.405 -135.835 ;
        RECT 165.075 -137.525 165.405 -137.195 ;
        RECT 165.075 -138.885 165.405 -138.555 ;
        RECT 165.075 -140.245 165.405 -139.915 ;
        RECT 165.075 -141.605 165.405 -141.275 ;
        RECT 165.075 -142.965 165.405 -142.635 ;
        RECT 165.075 -144.325 165.405 -143.995 ;
        RECT 165.075 -145.685 165.405 -145.355 ;
        RECT 165.075 -147.045 165.405 -146.715 ;
        RECT 165.075 -148.405 165.405 -148.075 ;
        RECT 165.075 -149.765 165.405 -149.435 ;
        RECT 165.075 -151.125 165.405 -150.795 ;
        RECT 165.075 -152.485 165.405 -152.155 ;
        RECT 165.075 -153.845 165.405 -153.515 ;
        RECT 165.075 -155.205 165.405 -154.875 ;
        RECT 165.075 -156.565 165.405 -156.235 ;
        RECT 165.075 -157.925 165.405 -157.595 ;
        RECT 165.075 -159.285 165.405 -158.955 ;
        RECT 165.075 -160.645 165.405 -160.315 ;
        RECT 165.075 -162.005 165.405 -161.675 ;
        RECT 165.075 -163.365 165.405 -163.035 ;
        RECT 165.075 -164.725 165.405 -164.395 ;
        RECT 165.075 -166.085 165.405 -165.755 ;
        RECT 165.075 -167.445 165.405 -167.115 ;
        RECT 165.075 -168.805 165.405 -168.475 ;
        RECT 165.075 -170.165 165.405 -169.835 ;
        RECT 165.075 -171.525 165.405 -171.195 ;
        RECT 165.075 -172.885 165.405 -172.555 ;
        RECT 165.075 -174.245 165.405 -173.915 ;
        RECT 165.075 -175.605 165.405 -175.275 ;
        RECT 165.075 -176.965 165.405 -176.635 ;
        RECT 165.075 -178.325 165.405 -177.995 ;
        RECT 165.075 -179.685 165.405 -179.355 ;
        RECT 165.075 -181.93 165.405 -180.8 ;
        RECT 165.08 -182.045 165.4 -95.035 ;
        RECT 165.075 -95.365 165.405 -95.035 ;
        RECT 165.075 -96.725 165.405 -96.395 ;
        RECT 165.075 -98.085 165.405 -97.755 ;
        RECT 165.075 -99.445 165.405 -99.115 ;
        RECT 165.075 -100.805 165.405 -100.475 ;
        RECT 165.075 -102.165 165.405 -101.835 ;
        RECT 165.075 -103.525 165.405 -103.195 ;
        RECT 165.075 -104.885 165.405 -104.555 ;
        RECT 165.075 -106.245 165.405 -105.915 ;
        RECT 165.075 -107.605 165.405 -107.275 ;
        RECT 165.075 -108.965 165.405 -108.635 ;
        RECT 165.075 -110.325 165.405 -109.995 ;
        RECT 165.075 -111.685 165.405 -111.355 ;
        RECT 165.075 -113.045 165.405 -112.715 ;
        RECT 165.075 -114.405 165.405 -114.075 ;
        RECT 165.075 -115.765 165.405 -115.435 ;
        RECT 165.075 -117.125 165.405 -116.795 ;
        RECT 165.075 -118.485 165.405 -118.155 ;
        RECT 165.075 -119.845 165.405 -119.515 ;
        RECT 165.075 -121.205 165.405 -120.875 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 241.32 119.165 242.45 ;
        RECT 118.835 239.195 119.165 239.525 ;
        RECT 118.835 237.835 119.165 238.165 ;
        RECT 118.84 237.16 119.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 -1.525 119.165 -1.195 ;
        RECT 118.835 -2.885 119.165 -2.555 ;
        RECT 118.84 -3.56 119.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 118.835 -95.365 119.165 -95.035 ;
        RECT 118.835 -96.725 119.165 -96.395 ;
        RECT 118.835 -98.085 119.165 -97.755 ;
        RECT 118.835 -99.445 119.165 -99.115 ;
        RECT 118.835 -100.805 119.165 -100.475 ;
        RECT 118.835 -102.165 119.165 -101.835 ;
        RECT 118.835 -103.525 119.165 -103.195 ;
        RECT 118.835 -104.885 119.165 -104.555 ;
        RECT 118.835 -106.245 119.165 -105.915 ;
        RECT 118.835 -107.605 119.165 -107.275 ;
        RECT 118.835 -108.965 119.165 -108.635 ;
        RECT 118.835 -110.325 119.165 -109.995 ;
        RECT 118.835 -111.685 119.165 -111.355 ;
        RECT 118.835 -113.045 119.165 -112.715 ;
        RECT 118.835 -114.405 119.165 -114.075 ;
        RECT 118.835 -115.765 119.165 -115.435 ;
        RECT 118.835 -117.125 119.165 -116.795 ;
        RECT 118.835 -118.485 119.165 -118.155 ;
        RECT 118.835 -119.845 119.165 -119.515 ;
        RECT 118.835 -121.205 119.165 -120.875 ;
        RECT 118.835 -122.565 119.165 -122.235 ;
        RECT 118.835 -123.925 119.165 -123.595 ;
        RECT 118.835 -125.285 119.165 -124.955 ;
        RECT 118.835 -126.645 119.165 -126.315 ;
        RECT 118.835 -128.005 119.165 -127.675 ;
        RECT 118.835 -129.365 119.165 -129.035 ;
        RECT 118.835 -130.725 119.165 -130.395 ;
        RECT 118.835 -132.085 119.165 -131.755 ;
        RECT 118.835 -133.445 119.165 -133.115 ;
        RECT 118.835 -134.805 119.165 -134.475 ;
        RECT 118.835 -136.165 119.165 -135.835 ;
        RECT 118.835 -137.525 119.165 -137.195 ;
        RECT 118.835 -138.885 119.165 -138.555 ;
        RECT 118.835 -140.245 119.165 -139.915 ;
        RECT 118.835 -141.605 119.165 -141.275 ;
        RECT 118.835 -142.965 119.165 -142.635 ;
        RECT 118.835 -144.325 119.165 -143.995 ;
        RECT 118.835 -145.685 119.165 -145.355 ;
        RECT 118.835 -147.045 119.165 -146.715 ;
        RECT 118.835 -148.405 119.165 -148.075 ;
        RECT 118.835 -149.765 119.165 -149.435 ;
        RECT 118.835 -151.125 119.165 -150.795 ;
        RECT 118.835 -152.485 119.165 -152.155 ;
        RECT 118.835 -153.845 119.165 -153.515 ;
        RECT 118.835 -155.205 119.165 -154.875 ;
        RECT 118.835 -156.565 119.165 -156.235 ;
        RECT 118.835 -157.925 119.165 -157.595 ;
        RECT 118.835 -159.285 119.165 -158.955 ;
        RECT 118.835 -160.645 119.165 -160.315 ;
        RECT 118.835 -162.005 119.165 -161.675 ;
        RECT 118.835 -163.365 119.165 -163.035 ;
        RECT 118.835 -164.725 119.165 -164.395 ;
        RECT 118.835 -166.085 119.165 -165.755 ;
        RECT 118.835 -167.445 119.165 -167.115 ;
        RECT 118.835 -168.805 119.165 -168.475 ;
        RECT 118.835 -170.165 119.165 -169.835 ;
        RECT 118.835 -171.525 119.165 -171.195 ;
        RECT 118.835 -172.885 119.165 -172.555 ;
        RECT 118.835 -174.245 119.165 -173.915 ;
        RECT 118.835 -175.605 119.165 -175.275 ;
        RECT 118.835 -176.965 119.165 -176.635 ;
        RECT 118.835 -178.325 119.165 -177.995 ;
        RECT 118.835 -179.685 119.165 -179.355 ;
        RECT 118.835 -181.93 119.165 -180.8 ;
        RECT 118.84 -182.045 119.16 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 241.32 120.525 242.45 ;
        RECT 120.195 239.195 120.525 239.525 ;
        RECT 120.195 237.835 120.525 238.165 ;
        RECT 120.2 237.16 120.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 -1.525 120.525 -1.195 ;
        RECT 120.195 -2.885 120.525 -2.555 ;
        RECT 120.2 -3.56 120.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 120.195 -95.365 120.525 -95.035 ;
        RECT 120.195 -96.725 120.525 -96.395 ;
        RECT 120.195 -98.085 120.525 -97.755 ;
        RECT 120.195 -99.445 120.525 -99.115 ;
        RECT 120.195 -100.805 120.525 -100.475 ;
        RECT 120.195 -102.165 120.525 -101.835 ;
        RECT 120.195 -103.525 120.525 -103.195 ;
        RECT 120.195 -104.885 120.525 -104.555 ;
        RECT 120.195 -106.245 120.525 -105.915 ;
        RECT 120.195 -107.605 120.525 -107.275 ;
        RECT 120.195 -108.965 120.525 -108.635 ;
        RECT 120.195 -110.325 120.525 -109.995 ;
        RECT 120.195 -111.685 120.525 -111.355 ;
        RECT 120.195 -113.045 120.525 -112.715 ;
        RECT 120.195 -114.405 120.525 -114.075 ;
        RECT 120.195 -115.765 120.525 -115.435 ;
        RECT 120.195 -117.125 120.525 -116.795 ;
        RECT 120.195 -118.485 120.525 -118.155 ;
        RECT 120.195 -119.845 120.525 -119.515 ;
        RECT 120.195 -121.205 120.525 -120.875 ;
        RECT 120.195 -122.565 120.525 -122.235 ;
        RECT 120.195 -123.925 120.525 -123.595 ;
        RECT 120.195 -125.285 120.525 -124.955 ;
        RECT 120.195 -126.645 120.525 -126.315 ;
        RECT 120.195 -128.005 120.525 -127.675 ;
        RECT 120.195 -129.365 120.525 -129.035 ;
        RECT 120.195 -130.725 120.525 -130.395 ;
        RECT 120.195 -132.085 120.525 -131.755 ;
        RECT 120.195 -133.445 120.525 -133.115 ;
        RECT 120.195 -134.805 120.525 -134.475 ;
        RECT 120.195 -136.165 120.525 -135.835 ;
        RECT 120.195 -137.525 120.525 -137.195 ;
        RECT 120.195 -138.885 120.525 -138.555 ;
        RECT 120.195 -140.245 120.525 -139.915 ;
        RECT 120.195 -141.605 120.525 -141.275 ;
        RECT 120.195 -142.965 120.525 -142.635 ;
        RECT 120.195 -144.325 120.525 -143.995 ;
        RECT 120.195 -145.685 120.525 -145.355 ;
        RECT 120.195 -147.045 120.525 -146.715 ;
        RECT 120.195 -148.405 120.525 -148.075 ;
        RECT 120.195 -149.765 120.525 -149.435 ;
        RECT 120.195 -151.125 120.525 -150.795 ;
        RECT 120.195 -152.485 120.525 -152.155 ;
        RECT 120.195 -153.845 120.525 -153.515 ;
        RECT 120.195 -155.205 120.525 -154.875 ;
        RECT 120.195 -156.565 120.525 -156.235 ;
        RECT 120.195 -157.925 120.525 -157.595 ;
        RECT 120.195 -159.285 120.525 -158.955 ;
        RECT 120.195 -160.645 120.525 -160.315 ;
        RECT 120.195 -162.005 120.525 -161.675 ;
        RECT 120.195 -163.365 120.525 -163.035 ;
        RECT 120.195 -164.725 120.525 -164.395 ;
        RECT 120.195 -166.085 120.525 -165.755 ;
        RECT 120.195 -167.445 120.525 -167.115 ;
        RECT 120.195 -168.805 120.525 -168.475 ;
        RECT 120.195 -170.165 120.525 -169.835 ;
        RECT 120.195 -171.525 120.525 -171.195 ;
        RECT 120.195 -172.885 120.525 -172.555 ;
        RECT 120.195 -174.245 120.525 -173.915 ;
        RECT 120.195 -175.605 120.525 -175.275 ;
        RECT 120.195 -176.965 120.525 -176.635 ;
        RECT 120.195 -178.325 120.525 -177.995 ;
        RECT 120.195 -179.685 120.525 -179.355 ;
        RECT 120.195 -181.93 120.525 -180.8 ;
        RECT 120.2 -182.045 120.52 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 241.32 121.885 242.45 ;
        RECT 121.555 239.195 121.885 239.525 ;
        RECT 121.555 237.835 121.885 238.165 ;
        RECT 121.56 237.16 121.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 -1.525 121.885 -1.195 ;
        RECT 121.555 -2.885 121.885 -2.555 ;
        RECT 121.56 -3.56 121.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 121.555 -95.365 121.885 -95.035 ;
        RECT 121.555 -96.725 121.885 -96.395 ;
        RECT 121.555 -98.085 121.885 -97.755 ;
        RECT 121.555 -99.445 121.885 -99.115 ;
        RECT 121.555 -100.805 121.885 -100.475 ;
        RECT 121.555 -102.165 121.885 -101.835 ;
        RECT 121.555 -103.525 121.885 -103.195 ;
        RECT 121.555 -104.885 121.885 -104.555 ;
        RECT 121.555 -106.245 121.885 -105.915 ;
        RECT 121.555 -107.605 121.885 -107.275 ;
        RECT 121.555 -108.965 121.885 -108.635 ;
        RECT 121.555 -110.325 121.885 -109.995 ;
        RECT 121.555 -111.685 121.885 -111.355 ;
        RECT 121.555 -113.045 121.885 -112.715 ;
        RECT 121.555 -114.405 121.885 -114.075 ;
        RECT 121.555 -115.765 121.885 -115.435 ;
        RECT 121.555 -117.125 121.885 -116.795 ;
        RECT 121.555 -118.485 121.885 -118.155 ;
        RECT 121.555 -119.845 121.885 -119.515 ;
        RECT 121.555 -121.205 121.885 -120.875 ;
        RECT 121.555 -122.565 121.885 -122.235 ;
        RECT 121.555 -123.925 121.885 -123.595 ;
        RECT 121.555 -125.285 121.885 -124.955 ;
        RECT 121.555 -126.645 121.885 -126.315 ;
        RECT 121.555 -128.005 121.885 -127.675 ;
        RECT 121.555 -129.365 121.885 -129.035 ;
        RECT 121.555 -130.725 121.885 -130.395 ;
        RECT 121.555 -132.085 121.885 -131.755 ;
        RECT 121.555 -133.445 121.885 -133.115 ;
        RECT 121.555 -134.805 121.885 -134.475 ;
        RECT 121.555 -136.165 121.885 -135.835 ;
        RECT 121.555 -137.525 121.885 -137.195 ;
        RECT 121.555 -138.885 121.885 -138.555 ;
        RECT 121.555 -140.245 121.885 -139.915 ;
        RECT 121.555 -141.605 121.885 -141.275 ;
        RECT 121.555 -142.965 121.885 -142.635 ;
        RECT 121.555 -144.325 121.885 -143.995 ;
        RECT 121.555 -145.685 121.885 -145.355 ;
        RECT 121.555 -147.045 121.885 -146.715 ;
        RECT 121.555 -148.405 121.885 -148.075 ;
        RECT 121.555 -149.765 121.885 -149.435 ;
        RECT 121.555 -151.125 121.885 -150.795 ;
        RECT 121.555 -152.485 121.885 -152.155 ;
        RECT 121.555 -153.845 121.885 -153.515 ;
        RECT 121.555 -155.205 121.885 -154.875 ;
        RECT 121.555 -156.565 121.885 -156.235 ;
        RECT 121.555 -157.925 121.885 -157.595 ;
        RECT 121.555 -159.285 121.885 -158.955 ;
        RECT 121.555 -160.645 121.885 -160.315 ;
        RECT 121.555 -162.005 121.885 -161.675 ;
        RECT 121.555 -163.365 121.885 -163.035 ;
        RECT 121.555 -164.725 121.885 -164.395 ;
        RECT 121.555 -166.085 121.885 -165.755 ;
        RECT 121.555 -167.445 121.885 -167.115 ;
        RECT 121.555 -168.805 121.885 -168.475 ;
        RECT 121.555 -170.165 121.885 -169.835 ;
        RECT 121.555 -171.525 121.885 -171.195 ;
        RECT 121.555 -172.885 121.885 -172.555 ;
        RECT 121.555 -174.245 121.885 -173.915 ;
        RECT 121.555 -175.605 121.885 -175.275 ;
        RECT 121.555 -176.965 121.885 -176.635 ;
        RECT 121.555 -178.325 121.885 -177.995 ;
        RECT 121.555 -179.685 121.885 -179.355 ;
        RECT 121.555 -181.93 121.885 -180.8 ;
        RECT 121.56 -182.045 121.88 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 241.32 123.245 242.45 ;
        RECT 122.915 239.195 123.245 239.525 ;
        RECT 122.915 237.835 123.245 238.165 ;
        RECT 122.92 237.16 123.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.915 -99.445 123.245 -99.115 ;
        RECT 122.915 -100.805 123.245 -100.475 ;
        RECT 122.915 -102.165 123.245 -101.835 ;
        RECT 122.915 -103.525 123.245 -103.195 ;
        RECT 122.915 -104.885 123.245 -104.555 ;
        RECT 122.915 -106.245 123.245 -105.915 ;
        RECT 122.915 -107.605 123.245 -107.275 ;
        RECT 122.915 -108.965 123.245 -108.635 ;
        RECT 122.915 -110.325 123.245 -109.995 ;
        RECT 122.915 -111.685 123.245 -111.355 ;
        RECT 122.915 -113.045 123.245 -112.715 ;
        RECT 122.915 -114.405 123.245 -114.075 ;
        RECT 122.915 -115.765 123.245 -115.435 ;
        RECT 122.915 -117.125 123.245 -116.795 ;
        RECT 122.915 -118.485 123.245 -118.155 ;
        RECT 122.915 -119.845 123.245 -119.515 ;
        RECT 122.915 -121.205 123.245 -120.875 ;
        RECT 122.915 -122.565 123.245 -122.235 ;
        RECT 122.915 -123.925 123.245 -123.595 ;
        RECT 122.915 -125.285 123.245 -124.955 ;
        RECT 122.915 -126.645 123.245 -126.315 ;
        RECT 122.915 -128.005 123.245 -127.675 ;
        RECT 122.915 -129.365 123.245 -129.035 ;
        RECT 122.915 -130.725 123.245 -130.395 ;
        RECT 122.915 -132.085 123.245 -131.755 ;
        RECT 122.915 -133.445 123.245 -133.115 ;
        RECT 122.915 -134.805 123.245 -134.475 ;
        RECT 122.915 -136.165 123.245 -135.835 ;
        RECT 122.915 -137.525 123.245 -137.195 ;
        RECT 122.915 -138.885 123.245 -138.555 ;
        RECT 122.915 -140.245 123.245 -139.915 ;
        RECT 122.915 -141.605 123.245 -141.275 ;
        RECT 122.915 -142.965 123.245 -142.635 ;
        RECT 122.915 -144.325 123.245 -143.995 ;
        RECT 122.915 -145.685 123.245 -145.355 ;
        RECT 122.915 -147.045 123.245 -146.715 ;
        RECT 122.915 -148.405 123.245 -148.075 ;
        RECT 122.915 -149.765 123.245 -149.435 ;
        RECT 122.915 -151.125 123.245 -150.795 ;
        RECT 122.915 -152.485 123.245 -152.155 ;
        RECT 122.915 -153.845 123.245 -153.515 ;
        RECT 122.915 -155.205 123.245 -154.875 ;
        RECT 122.915 -156.565 123.245 -156.235 ;
        RECT 122.915 -157.925 123.245 -157.595 ;
        RECT 122.915 -159.285 123.245 -158.955 ;
        RECT 122.915 -160.645 123.245 -160.315 ;
        RECT 122.915 -162.005 123.245 -161.675 ;
        RECT 122.915 -163.365 123.245 -163.035 ;
        RECT 122.915 -164.725 123.245 -164.395 ;
        RECT 122.915 -166.085 123.245 -165.755 ;
        RECT 122.915 -167.445 123.245 -167.115 ;
        RECT 122.915 -168.805 123.245 -168.475 ;
        RECT 122.915 -170.165 123.245 -169.835 ;
        RECT 122.915 -171.525 123.245 -171.195 ;
        RECT 122.915 -172.885 123.245 -172.555 ;
        RECT 122.915 -174.245 123.245 -173.915 ;
        RECT 122.915 -175.605 123.245 -175.275 ;
        RECT 122.915 -176.965 123.245 -176.635 ;
        RECT 122.915 -178.325 123.245 -177.995 ;
        RECT 122.915 -179.685 123.245 -179.355 ;
        RECT 122.915 -181.93 123.245 -180.8 ;
        RECT 122.92 -182.045 123.24 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.21 -98.075 123.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 241.32 124.605 242.45 ;
        RECT 124.275 239.195 124.605 239.525 ;
        RECT 124.275 237.835 124.605 238.165 ;
        RECT 124.28 237.16 124.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 124.275 -1.525 124.605 -1.195 ;
        RECT 124.275 -2.885 124.605 -2.555 ;
        RECT 124.28 -3.56 124.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.635 241.32 125.965 242.45 ;
        RECT 125.635 239.195 125.965 239.525 ;
        RECT 125.635 237.835 125.965 238.165 ;
        RECT 125.64 237.16 125.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.635 -1.525 125.965 -1.195 ;
        RECT 125.635 -2.885 125.965 -2.555 ;
        RECT 125.64 -3.56 125.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 241.32 127.325 242.45 ;
        RECT 126.995 239.195 127.325 239.525 ;
        RECT 126.995 237.835 127.325 238.165 ;
        RECT 127 237.16 127.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 -1.525 127.325 -1.195 ;
        RECT 126.995 -2.885 127.325 -2.555 ;
        RECT 127 -3.56 127.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 126.995 -95.365 127.325 -95.035 ;
        RECT 126.995 -96.725 127.325 -96.395 ;
        RECT 126.995 -98.085 127.325 -97.755 ;
        RECT 126.995 -99.445 127.325 -99.115 ;
        RECT 126.995 -100.805 127.325 -100.475 ;
        RECT 126.995 -102.165 127.325 -101.835 ;
        RECT 126.995 -103.525 127.325 -103.195 ;
        RECT 126.995 -104.885 127.325 -104.555 ;
        RECT 126.995 -106.245 127.325 -105.915 ;
        RECT 126.995 -107.605 127.325 -107.275 ;
        RECT 126.995 -108.965 127.325 -108.635 ;
        RECT 126.995 -110.325 127.325 -109.995 ;
        RECT 126.995 -111.685 127.325 -111.355 ;
        RECT 126.995 -113.045 127.325 -112.715 ;
        RECT 126.995 -114.405 127.325 -114.075 ;
        RECT 126.995 -115.765 127.325 -115.435 ;
        RECT 126.995 -117.125 127.325 -116.795 ;
        RECT 126.995 -118.485 127.325 -118.155 ;
        RECT 126.995 -119.845 127.325 -119.515 ;
        RECT 126.995 -121.205 127.325 -120.875 ;
        RECT 126.995 -122.565 127.325 -122.235 ;
        RECT 126.995 -123.925 127.325 -123.595 ;
        RECT 126.995 -125.285 127.325 -124.955 ;
        RECT 126.995 -126.645 127.325 -126.315 ;
        RECT 126.995 -128.005 127.325 -127.675 ;
        RECT 126.995 -129.365 127.325 -129.035 ;
        RECT 126.995 -130.725 127.325 -130.395 ;
        RECT 126.995 -132.085 127.325 -131.755 ;
        RECT 126.995 -133.445 127.325 -133.115 ;
        RECT 126.995 -134.805 127.325 -134.475 ;
        RECT 126.995 -136.165 127.325 -135.835 ;
        RECT 126.995 -137.525 127.325 -137.195 ;
        RECT 126.995 -138.885 127.325 -138.555 ;
        RECT 126.995 -140.245 127.325 -139.915 ;
        RECT 126.995 -141.605 127.325 -141.275 ;
        RECT 126.995 -142.965 127.325 -142.635 ;
        RECT 126.995 -144.325 127.325 -143.995 ;
        RECT 126.995 -145.685 127.325 -145.355 ;
        RECT 126.995 -147.045 127.325 -146.715 ;
        RECT 126.995 -148.405 127.325 -148.075 ;
        RECT 126.995 -149.765 127.325 -149.435 ;
        RECT 126.995 -151.125 127.325 -150.795 ;
        RECT 126.995 -152.485 127.325 -152.155 ;
        RECT 126.995 -153.845 127.325 -153.515 ;
        RECT 126.995 -155.205 127.325 -154.875 ;
        RECT 126.995 -156.565 127.325 -156.235 ;
        RECT 126.995 -157.925 127.325 -157.595 ;
        RECT 126.995 -159.285 127.325 -158.955 ;
        RECT 126.995 -160.645 127.325 -160.315 ;
        RECT 126.995 -162.005 127.325 -161.675 ;
        RECT 126.995 -163.365 127.325 -163.035 ;
        RECT 126.995 -164.725 127.325 -164.395 ;
        RECT 126.995 -166.085 127.325 -165.755 ;
        RECT 126.995 -167.445 127.325 -167.115 ;
        RECT 126.995 -168.805 127.325 -168.475 ;
        RECT 126.995 -170.165 127.325 -169.835 ;
        RECT 126.995 -171.525 127.325 -171.195 ;
        RECT 126.995 -172.885 127.325 -172.555 ;
        RECT 126.995 -174.245 127.325 -173.915 ;
        RECT 126.995 -175.605 127.325 -175.275 ;
        RECT 126.995 -176.965 127.325 -176.635 ;
        RECT 126.995 -178.325 127.325 -177.995 ;
        RECT 126.995 -179.685 127.325 -179.355 ;
        RECT 126.995 -181.93 127.325 -180.8 ;
        RECT 127 -182.045 127.32 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 241.32 128.685 242.45 ;
        RECT 128.355 239.195 128.685 239.525 ;
        RECT 128.355 237.835 128.685 238.165 ;
        RECT 128.36 237.16 128.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 -1.525 128.685 -1.195 ;
        RECT 128.355 -2.885 128.685 -2.555 ;
        RECT 128.36 -3.56 128.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 128.355 -95.365 128.685 -95.035 ;
        RECT 128.355 -96.725 128.685 -96.395 ;
        RECT 128.355 -98.085 128.685 -97.755 ;
        RECT 128.355 -99.445 128.685 -99.115 ;
        RECT 128.355 -100.805 128.685 -100.475 ;
        RECT 128.355 -102.165 128.685 -101.835 ;
        RECT 128.355 -103.525 128.685 -103.195 ;
        RECT 128.355 -104.885 128.685 -104.555 ;
        RECT 128.355 -106.245 128.685 -105.915 ;
        RECT 128.355 -107.605 128.685 -107.275 ;
        RECT 128.355 -108.965 128.685 -108.635 ;
        RECT 128.355 -110.325 128.685 -109.995 ;
        RECT 128.355 -111.685 128.685 -111.355 ;
        RECT 128.355 -113.045 128.685 -112.715 ;
        RECT 128.355 -114.405 128.685 -114.075 ;
        RECT 128.355 -115.765 128.685 -115.435 ;
        RECT 128.355 -117.125 128.685 -116.795 ;
        RECT 128.355 -118.485 128.685 -118.155 ;
        RECT 128.355 -119.845 128.685 -119.515 ;
        RECT 128.355 -121.205 128.685 -120.875 ;
        RECT 128.355 -122.565 128.685 -122.235 ;
        RECT 128.355 -123.925 128.685 -123.595 ;
        RECT 128.355 -125.285 128.685 -124.955 ;
        RECT 128.355 -126.645 128.685 -126.315 ;
        RECT 128.355 -128.005 128.685 -127.675 ;
        RECT 128.355 -129.365 128.685 -129.035 ;
        RECT 128.355 -130.725 128.685 -130.395 ;
        RECT 128.355 -132.085 128.685 -131.755 ;
        RECT 128.355 -133.445 128.685 -133.115 ;
        RECT 128.355 -134.805 128.685 -134.475 ;
        RECT 128.355 -136.165 128.685 -135.835 ;
        RECT 128.355 -137.525 128.685 -137.195 ;
        RECT 128.355 -138.885 128.685 -138.555 ;
        RECT 128.355 -140.245 128.685 -139.915 ;
        RECT 128.355 -141.605 128.685 -141.275 ;
        RECT 128.355 -142.965 128.685 -142.635 ;
        RECT 128.355 -144.325 128.685 -143.995 ;
        RECT 128.355 -145.685 128.685 -145.355 ;
        RECT 128.355 -147.045 128.685 -146.715 ;
        RECT 128.355 -148.405 128.685 -148.075 ;
        RECT 128.355 -149.765 128.685 -149.435 ;
        RECT 128.355 -151.125 128.685 -150.795 ;
        RECT 128.355 -152.485 128.685 -152.155 ;
        RECT 128.355 -153.845 128.685 -153.515 ;
        RECT 128.355 -155.205 128.685 -154.875 ;
        RECT 128.355 -156.565 128.685 -156.235 ;
        RECT 128.355 -157.925 128.685 -157.595 ;
        RECT 128.355 -159.285 128.685 -158.955 ;
        RECT 128.355 -160.645 128.685 -160.315 ;
        RECT 128.355 -162.005 128.685 -161.675 ;
        RECT 128.355 -163.365 128.685 -163.035 ;
        RECT 128.355 -164.725 128.685 -164.395 ;
        RECT 128.355 -166.085 128.685 -165.755 ;
        RECT 128.355 -167.445 128.685 -167.115 ;
        RECT 128.355 -168.805 128.685 -168.475 ;
        RECT 128.355 -170.165 128.685 -169.835 ;
        RECT 128.355 -171.525 128.685 -171.195 ;
        RECT 128.355 -172.885 128.685 -172.555 ;
        RECT 128.355 -174.245 128.685 -173.915 ;
        RECT 128.355 -175.605 128.685 -175.275 ;
        RECT 128.355 -176.965 128.685 -176.635 ;
        RECT 128.355 -178.325 128.685 -177.995 ;
        RECT 128.355 -179.685 128.685 -179.355 ;
        RECT 128.355 -181.93 128.685 -180.8 ;
        RECT 128.36 -182.045 128.68 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 241.32 130.045 242.45 ;
        RECT 129.715 239.195 130.045 239.525 ;
        RECT 129.715 237.835 130.045 238.165 ;
        RECT 129.72 237.16 130.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 -1.525 130.045 -1.195 ;
        RECT 129.715 -2.885 130.045 -2.555 ;
        RECT 129.72 -3.56 130.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.715 -95.365 130.045 -95.035 ;
        RECT 129.715 -96.725 130.045 -96.395 ;
        RECT 129.715 -98.085 130.045 -97.755 ;
        RECT 129.715 -99.445 130.045 -99.115 ;
        RECT 129.715 -100.805 130.045 -100.475 ;
        RECT 129.715 -102.165 130.045 -101.835 ;
        RECT 129.715 -103.525 130.045 -103.195 ;
        RECT 129.715 -104.885 130.045 -104.555 ;
        RECT 129.715 -106.245 130.045 -105.915 ;
        RECT 129.715 -107.605 130.045 -107.275 ;
        RECT 129.715 -108.965 130.045 -108.635 ;
        RECT 129.715 -110.325 130.045 -109.995 ;
        RECT 129.715 -111.685 130.045 -111.355 ;
        RECT 129.715 -113.045 130.045 -112.715 ;
        RECT 129.715 -114.405 130.045 -114.075 ;
        RECT 129.715 -115.765 130.045 -115.435 ;
        RECT 129.715 -117.125 130.045 -116.795 ;
        RECT 129.715 -118.485 130.045 -118.155 ;
        RECT 129.715 -119.845 130.045 -119.515 ;
        RECT 129.715 -121.205 130.045 -120.875 ;
        RECT 129.715 -122.565 130.045 -122.235 ;
        RECT 129.715 -123.925 130.045 -123.595 ;
        RECT 129.715 -125.285 130.045 -124.955 ;
        RECT 129.715 -126.645 130.045 -126.315 ;
        RECT 129.715 -128.005 130.045 -127.675 ;
        RECT 129.715 -129.365 130.045 -129.035 ;
        RECT 129.715 -130.725 130.045 -130.395 ;
        RECT 129.715 -132.085 130.045 -131.755 ;
        RECT 129.715 -133.445 130.045 -133.115 ;
        RECT 129.715 -134.805 130.045 -134.475 ;
        RECT 129.715 -136.165 130.045 -135.835 ;
        RECT 129.715 -137.525 130.045 -137.195 ;
        RECT 129.715 -138.885 130.045 -138.555 ;
        RECT 129.715 -140.245 130.045 -139.915 ;
        RECT 129.715 -141.605 130.045 -141.275 ;
        RECT 129.715 -142.965 130.045 -142.635 ;
        RECT 129.715 -144.325 130.045 -143.995 ;
        RECT 129.715 -145.685 130.045 -145.355 ;
        RECT 129.715 -147.045 130.045 -146.715 ;
        RECT 129.715 -148.405 130.045 -148.075 ;
        RECT 129.715 -149.765 130.045 -149.435 ;
        RECT 129.715 -151.125 130.045 -150.795 ;
        RECT 129.715 -152.485 130.045 -152.155 ;
        RECT 129.715 -153.845 130.045 -153.515 ;
        RECT 129.715 -155.205 130.045 -154.875 ;
        RECT 129.715 -156.565 130.045 -156.235 ;
        RECT 129.715 -157.925 130.045 -157.595 ;
        RECT 129.715 -159.285 130.045 -158.955 ;
        RECT 129.715 -160.645 130.045 -160.315 ;
        RECT 129.715 -162.005 130.045 -161.675 ;
        RECT 129.715 -163.365 130.045 -163.035 ;
        RECT 129.715 -164.725 130.045 -164.395 ;
        RECT 129.715 -166.085 130.045 -165.755 ;
        RECT 129.715 -167.445 130.045 -167.115 ;
        RECT 129.715 -168.805 130.045 -168.475 ;
        RECT 129.715 -170.165 130.045 -169.835 ;
        RECT 129.715 -171.525 130.045 -171.195 ;
        RECT 129.715 -172.885 130.045 -172.555 ;
        RECT 129.715 -174.245 130.045 -173.915 ;
        RECT 129.715 -175.605 130.045 -175.275 ;
        RECT 129.715 -176.965 130.045 -176.635 ;
        RECT 129.715 -178.325 130.045 -177.995 ;
        RECT 129.715 -179.685 130.045 -179.355 ;
        RECT 129.715 -181.93 130.045 -180.8 ;
        RECT 129.72 -182.045 130.04 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 241.32 131.405 242.45 ;
        RECT 131.075 239.195 131.405 239.525 ;
        RECT 131.075 237.835 131.405 238.165 ;
        RECT 131.08 237.16 131.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 -1.525 131.405 -1.195 ;
        RECT 131.075 -2.885 131.405 -2.555 ;
        RECT 131.08 -3.56 131.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.075 -95.365 131.405 -95.035 ;
        RECT 131.075 -96.725 131.405 -96.395 ;
        RECT 131.075 -98.085 131.405 -97.755 ;
        RECT 131.075 -99.445 131.405 -99.115 ;
        RECT 131.075 -100.805 131.405 -100.475 ;
        RECT 131.075 -102.165 131.405 -101.835 ;
        RECT 131.075 -103.525 131.405 -103.195 ;
        RECT 131.075 -104.885 131.405 -104.555 ;
        RECT 131.075 -106.245 131.405 -105.915 ;
        RECT 131.075 -107.605 131.405 -107.275 ;
        RECT 131.075 -108.965 131.405 -108.635 ;
        RECT 131.075 -110.325 131.405 -109.995 ;
        RECT 131.075 -111.685 131.405 -111.355 ;
        RECT 131.075 -113.045 131.405 -112.715 ;
        RECT 131.075 -114.405 131.405 -114.075 ;
        RECT 131.075 -115.765 131.405 -115.435 ;
        RECT 131.075 -117.125 131.405 -116.795 ;
        RECT 131.075 -118.485 131.405 -118.155 ;
        RECT 131.075 -119.845 131.405 -119.515 ;
        RECT 131.075 -121.205 131.405 -120.875 ;
        RECT 131.075 -122.565 131.405 -122.235 ;
        RECT 131.075 -123.925 131.405 -123.595 ;
        RECT 131.075 -125.285 131.405 -124.955 ;
        RECT 131.075 -126.645 131.405 -126.315 ;
        RECT 131.075 -128.005 131.405 -127.675 ;
        RECT 131.075 -129.365 131.405 -129.035 ;
        RECT 131.075 -130.725 131.405 -130.395 ;
        RECT 131.075 -132.085 131.405 -131.755 ;
        RECT 131.075 -133.445 131.405 -133.115 ;
        RECT 131.075 -134.805 131.405 -134.475 ;
        RECT 131.075 -136.165 131.405 -135.835 ;
        RECT 131.075 -137.525 131.405 -137.195 ;
        RECT 131.075 -138.885 131.405 -138.555 ;
        RECT 131.075 -140.245 131.405 -139.915 ;
        RECT 131.075 -141.605 131.405 -141.275 ;
        RECT 131.075 -142.965 131.405 -142.635 ;
        RECT 131.075 -144.325 131.405 -143.995 ;
        RECT 131.075 -145.685 131.405 -145.355 ;
        RECT 131.075 -147.045 131.405 -146.715 ;
        RECT 131.075 -148.405 131.405 -148.075 ;
        RECT 131.075 -149.765 131.405 -149.435 ;
        RECT 131.075 -151.125 131.405 -150.795 ;
        RECT 131.075 -152.485 131.405 -152.155 ;
        RECT 131.075 -153.845 131.405 -153.515 ;
        RECT 131.075 -155.205 131.405 -154.875 ;
        RECT 131.075 -156.565 131.405 -156.235 ;
        RECT 131.075 -157.925 131.405 -157.595 ;
        RECT 131.075 -159.285 131.405 -158.955 ;
        RECT 131.075 -160.645 131.405 -160.315 ;
        RECT 131.075 -162.005 131.405 -161.675 ;
        RECT 131.075 -163.365 131.405 -163.035 ;
        RECT 131.075 -164.725 131.405 -164.395 ;
        RECT 131.075 -166.085 131.405 -165.755 ;
        RECT 131.075 -167.445 131.405 -167.115 ;
        RECT 131.075 -168.805 131.405 -168.475 ;
        RECT 131.075 -170.165 131.405 -169.835 ;
        RECT 131.075 -171.525 131.405 -171.195 ;
        RECT 131.075 -172.885 131.405 -172.555 ;
        RECT 131.075 -174.245 131.405 -173.915 ;
        RECT 131.075 -175.605 131.405 -175.275 ;
        RECT 131.075 -176.965 131.405 -176.635 ;
        RECT 131.075 -178.325 131.405 -177.995 ;
        RECT 131.075 -179.685 131.405 -179.355 ;
        RECT 131.075 -181.93 131.405 -180.8 ;
        RECT 131.08 -182.045 131.4 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 241.32 132.765 242.45 ;
        RECT 132.435 239.195 132.765 239.525 ;
        RECT 132.435 237.835 132.765 238.165 ;
        RECT 132.44 237.16 132.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 -1.525 132.765 -1.195 ;
        RECT 132.435 -2.885 132.765 -2.555 ;
        RECT 132.44 -3.56 132.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 132.435 -95.365 132.765 -95.035 ;
        RECT 132.435 -96.725 132.765 -96.395 ;
        RECT 132.435 -98.085 132.765 -97.755 ;
        RECT 132.435 -99.445 132.765 -99.115 ;
        RECT 132.435 -100.805 132.765 -100.475 ;
        RECT 132.435 -102.165 132.765 -101.835 ;
        RECT 132.435 -103.525 132.765 -103.195 ;
        RECT 132.435 -104.885 132.765 -104.555 ;
        RECT 132.435 -106.245 132.765 -105.915 ;
        RECT 132.435 -107.605 132.765 -107.275 ;
        RECT 132.435 -108.965 132.765 -108.635 ;
        RECT 132.435 -110.325 132.765 -109.995 ;
        RECT 132.435 -111.685 132.765 -111.355 ;
        RECT 132.435 -113.045 132.765 -112.715 ;
        RECT 132.435 -114.405 132.765 -114.075 ;
        RECT 132.435 -115.765 132.765 -115.435 ;
        RECT 132.435 -117.125 132.765 -116.795 ;
        RECT 132.435 -118.485 132.765 -118.155 ;
        RECT 132.435 -119.845 132.765 -119.515 ;
        RECT 132.435 -121.205 132.765 -120.875 ;
        RECT 132.435 -122.565 132.765 -122.235 ;
        RECT 132.435 -123.925 132.765 -123.595 ;
        RECT 132.435 -125.285 132.765 -124.955 ;
        RECT 132.435 -126.645 132.765 -126.315 ;
        RECT 132.435 -128.005 132.765 -127.675 ;
        RECT 132.435 -129.365 132.765 -129.035 ;
        RECT 132.435 -130.725 132.765 -130.395 ;
        RECT 132.435 -132.085 132.765 -131.755 ;
        RECT 132.435 -133.445 132.765 -133.115 ;
        RECT 132.435 -134.805 132.765 -134.475 ;
        RECT 132.435 -136.165 132.765 -135.835 ;
        RECT 132.435 -137.525 132.765 -137.195 ;
        RECT 132.435 -138.885 132.765 -138.555 ;
        RECT 132.435 -140.245 132.765 -139.915 ;
        RECT 132.435 -141.605 132.765 -141.275 ;
        RECT 132.435 -142.965 132.765 -142.635 ;
        RECT 132.435 -144.325 132.765 -143.995 ;
        RECT 132.435 -145.685 132.765 -145.355 ;
        RECT 132.435 -147.045 132.765 -146.715 ;
        RECT 132.435 -148.405 132.765 -148.075 ;
        RECT 132.435 -149.765 132.765 -149.435 ;
        RECT 132.435 -151.125 132.765 -150.795 ;
        RECT 132.435 -152.485 132.765 -152.155 ;
        RECT 132.435 -153.845 132.765 -153.515 ;
        RECT 132.435 -155.205 132.765 -154.875 ;
        RECT 132.435 -156.565 132.765 -156.235 ;
        RECT 132.435 -157.925 132.765 -157.595 ;
        RECT 132.435 -159.285 132.765 -158.955 ;
        RECT 132.435 -160.645 132.765 -160.315 ;
        RECT 132.435 -162.005 132.765 -161.675 ;
        RECT 132.435 -163.365 132.765 -163.035 ;
        RECT 132.435 -164.725 132.765 -164.395 ;
        RECT 132.435 -166.085 132.765 -165.755 ;
        RECT 132.435 -167.445 132.765 -167.115 ;
        RECT 132.435 -168.805 132.765 -168.475 ;
        RECT 132.435 -170.165 132.765 -169.835 ;
        RECT 132.435 -171.525 132.765 -171.195 ;
        RECT 132.435 -172.885 132.765 -172.555 ;
        RECT 132.435 -174.245 132.765 -173.915 ;
        RECT 132.435 -175.605 132.765 -175.275 ;
        RECT 132.435 -176.965 132.765 -176.635 ;
        RECT 132.435 -178.325 132.765 -177.995 ;
        RECT 132.435 -179.685 132.765 -179.355 ;
        RECT 132.435 -181.93 132.765 -180.8 ;
        RECT 132.44 -182.045 132.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 241.32 134.125 242.45 ;
        RECT 133.795 239.195 134.125 239.525 ;
        RECT 133.795 237.835 134.125 238.165 ;
        RECT 133.8 237.16 134.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.795 -99.445 134.125 -99.115 ;
        RECT 133.795 -100.805 134.125 -100.475 ;
        RECT 133.795 -102.165 134.125 -101.835 ;
        RECT 133.795 -103.525 134.125 -103.195 ;
        RECT 133.795 -104.885 134.125 -104.555 ;
        RECT 133.795 -106.245 134.125 -105.915 ;
        RECT 133.795 -107.605 134.125 -107.275 ;
        RECT 133.795 -108.965 134.125 -108.635 ;
        RECT 133.795 -110.325 134.125 -109.995 ;
        RECT 133.795 -111.685 134.125 -111.355 ;
        RECT 133.795 -113.045 134.125 -112.715 ;
        RECT 133.795 -114.405 134.125 -114.075 ;
        RECT 133.795 -115.765 134.125 -115.435 ;
        RECT 133.795 -117.125 134.125 -116.795 ;
        RECT 133.795 -118.485 134.125 -118.155 ;
        RECT 133.795 -119.845 134.125 -119.515 ;
        RECT 133.795 -121.205 134.125 -120.875 ;
        RECT 133.795 -122.565 134.125 -122.235 ;
        RECT 133.795 -123.925 134.125 -123.595 ;
        RECT 133.795 -125.285 134.125 -124.955 ;
        RECT 133.795 -126.645 134.125 -126.315 ;
        RECT 133.795 -128.005 134.125 -127.675 ;
        RECT 133.795 -129.365 134.125 -129.035 ;
        RECT 133.795 -130.725 134.125 -130.395 ;
        RECT 133.795 -132.085 134.125 -131.755 ;
        RECT 133.795 -133.445 134.125 -133.115 ;
        RECT 133.795 -134.805 134.125 -134.475 ;
        RECT 133.795 -136.165 134.125 -135.835 ;
        RECT 133.795 -137.525 134.125 -137.195 ;
        RECT 133.795 -138.885 134.125 -138.555 ;
        RECT 133.795 -140.245 134.125 -139.915 ;
        RECT 133.795 -141.605 134.125 -141.275 ;
        RECT 133.795 -142.965 134.125 -142.635 ;
        RECT 133.795 -144.325 134.125 -143.995 ;
        RECT 133.795 -145.685 134.125 -145.355 ;
        RECT 133.795 -147.045 134.125 -146.715 ;
        RECT 133.795 -148.405 134.125 -148.075 ;
        RECT 133.795 -149.765 134.125 -149.435 ;
        RECT 133.795 -151.125 134.125 -150.795 ;
        RECT 133.795 -152.485 134.125 -152.155 ;
        RECT 133.795 -153.845 134.125 -153.515 ;
        RECT 133.795 -155.205 134.125 -154.875 ;
        RECT 133.795 -156.565 134.125 -156.235 ;
        RECT 133.795 -157.925 134.125 -157.595 ;
        RECT 133.795 -159.285 134.125 -158.955 ;
        RECT 133.795 -160.645 134.125 -160.315 ;
        RECT 133.795 -162.005 134.125 -161.675 ;
        RECT 133.795 -163.365 134.125 -163.035 ;
        RECT 133.795 -164.725 134.125 -164.395 ;
        RECT 133.795 -166.085 134.125 -165.755 ;
        RECT 133.795 -167.445 134.125 -167.115 ;
        RECT 133.795 -168.805 134.125 -168.475 ;
        RECT 133.795 -170.165 134.125 -169.835 ;
        RECT 133.795 -171.525 134.125 -171.195 ;
        RECT 133.795 -172.885 134.125 -172.555 ;
        RECT 133.795 -174.245 134.125 -173.915 ;
        RECT 133.795 -175.605 134.125 -175.275 ;
        RECT 133.795 -176.965 134.125 -176.635 ;
        RECT 133.795 -178.325 134.125 -177.995 ;
        RECT 133.795 -179.685 134.125 -179.355 ;
        RECT 133.795 -181.93 134.125 -180.8 ;
        RECT 133.8 -182.045 134.12 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 134.11 -98.075 134.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 241.32 135.485 242.45 ;
        RECT 135.155 239.195 135.485 239.525 ;
        RECT 135.155 237.835 135.485 238.165 ;
        RECT 135.16 237.16 135.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 135.155 -1.525 135.485 -1.195 ;
        RECT 135.155 -2.885 135.485 -2.555 ;
        RECT 135.16 -3.56 135.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 241.32 136.845 242.45 ;
        RECT 136.515 239.195 136.845 239.525 ;
        RECT 136.515 237.835 136.845 238.165 ;
        RECT 136.52 237.16 136.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 136.515 -1.525 136.845 -1.195 ;
        RECT 136.515 -2.885 136.845 -2.555 ;
        RECT 136.52 -3.56 136.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.875 241.32 138.205 242.45 ;
        RECT 137.875 239.195 138.205 239.525 ;
        RECT 137.875 237.835 138.205 238.165 ;
        RECT 137.88 237.16 138.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.875 -1.525 138.205 -1.195 ;
        RECT 137.875 -2.885 138.205 -2.555 ;
        RECT 137.88 -3.56 138.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 137.875 -95.365 138.205 -95.035 ;
        RECT 137.875 -96.725 138.205 -96.395 ;
        RECT 137.875 -98.085 138.205 -97.755 ;
        RECT 137.875 -99.445 138.205 -99.115 ;
        RECT 137.875 -100.805 138.205 -100.475 ;
        RECT 137.875 -102.165 138.205 -101.835 ;
        RECT 137.875 -103.525 138.205 -103.195 ;
        RECT 137.875 -104.885 138.205 -104.555 ;
        RECT 137.875 -106.245 138.205 -105.915 ;
        RECT 137.875 -107.605 138.205 -107.275 ;
        RECT 137.875 -108.965 138.205 -108.635 ;
        RECT 137.875 -110.325 138.205 -109.995 ;
        RECT 137.875 -111.685 138.205 -111.355 ;
        RECT 137.875 -113.045 138.205 -112.715 ;
        RECT 137.875 -114.405 138.205 -114.075 ;
        RECT 137.875 -115.765 138.205 -115.435 ;
        RECT 137.875 -117.125 138.205 -116.795 ;
        RECT 137.875 -118.485 138.205 -118.155 ;
        RECT 137.875 -119.845 138.205 -119.515 ;
        RECT 137.875 -121.205 138.205 -120.875 ;
        RECT 137.875 -122.565 138.205 -122.235 ;
        RECT 137.875 -123.925 138.205 -123.595 ;
        RECT 137.875 -125.285 138.205 -124.955 ;
        RECT 137.875 -126.645 138.205 -126.315 ;
        RECT 137.875 -128.005 138.205 -127.675 ;
        RECT 137.875 -129.365 138.205 -129.035 ;
        RECT 137.875 -130.725 138.205 -130.395 ;
        RECT 137.875 -132.085 138.205 -131.755 ;
        RECT 137.875 -133.445 138.205 -133.115 ;
        RECT 137.875 -134.805 138.205 -134.475 ;
        RECT 137.875 -136.165 138.205 -135.835 ;
        RECT 137.875 -137.525 138.205 -137.195 ;
        RECT 137.875 -138.885 138.205 -138.555 ;
        RECT 137.875 -140.245 138.205 -139.915 ;
        RECT 137.875 -141.605 138.205 -141.275 ;
        RECT 137.875 -142.965 138.205 -142.635 ;
        RECT 137.875 -144.325 138.205 -143.995 ;
        RECT 137.875 -145.685 138.205 -145.355 ;
        RECT 137.875 -147.045 138.205 -146.715 ;
        RECT 137.875 -148.405 138.205 -148.075 ;
        RECT 137.875 -149.765 138.205 -149.435 ;
        RECT 137.875 -151.125 138.205 -150.795 ;
        RECT 137.875 -152.485 138.205 -152.155 ;
        RECT 137.875 -153.845 138.205 -153.515 ;
        RECT 137.875 -155.205 138.205 -154.875 ;
        RECT 137.875 -156.565 138.205 -156.235 ;
        RECT 137.875 -157.925 138.205 -157.595 ;
        RECT 137.875 -159.285 138.205 -158.955 ;
        RECT 137.875 -160.645 138.205 -160.315 ;
        RECT 137.875 -162.005 138.205 -161.675 ;
        RECT 137.875 -163.365 138.205 -163.035 ;
        RECT 137.875 -164.725 138.205 -164.395 ;
        RECT 137.875 -166.085 138.205 -165.755 ;
        RECT 137.875 -167.445 138.205 -167.115 ;
        RECT 137.875 -168.805 138.205 -168.475 ;
        RECT 137.875 -170.165 138.205 -169.835 ;
        RECT 137.875 -171.525 138.205 -171.195 ;
        RECT 137.875 -172.885 138.205 -172.555 ;
        RECT 137.875 -174.245 138.205 -173.915 ;
        RECT 137.875 -175.605 138.205 -175.275 ;
        RECT 137.875 -176.965 138.205 -176.635 ;
        RECT 137.875 -178.325 138.205 -177.995 ;
        RECT 137.875 -179.685 138.205 -179.355 ;
        RECT 137.875 -181.93 138.205 -180.8 ;
        RECT 137.88 -182.045 138.2 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 241.32 139.565 242.45 ;
        RECT 139.235 239.195 139.565 239.525 ;
        RECT 139.235 237.835 139.565 238.165 ;
        RECT 139.24 237.16 139.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 -1.525 139.565 -1.195 ;
        RECT 139.235 -2.885 139.565 -2.555 ;
        RECT 139.24 -3.56 139.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 139.235 -95.365 139.565 -95.035 ;
        RECT 139.235 -96.725 139.565 -96.395 ;
        RECT 139.235 -98.085 139.565 -97.755 ;
        RECT 139.235 -99.445 139.565 -99.115 ;
        RECT 139.235 -100.805 139.565 -100.475 ;
        RECT 139.235 -102.165 139.565 -101.835 ;
        RECT 139.235 -103.525 139.565 -103.195 ;
        RECT 139.235 -104.885 139.565 -104.555 ;
        RECT 139.235 -106.245 139.565 -105.915 ;
        RECT 139.235 -107.605 139.565 -107.275 ;
        RECT 139.235 -108.965 139.565 -108.635 ;
        RECT 139.235 -110.325 139.565 -109.995 ;
        RECT 139.235 -111.685 139.565 -111.355 ;
        RECT 139.235 -113.045 139.565 -112.715 ;
        RECT 139.235 -114.405 139.565 -114.075 ;
        RECT 139.235 -115.765 139.565 -115.435 ;
        RECT 139.235 -117.125 139.565 -116.795 ;
        RECT 139.235 -118.485 139.565 -118.155 ;
        RECT 139.235 -119.845 139.565 -119.515 ;
        RECT 139.235 -121.205 139.565 -120.875 ;
        RECT 139.235 -122.565 139.565 -122.235 ;
        RECT 139.235 -123.925 139.565 -123.595 ;
        RECT 139.235 -125.285 139.565 -124.955 ;
        RECT 139.235 -126.645 139.565 -126.315 ;
        RECT 139.235 -128.005 139.565 -127.675 ;
        RECT 139.235 -129.365 139.565 -129.035 ;
        RECT 139.235 -130.725 139.565 -130.395 ;
        RECT 139.235 -132.085 139.565 -131.755 ;
        RECT 139.235 -133.445 139.565 -133.115 ;
        RECT 139.235 -134.805 139.565 -134.475 ;
        RECT 139.235 -136.165 139.565 -135.835 ;
        RECT 139.235 -137.525 139.565 -137.195 ;
        RECT 139.235 -138.885 139.565 -138.555 ;
        RECT 139.235 -140.245 139.565 -139.915 ;
        RECT 139.235 -141.605 139.565 -141.275 ;
        RECT 139.235 -142.965 139.565 -142.635 ;
        RECT 139.235 -144.325 139.565 -143.995 ;
        RECT 139.235 -145.685 139.565 -145.355 ;
        RECT 139.235 -147.045 139.565 -146.715 ;
        RECT 139.235 -148.405 139.565 -148.075 ;
        RECT 139.235 -149.765 139.565 -149.435 ;
        RECT 139.235 -151.125 139.565 -150.795 ;
        RECT 139.235 -152.485 139.565 -152.155 ;
        RECT 139.235 -153.845 139.565 -153.515 ;
        RECT 139.235 -155.205 139.565 -154.875 ;
        RECT 139.235 -156.565 139.565 -156.235 ;
        RECT 139.235 -157.925 139.565 -157.595 ;
        RECT 139.235 -159.285 139.565 -158.955 ;
        RECT 139.235 -160.645 139.565 -160.315 ;
        RECT 139.235 -162.005 139.565 -161.675 ;
        RECT 139.235 -163.365 139.565 -163.035 ;
        RECT 139.235 -164.725 139.565 -164.395 ;
        RECT 139.235 -166.085 139.565 -165.755 ;
        RECT 139.235 -167.445 139.565 -167.115 ;
        RECT 139.235 -168.805 139.565 -168.475 ;
        RECT 139.235 -170.165 139.565 -169.835 ;
        RECT 139.235 -171.525 139.565 -171.195 ;
        RECT 139.235 -172.885 139.565 -172.555 ;
        RECT 139.235 -174.245 139.565 -173.915 ;
        RECT 139.235 -175.605 139.565 -175.275 ;
        RECT 139.235 -176.965 139.565 -176.635 ;
        RECT 139.235 -178.325 139.565 -177.995 ;
        RECT 139.235 -179.685 139.565 -179.355 ;
        RECT 139.235 -181.93 139.565 -180.8 ;
        RECT 139.24 -182.045 139.56 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 241.32 140.925 242.45 ;
        RECT 140.595 239.195 140.925 239.525 ;
        RECT 140.595 237.835 140.925 238.165 ;
        RECT 140.6 237.16 140.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 -1.525 140.925 -1.195 ;
        RECT 140.595 -2.885 140.925 -2.555 ;
        RECT 140.6 -3.56 140.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 140.595 -95.365 140.925 -95.035 ;
        RECT 140.595 -96.725 140.925 -96.395 ;
        RECT 140.595 -98.085 140.925 -97.755 ;
        RECT 140.595 -99.445 140.925 -99.115 ;
        RECT 140.595 -100.805 140.925 -100.475 ;
        RECT 140.595 -102.165 140.925 -101.835 ;
        RECT 140.595 -103.525 140.925 -103.195 ;
        RECT 140.595 -104.885 140.925 -104.555 ;
        RECT 140.595 -106.245 140.925 -105.915 ;
        RECT 140.595 -107.605 140.925 -107.275 ;
        RECT 140.595 -108.965 140.925 -108.635 ;
        RECT 140.595 -110.325 140.925 -109.995 ;
        RECT 140.595 -111.685 140.925 -111.355 ;
        RECT 140.595 -113.045 140.925 -112.715 ;
        RECT 140.595 -114.405 140.925 -114.075 ;
        RECT 140.595 -115.765 140.925 -115.435 ;
        RECT 140.595 -117.125 140.925 -116.795 ;
        RECT 140.595 -118.485 140.925 -118.155 ;
        RECT 140.595 -119.845 140.925 -119.515 ;
        RECT 140.595 -121.205 140.925 -120.875 ;
        RECT 140.595 -122.565 140.925 -122.235 ;
        RECT 140.595 -123.925 140.925 -123.595 ;
        RECT 140.595 -125.285 140.925 -124.955 ;
        RECT 140.595 -126.645 140.925 -126.315 ;
        RECT 140.595 -128.005 140.925 -127.675 ;
        RECT 140.595 -129.365 140.925 -129.035 ;
        RECT 140.595 -130.725 140.925 -130.395 ;
        RECT 140.595 -132.085 140.925 -131.755 ;
        RECT 140.595 -133.445 140.925 -133.115 ;
        RECT 140.595 -134.805 140.925 -134.475 ;
        RECT 140.595 -136.165 140.925 -135.835 ;
        RECT 140.595 -137.525 140.925 -137.195 ;
        RECT 140.595 -138.885 140.925 -138.555 ;
        RECT 140.595 -140.245 140.925 -139.915 ;
        RECT 140.595 -141.605 140.925 -141.275 ;
        RECT 140.595 -142.965 140.925 -142.635 ;
        RECT 140.595 -144.325 140.925 -143.995 ;
        RECT 140.595 -145.685 140.925 -145.355 ;
        RECT 140.595 -147.045 140.925 -146.715 ;
        RECT 140.595 -148.405 140.925 -148.075 ;
        RECT 140.595 -149.765 140.925 -149.435 ;
        RECT 140.595 -151.125 140.925 -150.795 ;
        RECT 140.595 -152.485 140.925 -152.155 ;
        RECT 140.595 -153.845 140.925 -153.515 ;
        RECT 140.595 -155.205 140.925 -154.875 ;
        RECT 140.595 -156.565 140.925 -156.235 ;
        RECT 140.595 -157.925 140.925 -157.595 ;
        RECT 140.595 -159.285 140.925 -158.955 ;
        RECT 140.595 -160.645 140.925 -160.315 ;
        RECT 140.595 -162.005 140.925 -161.675 ;
        RECT 140.595 -163.365 140.925 -163.035 ;
        RECT 140.595 -164.725 140.925 -164.395 ;
        RECT 140.595 -166.085 140.925 -165.755 ;
        RECT 140.595 -167.445 140.925 -167.115 ;
        RECT 140.595 -168.805 140.925 -168.475 ;
        RECT 140.595 -170.165 140.925 -169.835 ;
        RECT 140.595 -171.525 140.925 -171.195 ;
        RECT 140.595 -172.885 140.925 -172.555 ;
        RECT 140.595 -174.245 140.925 -173.915 ;
        RECT 140.595 -175.605 140.925 -175.275 ;
        RECT 140.595 -176.965 140.925 -176.635 ;
        RECT 140.595 -178.325 140.925 -177.995 ;
        RECT 140.595 -179.685 140.925 -179.355 ;
        RECT 140.595 -181.93 140.925 -180.8 ;
        RECT 140.6 -182.045 140.92 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 241.32 142.285 242.45 ;
        RECT 141.955 239.195 142.285 239.525 ;
        RECT 141.955 237.835 142.285 238.165 ;
        RECT 141.96 237.16 142.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 141.955 -2.885 142.285 -2.555 ;
        RECT 141.96 -3.56 142.28 -0.52 ;
        RECT 141.955 -1.525 142.285 -1.195 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 241.32 91.965 242.45 ;
        RECT 91.635 239.195 91.965 239.525 ;
        RECT 91.635 237.835 91.965 238.165 ;
        RECT 91.64 237.16 91.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 91.635 -1.525 91.965 -1.195 ;
        RECT 91.635 -2.885 91.965 -2.555 ;
        RECT 91.64 -3.56 91.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 241.32 93.325 242.45 ;
        RECT 92.995 239.195 93.325 239.525 ;
        RECT 92.995 237.835 93.325 238.165 ;
        RECT 93 237.16 93.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 92.995 -1.525 93.325 -1.195 ;
        RECT 92.995 -2.885 93.325 -2.555 ;
        RECT 93 -3.56 93.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 241.32 94.685 242.45 ;
        RECT 94.355 239.195 94.685 239.525 ;
        RECT 94.355 237.835 94.685 238.165 ;
        RECT 94.36 237.16 94.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 -1.525 94.685 -1.195 ;
        RECT 94.355 -2.885 94.685 -2.555 ;
        RECT 94.36 -3.56 94.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 94.355 -95.365 94.685 -95.035 ;
        RECT 94.355 -96.725 94.685 -96.395 ;
        RECT 94.355 -98.085 94.685 -97.755 ;
        RECT 94.355 -99.445 94.685 -99.115 ;
        RECT 94.355 -100.805 94.685 -100.475 ;
        RECT 94.355 -102.165 94.685 -101.835 ;
        RECT 94.355 -103.525 94.685 -103.195 ;
        RECT 94.355 -104.885 94.685 -104.555 ;
        RECT 94.355 -106.245 94.685 -105.915 ;
        RECT 94.355 -107.605 94.685 -107.275 ;
        RECT 94.355 -108.965 94.685 -108.635 ;
        RECT 94.355 -110.325 94.685 -109.995 ;
        RECT 94.355 -111.685 94.685 -111.355 ;
        RECT 94.355 -113.045 94.685 -112.715 ;
        RECT 94.355 -114.405 94.685 -114.075 ;
        RECT 94.355 -115.765 94.685 -115.435 ;
        RECT 94.355 -117.125 94.685 -116.795 ;
        RECT 94.355 -118.485 94.685 -118.155 ;
        RECT 94.355 -119.845 94.685 -119.515 ;
        RECT 94.355 -121.205 94.685 -120.875 ;
        RECT 94.355 -122.565 94.685 -122.235 ;
        RECT 94.355 -123.925 94.685 -123.595 ;
        RECT 94.355 -125.285 94.685 -124.955 ;
        RECT 94.355 -126.645 94.685 -126.315 ;
        RECT 94.355 -128.005 94.685 -127.675 ;
        RECT 94.355 -129.365 94.685 -129.035 ;
        RECT 94.355 -130.725 94.685 -130.395 ;
        RECT 94.355 -132.085 94.685 -131.755 ;
        RECT 94.355 -133.445 94.685 -133.115 ;
        RECT 94.355 -134.805 94.685 -134.475 ;
        RECT 94.355 -136.165 94.685 -135.835 ;
        RECT 94.355 -137.525 94.685 -137.195 ;
        RECT 94.355 -138.885 94.685 -138.555 ;
        RECT 94.355 -140.245 94.685 -139.915 ;
        RECT 94.355 -141.605 94.685 -141.275 ;
        RECT 94.355 -142.965 94.685 -142.635 ;
        RECT 94.355 -144.325 94.685 -143.995 ;
        RECT 94.355 -145.685 94.685 -145.355 ;
        RECT 94.355 -147.045 94.685 -146.715 ;
        RECT 94.355 -148.405 94.685 -148.075 ;
        RECT 94.355 -149.765 94.685 -149.435 ;
        RECT 94.355 -151.125 94.685 -150.795 ;
        RECT 94.355 -152.485 94.685 -152.155 ;
        RECT 94.355 -153.845 94.685 -153.515 ;
        RECT 94.355 -155.205 94.685 -154.875 ;
        RECT 94.355 -156.565 94.685 -156.235 ;
        RECT 94.355 -157.925 94.685 -157.595 ;
        RECT 94.355 -159.285 94.685 -158.955 ;
        RECT 94.355 -160.645 94.685 -160.315 ;
        RECT 94.355 -162.005 94.685 -161.675 ;
        RECT 94.355 -163.365 94.685 -163.035 ;
        RECT 94.355 -164.725 94.685 -164.395 ;
        RECT 94.355 -166.085 94.685 -165.755 ;
        RECT 94.355 -167.445 94.685 -167.115 ;
        RECT 94.355 -168.805 94.685 -168.475 ;
        RECT 94.355 -170.165 94.685 -169.835 ;
        RECT 94.355 -171.525 94.685 -171.195 ;
        RECT 94.355 -172.885 94.685 -172.555 ;
        RECT 94.355 -174.245 94.685 -173.915 ;
        RECT 94.355 -175.605 94.685 -175.275 ;
        RECT 94.355 -176.965 94.685 -176.635 ;
        RECT 94.355 -178.325 94.685 -177.995 ;
        RECT 94.355 -179.685 94.685 -179.355 ;
        RECT 94.355 -181.93 94.685 -180.8 ;
        RECT 94.36 -182.045 94.68 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 241.32 96.045 242.45 ;
        RECT 95.715 239.195 96.045 239.525 ;
        RECT 95.715 237.835 96.045 238.165 ;
        RECT 95.72 237.16 96.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 -1.525 96.045 -1.195 ;
        RECT 95.715 -2.885 96.045 -2.555 ;
        RECT 95.72 -3.56 96.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 95.715 -95.365 96.045 -95.035 ;
        RECT 95.715 -96.725 96.045 -96.395 ;
        RECT 95.715 -98.085 96.045 -97.755 ;
        RECT 95.715 -99.445 96.045 -99.115 ;
        RECT 95.715 -100.805 96.045 -100.475 ;
        RECT 95.715 -102.165 96.045 -101.835 ;
        RECT 95.715 -103.525 96.045 -103.195 ;
        RECT 95.715 -104.885 96.045 -104.555 ;
        RECT 95.715 -106.245 96.045 -105.915 ;
        RECT 95.715 -107.605 96.045 -107.275 ;
        RECT 95.715 -108.965 96.045 -108.635 ;
        RECT 95.715 -110.325 96.045 -109.995 ;
        RECT 95.715 -111.685 96.045 -111.355 ;
        RECT 95.715 -113.045 96.045 -112.715 ;
        RECT 95.715 -114.405 96.045 -114.075 ;
        RECT 95.715 -115.765 96.045 -115.435 ;
        RECT 95.715 -117.125 96.045 -116.795 ;
        RECT 95.715 -118.485 96.045 -118.155 ;
        RECT 95.715 -119.845 96.045 -119.515 ;
        RECT 95.715 -121.205 96.045 -120.875 ;
        RECT 95.715 -122.565 96.045 -122.235 ;
        RECT 95.715 -123.925 96.045 -123.595 ;
        RECT 95.715 -125.285 96.045 -124.955 ;
        RECT 95.715 -126.645 96.045 -126.315 ;
        RECT 95.715 -128.005 96.045 -127.675 ;
        RECT 95.715 -129.365 96.045 -129.035 ;
        RECT 95.715 -130.725 96.045 -130.395 ;
        RECT 95.715 -132.085 96.045 -131.755 ;
        RECT 95.715 -133.445 96.045 -133.115 ;
        RECT 95.715 -134.805 96.045 -134.475 ;
        RECT 95.715 -136.165 96.045 -135.835 ;
        RECT 95.715 -137.525 96.045 -137.195 ;
        RECT 95.715 -138.885 96.045 -138.555 ;
        RECT 95.715 -140.245 96.045 -139.915 ;
        RECT 95.715 -141.605 96.045 -141.275 ;
        RECT 95.715 -142.965 96.045 -142.635 ;
        RECT 95.715 -144.325 96.045 -143.995 ;
        RECT 95.715 -145.685 96.045 -145.355 ;
        RECT 95.715 -147.045 96.045 -146.715 ;
        RECT 95.715 -148.405 96.045 -148.075 ;
        RECT 95.715 -149.765 96.045 -149.435 ;
        RECT 95.715 -151.125 96.045 -150.795 ;
        RECT 95.715 -152.485 96.045 -152.155 ;
        RECT 95.715 -153.845 96.045 -153.515 ;
        RECT 95.715 -155.205 96.045 -154.875 ;
        RECT 95.715 -156.565 96.045 -156.235 ;
        RECT 95.715 -157.925 96.045 -157.595 ;
        RECT 95.715 -159.285 96.045 -158.955 ;
        RECT 95.715 -160.645 96.045 -160.315 ;
        RECT 95.715 -162.005 96.045 -161.675 ;
        RECT 95.715 -163.365 96.045 -163.035 ;
        RECT 95.715 -164.725 96.045 -164.395 ;
        RECT 95.715 -166.085 96.045 -165.755 ;
        RECT 95.715 -167.445 96.045 -167.115 ;
        RECT 95.715 -168.805 96.045 -168.475 ;
        RECT 95.715 -170.165 96.045 -169.835 ;
        RECT 95.715 -171.525 96.045 -171.195 ;
        RECT 95.715 -172.885 96.045 -172.555 ;
        RECT 95.715 -174.245 96.045 -173.915 ;
        RECT 95.715 -175.605 96.045 -175.275 ;
        RECT 95.715 -176.965 96.045 -176.635 ;
        RECT 95.715 -178.325 96.045 -177.995 ;
        RECT 95.715 -179.685 96.045 -179.355 ;
        RECT 95.715 -181.93 96.045 -180.8 ;
        RECT 95.72 -182.045 96.04 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 241.32 97.405 242.45 ;
        RECT 97.075 239.195 97.405 239.525 ;
        RECT 97.075 237.835 97.405 238.165 ;
        RECT 97.08 237.16 97.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 -1.525 97.405 -1.195 ;
        RECT 97.075 -2.885 97.405 -2.555 ;
        RECT 97.08 -3.56 97.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 97.075 -95.365 97.405 -95.035 ;
        RECT 97.075 -96.725 97.405 -96.395 ;
        RECT 97.075 -98.085 97.405 -97.755 ;
        RECT 97.075 -99.445 97.405 -99.115 ;
        RECT 97.075 -100.805 97.405 -100.475 ;
        RECT 97.075 -102.165 97.405 -101.835 ;
        RECT 97.075 -103.525 97.405 -103.195 ;
        RECT 97.075 -104.885 97.405 -104.555 ;
        RECT 97.075 -106.245 97.405 -105.915 ;
        RECT 97.075 -107.605 97.405 -107.275 ;
        RECT 97.075 -108.965 97.405 -108.635 ;
        RECT 97.075 -110.325 97.405 -109.995 ;
        RECT 97.075 -111.685 97.405 -111.355 ;
        RECT 97.075 -113.045 97.405 -112.715 ;
        RECT 97.075 -114.405 97.405 -114.075 ;
        RECT 97.075 -115.765 97.405 -115.435 ;
        RECT 97.075 -117.125 97.405 -116.795 ;
        RECT 97.075 -118.485 97.405 -118.155 ;
        RECT 97.075 -119.845 97.405 -119.515 ;
        RECT 97.075 -121.205 97.405 -120.875 ;
        RECT 97.075 -122.565 97.405 -122.235 ;
        RECT 97.075 -123.925 97.405 -123.595 ;
        RECT 97.075 -125.285 97.405 -124.955 ;
        RECT 97.075 -126.645 97.405 -126.315 ;
        RECT 97.075 -128.005 97.405 -127.675 ;
        RECT 97.075 -129.365 97.405 -129.035 ;
        RECT 97.075 -130.725 97.405 -130.395 ;
        RECT 97.075 -132.085 97.405 -131.755 ;
        RECT 97.075 -133.445 97.405 -133.115 ;
        RECT 97.075 -134.805 97.405 -134.475 ;
        RECT 97.075 -136.165 97.405 -135.835 ;
        RECT 97.075 -137.525 97.405 -137.195 ;
        RECT 97.075 -138.885 97.405 -138.555 ;
        RECT 97.075 -140.245 97.405 -139.915 ;
        RECT 97.075 -141.605 97.405 -141.275 ;
        RECT 97.075 -142.965 97.405 -142.635 ;
        RECT 97.075 -144.325 97.405 -143.995 ;
        RECT 97.075 -145.685 97.405 -145.355 ;
        RECT 97.075 -147.045 97.405 -146.715 ;
        RECT 97.075 -148.405 97.405 -148.075 ;
        RECT 97.075 -149.765 97.405 -149.435 ;
        RECT 97.075 -151.125 97.405 -150.795 ;
        RECT 97.075 -152.485 97.405 -152.155 ;
        RECT 97.075 -153.845 97.405 -153.515 ;
        RECT 97.075 -155.205 97.405 -154.875 ;
        RECT 97.075 -156.565 97.405 -156.235 ;
        RECT 97.075 -157.925 97.405 -157.595 ;
        RECT 97.075 -159.285 97.405 -158.955 ;
        RECT 97.075 -160.645 97.405 -160.315 ;
        RECT 97.075 -162.005 97.405 -161.675 ;
        RECT 97.075 -163.365 97.405 -163.035 ;
        RECT 97.075 -164.725 97.405 -164.395 ;
        RECT 97.075 -166.085 97.405 -165.755 ;
        RECT 97.075 -167.445 97.405 -167.115 ;
        RECT 97.075 -168.805 97.405 -168.475 ;
        RECT 97.075 -170.165 97.405 -169.835 ;
        RECT 97.075 -171.525 97.405 -171.195 ;
        RECT 97.075 -172.885 97.405 -172.555 ;
        RECT 97.075 -174.245 97.405 -173.915 ;
        RECT 97.075 -175.605 97.405 -175.275 ;
        RECT 97.075 -176.965 97.405 -176.635 ;
        RECT 97.075 -178.325 97.405 -177.995 ;
        RECT 97.075 -179.685 97.405 -179.355 ;
        RECT 97.075 -181.93 97.405 -180.8 ;
        RECT 97.08 -182.045 97.4 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 241.32 98.765 242.45 ;
        RECT 98.435 239.195 98.765 239.525 ;
        RECT 98.435 237.835 98.765 238.165 ;
        RECT 98.44 237.16 98.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 -1.525 98.765 -1.195 ;
        RECT 98.435 -2.885 98.765 -2.555 ;
        RECT 98.44 -3.56 98.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 98.435 -95.365 98.765 -95.035 ;
        RECT 98.435 -96.725 98.765 -96.395 ;
        RECT 98.435 -98.085 98.765 -97.755 ;
        RECT 98.435 -99.445 98.765 -99.115 ;
        RECT 98.435 -100.805 98.765 -100.475 ;
        RECT 98.435 -102.165 98.765 -101.835 ;
        RECT 98.435 -103.525 98.765 -103.195 ;
        RECT 98.435 -104.885 98.765 -104.555 ;
        RECT 98.435 -106.245 98.765 -105.915 ;
        RECT 98.435 -107.605 98.765 -107.275 ;
        RECT 98.435 -108.965 98.765 -108.635 ;
        RECT 98.435 -110.325 98.765 -109.995 ;
        RECT 98.435 -111.685 98.765 -111.355 ;
        RECT 98.435 -113.045 98.765 -112.715 ;
        RECT 98.435 -114.405 98.765 -114.075 ;
        RECT 98.435 -115.765 98.765 -115.435 ;
        RECT 98.435 -117.125 98.765 -116.795 ;
        RECT 98.435 -118.485 98.765 -118.155 ;
        RECT 98.435 -119.845 98.765 -119.515 ;
        RECT 98.435 -121.205 98.765 -120.875 ;
        RECT 98.435 -122.565 98.765 -122.235 ;
        RECT 98.435 -123.925 98.765 -123.595 ;
        RECT 98.435 -125.285 98.765 -124.955 ;
        RECT 98.435 -126.645 98.765 -126.315 ;
        RECT 98.435 -128.005 98.765 -127.675 ;
        RECT 98.435 -129.365 98.765 -129.035 ;
        RECT 98.435 -130.725 98.765 -130.395 ;
        RECT 98.435 -132.085 98.765 -131.755 ;
        RECT 98.435 -133.445 98.765 -133.115 ;
        RECT 98.435 -134.805 98.765 -134.475 ;
        RECT 98.435 -136.165 98.765 -135.835 ;
        RECT 98.435 -137.525 98.765 -137.195 ;
        RECT 98.435 -138.885 98.765 -138.555 ;
        RECT 98.435 -140.245 98.765 -139.915 ;
        RECT 98.435 -141.605 98.765 -141.275 ;
        RECT 98.435 -142.965 98.765 -142.635 ;
        RECT 98.435 -144.325 98.765 -143.995 ;
        RECT 98.435 -145.685 98.765 -145.355 ;
        RECT 98.435 -147.045 98.765 -146.715 ;
        RECT 98.435 -148.405 98.765 -148.075 ;
        RECT 98.435 -149.765 98.765 -149.435 ;
        RECT 98.435 -151.125 98.765 -150.795 ;
        RECT 98.435 -152.485 98.765 -152.155 ;
        RECT 98.435 -153.845 98.765 -153.515 ;
        RECT 98.435 -155.205 98.765 -154.875 ;
        RECT 98.435 -156.565 98.765 -156.235 ;
        RECT 98.435 -157.925 98.765 -157.595 ;
        RECT 98.435 -159.285 98.765 -158.955 ;
        RECT 98.435 -160.645 98.765 -160.315 ;
        RECT 98.435 -162.005 98.765 -161.675 ;
        RECT 98.435 -163.365 98.765 -163.035 ;
        RECT 98.435 -164.725 98.765 -164.395 ;
        RECT 98.435 -166.085 98.765 -165.755 ;
        RECT 98.435 -167.445 98.765 -167.115 ;
        RECT 98.435 -168.805 98.765 -168.475 ;
        RECT 98.435 -170.165 98.765 -169.835 ;
        RECT 98.435 -171.525 98.765 -171.195 ;
        RECT 98.435 -172.885 98.765 -172.555 ;
        RECT 98.435 -174.245 98.765 -173.915 ;
        RECT 98.435 -175.605 98.765 -175.275 ;
        RECT 98.435 -176.965 98.765 -176.635 ;
        RECT 98.435 -178.325 98.765 -177.995 ;
        RECT 98.435 -179.685 98.765 -179.355 ;
        RECT 98.435 -181.93 98.765 -180.8 ;
        RECT 98.44 -182.045 98.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 241.32 100.125 242.45 ;
        RECT 99.795 239.195 100.125 239.525 ;
        RECT 99.795 237.835 100.125 238.165 ;
        RECT 99.8 237.16 100.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 -1.525 100.125 -1.195 ;
        RECT 99.795 -2.885 100.125 -2.555 ;
        RECT 99.8 -3.56 100.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 99.795 -95.365 100.125 -95.035 ;
        RECT 99.795 -96.725 100.125 -96.395 ;
        RECT 99.795 -98.085 100.125 -97.755 ;
        RECT 99.795 -99.445 100.125 -99.115 ;
        RECT 99.795 -100.805 100.125 -100.475 ;
        RECT 99.795 -102.165 100.125 -101.835 ;
        RECT 99.795 -103.525 100.125 -103.195 ;
        RECT 99.795 -104.885 100.125 -104.555 ;
        RECT 99.795 -106.245 100.125 -105.915 ;
        RECT 99.795 -107.605 100.125 -107.275 ;
        RECT 99.795 -108.965 100.125 -108.635 ;
        RECT 99.795 -110.325 100.125 -109.995 ;
        RECT 99.795 -111.685 100.125 -111.355 ;
        RECT 99.795 -113.045 100.125 -112.715 ;
        RECT 99.795 -114.405 100.125 -114.075 ;
        RECT 99.795 -115.765 100.125 -115.435 ;
        RECT 99.795 -117.125 100.125 -116.795 ;
        RECT 99.795 -118.485 100.125 -118.155 ;
        RECT 99.795 -119.845 100.125 -119.515 ;
        RECT 99.795 -121.205 100.125 -120.875 ;
        RECT 99.795 -122.565 100.125 -122.235 ;
        RECT 99.795 -123.925 100.125 -123.595 ;
        RECT 99.795 -125.285 100.125 -124.955 ;
        RECT 99.795 -126.645 100.125 -126.315 ;
        RECT 99.795 -128.005 100.125 -127.675 ;
        RECT 99.795 -129.365 100.125 -129.035 ;
        RECT 99.795 -130.725 100.125 -130.395 ;
        RECT 99.795 -132.085 100.125 -131.755 ;
        RECT 99.795 -133.445 100.125 -133.115 ;
        RECT 99.795 -134.805 100.125 -134.475 ;
        RECT 99.795 -136.165 100.125 -135.835 ;
        RECT 99.795 -137.525 100.125 -137.195 ;
        RECT 99.795 -138.885 100.125 -138.555 ;
        RECT 99.795 -140.245 100.125 -139.915 ;
        RECT 99.795 -141.605 100.125 -141.275 ;
        RECT 99.795 -142.965 100.125 -142.635 ;
        RECT 99.795 -144.325 100.125 -143.995 ;
        RECT 99.795 -145.685 100.125 -145.355 ;
        RECT 99.795 -147.045 100.125 -146.715 ;
        RECT 99.795 -148.405 100.125 -148.075 ;
        RECT 99.795 -149.765 100.125 -149.435 ;
        RECT 99.795 -151.125 100.125 -150.795 ;
        RECT 99.795 -152.485 100.125 -152.155 ;
        RECT 99.795 -153.845 100.125 -153.515 ;
        RECT 99.795 -155.205 100.125 -154.875 ;
        RECT 99.795 -156.565 100.125 -156.235 ;
        RECT 99.795 -157.925 100.125 -157.595 ;
        RECT 99.795 -159.285 100.125 -158.955 ;
        RECT 99.795 -160.645 100.125 -160.315 ;
        RECT 99.795 -162.005 100.125 -161.675 ;
        RECT 99.795 -163.365 100.125 -163.035 ;
        RECT 99.795 -164.725 100.125 -164.395 ;
        RECT 99.795 -166.085 100.125 -165.755 ;
        RECT 99.795 -167.445 100.125 -167.115 ;
        RECT 99.795 -168.805 100.125 -168.475 ;
        RECT 99.795 -170.165 100.125 -169.835 ;
        RECT 99.795 -171.525 100.125 -171.195 ;
        RECT 99.795 -172.885 100.125 -172.555 ;
        RECT 99.795 -174.245 100.125 -173.915 ;
        RECT 99.795 -175.605 100.125 -175.275 ;
        RECT 99.795 -176.965 100.125 -176.635 ;
        RECT 99.795 -178.325 100.125 -177.995 ;
        RECT 99.795 -179.685 100.125 -179.355 ;
        RECT 99.795 -181.93 100.125 -180.8 ;
        RECT 99.8 -182.045 100.12 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.155 241.32 101.485 242.45 ;
        RECT 101.155 239.195 101.485 239.525 ;
        RECT 101.155 237.835 101.485 238.165 ;
        RECT 101.16 237.16 101.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.155 -99.445 101.485 -99.115 ;
        RECT 101.155 -100.805 101.485 -100.475 ;
        RECT 101.155 -102.165 101.485 -101.835 ;
        RECT 101.155 -103.525 101.485 -103.195 ;
        RECT 101.155 -104.885 101.485 -104.555 ;
        RECT 101.155 -106.245 101.485 -105.915 ;
        RECT 101.155 -107.605 101.485 -107.275 ;
        RECT 101.155 -108.965 101.485 -108.635 ;
        RECT 101.155 -110.325 101.485 -109.995 ;
        RECT 101.155 -111.685 101.485 -111.355 ;
        RECT 101.155 -113.045 101.485 -112.715 ;
        RECT 101.155 -114.405 101.485 -114.075 ;
        RECT 101.155 -115.765 101.485 -115.435 ;
        RECT 101.155 -117.125 101.485 -116.795 ;
        RECT 101.155 -118.485 101.485 -118.155 ;
        RECT 101.155 -119.845 101.485 -119.515 ;
        RECT 101.155 -121.205 101.485 -120.875 ;
        RECT 101.155 -122.565 101.485 -122.235 ;
        RECT 101.155 -123.925 101.485 -123.595 ;
        RECT 101.155 -125.285 101.485 -124.955 ;
        RECT 101.155 -126.645 101.485 -126.315 ;
        RECT 101.155 -128.005 101.485 -127.675 ;
        RECT 101.155 -129.365 101.485 -129.035 ;
        RECT 101.155 -130.725 101.485 -130.395 ;
        RECT 101.155 -132.085 101.485 -131.755 ;
        RECT 101.155 -133.445 101.485 -133.115 ;
        RECT 101.155 -134.805 101.485 -134.475 ;
        RECT 101.155 -136.165 101.485 -135.835 ;
        RECT 101.155 -137.525 101.485 -137.195 ;
        RECT 101.155 -138.885 101.485 -138.555 ;
        RECT 101.155 -140.245 101.485 -139.915 ;
        RECT 101.155 -141.605 101.485 -141.275 ;
        RECT 101.155 -142.965 101.485 -142.635 ;
        RECT 101.155 -144.325 101.485 -143.995 ;
        RECT 101.155 -145.685 101.485 -145.355 ;
        RECT 101.155 -147.045 101.485 -146.715 ;
        RECT 101.155 -148.405 101.485 -148.075 ;
        RECT 101.155 -149.765 101.485 -149.435 ;
        RECT 101.155 -151.125 101.485 -150.795 ;
        RECT 101.155 -152.485 101.485 -152.155 ;
        RECT 101.155 -153.845 101.485 -153.515 ;
        RECT 101.155 -155.205 101.485 -154.875 ;
        RECT 101.155 -156.565 101.485 -156.235 ;
        RECT 101.155 -157.925 101.485 -157.595 ;
        RECT 101.155 -159.285 101.485 -158.955 ;
        RECT 101.155 -160.645 101.485 -160.315 ;
        RECT 101.155 -162.005 101.485 -161.675 ;
        RECT 101.155 -163.365 101.485 -163.035 ;
        RECT 101.155 -164.725 101.485 -164.395 ;
        RECT 101.155 -166.085 101.485 -165.755 ;
        RECT 101.155 -167.445 101.485 -167.115 ;
        RECT 101.155 -168.805 101.485 -168.475 ;
        RECT 101.155 -170.165 101.485 -169.835 ;
        RECT 101.155 -171.525 101.485 -171.195 ;
        RECT 101.155 -172.885 101.485 -172.555 ;
        RECT 101.155 -174.245 101.485 -173.915 ;
        RECT 101.155 -175.605 101.485 -175.275 ;
        RECT 101.155 -176.965 101.485 -176.635 ;
        RECT 101.155 -178.325 101.485 -177.995 ;
        RECT 101.155 -179.685 101.485 -179.355 ;
        RECT 101.155 -181.93 101.485 -180.8 ;
        RECT 101.16 -182.045 101.48 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 101.41 -98.075 101.74 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 241.32 102.845 242.45 ;
        RECT 102.515 239.195 102.845 239.525 ;
        RECT 102.515 237.835 102.845 238.165 ;
        RECT 102.52 237.16 102.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 102.515 -1.525 102.845 -1.195 ;
        RECT 102.515 -2.885 102.845 -2.555 ;
        RECT 102.52 -3.56 102.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 241.32 104.205 242.45 ;
        RECT 103.875 239.195 104.205 239.525 ;
        RECT 103.875 237.835 104.205 238.165 ;
        RECT 103.88 237.16 104.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 103.875 -1.525 104.205 -1.195 ;
        RECT 103.875 -2.885 104.205 -2.555 ;
        RECT 103.88 -3.56 104.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 241.32 105.565 242.45 ;
        RECT 105.235 239.195 105.565 239.525 ;
        RECT 105.235 237.835 105.565 238.165 ;
        RECT 105.24 237.16 105.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 -1.525 105.565 -1.195 ;
        RECT 105.235 -2.885 105.565 -2.555 ;
        RECT 105.24 -3.56 105.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 105.235 -95.365 105.565 -95.035 ;
        RECT 105.235 -96.725 105.565 -96.395 ;
        RECT 105.235 -98.085 105.565 -97.755 ;
        RECT 105.235 -99.445 105.565 -99.115 ;
        RECT 105.235 -100.805 105.565 -100.475 ;
        RECT 105.235 -102.165 105.565 -101.835 ;
        RECT 105.235 -103.525 105.565 -103.195 ;
        RECT 105.235 -104.885 105.565 -104.555 ;
        RECT 105.235 -106.245 105.565 -105.915 ;
        RECT 105.235 -107.605 105.565 -107.275 ;
        RECT 105.235 -108.965 105.565 -108.635 ;
        RECT 105.235 -110.325 105.565 -109.995 ;
        RECT 105.235 -111.685 105.565 -111.355 ;
        RECT 105.235 -113.045 105.565 -112.715 ;
        RECT 105.235 -114.405 105.565 -114.075 ;
        RECT 105.235 -115.765 105.565 -115.435 ;
        RECT 105.235 -117.125 105.565 -116.795 ;
        RECT 105.235 -118.485 105.565 -118.155 ;
        RECT 105.235 -119.845 105.565 -119.515 ;
        RECT 105.235 -121.205 105.565 -120.875 ;
        RECT 105.235 -122.565 105.565 -122.235 ;
        RECT 105.235 -123.925 105.565 -123.595 ;
        RECT 105.235 -125.285 105.565 -124.955 ;
        RECT 105.235 -126.645 105.565 -126.315 ;
        RECT 105.235 -128.005 105.565 -127.675 ;
        RECT 105.235 -129.365 105.565 -129.035 ;
        RECT 105.235 -130.725 105.565 -130.395 ;
        RECT 105.235 -132.085 105.565 -131.755 ;
        RECT 105.235 -133.445 105.565 -133.115 ;
        RECT 105.235 -134.805 105.565 -134.475 ;
        RECT 105.235 -136.165 105.565 -135.835 ;
        RECT 105.235 -137.525 105.565 -137.195 ;
        RECT 105.235 -138.885 105.565 -138.555 ;
        RECT 105.235 -140.245 105.565 -139.915 ;
        RECT 105.235 -141.605 105.565 -141.275 ;
        RECT 105.235 -142.965 105.565 -142.635 ;
        RECT 105.235 -144.325 105.565 -143.995 ;
        RECT 105.235 -145.685 105.565 -145.355 ;
        RECT 105.235 -147.045 105.565 -146.715 ;
        RECT 105.235 -148.405 105.565 -148.075 ;
        RECT 105.235 -149.765 105.565 -149.435 ;
        RECT 105.235 -151.125 105.565 -150.795 ;
        RECT 105.235 -152.485 105.565 -152.155 ;
        RECT 105.235 -153.845 105.565 -153.515 ;
        RECT 105.235 -155.205 105.565 -154.875 ;
        RECT 105.235 -156.565 105.565 -156.235 ;
        RECT 105.235 -157.925 105.565 -157.595 ;
        RECT 105.235 -159.285 105.565 -158.955 ;
        RECT 105.235 -160.645 105.565 -160.315 ;
        RECT 105.235 -162.005 105.565 -161.675 ;
        RECT 105.235 -163.365 105.565 -163.035 ;
        RECT 105.235 -164.725 105.565 -164.395 ;
        RECT 105.235 -166.085 105.565 -165.755 ;
        RECT 105.235 -167.445 105.565 -167.115 ;
        RECT 105.235 -168.805 105.565 -168.475 ;
        RECT 105.235 -170.165 105.565 -169.835 ;
        RECT 105.235 -171.525 105.565 -171.195 ;
        RECT 105.235 -172.885 105.565 -172.555 ;
        RECT 105.235 -174.245 105.565 -173.915 ;
        RECT 105.235 -175.605 105.565 -175.275 ;
        RECT 105.235 -176.965 105.565 -176.635 ;
        RECT 105.235 -178.325 105.565 -177.995 ;
        RECT 105.235 -179.685 105.565 -179.355 ;
        RECT 105.235 -181.93 105.565 -180.8 ;
        RECT 105.24 -182.045 105.56 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 241.32 106.925 242.45 ;
        RECT 106.595 239.195 106.925 239.525 ;
        RECT 106.595 237.835 106.925 238.165 ;
        RECT 106.6 237.16 106.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 -1.525 106.925 -1.195 ;
        RECT 106.595 -2.885 106.925 -2.555 ;
        RECT 106.6 -3.56 106.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 106.595 -95.365 106.925 -95.035 ;
        RECT 106.595 -96.725 106.925 -96.395 ;
        RECT 106.595 -98.085 106.925 -97.755 ;
        RECT 106.595 -99.445 106.925 -99.115 ;
        RECT 106.595 -100.805 106.925 -100.475 ;
        RECT 106.595 -102.165 106.925 -101.835 ;
        RECT 106.595 -103.525 106.925 -103.195 ;
        RECT 106.595 -104.885 106.925 -104.555 ;
        RECT 106.595 -106.245 106.925 -105.915 ;
        RECT 106.595 -107.605 106.925 -107.275 ;
        RECT 106.595 -108.965 106.925 -108.635 ;
        RECT 106.595 -110.325 106.925 -109.995 ;
        RECT 106.595 -111.685 106.925 -111.355 ;
        RECT 106.595 -113.045 106.925 -112.715 ;
        RECT 106.595 -114.405 106.925 -114.075 ;
        RECT 106.595 -115.765 106.925 -115.435 ;
        RECT 106.595 -117.125 106.925 -116.795 ;
        RECT 106.595 -118.485 106.925 -118.155 ;
        RECT 106.595 -119.845 106.925 -119.515 ;
        RECT 106.595 -121.205 106.925 -120.875 ;
        RECT 106.595 -122.565 106.925 -122.235 ;
        RECT 106.595 -123.925 106.925 -123.595 ;
        RECT 106.595 -125.285 106.925 -124.955 ;
        RECT 106.595 -126.645 106.925 -126.315 ;
        RECT 106.595 -128.005 106.925 -127.675 ;
        RECT 106.595 -129.365 106.925 -129.035 ;
        RECT 106.595 -130.725 106.925 -130.395 ;
        RECT 106.595 -132.085 106.925 -131.755 ;
        RECT 106.595 -133.445 106.925 -133.115 ;
        RECT 106.595 -134.805 106.925 -134.475 ;
        RECT 106.595 -136.165 106.925 -135.835 ;
        RECT 106.595 -137.525 106.925 -137.195 ;
        RECT 106.595 -138.885 106.925 -138.555 ;
        RECT 106.595 -140.245 106.925 -139.915 ;
        RECT 106.595 -141.605 106.925 -141.275 ;
        RECT 106.595 -142.965 106.925 -142.635 ;
        RECT 106.595 -144.325 106.925 -143.995 ;
        RECT 106.595 -145.685 106.925 -145.355 ;
        RECT 106.595 -147.045 106.925 -146.715 ;
        RECT 106.595 -148.405 106.925 -148.075 ;
        RECT 106.595 -149.765 106.925 -149.435 ;
        RECT 106.595 -151.125 106.925 -150.795 ;
        RECT 106.595 -152.485 106.925 -152.155 ;
        RECT 106.595 -153.845 106.925 -153.515 ;
        RECT 106.595 -155.205 106.925 -154.875 ;
        RECT 106.595 -156.565 106.925 -156.235 ;
        RECT 106.595 -157.925 106.925 -157.595 ;
        RECT 106.595 -159.285 106.925 -158.955 ;
        RECT 106.595 -160.645 106.925 -160.315 ;
        RECT 106.595 -162.005 106.925 -161.675 ;
        RECT 106.595 -163.365 106.925 -163.035 ;
        RECT 106.595 -164.725 106.925 -164.395 ;
        RECT 106.595 -166.085 106.925 -165.755 ;
        RECT 106.595 -167.445 106.925 -167.115 ;
        RECT 106.595 -168.805 106.925 -168.475 ;
        RECT 106.595 -170.165 106.925 -169.835 ;
        RECT 106.595 -171.525 106.925 -171.195 ;
        RECT 106.595 -172.885 106.925 -172.555 ;
        RECT 106.595 -174.245 106.925 -173.915 ;
        RECT 106.595 -175.605 106.925 -175.275 ;
        RECT 106.595 -176.965 106.925 -176.635 ;
        RECT 106.595 -178.325 106.925 -177.995 ;
        RECT 106.595 -179.685 106.925 -179.355 ;
        RECT 106.595 -181.93 106.925 -180.8 ;
        RECT 106.6 -182.045 106.92 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 241.32 108.285 242.45 ;
        RECT 107.955 239.195 108.285 239.525 ;
        RECT 107.955 237.835 108.285 238.165 ;
        RECT 107.96 237.16 108.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 -1.525 108.285 -1.195 ;
        RECT 107.955 -2.885 108.285 -2.555 ;
        RECT 107.96 -3.56 108.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 107.955 -95.365 108.285 -95.035 ;
        RECT 107.955 -96.725 108.285 -96.395 ;
        RECT 107.955 -98.085 108.285 -97.755 ;
        RECT 107.955 -99.445 108.285 -99.115 ;
        RECT 107.955 -100.805 108.285 -100.475 ;
        RECT 107.955 -102.165 108.285 -101.835 ;
        RECT 107.955 -103.525 108.285 -103.195 ;
        RECT 107.955 -104.885 108.285 -104.555 ;
        RECT 107.955 -106.245 108.285 -105.915 ;
        RECT 107.955 -107.605 108.285 -107.275 ;
        RECT 107.955 -108.965 108.285 -108.635 ;
        RECT 107.955 -110.325 108.285 -109.995 ;
        RECT 107.955 -111.685 108.285 -111.355 ;
        RECT 107.955 -113.045 108.285 -112.715 ;
        RECT 107.955 -114.405 108.285 -114.075 ;
        RECT 107.955 -115.765 108.285 -115.435 ;
        RECT 107.955 -117.125 108.285 -116.795 ;
        RECT 107.955 -118.485 108.285 -118.155 ;
        RECT 107.955 -119.845 108.285 -119.515 ;
        RECT 107.955 -121.205 108.285 -120.875 ;
        RECT 107.955 -122.565 108.285 -122.235 ;
        RECT 107.955 -123.925 108.285 -123.595 ;
        RECT 107.955 -125.285 108.285 -124.955 ;
        RECT 107.955 -126.645 108.285 -126.315 ;
        RECT 107.955 -128.005 108.285 -127.675 ;
        RECT 107.955 -129.365 108.285 -129.035 ;
        RECT 107.955 -130.725 108.285 -130.395 ;
        RECT 107.955 -132.085 108.285 -131.755 ;
        RECT 107.955 -133.445 108.285 -133.115 ;
        RECT 107.955 -134.805 108.285 -134.475 ;
        RECT 107.955 -136.165 108.285 -135.835 ;
        RECT 107.955 -137.525 108.285 -137.195 ;
        RECT 107.955 -138.885 108.285 -138.555 ;
        RECT 107.955 -140.245 108.285 -139.915 ;
        RECT 107.955 -141.605 108.285 -141.275 ;
        RECT 107.955 -142.965 108.285 -142.635 ;
        RECT 107.955 -144.325 108.285 -143.995 ;
        RECT 107.955 -145.685 108.285 -145.355 ;
        RECT 107.955 -147.045 108.285 -146.715 ;
        RECT 107.955 -148.405 108.285 -148.075 ;
        RECT 107.955 -149.765 108.285 -149.435 ;
        RECT 107.955 -151.125 108.285 -150.795 ;
        RECT 107.955 -152.485 108.285 -152.155 ;
        RECT 107.955 -153.845 108.285 -153.515 ;
        RECT 107.955 -155.205 108.285 -154.875 ;
        RECT 107.955 -156.565 108.285 -156.235 ;
        RECT 107.955 -157.925 108.285 -157.595 ;
        RECT 107.955 -159.285 108.285 -158.955 ;
        RECT 107.955 -160.645 108.285 -160.315 ;
        RECT 107.955 -162.005 108.285 -161.675 ;
        RECT 107.955 -163.365 108.285 -163.035 ;
        RECT 107.955 -164.725 108.285 -164.395 ;
        RECT 107.955 -166.085 108.285 -165.755 ;
        RECT 107.955 -167.445 108.285 -167.115 ;
        RECT 107.955 -168.805 108.285 -168.475 ;
        RECT 107.955 -170.165 108.285 -169.835 ;
        RECT 107.955 -171.525 108.285 -171.195 ;
        RECT 107.955 -172.885 108.285 -172.555 ;
        RECT 107.955 -174.245 108.285 -173.915 ;
        RECT 107.955 -175.605 108.285 -175.275 ;
        RECT 107.955 -176.965 108.285 -176.635 ;
        RECT 107.955 -178.325 108.285 -177.995 ;
        RECT 107.955 -179.685 108.285 -179.355 ;
        RECT 107.955 -181.93 108.285 -180.8 ;
        RECT 107.96 -182.045 108.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 241.32 109.645 242.45 ;
        RECT 109.315 239.195 109.645 239.525 ;
        RECT 109.315 237.835 109.645 238.165 ;
        RECT 109.32 237.16 109.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 -1.525 109.645 -1.195 ;
        RECT 109.315 -2.885 109.645 -2.555 ;
        RECT 109.32 -3.56 109.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 109.315 -95.365 109.645 -95.035 ;
        RECT 109.315 -96.725 109.645 -96.395 ;
        RECT 109.315 -98.085 109.645 -97.755 ;
        RECT 109.315 -99.445 109.645 -99.115 ;
        RECT 109.315 -100.805 109.645 -100.475 ;
        RECT 109.315 -102.165 109.645 -101.835 ;
        RECT 109.315 -103.525 109.645 -103.195 ;
        RECT 109.315 -104.885 109.645 -104.555 ;
        RECT 109.315 -106.245 109.645 -105.915 ;
        RECT 109.315 -107.605 109.645 -107.275 ;
        RECT 109.315 -108.965 109.645 -108.635 ;
        RECT 109.315 -110.325 109.645 -109.995 ;
        RECT 109.315 -111.685 109.645 -111.355 ;
        RECT 109.315 -113.045 109.645 -112.715 ;
        RECT 109.315 -114.405 109.645 -114.075 ;
        RECT 109.315 -115.765 109.645 -115.435 ;
        RECT 109.315 -117.125 109.645 -116.795 ;
        RECT 109.315 -118.485 109.645 -118.155 ;
        RECT 109.315 -119.845 109.645 -119.515 ;
        RECT 109.315 -121.205 109.645 -120.875 ;
        RECT 109.315 -122.565 109.645 -122.235 ;
        RECT 109.315 -123.925 109.645 -123.595 ;
        RECT 109.315 -125.285 109.645 -124.955 ;
        RECT 109.315 -126.645 109.645 -126.315 ;
        RECT 109.315 -128.005 109.645 -127.675 ;
        RECT 109.315 -129.365 109.645 -129.035 ;
        RECT 109.315 -130.725 109.645 -130.395 ;
        RECT 109.315 -132.085 109.645 -131.755 ;
        RECT 109.315 -133.445 109.645 -133.115 ;
        RECT 109.315 -134.805 109.645 -134.475 ;
        RECT 109.315 -136.165 109.645 -135.835 ;
        RECT 109.315 -137.525 109.645 -137.195 ;
        RECT 109.315 -138.885 109.645 -138.555 ;
        RECT 109.315 -140.245 109.645 -139.915 ;
        RECT 109.315 -141.605 109.645 -141.275 ;
        RECT 109.315 -142.965 109.645 -142.635 ;
        RECT 109.315 -144.325 109.645 -143.995 ;
        RECT 109.315 -145.685 109.645 -145.355 ;
        RECT 109.315 -147.045 109.645 -146.715 ;
        RECT 109.315 -148.405 109.645 -148.075 ;
        RECT 109.315 -149.765 109.645 -149.435 ;
        RECT 109.315 -151.125 109.645 -150.795 ;
        RECT 109.315 -152.485 109.645 -152.155 ;
        RECT 109.315 -153.845 109.645 -153.515 ;
        RECT 109.315 -155.205 109.645 -154.875 ;
        RECT 109.315 -156.565 109.645 -156.235 ;
        RECT 109.315 -157.925 109.645 -157.595 ;
        RECT 109.315 -159.285 109.645 -158.955 ;
        RECT 109.315 -160.645 109.645 -160.315 ;
        RECT 109.315 -162.005 109.645 -161.675 ;
        RECT 109.315 -163.365 109.645 -163.035 ;
        RECT 109.315 -164.725 109.645 -164.395 ;
        RECT 109.315 -166.085 109.645 -165.755 ;
        RECT 109.315 -167.445 109.645 -167.115 ;
        RECT 109.315 -168.805 109.645 -168.475 ;
        RECT 109.315 -170.165 109.645 -169.835 ;
        RECT 109.315 -171.525 109.645 -171.195 ;
        RECT 109.315 -172.885 109.645 -172.555 ;
        RECT 109.315 -174.245 109.645 -173.915 ;
        RECT 109.315 -175.605 109.645 -175.275 ;
        RECT 109.315 -176.965 109.645 -176.635 ;
        RECT 109.315 -178.325 109.645 -177.995 ;
        RECT 109.315 -179.685 109.645 -179.355 ;
        RECT 109.315 -181.93 109.645 -180.8 ;
        RECT 109.32 -182.045 109.64 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 241.32 111.005 242.45 ;
        RECT 110.675 239.195 111.005 239.525 ;
        RECT 110.675 237.835 111.005 238.165 ;
        RECT 110.68 237.16 111 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 -1.525 111.005 -1.195 ;
        RECT 110.675 -2.885 111.005 -2.555 ;
        RECT 110.68 -3.56 111 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 110.675 -95.365 111.005 -95.035 ;
        RECT 110.675 -96.725 111.005 -96.395 ;
        RECT 110.675 -98.085 111.005 -97.755 ;
        RECT 110.675 -99.445 111.005 -99.115 ;
        RECT 110.675 -100.805 111.005 -100.475 ;
        RECT 110.675 -102.165 111.005 -101.835 ;
        RECT 110.675 -103.525 111.005 -103.195 ;
        RECT 110.675 -104.885 111.005 -104.555 ;
        RECT 110.675 -106.245 111.005 -105.915 ;
        RECT 110.675 -107.605 111.005 -107.275 ;
        RECT 110.675 -108.965 111.005 -108.635 ;
        RECT 110.675 -110.325 111.005 -109.995 ;
        RECT 110.675 -111.685 111.005 -111.355 ;
        RECT 110.675 -113.045 111.005 -112.715 ;
        RECT 110.675 -114.405 111.005 -114.075 ;
        RECT 110.675 -115.765 111.005 -115.435 ;
        RECT 110.675 -117.125 111.005 -116.795 ;
        RECT 110.675 -118.485 111.005 -118.155 ;
        RECT 110.675 -119.845 111.005 -119.515 ;
        RECT 110.675 -121.205 111.005 -120.875 ;
        RECT 110.675 -122.565 111.005 -122.235 ;
        RECT 110.675 -123.925 111.005 -123.595 ;
        RECT 110.675 -125.285 111.005 -124.955 ;
        RECT 110.675 -126.645 111.005 -126.315 ;
        RECT 110.675 -128.005 111.005 -127.675 ;
        RECT 110.675 -129.365 111.005 -129.035 ;
        RECT 110.675 -130.725 111.005 -130.395 ;
        RECT 110.675 -132.085 111.005 -131.755 ;
        RECT 110.675 -133.445 111.005 -133.115 ;
        RECT 110.675 -134.805 111.005 -134.475 ;
        RECT 110.675 -136.165 111.005 -135.835 ;
        RECT 110.675 -137.525 111.005 -137.195 ;
        RECT 110.675 -138.885 111.005 -138.555 ;
        RECT 110.675 -140.245 111.005 -139.915 ;
        RECT 110.675 -141.605 111.005 -141.275 ;
        RECT 110.675 -142.965 111.005 -142.635 ;
        RECT 110.675 -144.325 111.005 -143.995 ;
        RECT 110.675 -145.685 111.005 -145.355 ;
        RECT 110.675 -147.045 111.005 -146.715 ;
        RECT 110.675 -148.405 111.005 -148.075 ;
        RECT 110.675 -149.765 111.005 -149.435 ;
        RECT 110.675 -151.125 111.005 -150.795 ;
        RECT 110.675 -152.485 111.005 -152.155 ;
        RECT 110.675 -153.845 111.005 -153.515 ;
        RECT 110.675 -155.205 111.005 -154.875 ;
        RECT 110.675 -156.565 111.005 -156.235 ;
        RECT 110.675 -157.925 111.005 -157.595 ;
        RECT 110.675 -159.285 111.005 -158.955 ;
        RECT 110.675 -160.645 111.005 -160.315 ;
        RECT 110.675 -162.005 111.005 -161.675 ;
        RECT 110.675 -163.365 111.005 -163.035 ;
        RECT 110.675 -164.725 111.005 -164.395 ;
        RECT 110.675 -166.085 111.005 -165.755 ;
        RECT 110.675 -167.445 111.005 -167.115 ;
        RECT 110.675 -168.805 111.005 -168.475 ;
        RECT 110.675 -170.165 111.005 -169.835 ;
        RECT 110.675 -171.525 111.005 -171.195 ;
        RECT 110.675 -172.885 111.005 -172.555 ;
        RECT 110.675 -174.245 111.005 -173.915 ;
        RECT 110.675 -175.605 111.005 -175.275 ;
        RECT 110.675 -176.965 111.005 -176.635 ;
        RECT 110.675 -178.325 111.005 -177.995 ;
        RECT 110.675 -179.685 111.005 -179.355 ;
        RECT 110.675 -181.93 111.005 -180.8 ;
        RECT 110.68 -182.045 111 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 241.32 112.365 242.45 ;
        RECT 112.035 239.195 112.365 239.525 ;
        RECT 112.035 237.835 112.365 238.165 ;
        RECT 112.04 237.16 112.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.035 -99.445 112.365 -99.115 ;
        RECT 112.035 -100.805 112.365 -100.475 ;
        RECT 112.035 -102.165 112.365 -101.835 ;
        RECT 112.035 -103.525 112.365 -103.195 ;
        RECT 112.035 -104.885 112.365 -104.555 ;
        RECT 112.035 -106.245 112.365 -105.915 ;
        RECT 112.035 -107.605 112.365 -107.275 ;
        RECT 112.035 -108.965 112.365 -108.635 ;
        RECT 112.035 -110.325 112.365 -109.995 ;
        RECT 112.035 -111.685 112.365 -111.355 ;
        RECT 112.035 -113.045 112.365 -112.715 ;
        RECT 112.035 -114.405 112.365 -114.075 ;
        RECT 112.035 -115.765 112.365 -115.435 ;
        RECT 112.035 -117.125 112.365 -116.795 ;
        RECT 112.035 -118.485 112.365 -118.155 ;
        RECT 112.035 -119.845 112.365 -119.515 ;
        RECT 112.035 -121.205 112.365 -120.875 ;
        RECT 112.035 -122.565 112.365 -122.235 ;
        RECT 112.035 -123.925 112.365 -123.595 ;
        RECT 112.035 -125.285 112.365 -124.955 ;
        RECT 112.035 -126.645 112.365 -126.315 ;
        RECT 112.035 -128.005 112.365 -127.675 ;
        RECT 112.035 -129.365 112.365 -129.035 ;
        RECT 112.035 -130.725 112.365 -130.395 ;
        RECT 112.035 -132.085 112.365 -131.755 ;
        RECT 112.035 -133.445 112.365 -133.115 ;
        RECT 112.035 -134.805 112.365 -134.475 ;
        RECT 112.035 -136.165 112.365 -135.835 ;
        RECT 112.035 -137.525 112.365 -137.195 ;
        RECT 112.035 -138.885 112.365 -138.555 ;
        RECT 112.035 -140.245 112.365 -139.915 ;
        RECT 112.035 -141.605 112.365 -141.275 ;
        RECT 112.035 -142.965 112.365 -142.635 ;
        RECT 112.035 -144.325 112.365 -143.995 ;
        RECT 112.035 -145.685 112.365 -145.355 ;
        RECT 112.035 -147.045 112.365 -146.715 ;
        RECT 112.035 -148.405 112.365 -148.075 ;
        RECT 112.035 -149.765 112.365 -149.435 ;
        RECT 112.035 -151.125 112.365 -150.795 ;
        RECT 112.035 -152.485 112.365 -152.155 ;
        RECT 112.035 -153.845 112.365 -153.515 ;
        RECT 112.035 -155.205 112.365 -154.875 ;
        RECT 112.035 -156.565 112.365 -156.235 ;
        RECT 112.035 -157.925 112.365 -157.595 ;
        RECT 112.035 -159.285 112.365 -158.955 ;
        RECT 112.035 -160.645 112.365 -160.315 ;
        RECT 112.035 -162.005 112.365 -161.675 ;
        RECT 112.035 -163.365 112.365 -163.035 ;
        RECT 112.035 -164.725 112.365 -164.395 ;
        RECT 112.035 -166.085 112.365 -165.755 ;
        RECT 112.035 -167.445 112.365 -167.115 ;
        RECT 112.035 -168.805 112.365 -168.475 ;
        RECT 112.035 -170.165 112.365 -169.835 ;
        RECT 112.035 -171.525 112.365 -171.195 ;
        RECT 112.035 -172.885 112.365 -172.555 ;
        RECT 112.035 -174.245 112.365 -173.915 ;
        RECT 112.035 -175.605 112.365 -175.275 ;
        RECT 112.035 -176.965 112.365 -176.635 ;
        RECT 112.035 -178.325 112.365 -177.995 ;
        RECT 112.035 -179.685 112.365 -179.355 ;
        RECT 112.035 -181.93 112.365 -180.8 ;
        RECT 112.04 -182.045 112.36 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 112.31 -98.075 112.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.395 241.32 113.725 242.45 ;
        RECT 113.395 239.195 113.725 239.525 ;
        RECT 113.395 237.835 113.725 238.165 ;
        RECT 113.4 237.16 113.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 113.395 -1.525 113.725 -1.195 ;
        RECT 113.395 -2.885 113.725 -2.555 ;
        RECT 113.4 -3.56 113.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 241.32 115.085 242.45 ;
        RECT 114.755 239.195 115.085 239.525 ;
        RECT 114.755 237.835 115.085 238.165 ;
        RECT 114.76 237.16 115.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 114.755 -1.525 115.085 -1.195 ;
        RECT 114.755 -2.885 115.085 -2.555 ;
        RECT 114.76 -3.56 115.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 241.32 116.445 242.45 ;
        RECT 116.115 239.195 116.445 239.525 ;
        RECT 116.115 237.835 116.445 238.165 ;
        RECT 116.12 237.16 116.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 -1.525 116.445 -1.195 ;
        RECT 116.115 -2.885 116.445 -2.555 ;
        RECT 116.12 -3.56 116.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 116.115 -95.365 116.445 -95.035 ;
        RECT 116.115 -96.725 116.445 -96.395 ;
        RECT 116.115 -98.085 116.445 -97.755 ;
        RECT 116.115 -99.445 116.445 -99.115 ;
        RECT 116.115 -100.805 116.445 -100.475 ;
        RECT 116.115 -102.165 116.445 -101.835 ;
        RECT 116.115 -103.525 116.445 -103.195 ;
        RECT 116.115 -104.885 116.445 -104.555 ;
        RECT 116.115 -106.245 116.445 -105.915 ;
        RECT 116.115 -107.605 116.445 -107.275 ;
        RECT 116.115 -108.965 116.445 -108.635 ;
        RECT 116.115 -110.325 116.445 -109.995 ;
        RECT 116.115 -111.685 116.445 -111.355 ;
        RECT 116.115 -113.045 116.445 -112.715 ;
        RECT 116.115 -114.405 116.445 -114.075 ;
        RECT 116.115 -115.765 116.445 -115.435 ;
        RECT 116.115 -117.125 116.445 -116.795 ;
        RECT 116.115 -118.485 116.445 -118.155 ;
        RECT 116.115 -119.845 116.445 -119.515 ;
        RECT 116.115 -121.205 116.445 -120.875 ;
        RECT 116.115 -122.565 116.445 -122.235 ;
        RECT 116.115 -123.925 116.445 -123.595 ;
        RECT 116.115 -125.285 116.445 -124.955 ;
        RECT 116.115 -126.645 116.445 -126.315 ;
        RECT 116.115 -128.005 116.445 -127.675 ;
        RECT 116.115 -129.365 116.445 -129.035 ;
        RECT 116.115 -130.725 116.445 -130.395 ;
        RECT 116.115 -132.085 116.445 -131.755 ;
        RECT 116.115 -133.445 116.445 -133.115 ;
        RECT 116.115 -134.805 116.445 -134.475 ;
        RECT 116.115 -136.165 116.445 -135.835 ;
        RECT 116.115 -137.525 116.445 -137.195 ;
        RECT 116.115 -138.885 116.445 -138.555 ;
        RECT 116.115 -140.245 116.445 -139.915 ;
        RECT 116.115 -141.605 116.445 -141.275 ;
        RECT 116.115 -142.965 116.445 -142.635 ;
        RECT 116.115 -144.325 116.445 -143.995 ;
        RECT 116.115 -145.685 116.445 -145.355 ;
        RECT 116.115 -147.045 116.445 -146.715 ;
        RECT 116.115 -148.405 116.445 -148.075 ;
        RECT 116.115 -149.765 116.445 -149.435 ;
        RECT 116.115 -151.125 116.445 -150.795 ;
        RECT 116.115 -152.485 116.445 -152.155 ;
        RECT 116.115 -153.845 116.445 -153.515 ;
        RECT 116.115 -155.205 116.445 -154.875 ;
        RECT 116.115 -156.565 116.445 -156.235 ;
        RECT 116.115 -157.925 116.445 -157.595 ;
        RECT 116.115 -159.285 116.445 -158.955 ;
        RECT 116.115 -160.645 116.445 -160.315 ;
        RECT 116.115 -162.005 116.445 -161.675 ;
        RECT 116.115 -163.365 116.445 -163.035 ;
        RECT 116.115 -164.725 116.445 -164.395 ;
        RECT 116.115 -166.085 116.445 -165.755 ;
        RECT 116.115 -167.445 116.445 -167.115 ;
        RECT 116.115 -168.805 116.445 -168.475 ;
        RECT 116.115 -170.165 116.445 -169.835 ;
        RECT 116.115 -171.525 116.445 -171.195 ;
        RECT 116.115 -172.885 116.445 -172.555 ;
        RECT 116.115 -174.245 116.445 -173.915 ;
        RECT 116.115 -175.605 116.445 -175.275 ;
        RECT 116.115 -176.965 116.445 -176.635 ;
        RECT 116.115 -178.325 116.445 -177.995 ;
        RECT 116.115 -179.685 116.445 -179.355 ;
        RECT 116.115 -181.93 116.445 -180.8 ;
        RECT 116.12 -182.045 116.44 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 241.32 117.805 242.45 ;
        RECT 117.475 239.195 117.805 239.525 ;
        RECT 117.475 237.835 117.805 238.165 ;
        RECT 117.48 237.16 117.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 -1.525 117.805 -1.195 ;
        RECT 117.475 -2.885 117.805 -2.555 ;
        RECT 117.48 -3.56 117.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 117.475 -149.765 117.805 -149.435 ;
        RECT 117.475 -151.125 117.805 -150.795 ;
        RECT 117.475 -152.485 117.805 -152.155 ;
        RECT 117.475 -153.845 117.805 -153.515 ;
        RECT 117.475 -155.205 117.805 -154.875 ;
        RECT 117.475 -156.565 117.805 -156.235 ;
        RECT 117.475 -157.925 117.805 -157.595 ;
        RECT 117.475 -159.285 117.805 -158.955 ;
        RECT 117.475 -160.645 117.805 -160.315 ;
        RECT 117.475 -162.005 117.805 -161.675 ;
        RECT 117.475 -163.365 117.805 -163.035 ;
        RECT 117.475 -164.725 117.805 -164.395 ;
        RECT 117.475 -166.085 117.805 -165.755 ;
        RECT 117.475 -167.445 117.805 -167.115 ;
        RECT 117.475 -168.805 117.805 -168.475 ;
        RECT 117.475 -170.165 117.805 -169.835 ;
        RECT 117.475 -171.525 117.805 -171.195 ;
        RECT 117.475 -172.885 117.805 -172.555 ;
        RECT 117.475 -174.245 117.805 -173.915 ;
        RECT 117.475 -175.605 117.805 -175.275 ;
        RECT 117.475 -176.965 117.805 -176.635 ;
        RECT 117.475 -178.325 117.805 -177.995 ;
        RECT 117.475 -179.685 117.805 -179.355 ;
        RECT 117.475 -181.93 117.805 -180.8 ;
        RECT 117.48 -182.045 117.8 -95.035 ;
        RECT 117.475 -95.365 117.805 -95.035 ;
        RECT 117.475 -96.725 117.805 -96.395 ;
        RECT 117.475 -98.085 117.805 -97.755 ;
        RECT 117.475 -99.445 117.805 -99.115 ;
        RECT 117.475 -100.805 117.805 -100.475 ;
        RECT 117.475 -102.165 117.805 -101.835 ;
        RECT 117.475 -103.525 117.805 -103.195 ;
        RECT 117.475 -104.885 117.805 -104.555 ;
        RECT 117.475 -106.245 117.805 -105.915 ;
        RECT 117.475 -107.605 117.805 -107.275 ;
        RECT 117.475 -108.965 117.805 -108.635 ;
        RECT 117.475 -110.325 117.805 -109.995 ;
        RECT 117.475 -111.685 117.805 -111.355 ;
        RECT 117.475 -113.045 117.805 -112.715 ;
        RECT 117.475 -114.405 117.805 -114.075 ;
        RECT 117.475 -115.765 117.805 -115.435 ;
        RECT 117.475 -117.125 117.805 -116.795 ;
        RECT 117.475 -118.485 117.805 -118.155 ;
        RECT 117.475 -119.845 117.805 -119.515 ;
        RECT 117.475 -121.205 117.805 -120.875 ;
        RECT 117.475 -122.565 117.805 -122.235 ;
        RECT 117.475 -123.925 117.805 -123.595 ;
        RECT 117.475 -125.285 117.805 -124.955 ;
        RECT 117.475 -126.645 117.805 -126.315 ;
        RECT 117.475 -128.005 117.805 -127.675 ;
        RECT 117.475 -129.365 117.805 -129.035 ;
        RECT 117.475 -130.725 117.805 -130.395 ;
        RECT 117.475 -132.085 117.805 -131.755 ;
        RECT 117.475 -133.445 117.805 -133.115 ;
        RECT 117.475 -134.805 117.805 -134.475 ;
        RECT 117.475 -136.165 117.805 -135.835 ;
        RECT 117.475 -137.525 117.805 -137.195 ;
        RECT 117.475 -138.885 117.805 -138.555 ;
        RECT 117.475 -140.245 117.805 -139.915 ;
        RECT 117.475 -141.605 117.805 -141.275 ;
        RECT 117.475 -142.965 117.805 -142.635 ;
        RECT 117.475 -144.325 117.805 -143.995 ;
        RECT 117.475 -145.685 117.805 -145.355 ;
        RECT 117.475 -147.045 117.805 -146.715 ;
        RECT 117.475 -148.405 117.805 -148.075 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 241.32 68.845 242.45 ;
        RECT 68.515 239.195 68.845 239.525 ;
        RECT 68.515 237.835 68.845 238.165 ;
        RECT 68.52 237.16 68.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.515 -99.445 68.845 -99.115 ;
        RECT 68.515 -100.805 68.845 -100.475 ;
        RECT 68.515 -102.165 68.845 -101.835 ;
        RECT 68.515 -103.525 68.845 -103.195 ;
        RECT 68.515 -104.885 68.845 -104.555 ;
        RECT 68.515 -106.245 68.845 -105.915 ;
        RECT 68.515 -107.605 68.845 -107.275 ;
        RECT 68.515 -108.965 68.845 -108.635 ;
        RECT 68.515 -110.325 68.845 -109.995 ;
        RECT 68.515 -111.685 68.845 -111.355 ;
        RECT 68.515 -113.045 68.845 -112.715 ;
        RECT 68.515 -114.405 68.845 -114.075 ;
        RECT 68.515 -115.765 68.845 -115.435 ;
        RECT 68.515 -117.125 68.845 -116.795 ;
        RECT 68.515 -118.485 68.845 -118.155 ;
        RECT 68.515 -119.845 68.845 -119.515 ;
        RECT 68.515 -121.205 68.845 -120.875 ;
        RECT 68.515 -122.565 68.845 -122.235 ;
        RECT 68.515 -123.925 68.845 -123.595 ;
        RECT 68.515 -125.285 68.845 -124.955 ;
        RECT 68.515 -126.645 68.845 -126.315 ;
        RECT 68.515 -128.005 68.845 -127.675 ;
        RECT 68.515 -129.365 68.845 -129.035 ;
        RECT 68.515 -130.725 68.845 -130.395 ;
        RECT 68.515 -132.085 68.845 -131.755 ;
        RECT 68.515 -133.445 68.845 -133.115 ;
        RECT 68.515 -134.805 68.845 -134.475 ;
        RECT 68.515 -136.165 68.845 -135.835 ;
        RECT 68.515 -137.525 68.845 -137.195 ;
        RECT 68.515 -138.885 68.845 -138.555 ;
        RECT 68.515 -140.245 68.845 -139.915 ;
        RECT 68.515 -141.605 68.845 -141.275 ;
        RECT 68.515 -142.965 68.845 -142.635 ;
        RECT 68.515 -144.325 68.845 -143.995 ;
        RECT 68.515 -145.685 68.845 -145.355 ;
        RECT 68.515 -147.045 68.845 -146.715 ;
        RECT 68.515 -148.405 68.845 -148.075 ;
        RECT 68.515 -149.765 68.845 -149.435 ;
        RECT 68.515 -151.125 68.845 -150.795 ;
        RECT 68.515 -152.485 68.845 -152.155 ;
        RECT 68.515 -153.845 68.845 -153.515 ;
        RECT 68.515 -155.205 68.845 -154.875 ;
        RECT 68.515 -156.565 68.845 -156.235 ;
        RECT 68.515 -157.925 68.845 -157.595 ;
        RECT 68.515 -159.285 68.845 -158.955 ;
        RECT 68.515 -160.645 68.845 -160.315 ;
        RECT 68.515 -162.005 68.845 -161.675 ;
        RECT 68.515 -163.365 68.845 -163.035 ;
        RECT 68.515 -164.725 68.845 -164.395 ;
        RECT 68.515 -166.085 68.845 -165.755 ;
        RECT 68.515 -167.445 68.845 -167.115 ;
        RECT 68.515 -168.805 68.845 -168.475 ;
        RECT 68.515 -170.165 68.845 -169.835 ;
        RECT 68.515 -171.525 68.845 -171.195 ;
        RECT 68.515 -172.885 68.845 -172.555 ;
        RECT 68.515 -174.245 68.845 -173.915 ;
        RECT 68.515 -175.605 68.845 -175.275 ;
        RECT 68.515 -176.965 68.845 -176.635 ;
        RECT 68.515 -178.325 68.845 -177.995 ;
        RECT 68.515 -179.685 68.845 -179.355 ;
        RECT 68.515 -181.93 68.845 -180.8 ;
        RECT 68.52 -182.045 68.84 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 68.71 -98.075 69.04 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 241.32 70.205 242.45 ;
        RECT 69.875 239.195 70.205 239.525 ;
        RECT 69.875 237.835 70.205 238.165 ;
        RECT 69.88 237.16 70.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 69.875 -1.525 70.205 -1.195 ;
        RECT 69.875 -2.885 70.205 -2.555 ;
        RECT 69.88 -3.56 70.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 241.32 71.565 242.45 ;
        RECT 71.235 239.195 71.565 239.525 ;
        RECT 71.235 237.835 71.565 238.165 ;
        RECT 71.24 237.16 71.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 71.235 -1.525 71.565 -1.195 ;
        RECT 71.235 -2.885 71.565 -2.555 ;
        RECT 71.24 -3.56 71.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 241.32 72.925 242.45 ;
        RECT 72.595 239.195 72.925 239.525 ;
        RECT 72.595 237.835 72.925 238.165 ;
        RECT 72.6 237.16 72.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 -1.525 72.925 -1.195 ;
        RECT 72.595 -2.885 72.925 -2.555 ;
        RECT 72.6 -3.56 72.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 72.595 -95.365 72.925 -95.035 ;
        RECT 72.595 -96.725 72.925 -96.395 ;
        RECT 72.595 -98.085 72.925 -97.755 ;
        RECT 72.595 -99.445 72.925 -99.115 ;
        RECT 72.595 -100.805 72.925 -100.475 ;
        RECT 72.595 -102.165 72.925 -101.835 ;
        RECT 72.595 -103.525 72.925 -103.195 ;
        RECT 72.595 -104.885 72.925 -104.555 ;
        RECT 72.595 -106.245 72.925 -105.915 ;
        RECT 72.595 -107.605 72.925 -107.275 ;
        RECT 72.595 -108.965 72.925 -108.635 ;
        RECT 72.595 -110.325 72.925 -109.995 ;
        RECT 72.595 -111.685 72.925 -111.355 ;
        RECT 72.595 -113.045 72.925 -112.715 ;
        RECT 72.595 -114.405 72.925 -114.075 ;
        RECT 72.595 -115.765 72.925 -115.435 ;
        RECT 72.595 -117.125 72.925 -116.795 ;
        RECT 72.595 -118.485 72.925 -118.155 ;
        RECT 72.595 -119.845 72.925 -119.515 ;
        RECT 72.595 -121.205 72.925 -120.875 ;
        RECT 72.595 -122.565 72.925 -122.235 ;
        RECT 72.595 -123.925 72.925 -123.595 ;
        RECT 72.595 -125.285 72.925 -124.955 ;
        RECT 72.595 -126.645 72.925 -126.315 ;
        RECT 72.595 -128.005 72.925 -127.675 ;
        RECT 72.595 -129.365 72.925 -129.035 ;
        RECT 72.595 -130.725 72.925 -130.395 ;
        RECT 72.595 -132.085 72.925 -131.755 ;
        RECT 72.595 -133.445 72.925 -133.115 ;
        RECT 72.595 -134.805 72.925 -134.475 ;
        RECT 72.595 -136.165 72.925 -135.835 ;
        RECT 72.595 -137.525 72.925 -137.195 ;
        RECT 72.595 -138.885 72.925 -138.555 ;
        RECT 72.595 -140.245 72.925 -139.915 ;
        RECT 72.595 -141.605 72.925 -141.275 ;
        RECT 72.595 -142.965 72.925 -142.635 ;
        RECT 72.595 -144.325 72.925 -143.995 ;
        RECT 72.595 -145.685 72.925 -145.355 ;
        RECT 72.595 -147.045 72.925 -146.715 ;
        RECT 72.595 -148.405 72.925 -148.075 ;
        RECT 72.595 -149.765 72.925 -149.435 ;
        RECT 72.595 -151.125 72.925 -150.795 ;
        RECT 72.595 -152.485 72.925 -152.155 ;
        RECT 72.595 -153.845 72.925 -153.515 ;
        RECT 72.595 -155.205 72.925 -154.875 ;
        RECT 72.595 -156.565 72.925 -156.235 ;
        RECT 72.595 -157.925 72.925 -157.595 ;
        RECT 72.595 -159.285 72.925 -158.955 ;
        RECT 72.595 -160.645 72.925 -160.315 ;
        RECT 72.595 -162.005 72.925 -161.675 ;
        RECT 72.595 -163.365 72.925 -163.035 ;
        RECT 72.595 -164.725 72.925 -164.395 ;
        RECT 72.595 -166.085 72.925 -165.755 ;
        RECT 72.595 -167.445 72.925 -167.115 ;
        RECT 72.595 -168.805 72.925 -168.475 ;
        RECT 72.595 -170.165 72.925 -169.835 ;
        RECT 72.595 -171.525 72.925 -171.195 ;
        RECT 72.595 -172.885 72.925 -172.555 ;
        RECT 72.595 -174.245 72.925 -173.915 ;
        RECT 72.595 -175.605 72.925 -175.275 ;
        RECT 72.595 -176.965 72.925 -176.635 ;
        RECT 72.595 -178.325 72.925 -177.995 ;
        RECT 72.595 -179.685 72.925 -179.355 ;
        RECT 72.595 -181.93 72.925 -180.8 ;
        RECT 72.6 -182.045 72.92 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 241.32 74.285 242.45 ;
        RECT 73.955 239.195 74.285 239.525 ;
        RECT 73.955 237.835 74.285 238.165 ;
        RECT 73.96 237.16 74.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 -1.525 74.285 -1.195 ;
        RECT 73.955 -2.885 74.285 -2.555 ;
        RECT 73.96 -3.56 74.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 73.955 -95.365 74.285 -95.035 ;
        RECT 73.955 -96.725 74.285 -96.395 ;
        RECT 73.955 -98.085 74.285 -97.755 ;
        RECT 73.955 -99.445 74.285 -99.115 ;
        RECT 73.955 -100.805 74.285 -100.475 ;
        RECT 73.955 -102.165 74.285 -101.835 ;
        RECT 73.955 -103.525 74.285 -103.195 ;
        RECT 73.955 -104.885 74.285 -104.555 ;
        RECT 73.955 -106.245 74.285 -105.915 ;
        RECT 73.955 -107.605 74.285 -107.275 ;
        RECT 73.955 -108.965 74.285 -108.635 ;
        RECT 73.955 -110.325 74.285 -109.995 ;
        RECT 73.955 -111.685 74.285 -111.355 ;
        RECT 73.955 -113.045 74.285 -112.715 ;
        RECT 73.955 -114.405 74.285 -114.075 ;
        RECT 73.955 -115.765 74.285 -115.435 ;
        RECT 73.955 -117.125 74.285 -116.795 ;
        RECT 73.955 -118.485 74.285 -118.155 ;
        RECT 73.955 -119.845 74.285 -119.515 ;
        RECT 73.955 -121.205 74.285 -120.875 ;
        RECT 73.955 -122.565 74.285 -122.235 ;
        RECT 73.955 -123.925 74.285 -123.595 ;
        RECT 73.955 -125.285 74.285 -124.955 ;
        RECT 73.955 -126.645 74.285 -126.315 ;
        RECT 73.955 -128.005 74.285 -127.675 ;
        RECT 73.955 -129.365 74.285 -129.035 ;
        RECT 73.955 -130.725 74.285 -130.395 ;
        RECT 73.955 -132.085 74.285 -131.755 ;
        RECT 73.955 -133.445 74.285 -133.115 ;
        RECT 73.955 -134.805 74.285 -134.475 ;
        RECT 73.955 -136.165 74.285 -135.835 ;
        RECT 73.955 -137.525 74.285 -137.195 ;
        RECT 73.955 -138.885 74.285 -138.555 ;
        RECT 73.955 -140.245 74.285 -139.915 ;
        RECT 73.955 -141.605 74.285 -141.275 ;
        RECT 73.955 -142.965 74.285 -142.635 ;
        RECT 73.955 -144.325 74.285 -143.995 ;
        RECT 73.955 -145.685 74.285 -145.355 ;
        RECT 73.955 -147.045 74.285 -146.715 ;
        RECT 73.955 -148.405 74.285 -148.075 ;
        RECT 73.955 -149.765 74.285 -149.435 ;
        RECT 73.955 -151.125 74.285 -150.795 ;
        RECT 73.955 -152.485 74.285 -152.155 ;
        RECT 73.955 -153.845 74.285 -153.515 ;
        RECT 73.955 -155.205 74.285 -154.875 ;
        RECT 73.955 -156.565 74.285 -156.235 ;
        RECT 73.955 -157.925 74.285 -157.595 ;
        RECT 73.955 -159.285 74.285 -158.955 ;
        RECT 73.955 -160.645 74.285 -160.315 ;
        RECT 73.955 -162.005 74.285 -161.675 ;
        RECT 73.955 -163.365 74.285 -163.035 ;
        RECT 73.955 -164.725 74.285 -164.395 ;
        RECT 73.955 -166.085 74.285 -165.755 ;
        RECT 73.955 -167.445 74.285 -167.115 ;
        RECT 73.955 -168.805 74.285 -168.475 ;
        RECT 73.955 -170.165 74.285 -169.835 ;
        RECT 73.955 -171.525 74.285 -171.195 ;
        RECT 73.955 -172.885 74.285 -172.555 ;
        RECT 73.955 -174.245 74.285 -173.915 ;
        RECT 73.955 -175.605 74.285 -175.275 ;
        RECT 73.955 -176.965 74.285 -176.635 ;
        RECT 73.955 -178.325 74.285 -177.995 ;
        RECT 73.955 -179.685 74.285 -179.355 ;
        RECT 73.955 -181.93 74.285 -180.8 ;
        RECT 73.96 -182.045 74.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 241.32 75.645 242.45 ;
        RECT 75.315 239.195 75.645 239.525 ;
        RECT 75.315 237.835 75.645 238.165 ;
        RECT 75.32 237.16 75.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 -1.525 75.645 -1.195 ;
        RECT 75.315 -2.885 75.645 -2.555 ;
        RECT 75.32 -3.56 75.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 75.315 -95.365 75.645 -95.035 ;
        RECT 75.315 -96.725 75.645 -96.395 ;
        RECT 75.315 -98.085 75.645 -97.755 ;
        RECT 75.315 -99.445 75.645 -99.115 ;
        RECT 75.315 -100.805 75.645 -100.475 ;
        RECT 75.315 -102.165 75.645 -101.835 ;
        RECT 75.315 -103.525 75.645 -103.195 ;
        RECT 75.315 -104.885 75.645 -104.555 ;
        RECT 75.315 -106.245 75.645 -105.915 ;
        RECT 75.315 -107.605 75.645 -107.275 ;
        RECT 75.315 -108.965 75.645 -108.635 ;
        RECT 75.315 -110.325 75.645 -109.995 ;
        RECT 75.315 -111.685 75.645 -111.355 ;
        RECT 75.315 -113.045 75.645 -112.715 ;
        RECT 75.315 -114.405 75.645 -114.075 ;
        RECT 75.315 -115.765 75.645 -115.435 ;
        RECT 75.315 -117.125 75.645 -116.795 ;
        RECT 75.315 -118.485 75.645 -118.155 ;
        RECT 75.315 -119.845 75.645 -119.515 ;
        RECT 75.315 -121.205 75.645 -120.875 ;
        RECT 75.315 -122.565 75.645 -122.235 ;
        RECT 75.315 -123.925 75.645 -123.595 ;
        RECT 75.315 -125.285 75.645 -124.955 ;
        RECT 75.315 -126.645 75.645 -126.315 ;
        RECT 75.315 -128.005 75.645 -127.675 ;
        RECT 75.315 -129.365 75.645 -129.035 ;
        RECT 75.315 -130.725 75.645 -130.395 ;
        RECT 75.315 -132.085 75.645 -131.755 ;
        RECT 75.315 -133.445 75.645 -133.115 ;
        RECT 75.315 -134.805 75.645 -134.475 ;
        RECT 75.315 -136.165 75.645 -135.835 ;
        RECT 75.315 -137.525 75.645 -137.195 ;
        RECT 75.315 -138.885 75.645 -138.555 ;
        RECT 75.315 -140.245 75.645 -139.915 ;
        RECT 75.315 -141.605 75.645 -141.275 ;
        RECT 75.315 -142.965 75.645 -142.635 ;
        RECT 75.315 -144.325 75.645 -143.995 ;
        RECT 75.315 -145.685 75.645 -145.355 ;
        RECT 75.315 -147.045 75.645 -146.715 ;
        RECT 75.315 -148.405 75.645 -148.075 ;
        RECT 75.315 -149.765 75.645 -149.435 ;
        RECT 75.315 -151.125 75.645 -150.795 ;
        RECT 75.315 -152.485 75.645 -152.155 ;
        RECT 75.315 -153.845 75.645 -153.515 ;
        RECT 75.315 -155.205 75.645 -154.875 ;
        RECT 75.315 -156.565 75.645 -156.235 ;
        RECT 75.315 -157.925 75.645 -157.595 ;
        RECT 75.315 -159.285 75.645 -158.955 ;
        RECT 75.315 -160.645 75.645 -160.315 ;
        RECT 75.315 -162.005 75.645 -161.675 ;
        RECT 75.315 -163.365 75.645 -163.035 ;
        RECT 75.315 -164.725 75.645 -164.395 ;
        RECT 75.315 -166.085 75.645 -165.755 ;
        RECT 75.315 -167.445 75.645 -167.115 ;
        RECT 75.315 -168.805 75.645 -168.475 ;
        RECT 75.315 -170.165 75.645 -169.835 ;
        RECT 75.315 -171.525 75.645 -171.195 ;
        RECT 75.315 -172.885 75.645 -172.555 ;
        RECT 75.315 -174.245 75.645 -173.915 ;
        RECT 75.315 -175.605 75.645 -175.275 ;
        RECT 75.315 -176.965 75.645 -176.635 ;
        RECT 75.315 -178.325 75.645 -177.995 ;
        RECT 75.315 -179.685 75.645 -179.355 ;
        RECT 75.315 -181.93 75.645 -180.8 ;
        RECT 75.32 -182.045 75.64 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.675 241.32 77.005 242.45 ;
        RECT 76.675 239.195 77.005 239.525 ;
        RECT 76.675 237.835 77.005 238.165 ;
        RECT 76.68 237.16 77 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.675 -1.525 77.005 -1.195 ;
        RECT 76.675 -2.885 77.005 -2.555 ;
        RECT 76.68 -3.56 77 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 76.675 -95.365 77.005 -95.035 ;
        RECT 76.675 -96.725 77.005 -96.395 ;
        RECT 76.675 -98.085 77.005 -97.755 ;
        RECT 76.675 -99.445 77.005 -99.115 ;
        RECT 76.675 -100.805 77.005 -100.475 ;
        RECT 76.675 -102.165 77.005 -101.835 ;
        RECT 76.675 -103.525 77.005 -103.195 ;
        RECT 76.675 -104.885 77.005 -104.555 ;
        RECT 76.675 -106.245 77.005 -105.915 ;
        RECT 76.675 -107.605 77.005 -107.275 ;
        RECT 76.675 -108.965 77.005 -108.635 ;
        RECT 76.675 -110.325 77.005 -109.995 ;
        RECT 76.675 -111.685 77.005 -111.355 ;
        RECT 76.675 -113.045 77.005 -112.715 ;
        RECT 76.675 -114.405 77.005 -114.075 ;
        RECT 76.675 -115.765 77.005 -115.435 ;
        RECT 76.675 -117.125 77.005 -116.795 ;
        RECT 76.675 -118.485 77.005 -118.155 ;
        RECT 76.675 -119.845 77.005 -119.515 ;
        RECT 76.675 -121.205 77.005 -120.875 ;
        RECT 76.675 -122.565 77.005 -122.235 ;
        RECT 76.675 -123.925 77.005 -123.595 ;
        RECT 76.675 -125.285 77.005 -124.955 ;
        RECT 76.675 -126.645 77.005 -126.315 ;
        RECT 76.675 -128.005 77.005 -127.675 ;
        RECT 76.675 -129.365 77.005 -129.035 ;
        RECT 76.675 -130.725 77.005 -130.395 ;
        RECT 76.675 -132.085 77.005 -131.755 ;
        RECT 76.675 -133.445 77.005 -133.115 ;
        RECT 76.675 -134.805 77.005 -134.475 ;
        RECT 76.675 -136.165 77.005 -135.835 ;
        RECT 76.675 -137.525 77.005 -137.195 ;
        RECT 76.675 -138.885 77.005 -138.555 ;
        RECT 76.675 -140.245 77.005 -139.915 ;
        RECT 76.675 -141.605 77.005 -141.275 ;
        RECT 76.675 -142.965 77.005 -142.635 ;
        RECT 76.675 -144.325 77.005 -143.995 ;
        RECT 76.675 -145.685 77.005 -145.355 ;
        RECT 76.675 -147.045 77.005 -146.715 ;
        RECT 76.675 -148.405 77.005 -148.075 ;
        RECT 76.675 -149.765 77.005 -149.435 ;
        RECT 76.675 -151.125 77.005 -150.795 ;
        RECT 76.675 -152.485 77.005 -152.155 ;
        RECT 76.675 -153.845 77.005 -153.515 ;
        RECT 76.675 -155.205 77.005 -154.875 ;
        RECT 76.675 -156.565 77.005 -156.235 ;
        RECT 76.675 -157.925 77.005 -157.595 ;
        RECT 76.675 -159.285 77.005 -158.955 ;
        RECT 76.675 -160.645 77.005 -160.315 ;
        RECT 76.675 -162.005 77.005 -161.675 ;
        RECT 76.675 -163.365 77.005 -163.035 ;
        RECT 76.675 -164.725 77.005 -164.395 ;
        RECT 76.675 -166.085 77.005 -165.755 ;
        RECT 76.675 -167.445 77.005 -167.115 ;
        RECT 76.675 -168.805 77.005 -168.475 ;
        RECT 76.675 -170.165 77.005 -169.835 ;
        RECT 76.675 -171.525 77.005 -171.195 ;
        RECT 76.675 -172.885 77.005 -172.555 ;
        RECT 76.675 -174.245 77.005 -173.915 ;
        RECT 76.675 -175.605 77.005 -175.275 ;
        RECT 76.675 -176.965 77.005 -176.635 ;
        RECT 76.675 -178.325 77.005 -177.995 ;
        RECT 76.675 -179.685 77.005 -179.355 ;
        RECT 76.675 -181.93 77.005 -180.8 ;
        RECT 76.68 -182.045 77 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 241.32 78.365 242.45 ;
        RECT 78.035 239.195 78.365 239.525 ;
        RECT 78.035 237.835 78.365 238.165 ;
        RECT 78.04 237.16 78.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 -1.525 78.365 -1.195 ;
        RECT 78.035 -2.885 78.365 -2.555 ;
        RECT 78.04 -3.56 78.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 78.035 -95.365 78.365 -95.035 ;
        RECT 78.035 -96.725 78.365 -96.395 ;
        RECT 78.035 -98.085 78.365 -97.755 ;
        RECT 78.035 -99.445 78.365 -99.115 ;
        RECT 78.035 -100.805 78.365 -100.475 ;
        RECT 78.035 -102.165 78.365 -101.835 ;
        RECT 78.035 -103.525 78.365 -103.195 ;
        RECT 78.035 -104.885 78.365 -104.555 ;
        RECT 78.035 -106.245 78.365 -105.915 ;
        RECT 78.035 -107.605 78.365 -107.275 ;
        RECT 78.035 -108.965 78.365 -108.635 ;
        RECT 78.035 -110.325 78.365 -109.995 ;
        RECT 78.035 -111.685 78.365 -111.355 ;
        RECT 78.035 -113.045 78.365 -112.715 ;
        RECT 78.035 -114.405 78.365 -114.075 ;
        RECT 78.035 -115.765 78.365 -115.435 ;
        RECT 78.035 -117.125 78.365 -116.795 ;
        RECT 78.035 -118.485 78.365 -118.155 ;
        RECT 78.035 -119.845 78.365 -119.515 ;
        RECT 78.035 -121.205 78.365 -120.875 ;
        RECT 78.035 -122.565 78.365 -122.235 ;
        RECT 78.035 -123.925 78.365 -123.595 ;
        RECT 78.035 -125.285 78.365 -124.955 ;
        RECT 78.035 -126.645 78.365 -126.315 ;
        RECT 78.035 -128.005 78.365 -127.675 ;
        RECT 78.035 -129.365 78.365 -129.035 ;
        RECT 78.035 -130.725 78.365 -130.395 ;
        RECT 78.035 -132.085 78.365 -131.755 ;
        RECT 78.035 -133.445 78.365 -133.115 ;
        RECT 78.035 -134.805 78.365 -134.475 ;
        RECT 78.035 -136.165 78.365 -135.835 ;
        RECT 78.035 -137.525 78.365 -137.195 ;
        RECT 78.035 -138.885 78.365 -138.555 ;
        RECT 78.035 -140.245 78.365 -139.915 ;
        RECT 78.035 -141.605 78.365 -141.275 ;
        RECT 78.035 -142.965 78.365 -142.635 ;
        RECT 78.035 -144.325 78.365 -143.995 ;
        RECT 78.035 -145.685 78.365 -145.355 ;
        RECT 78.035 -147.045 78.365 -146.715 ;
        RECT 78.035 -148.405 78.365 -148.075 ;
        RECT 78.035 -149.765 78.365 -149.435 ;
        RECT 78.035 -151.125 78.365 -150.795 ;
        RECT 78.035 -152.485 78.365 -152.155 ;
        RECT 78.035 -153.845 78.365 -153.515 ;
        RECT 78.035 -155.205 78.365 -154.875 ;
        RECT 78.035 -156.565 78.365 -156.235 ;
        RECT 78.035 -157.925 78.365 -157.595 ;
        RECT 78.035 -159.285 78.365 -158.955 ;
        RECT 78.035 -160.645 78.365 -160.315 ;
        RECT 78.035 -162.005 78.365 -161.675 ;
        RECT 78.035 -163.365 78.365 -163.035 ;
        RECT 78.035 -164.725 78.365 -164.395 ;
        RECT 78.035 -166.085 78.365 -165.755 ;
        RECT 78.035 -167.445 78.365 -167.115 ;
        RECT 78.035 -168.805 78.365 -168.475 ;
        RECT 78.035 -170.165 78.365 -169.835 ;
        RECT 78.035 -171.525 78.365 -171.195 ;
        RECT 78.035 -172.885 78.365 -172.555 ;
        RECT 78.035 -174.245 78.365 -173.915 ;
        RECT 78.035 -175.605 78.365 -175.275 ;
        RECT 78.035 -176.965 78.365 -176.635 ;
        RECT 78.035 -178.325 78.365 -177.995 ;
        RECT 78.035 -179.685 78.365 -179.355 ;
        RECT 78.035 -181.93 78.365 -180.8 ;
        RECT 78.04 -182.045 78.36 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 241.32 79.725 242.45 ;
        RECT 79.395 239.195 79.725 239.525 ;
        RECT 79.395 237.835 79.725 238.165 ;
        RECT 79.4 237.16 79.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.395 -99.445 79.725 -99.115 ;
        RECT 79.395 -100.805 79.725 -100.475 ;
        RECT 79.395 -102.165 79.725 -101.835 ;
        RECT 79.395 -103.525 79.725 -103.195 ;
        RECT 79.395 -104.885 79.725 -104.555 ;
        RECT 79.395 -106.245 79.725 -105.915 ;
        RECT 79.395 -107.605 79.725 -107.275 ;
        RECT 79.395 -108.965 79.725 -108.635 ;
        RECT 79.395 -110.325 79.725 -109.995 ;
        RECT 79.395 -111.685 79.725 -111.355 ;
        RECT 79.395 -113.045 79.725 -112.715 ;
        RECT 79.395 -114.405 79.725 -114.075 ;
        RECT 79.395 -115.765 79.725 -115.435 ;
        RECT 79.395 -117.125 79.725 -116.795 ;
        RECT 79.395 -118.485 79.725 -118.155 ;
        RECT 79.395 -119.845 79.725 -119.515 ;
        RECT 79.395 -121.205 79.725 -120.875 ;
        RECT 79.395 -122.565 79.725 -122.235 ;
        RECT 79.395 -123.925 79.725 -123.595 ;
        RECT 79.395 -125.285 79.725 -124.955 ;
        RECT 79.395 -126.645 79.725 -126.315 ;
        RECT 79.395 -128.005 79.725 -127.675 ;
        RECT 79.395 -129.365 79.725 -129.035 ;
        RECT 79.395 -130.725 79.725 -130.395 ;
        RECT 79.395 -132.085 79.725 -131.755 ;
        RECT 79.395 -133.445 79.725 -133.115 ;
        RECT 79.395 -134.805 79.725 -134.475 ;
        RECT 79.395 -136.165 79.725 -135.835 ;
        RECT 79.395 -137.525 79.725 -137.195 ;
        RECT 79.395 -138.885 79.725 -138.555 ;
        RECT 79.395 -140.245 79.725 -139.915 ;
        RECT 79.395 -141.605 79.725 -141.275 ;
        RECT 79.395 -142.965 79.725 -142.635 ;
        RECT 79.395 -144.325 79.725 -143.995 ;
        RECT 79.395 -145.685 79.725 -145.355 ;
        RECT 79.395 -147.045 79.725 -146.715 ;
        RECT 79.395 -148.405 79.725 -148.075 ;
        RECT 79.395 -149.765 79.725 -149.435 ;
        RECT 79.395 -151.125 79.725 -150.795 ;
        RECT 79.395 -152.485 79.725 -152.155 ;
        RECT 79.395 -153.845 79.725 -153.515 ;
        RECT 79.395 -155.205 79.725 -154.875 ;
        RECT 79.395 -156.565 79.725 -156.235 ;
        RECT 79.395 -157.925 79.725 -157.595 ;
        RECT 79.395 -159.285 79.725 -158.955 ;
        RECT 79.395 -160.645 79.725 -160.315 ;
        RECT 79.395 -162.005 79.725 -161.675 ;
        RECT 79.395 -163.365 79.725 -163.035 ;
        RECT 79.395 -164.725 79.725 -164.395 ;
        RECT 79.395 -166.085 79.725 -165.755 ;
        RECT 79.395 -167.445 79.725 -167.115 ;
        RECT 79.395 -168.805 79.725 -168.475 ;
        RECT 79.395 -170.165 79.725 -169.835 ;
        RECT 79.395 -171.525 79.725 -171.195 ;
        RECT 79.395 -172.885 79.725 -172.555 ;
        RECT 79.395 -174.245 79.725 -173.915 ;
        RECT 79.395 -175.605 79.725 -175.275 ;
        RECT 79.395 -176.965 79.725 -176.635 ;
        RECT 79.395 -178.325 79.725 -177.995 ;
        RECT 79.395 -179.685 79.725 -179.355 ;
        RECT 79.395 -181.93 79.725 -180.8 ;
        RECT 79.4 -182.045 79.72 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 79.61 -98.075 79.94 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 241.32 81.085 242.45 ;
        RECT 80.755 239.195 81.085 239.525 ;
        RECT 80.755 237.835 81.085 238.165 ;
        RECT 80.76 237.16 81.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 80.755 -1.525 81.085 -1.195 ;
        RECT 80.755 -2.885 81.085 -2.555 ;
        RECT 80.76 -3.56 81.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 241.32 82.445 242.45 ;
        RECT 82.115 239.195 82.445 239.525 ;
        RECT 82.115 237.835 82.445 238.165 ;
        RECT 82.12 237.16 82.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 82.115 -1.525 82.445 -1.195 ;
        RECT 82.115 -2.885 82.445 -2.555 ;
        RECT 82.12 -3.56 82.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 241.32 83.805 242.45 ;
        RECT 83.475 239.195 83.805 239.525 ;
        RECT 83.475 237.835 83.805 238.165 ;
        RECT 83.48 237.16 83.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 -1.525 83.805 -1.195 ;
        RECT 83.475 -2.885 83.805 -2.555 ;
        RECT 83.48 -3.56 83.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 83.475 -95.365 83.805 -95.035 ;
        RECT 83.475 -96.725 83.805 -96.395 ;
        RECT 83.475 -98.085 83.805 -97.755 ;
        RECT 83.475 -99.445 83.805 -99.115 ;
        RECT 83.475 -100.805 83.805 -100.475 ;
        RECT 83.475 -102.165 83.805 -101.835 ;
        RECT 83.475 -103.525 83.805 -103.195 ;
        RECT 83.475 -104.885 83.805 -104.555 ;
        RECT 83.475 -106.245 83.805 -105.915 ;
        RECT 83.475 -107.605 83.805 -107.275 ;
        RECT 83.475 -108.965 83.805 -108.635 ;
        RECT 83.475 -110.325 83.805 -109.995 ;
        RECT 83.475 -111.685 83.805 -111.355 ;
        RECT 83.475 -113.045 83.805 -112.715 ;
        RECT 83.475 -114.405 83.805 -114.075 ;
        RECT 83.475 -115.765 83.805 -115.435 ;
        RECT 83.475 -117.125 83.805 -116.795 ;
        RECT 83.475 -118.485 83.805 -118.155 ;
        RECT 83.475 -119.845 83.805 -119.515 ;
        RECT 83.475 -121.205 83.805 -120.875 ;
        RECT 83.475 -122.565 83.805 -122.235 ;
        RECT 83.475 -123.925 83.805 -123.595 ;
        RECT 83.475 -125.285 83.805 -124.955 ;
        RECT 83.475 -126.645 83.805 -126.315 ;
        RECT 83.475 -128.005 83.805 -127.675 ;
        RECT 83.475 -129.365 83.805 -129.035 ;
        RECT 83.475 -130.725 83.805 -130.395 ;
        RECT 83.475 -132.085 83.805 -131.755 ;
        RECT 83.475 -133.445 83.805 -133.115 ;
        RECT 83.475 -134.805 83.805 -134.475 ;
        RECT 83.475 -136.165 83.805 -135.835 ;
        RECT 83.475 -137.525 83.805 -137.195 ;
        RECT 83.475 -138.885 83.805 -138.555 ;
        RECT 83.475 -140.245 83.805 -139.915 ;
        RECT 83.475 -141.605 83.805 -141.275 ;
        RECT 83.475 -142.965 83.805 -142.635 ;
        RECT 83.475 -144.325 83.805 -143.995 ;
        RECT 83.475 -145.685 83.805 -145.355 ;
        RECT 83.475 -147.045 83.805 -146.715 ;
        RECT 83.475 -148.405 83.805 -148.075 ;
        RECT 83.475 -149.765 83.805 -149.435 ;
        RECT 83.475 -151.125 83.805 -150.795 ;
        RECT 83.475 -152.485 83.805 -152.155 ;
        RECT 83.475 -153.845 83.805 -153.515 ;
        RECT 83.475 -155.205 83.805 -154.875 ;
        RECT 83.475 -156.565 83.805 -156.235 ;
        RECT 83.475 -157.925 83.805 -157.595 ;
        RECT 83.475 -159.285 83.805 -158.955 ;
        RECT 83.475 -160.645 83.805 -160.315 ;
        RECT 83.475 -162.005 83.805 -161.675 ;
        RECT 83.475 -163.365 83.805 -163.035 ;
        RECT 83.475 -164.725 83.805 -164.395 ;
        RECT 83.475 -166.085 83.805 -165.755 ;
        RECT 83.475 -167.445 83.805 -167.115 ;
        RECT 83.475 -168.805 83.805 -168.475 ;
        RECT 83.475 -170.165 83.805 -169.835 ;
        RECT 83.475 -171.525 83.805 -171.195 ;
        RECT 83.475 -172.885 83.805 -172.555 ;
        RECT 83.475 -174.245 83.805 -173.915 ;
        RECT 83.475 -175.605 83.805 -175.275 ;
        RECT 83.475 -176.965 83.805 -176.635 ;
        RECT 83.475 -178.325 83.805 -177.995 ;
        RECT 83.475 -179.685 83.805 -179.355 ;
        RECT 83.475 -181.93 83.805 -180.8 ;
        RECT 83.48 -182.045 83.8 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 241.32 85.165 242.45 ;
        RECT 84.835 239.195 85.165 239.525 ;
        RECT 84.835 237.835 85.165 238.165 ;
        RECT 84.84 237.16 85.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 -1.525 85.165 -1.195 ;
        RECT 84.835 -2.885 85.165 -2.555 ;
        RECT 84.84 -3.56 85.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 84.835 -95.365 85.165 -95.035 ;
        RECT 84.835 -96.725 85.165 -96.395 ;
        RECT 84.835 -98.085 85.165 -97.755 ;
        RECT 84.835 -99.445 85.165 -99.115 ;
        RECT 84.835 -100.805 85.165 -100.475 ;
        RECT 84.835 -102.165 85.165 -101.835 ;
        RECT 84.835 -103.525 85.165 -103.195 ;
        RECT 84.835 -104.885 85.165 -104.555 ;
        RECT 84.835 -106.245 85.165 -105.915 ;
        RECT 84.835 -107.605 85.165 -107.275 ;
        RECT 84.835 -108.965 85.165 -108.635 ;
        RECT 84.835 -110.325 85.165 -109.995 ;
        RECT 84.835 -111.685 85.165 -111.355 ;
        RECT 84.835 -113.045 85.165 -112.715 ;
        RECT 84.835 -114.405 85.165 -114.075 ;
        RECT 84.835 -115.765 85.165 -115.435 ;
        RECT 84.835 -117.125 85.165 -116.795 ;
        RECT 84.835 -118.485 85.165 -118.155 ;
        RECT 84.835 -119.845 85.165 -119.515 ;
        RECT 84.835 -121.205 85.165 -120.875 ;
        RECT 84.835 -122.565 85.165 -122.235 ;
        RECT 84.835 -123.925 85.165 -123.595 ;
        RECT 84.835 -125.285 85.165 -124.955 ;
        RECT 84.835 -126.645 85.165 -126.315 ;
        RECT 84.835 -128.005 85.165 -127.675 ;
        RECT 84.835 -129.365 85.165 -129.035 ;
        RECT 84.835 -130.725 85.165 -130.395 ;
        RECT 84.835 -132.085 85.165 -131.755 ;
        RECT 84.835 -133.445 85.165 -133.115 ;
        RECT 84.835 -134.805 85.165 -134.475 ;
        RECT 84.835 -136.165 85.165 -135.835 ;
        RECT 84.835 -137.525 85.165 -137.195 ;
        RECT 84.835 -138.885 85.165 -138.555 ;
        RECT 84.835 -140.245 85.165 -139.915 ;
        RECT 84.835 -141.605 85.165 -141.275 ;
        RECT 84.835 -142.965 85.165 -142.635 ;
        RECT 84.835 -144.325 85.165 -143.995 ;
        RECT 84.835 -145.685 85.165 -145.355 ;
        RECT 84.835 -147.045 85.165 -146.715 ;
        RECT 84.835 -148.405 85.165 -148.075 ;
        RECT 84.835 -149.765 85.165 -149.435 ;
        RECT 84.835 -151.125 85.165 -150.795 ;
        RECT 84.835 -152.485 85.165 -152.155 ;
        RECT 84.835 -153.845 85.165 -153.515 ;
        RECT 84.835 -155.205 85.165 -154.875 ;
        RECT 84.835 -156.565 85.165 -156.235 ;
        RECT 84.835 -157.925 85.165 -157.595 ;
        RECT 84.835 -159.285 85.165 -158.955 ;
        RECT 84.835 -160.645 85.165 -160.315 ;
        RECT 84.835 -162.005 85.165 -161.675 ;
        RECT 84.835 -163.365 85.165 -163.035 ;
        RECT 84.835 -164.725 85.165 -164.395 ;
        RECT 84.835 -166.085 85.165 -165.755 ;
        RECT 84.835 -167.445 85.165 -167.115 ;
        RECT 84.835 -168.805 85.165 -168.475 ;
        RECT 84.835 -170.165 85.165 -169.835 ;
        RECT 84.835 -171.525 85.165 -171.195 ;
        RECT 84.835 -172.885 85.165 -172.555 ;
        RECT 84.835 -174.245 85.165 -173.915 ;
        RECT 84.835 -175.605 85.165 -175.275 ;
        RECT 84.835 -176.965 85.165 -176.635 ;
        RECT 84.835 -178.325 85.165 -177.995 ;
        RECT 84.835 -179.685 85.165 -179.355 ;
        RECT 84.835 -181.93 85.165 -180.8 ;
        RECT 84.84 -182.045 85.16 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 241.32 86.525 242.45 ;
        RECT 86.195 239.195 86.525 239.525 ;
        RECT 86.195 237.835 86.525 238.165 ;
        RECT 86.2 237.16 86.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 -1.525 86.525 -1.195 ;
        RECT 86.195 -2.885 86.525 -2.555 ;
        RECT 86.2 -3.56 86.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 86.195 -95.365 86.525 -95.035 ;
        RECT 86.195 -96.725 86.525 -96.395 ;
        RECT 86.195 -98.085 86.525 -97.755 ;
        RECT 86.195 -99.445 86.525 -99.115 ;
        RECT 86.195 -100.805 86.525 -100.475 ;
        RECT 86.195 -102.165 86.525 -101.835 ;
        RECT 86.195 -103.525 86.525 -103.195 ;
        RECT 86.195 -104.885 86.525 -104.555 ;
        RECT 86.195 -106.245 86.525 -105.915 ;
        RECT 86.195 -107.605 86.525 -107.275 ;
        RECT 86.195 -108.965 86.525 -108.635 ;
        RECT 86.195 -110.325 86.525 -109.995 ;
        RECT 86.195 -111.685 86.525 -111.355 ;
        RECT 86.195 -113.045 86.525 -112.715 ;
        RECT 86.195 -114.405 86.525 -114.075 ;
        RECT 86.195 -115.765 86.525 -115.435 ;
        RECT 86.195 -117.125 86.525 -116.795 ;
        RECT 86.195 -118.485 86.525 -118.155 ;
        RECT 86.195 -119.845 86.525 -119.515 ;
        RECT 86.195 -121.205 86.525 -120.875 ;
        RECT 86.195 -122.565 86.525 -122.235 ;
        RECT 86.195 -123.925 86.525 -123.595 ;
        RECT 86.195 -125.285 86.525 -124.955 ;
        RECT 86.195 -126.645 86.525 -126.315 ;
        RECT 86.195 -128.005 86.525 -127.675 ;
        RECT 86.195 -129.365 86.525 -129.035 ;
        RECT 86.195 -130.725 86.525 -130.395 ;
        RECT 86.195 -132.085 86.525 -131.755 ;
        RECT 86.195 -133.445 86.525 -133.115 ;
        RECT 86.195 -134.805 86.525 -134.475 ;
        RECT 86.195 -136.165 86.525 -135.835 ;
        RECT 86.195 -137.525 86.525 -137.195 ;
        RECT 86.195 -138.885 86.525 -138.555 ;
        RECT 86.195 -140.245 86.525 -139.915 ;
        RECT 86.195 -141.605 86.525 -141.275 ;
        RECT 86.195 -142.965 86.525 -142.635 ;
        RECT 86.195 -144.325 86.525 -143.995 ;
        RECT 86.195 -145.685 86.525 -145.355 ;
        RECT 86.195 -147.045 86.525 -146.715 ;
        RECT 86.195 -148.405 86.525 -148.075 ;
        RECT 86.195 -149.765 86.525 -149.435 ;
        RECT 86.195 -151.125 86.525 -150.795 ;
        RECT 86.195 -152.485 86.525 -152.155 ;
        RECT 86.195 -153.845 86.525 -153.515 ;
        RECT 86.195 -155.205 86.525 -154.875 ;
        RECT 86.195 -156.565 86.525 -156.235 ;
        RECT 86.195 -157.925 86.525 -157.595 ;
        RECT 86.195 -159.285 86.525 -158.955 ;
        RECT 86.195 -160.645 86.525 -160.315 ;
        RECT 86.195 -162.005 86.525 -161.675 ;
        RECT 86.195 -163.365 86.525 -163.035 ;
        RECT 86.195 -164.725 86.525 -164.395 ;
        RECT 86.195 -166.085 86.525 -165.755 ;
        RECT 86.195 -167.445 86.525 -167.115 ;
        RECT 86.195 -168.805 86.525 -168.475 ;
        RECT 86.195 -170.165 86.525 -169.835 ;
        RECT 86.195 -171.525 86.525 -171.195 ;
        RECT 86.195 -172.885 86.525 -172.555 ;
        RECT 86.195 -174.245 86.525 -173.915 ;
        RECT 86.195 -175.605 86.525 -175.275 ;
        RECT 86.195 -176.965 86.525 -176.635 ;
        RECT 86.195 -178.325 86.525 -177.995 ;
        RECT 86.195 -179.685 86.525 -179.355 ;
        RECT 86.195 -181.93 86.525 -180.8 ;
        RECT 86.2 -182.045 86.52 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 241.32 87.885 242.45 ;
        RECT 87.555 239.195 87.885 239.525 ;
        RECT 87.555 237.835 87.885 238.165 ;
        RECT 87.56 237.16 87.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 -1.525 87.885 -1.195 ;
        RECT 87.555 -2.885 87.885 -2.555 ;
        RECT 87.56 -3.56 87.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 87.555 -95.365 87.885 -95.035 ;
        RECT 87.555 -96.725 87.885 -96.395 ;
        RECT 87.555 -98.085 87.885 -97.755 ;
        RECT 87.555 -99.445 87.885 -99.115 ;
        RECT 87.555 -100.805 87.885 -100.475 ;
        RECT 87.555 -102.165 87.885 -101.835 ;
        RECT 87.555 -103.525 87.885 -103.195 ;
        RECT 87.555 -104.885 87.885 -104.555 ;
        RECT 87.555 -106.245 87.885 -105.915 ;
        RECT 87.555 -107.605 87.885 -107.275 ;
        RECT 87.555 -108.965 87.885 -108.635 ;
        RECT 87.555 -110.325 87.885 -109.995 ;
        RECT 87.555 -111.685 87.885 -111.355 ;
        RECT 87.555 -113.045 87.885 -112.715 ;
        RECT 87.555 -114.405 87.885 -114.075 ;
        RECT 87.555 -115.765 87.885 -115.435 ;
        RECT 87.555 -117.125 87.885 -116.795 ;
        RECT 87.555 -118.485 87.885 -118.155 ;
        RECT 87.555 -119.845 87.885 -119.515 ;
        RECT 87.555 -121.205 87.885 -120.875 ;
        RECT 87.555 -122.565 87.885 -122.235 ;
        RECT 87.555 -123.925 87.885 -123.595 ;
        RECT 87.555 -125.285 87.885 -124.955 ;
        RECT 87.555 -126.645 87.885 -126.315 ;
        RECT 87.555 -128.005 87.885 -127.675 ;
        RECT 87.555 -129.365 87.885 -129.035 ;
        RECT 87.555 -130.725 87.885 -130.395 ;
        RECT 87.555 -132.085 87.885 -131.755 ;
        RECT 87.555 -133.445 87.885 -133.115 ;
        RECT 87.555 -134.805 87.885 -134.475 ;
        RECT 87.555 -136.165 87.885 -135.835 ;
        RECT 87.555 -137.525 87.885 -137.195 ;
        RECT 87.555 -138.885 87.885 -138.555 ;
        RECT 87.555 -140.245 87.885 -139.915 ;
        RECT 87.555 -141.605 87.885 -141.275 ;
        RECT 87.555 -142.965 87.885 -142.635 ;
        RECT 87.555 -144.325 87.885 -143.995 ;
        RECT 87.555 -145.685 87.885 -145.355 ;
        RECT 87.555 -147.045 87.885 -146.715 ;
        RECT 87.555 -148.405 87.885 -148.075 ;
        RECT 87.555 -149.765 87.885 -149.435 ;
        RECT 87.555 -151.125 87.885 -150.795 ;
        RECT 87.555 -152.485 87.885 -152.155 ;
        RECT 87.555 -153.845 87.885 -153.515 ;
        RECT 87.555 -155.205 87.885 -154.875 ;
        RECT 87.555 -156.565 87.885 -156.235 ;
        RECT 87.555 -157.925 87.885 -157.595 ;
        RECT 87.555 -159.285 87.885 -158.955 ;
        RECT 87.555 -160.645 87.885 -160.315 ;
        RECT 87.555 -162.005 87.885 -161.675 ;
        RECT 87.555 -163.365 87.885 -163.035 ;
        RECT 87.555 -164.725 87.885 -164.395 ;
        RECT 87.555 -166.085 87.885 -165.755 ;
        RECT 87.555 -167.445 87.885 -167.115 ;
        RECT 87.555 -168.805 87.885 -168.475 ;
        RECT 87.555 -170.165 87.885 -169.835 ;
        RECT 87.555 -171.525 87.885 -171.195 ;
        RECT 87.555 -172.885 87.885 -172.555 ;
        RECT 87.555 -174.245 87.885 -173.915 ;
        RECT 87.555 -175.605 87.885 -175.275 ;
        RECT 87.555 -176.965 87.885 -176.635 ;
        RECT 87.555 -178.325 87.885 -177.995 ;
        RECT 87.555 -179.685 87.885 -179.355 ;
        RECT 87.555 -181.93 87.885 -180.8 ;
        RECT 87.56 -182.045 87.88 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.915 241.32 89.245 242.45 ;
        RECT 88.915 239.195 89.245 239.525 ;
        RECT 88.915 237.835 89.245 238.165 ;
        RECT 88.92 237.16 89.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.915 -1.525 89.245 -1.195 ;
        RECT 88.915 -2.885 89.245 -2.555 ;
        RECT 88.92 -3.56 89.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 88.915 -95.365 89.245 -95.035 ;
        RECT 88.915 -96.725 89.245 -96.395 ;
        RECT 88.915 -98.085 89.245 -97.755 ;
        RECT 88.915 -99.445 89.245 -99.115 ;
        RECT 88.915 -100.805 89.245 -100.475 ;
        RECT 88.915 -102.165 89.245 -101.835 ;
        RECT 88.915 -103.525 89.245 -103.195 ;
        RECT 88.915 -104.885 89.245 -104.555 ;
        RECT 88.915 -106.245 89.245 -105.915 ;
        RECT 88.915 -107.605 89.245 -107.275 ;
        RECT 88.915 -108.965 89.245 -108.635 ;
        RECT 88.915 -110.325 89.245 -109.995 ;
        RECT 88.915 -111.685 89.245 -111.355 ;
        RECT 88.915 -113.045 89.245 -112.715 ;
        RECT 88.915 -114.405 89.245 -114.075 ;
        RECT 88.915 -115.765 89.245 -115.435 ;
        RECT 88.915 -117.125 89.245 -116.795 ;
        RECT 88.915 -118.485 89.245 -118.155 ;
        RECT 88.915 -119.845 89.245 -119.515 ;
        RECT 88.915 -121.205 89.245 -120.875 ;
        RECT 88.915 -122.565 89.245 -122.235 ;
        RECT 88.915 -123.925 89.245 -123.595 ;
        RECT 88.915 -125.285 89.245 -124.955 ;
        RECT 88.915 -126.645 89.245 -126.315 ;
        RECT 88.915 -128.005 89.245 -127.675 ;
        RECT 88.915 -129.365 89.245 -129.035 ;
        RECT 88.915 -130.725 89.245 -130.395 ;
        RECT 88.915 -132.085 89.245 -131.755 ;
        RECT 88.915 -133.445 89.245 -133.115 ;
        RECT 88.915 -134.805 89.245 -134.475 ;
        RECT 88.915 -136.165 89.245 -135.835 ;
        RECT 88.915 -137.525 89.245 -137.195 ;
        RECT 88.915 -138.885 89.245 -138.555 ;
        RECT 88.915 -140.245 89.245 -139.915 ;
        RECT 88.915 -141.605 89.245 -141.275 ;
        RECT 88.915 -142.965 89.245 -142.635 ;
        RECT 88.915 -144.325 89.245 -143.995 ;
        RECT 88.915 -145.685 89.245 -145.355 ;
        RECT 88.915 -147.045 89.245 -146.715 ;
        RECT 88.915 -148.405 89.245 -148.075 ;
        RECT 88.915 -149.765 89.245 -149.435 ;
        RECT 88.915 -151.125 89.245 -150.795 ;
        RECT 88.915 -152.485 89.245 -152.155 ;
        RECT 88.915 -153.845 89.245 -153.515 ;
        RECT 88.915 -155.205 89.245 -154.875 ;
        RECT 88.915 -156.565 89.245 -156.235 ;
        RECT 88.915 -157.925 89.245 -157.595 ;
        RECT 88.915 -159.285 89.245 -158.955 ;
        RECT 88.915 -160.645 89.245 -160.315 ;
        RECT 88.915 -162.005 89.245 -161.675 ;
        RECT 88.915 -163.365 89.245 -163.035 ;
        RECT 88.915 -164.725 89.245 -164.395 ;
        RECT 88.915 -166.085 89.245 -165.755 ;
        RECT 88.915 -167.445 89.245 -167.115 ;
        RECT 88.915 -168.805 89.245 -168.475 ;
        RECT 88.915 -170.165 89.245 -169.835 ;
        RECT 88.915 -171.525 89.245 -171.195 ;
        RECT 88.915 -172.885 89.245 -172.555 ;
        RECT 88.915 -174.245 89.245 -173.915 ;
        RECT 88.915 -175.605 89.245 -175.275 ;
        RECT 88.915 -176.965 89.245 -176.635 ;
        RECT 88.915 -178.325 89.245 -177.995 ;
        RECT 88.915 -179.685 89.245 -179.355 ;
        RECT 88.915 -181.93 89.245 -180.8 ;
        RECT 88.92 -182.045 89.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 241.32 90.605 242.45 ;
        RECT 90.275 239.195 90.605 239.525 ;
        RECT 90.275 237.835 90.605 238.165 ;
        RECT 90.28 237.16 90.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.275 -99.445 90.605 -99.115 ;
        RECT 90.275 -100.805 90.605 -100.475 ;
        RECT 90.275 -102.165 90.605 -101.835 ;
        RECT 90.275 -103.525 90.605 -103.195 ;
        RECT 90.275 -104.885 90.605 -104.555 ;
        RECT 90.275 -106.245 90.605 -105.915 ;
        RECT 90.275 -107.605 90.605 -107.275 ;
        RECT 90.275 -108.965 90.605 -108.635 ;
        RECT 90.275 -110.325 90.605 -109.995 ;
        RECT 90.275 -111.685 90.605 -111.355 ;
        RECT 90.275 -113.045 90.605 -112.715 ;
        RECT 90.275 -114.405 90.605 -114.075 ;
        RECT 90.275 -115.765 90.605 -115.435 ;
        RECT 90.275 -117.125 90.605 -116.795 ;
        RECT 90.275 -118.485 90.605 -118.155 ;
        RECT 90.275 -119.845 90.605 -119.515 ;
        RECT 90.275 -121.205 90.605 -120.875 ;
        RECT 90.275 -122.565 90.605 -122.235 ;
        RECT 90.275 -123.925 90.605 -123.595 ;
        RECT 90.275 -125.285 90.605 -124.955 ;
        RECT 90.275 -126.645 90.605 -126.315 ;
        RECT 90.275 -128.005 90.605 -127.675 ;
        RECT 90.275 -129.365 90.605 -129.035 ;
        RECT 90.275 -130.725 90.605 -130.395 ;
        RECT 90.275 -132.085 90.605 -131.755 ;
        RECT 90.275 -133.445 90.605 -133.115 ;
        RECT 90.275 -134.805 90.605 -134.475 ;
        RECT 90.275 -136.165 90.605 -135.835 ;
        RECT 90.275 -137.525 90.605 -137.195 ;
        RECT 90.275 -138.885 90.605 -138.555 ;
        RECT 90.275 -140.245 90.605 -139.915 ;
        RECT 90.275 -141.605 90.605 -141.275 ;
        RECT 90.275 -142.965 90.605 -142.635 ;
        RECT 90.275 -144.325 90.605 -143.995 ;
        RECT 90.275 -145.685 90.605 -145.355 ;
        RECT 90.275 -147.045 90.605 -146.715 ;
        RECT 90.275 -148.405 90.605 -148.075 ;
        RECT 90.275 -149.765 90.605 -149.435 ;
        RECT 90.275 -151.125 90.605 -150.795 ;
        RECT 90.275 -152.485 90.605 -152.155 ;
        RECT 90.275 -153.845 90.605 -153.515 ;
        RECT 90.275 -155.205 90.605 -154.875 ;
        RECT 90.275 -156.565 90.605 -156.235 ;
        RECT 90.275 -157.925 90.605 -157.595 ;
        RECT 90.275 -159.285 90.605 -158.955 ;
        RECT 90.275 -160.645 90.605 -160.315 ;
        RECT 90.275 -162.005 90.605 -161.675 ;
        RECT 90.275 -163.365 90.605 -163.035 ;
        RECT 90.275 -164.725 90.605 -164.395 ;
        RECT 90.275 -166.085 90.605 -165.755 ;
        RECT 90.275 -167.445 90.605 -167.115 ;
        RECT 90.275 -168.805 90.605 -168.475 ;
        RECT 90.275 -170.165 90.605 -169.835 ;
        RECT 90.275 -171.525 90.605 -171.195 ;
        RECT 90.275 -172.885 90.605 -172.555 ;
        RECT 90.275 -174.245 90.605 -173.915 ;
        RECT 90.275 -175.605 90.605 -175.275 ;
        RECT 90.275 -176.965 90.605 -176.635 ;
        RECT 90.275 -178.325 90.605 -177.995 ;
        RECT 90.275 -179.685 90.605 -179.355 ;
        RECT 90.275 -181.93 90.605 -180.8 ;
        RECT 90.28 -182.045 90.6 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 90.51 -98.075 90.84 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 241.32 44.365 242.45 ;
        RECT 44.035 239.195 44.365 239.525 ;
        RECT 44.035 237.835 44.365 238.165 ;
        RECT 44.04 237.16 44.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 -1.525 44.365 -1.195 ;
        RECT 44.035 -2.885 44.365 -2.555 ;
        RECT 44.04 -3.56 44.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 44.035 -95.365 44.365 -95.035 ;
        RECT 44.035 -96.725 44.365 -96.395 ;
        RECT 44.035 -98.085 44.365 -97.755 ;
        RECT 44.035 -99.445 44.365 -99.115 ;
        RECT 44.035 -100.805 44.365 -100.475 ;
        RECT 44.035 -102.165 44.365 -101.835 ;
        RECT 44.035 -103.525 44.365 -103.195 ;
        RECT 44.035 -104.885 44.365 -104.555 ;
        RECT 44.035 -106.245 44.365 -105.915 ;
        RECT 44.035 -107.605 44.365 -107.275 ;
        RECT 44.035 -108.965 44.365 -108.635 ;
        RECT 44.035 -110.325 44.365 -109.995 ;
        RECT 44.035 -111.685 44.365 -111.355 ;
        RECT 44.035 -113.045 44.365 -112.715 ;
        RECT 44.035 -114.405 44.365 -114.075 ;
        RECT 44.035 -115.765 44.365 -115.435 ;
        RECT 44.035 -117.125 44.365 -116.795 ;
        RECT 44.035 -118.485 44.365 -118.155 ;
        RECT 44.035 -119.845 44.365 -119.515 ;
        RECT 44.035 -121.205 44.365 -120.875 ;
        RECT 44.035 -122.565 44.365 -122.235 ;
        RECT 44.035 -123.925 44.365 -123.595 ;
        RECT 44.035 -125.285 44.365 -124.955 ;
        RECT 44.035 -126.645 44.365 -126.315 ;
        RECT 44.035 -128.005 44.365 -127.675 ;
        RECT 44.035 -129.365 44.365 -129.035 ;
        RECT 44.035 -130.725 44.365 -130.395 ;
        RECT 44.035 -132.085 44.365 -131.755 ;
        RECT 44.035 -133.445 44.365 -133.115 ;
        RECT 44.035 -134.805 44.365 -134.475 ;
        RECT 44.035 -136.165 44.365 -135.835 ;
        RECT 44.035 -137.525 44.365 -137.195 ;
        RECT 44.035 -138.885 44.365 -138.555 ;
        RECT 44.035 -140.245 44.365 -139.915 ;
        RECT 44.035 -141.605 44.365 -141.275 ;
        RECT 44.035 -142.965 44.365 -142.635 ;
        RECT 44.035 -144.325 44.365 -143.995 ;
        RECT 44.035 -145.685 44.365 -145.355 ;
        RECT 44.035 -147.045 44.365 -146.715 ;
        RECT 44.035 -148.405 44.365 -148.075 ;
        RECT 44.035 -149.765 44.365 -149.435 ;
        RECT 44.035 -151.125 44.365 -150.795 ;
        RECT 44.035 -152.485 44.365 -152.155 ;
        RECT 44.035 -153.845 44.365 -153.515 ;
        RECT 44.035 -155.205 44.365 -154.875 ;
        RECT 44.035 -156.565 44.365 -156.235 ;
        RECT 44.035 -157.925 44.365 -157.595 ;
        RECT 44.035 -159.285 44.365 -158.955 ;
        RECT 44.035 -160.645 44.365 -160.315 ;
        RECT 44.035 -162.005 44.365 -161.675 ;
        RECT 44.035 -163.365 44.365 -163.035 ;
        RECT 44.035 -164.725 44.365 -164.395 ;
        RECT 44.035 -166.085 44.365 -165.755 ;
        RECT 44.035 -167.445 44.365 -167.115 ;
        RECT 44.035 -168.805 44.365 -168.475 ;
        RECT 44.035 -170.165 44.365 -169.835 ;
        RECT 44.035 -171.525 44.365 -171.195 ;
        RECT 44.035 -172.885 44.365 -172.555 ;
        RECT 44.035 -174.245 44.365 -173.915 ;
        RECT 44.035 -175.605 44.365 -175.275 ;
        RECT 44.035 -176.965 44.365 -176.635 ;
        RECT 44.035 -178.325 44.365 -177.995 ;
        RECT 44.035 -179.685 44.365 -179.355 ;
        RECT 44.035 -181.93 44.365 -180.8 ;
        RECT 44.04 -182.045 44.36 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 241.32 45.725 242.45 ;
        RECT 45.395 239.195 45.725 239.525 ;
        RECT 45.395 237.835 45.725 238.165 ;
        RECT 45.4 237.16 45.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 -1.525 45.725 -1.195 ;
        RECT 45.395 -2.885 45.725 -2.555 ;
        RECT 45.4 -3.56 45.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 45.395 -95.365 45.725 -95.035 ;
        RECT 45.395 -96.725 45.725 -96.395 ;
        RECT 45.395 -98.085 45.725 -97.755 ;
        RECT 45.395 -99.445 45.725 -99.115 ;
        RECT 45.395 -100.805 45.725 -100.475 ;
        RECT 45.395 -102.165 45.725 -101.835 ;
        RECT 45.395 -103.525 45.725 -103.195 ;
        RECT 45.395 -104.885 45.725 -104.555 ;
        RECT 45.395 -106.245 45.725 -105.915 ;
        RECT 45.395 -107.605 45.725 -107.275 ;
        RECT 45.395 -108.965 45.725 -108.635 ;
        RECT 45.395 -110.325 45.725 -109.995 ;
        RECT 45.395 -111.685 45.725 -111.355 ;
        RECT 45.395 -113.045 45.725 -112.715 ;
        RECT 45.395 -114.405 45.725 -114.075 ;
        RECT 45.395 -115.765 45.725 -115.435 ;
        RECT 45.395 -117.125 45.725 -116.795 ;
        RECT 45.395 -118.485 45.725 -118.155 ;
        RECT 45.395 -119.845 45.725 -119.515 ;
        RECT 45.395 -121.205 45.725 -120.875 ;
        RECT 45.395 -122.565 45.725 -122.235 ;
        RECT 45.395 -123.925 45.725 -123.595 ;
        RECT 45.395 -125.285 45.725 -124.955 ;
        RECT 45.395 -126.645 45.725 -126.315 ;
        RECT 45.395 -128.005 45.725 -127.675 ;
        RECT 45.395 -129.365 45.725 -129.035 ;
        RECT 45.395 -130.725 45.725 -130.395 ;
        RECT 45.395 -132.085 45.725 -131.755 ;
        RECT 45.395 -133.445 45.725 -133.115 ;
        RECT 45.395 -134.805 45.725 -134.475 ;
        RECT 45.395 -136.165 45.725 -135.835 ;
        RECT 45.395 -137.525 45.725 -137.195 ;
        RECT 45.395 -138.885 45.725 -138.555 ;
        RECT 45.395 -140.245 45.725 -139.915 ;
        RECT 45.395 -141.605 45.725 -141.275 ;
        RECT 45.395 -142.965 45.725 -142.635 ;
        RECT 45.395 -144.325 45.725 -143.995 ;
        RECT 45.395 -145.685 45.725 -145.355 ;
        RECT 45.395 -147.045 45.725 -146.715 ;
        RECT 45.395 -148.405 45.725 -148.075 ;
        RECT 45.395 -149.765 45.725 -149.435 ;
        RECT 45.395 -151.125 45.725 -150.795 ;
        RECT 45.395 -152.485 45.725 -152.155 ;
        RECT 45.395 -153.845 45.725 -153.515 ;
        RECT 45.395 -155.205 45.725 -154.875 ;
        RECT 45.395 -156.565 45.725 -156.235 ;
        RECT 45.395 -157.925 45.725 -157.595 ;
        RECT 45.395 -159.285 45.725 -158.955 ;
        RECT 45.395 -160.645 45.725 -160.315 ;
        RECT 45.395 -162.005 45.725 -161.675 ;
        RECT 45.395 -163.365 45.725 -163.035 ;
        RECT 45.395 -164.725 45.725 -164.395 ;
        RECT 45.395 -166.085 45.725 -165.755 ;
        RECT 45.395 -167.445 45.725 -167.115 ;
        RECT 45.395 -168.805 45.725 -168.475 ;
        RECT 45.395 -170.165 45.725 -169.835 ;
        RECT 45.395 -171.525 45.725 -171.195 ;
        RECT 45.395 -172.885 45.725 -172.555 ;
        RECT 45.395 -174.245 45.725 -173.915 ;
        RECT 45.395 -175.605 45.725 -175.275 ;
        RECT 45.395 -176.965 45.725 -176.635 ;
        RECT 45.395 -178.325 45.725 -177.995 ;
        RECT 45.395 -179.685 45.725 -179.355 ;
        RECT 45.395 -181.93 45.725 -180.8 ;
        RECT 45.4 -182.045 45.72 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 241.32 47.085 242.45 ;
        RECT 46.755 239.195 47.085 239.525 ;
        RECT 46.755 237.835 47.085 238.165 ;
        RECT 46.76 237.16 47.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.755 -99.445 47.085 -99.115 ;
        RECT 46.755 -100.805 47.085 -100.475 ;
        RECT 46.755 -102.165 47.085 -101.835 ;
        RECT 46.755 -103.525 47.085 -103.195 ;
        RECT 46.755 -104.885 47.085 -104.555 ;
        RECT 46.755 -106.245 47.085 -105.915 ;
        RECT 46.755 -107.605 47.085 -107.275 ;
        RECT 46.755 -108.965 47.085 -108.635 ;
        RECT 46.755 -110.325 47.085 -109.995 ;
        RECT 46.755 -111.685 47.085 -111.355 ;
        RECT 46.755 -113.045 47.085 -112.715 ;
        RECT 46.755 -114.405 47.085 -114.075 ;
        RECT 46.755 -115.765 47.085 -115.435 ;
        RECT 46.755 -117.125 47.085 -116.795 ;
        RECT 46.755 -118.485 47.085 -118.155 ;
        RECT 46.755 -119.845 47.085 -119.515 ;
        RECT 46.755 -121.205 47.085 -120.875 ;
        RECT 46.755 -122.565 47.085 -122.235 ;
        RECT 46.755 -123.925 47.085 -123.595 ;
        RECT 46.755 -125.285 47.085 -124.955 ;
        RECT 46.755 -126.645 47.085 -126.315 ;
        RECT 46.755 -128.005 47.085 -127.675 ;
        RECT 46.755 -129.365 47.085 -129.035 ;
        RECT 46.755 -130.725 47.085 -130.395 ;
        RECT 46.755 -132.085 47.085 -131.755 ;
        RECT 46.755 -133.445 47.085 -133.115 ;
        RECT 46.755 -134.805 47.085 -134.475 ;
        RECT 46.755 -136.165 47.085 -135.835 ;
        RECT 46.755 -137.525 47.085 -137.195 ;
        RECT 46.755 -138.885 47.085 -138.555 ;
        RECT 46.755 -140.245 47.085 -139.915 ;
        RECT 46.755 -141.605 47.085 -141.275 ;
        RECT 46.755 -142.965 47.085 -142.635 ;
        RECT 46.755 -144.325 47.085 -143.995 ;
        RECT 46.755 -145.685 47.085 -145.355 ;
        RECT 46.755 -147.045 47.085 -146.715 ;
        RECT 46.755 -148.405 47.085 -148.075 ;
        RECT 46.755 -149.765 47.085 -149.435 ;
        RECT 46.755 -151.125 47.085 -150.795 ;
        RECT 46.755 -152.485 47.085 -152.155 ;
        RECT 46.755 -153.845 47.085 -153.515 ;
        RECT 46.755 -155.205 47.085 -154.875 ;
        RECT 46.755 -156.565 47.085 -156.235 ;
        RECT 46.755 -157.925 47.085 -157.595 ;
        RECT 46.755 -159.285 47.085 -158.955 ;
        RECT 46.755 -160.645 47.085 -160.315 ;
        RECT 46.755 -162.005 47.085 -161.675 ;
        RECT 46.755 -163.365 47.085 -163.035 ;
        RECT 46.755 -164.725 47.085 -164.395 ;
        RECT 46.755 -166.085 47.085 -165.755 ;
        RECT 46.755 -167.445 47.085 -167.115 ;
        RECT 46.755 -168.805 47.085 -168.475 ;
        RECT 46.755 -170.165 47.085 -169.835 ;
        RECT 46.755 -171.525 47.085 -171.195 ;
        RECT 46.755 -172.885 47.085 -172.555 ;
        RECT 46.755 -174.245 47.085 -173.915 ;
        RECT 46.755 -175.605 47.085 -175.275 ;
        RECT 46.755 -176.965 47.085 -176.635 ;
        RECT 46.755 -178.325 47.085 -177.995 ;
        RECT 46.755 -179.685 47.085 -179.355 ;
        RECT 46.755 -181.93 47.085 -180.8 ;
        RECT 46.76 -182.045 47.08 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 46.91 -98.075 47.24 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 241.32 48.445 242.45 ;
        RECT 48.115 239.195 48.445 239.525 ;
        RECT 48.115 237.835 48.445 238.165 ;
        RECT 48.12 237.16 48.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 48.115 -1.525 48.445 -1.195 ;
        RECT 48.115 -2.885 48.445 -2.555 ;
        RECT 48.12 -3.56 48.44 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 241.32 49.805 242.45 ;
        RECT 49.475 239.195 49.805 239.525 ;
        RECT 49.475 237.835 49.805 238.165 ;
        RECT 49.48 237.16 49.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 49.475 -1.525 49.805 -1.195 ;
        RECT 49.475 -2.885 49.805 -2.555 ;
        RECT 49.48 -3.56 49.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 241.32 51.165 242.45 ;
        RECT 50.835 239.195 51.165 239.525 ;
        RECT 50.835 237.835 51.165 238.165 ;
        RECT 50.84 237.16 51.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 -1.525 51.165 -1.195 ;
        RECT 50.835 -2.885 51.165 -2.555 ;
        RECT 50.84 -3.56 51.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 50.835 -95.365 51.165 -95.035 ;
        RECT 50.835 -96.725 51.165 -96.395 ;
        RECT 50.835 -98.085 51.165 -97.755 ;
        RECT 50.835 -99.445 51.165 -99.115 ;
        RECT 50.835 -100.805 51.165 -100.475 ;
        RECT 50.835 -102.165 51.165 -101.835 ;
        RECT 50.835 -103.525 51.165 -103.195 ;
        RECT 50.835 -104.885 51.165 -104.555 ;
        RECT 50.835 -106.245 51.165 -105.915 ;
        RECT 50.835 -107.605 51.165 -107.275 ;
        RECT 50.835 -108.965 51.165 -108.635 ;
        RECT 50.835 -110.325 51.165 -109.995 ;
        RECT 50.835 -111.685 51.165 -111.355 ;
        RECT 50.835 -113.045 51.165 -112.715 ;
        RECT 50.835 -114.405 51.165 -114.075 ;
        RECT 50.835 -115.765 51.165 -115.435 ;
        RECT 50.835 -117.125 51.165 -116.795 ;
        RECT 50.835 -118.485 51.165 -118.155 ;
        RECT 50.835 -119.845 51.165 -119.515 ;
        RECT 50.835 -121.205 51.165 -120.875 ;
        RECT 50.835 -122.565 51.165 -122.235 ;
        RECT 50.835 -123.925 51.165 -123.595 ;
        RECT 50.835 -125.285 51.165 -124.955 ;
        RECT 50.835 -126.645 51.165 -126.315 ;
        RECT 50.835 -128.005 51.165 -127.675 ;
        RECT 50.835 -129.365 51.165 -129.035 ;
        RECT 50.835 -130.725 51.165 -130.395 ;
        RECT 50.835 -132.085 51.165 -131.755 ;
        RECT 50.835 -133.445 51.165 -133.115 ;
        RECT 50.835 -134.805 51.165 -134.475 ;
        RECT 50.835 -136.165 51.165 -135.835 ;
        RECT 50.835 -137.525 51.165 -137.195 ;
        RECT 50.835 -138.885 51.165 -138.555 ;
        RECT 50.835 -140.245 51.165 -139.915 ;
        RECT 50.835 -141.605 51.165 -141.275 ;
        RECT 50.835 -142.965 51.165 -142.635 ;
        RECT 50.835 -144.325 51.165 -143.995 ;
        RECT 50.835 -145.685 51.165 -145.355 ;
        RECT 50.835 -147.045 51.165 -146.715 ;
        RECT 50.835 -148.405 51.165 -148.075 ;
        RECT 50.835 -149.765 51.165 -149.435 ;
        RECT 50.835 -151.125 51.165 -150.795 ;
        RECT 50.835 -152.485 51.165 -152.155 ;
        RECT 50.835 -153.845 51.165 -153.515 ;
        RECT 50.835 -155.205 51.165 -154.875 ;
        RECT 50.835 -156.565 51.165 -156.235 ;
        RECT 50.835 -157.925 51.165 -157.595 ;
        RECT 50.835 -159.285 51.165 -158.955 ;
        RECT 50.835 -160.645 51.165 -160.315 ;
        RECT 50.835 -162.005 51.165 -161.675 ;
        RECT 50.835 -163.365 51.165 -163.035 ;
        RECT 50.835 -164.725 51.165 -164.395 ;
        RECT 50.835 -166.085 51.165 -165.755 ;
        RECT 50.835 -167.445 51.165 -167.115 ;
        RECT 50.835 -168.805 51.165 -168.475 ;
        RECT 50.835 -170.165 51.165 -169.835 ;
        RECT 50.835 -171.525 51.165 -171.195 ;
        RECT 50.835 -172.885 51.165 -172.555 ;
        RECT 50.835 -174.245 51.165 -173.915 ;
        RECT 50.835 -175.605 51.165 -175.275 ;
        RECT 50.835 -176.965 51.165 -176.635 ;
        RECT 50.835 -178.325 51.165 -177.995 ;
        RECT 50.835 -179.685 51.165 -179.355 ;
        RECT 50.835 -181.93 51.165 -180.8 ;
        RECT 50.84 -182.045 51.16 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.195 241.32 52.525 242.45 ;
        RECT 52.195 239.195 52.525 239.525 ;
        RECT 52.195 237.835 52.525 238.165 ;
        RECT 52.2 237.16 52.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.195 -1.525 52.525 -1.195 ;
        RECT 52.195 -2.885 52.525 -2.555 ;
        RECT 52.2 -3.56 52.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 52.195 -95.365 52.525 -95.035 ;
        RECT 52.195 -96.725 52.525 -96.395 ;
        RECT 52.195 -98.085 52.525 -97.755 ;
        RECT 52.195 -99.445 52.525 -99.115 ;
        RECT 52.195 -100.805 52.525 -100.475 ;
        RECT 52.195 -102.165 52.525 -101.835 ;
        RECT 52.195 -103.525 52.525 -103.195 ;
        RECT 52.195 -104.885 52.525 -104.555 ;
        RECT 52.195 -106.245 52.525 -105.915 ;
        RECT 52.195 -107.605 52.525 -107.275 ;
        RECT 52.195 -108.965 52.525 -108.635 ;
        RECT 52.195 -110.325 52.525 -109.995 ;
        RECT 52.195 -111.685 52.525 -111.355 ;
        RECT 52.195 -113.045 52.525 -112.715 ;
        RECT 52.195 -114.405 52.525 -114.075 ;
        RECT 52.195 -115.765 52.525 -115.435 ;
        RECT 52.195 -117.125 52.525 -116.795 ;
        RECT 52.195 -118.485 52.525 -118.155 ;
        RECT 52.195 -119.845 52.525 -119.515 ;
        RECT 52.195 -121.205 52.525 -120.875 ;
        RECT 52.195 -122.565 52.525 -122.235 ;
        RECT 52.195 -123.925 52.525 -123.595 ;
        RECT 52.195 -125.285 52.525 -124.955 ;
        RECT 52.195 -126.645 52.525 -126.315 ;
        RECT 52.195 -128.005 52.525 -127.675 ;
        RECT 52.195 -129.365 52.525 -129.035 ;
        RECT 52.195 -130.725 52.525 -130.395 ;
        RECT 52.195 -132.085 52.525 -131.755 ;
        RECT 52.195 -133.445 52.525 -133.115 ;
        RECT 52.195 -134.805 52.525 -134.475 ;
        RECT 52.195 -136.165 52.525 -135.835 ;
        RECT 52.195 -137.525 52.525 -137.195 ;
        RECT 52.195 -138.885 52.525 -138.555 ;
        RECT 52.195 -140.245 52.525 -139.915 ;
        RECT 52.195 -141.605 52.525 -141.275 ;
        RECT 52.195 -142.965 52.525 -142.635 ;
        RECT 52.195 -144.325 52.525 -143.995 ;
        RECT 52.195 -145.685 52.525 -145.355 ;
        RECT 52.195 -147.045 52.525 -146.715 ;
        RECT 52.195 -148.405 52.525 -148.075 ;
        RECT 52.195 -149.765 52.525 -149.435 ;
        RECT 52.195 -151.125 52.525 -150.795 ;
        RECT 52.195 -152.485 52.525 -152.155 ;
        RECT 52.195 -153.845 52.525 -153.515 ;
        RECT 52.195 -155.205 52.525 -154.875 ;
        RECT 52.195 -156.565 52.525 -156.235 ;
        RECT 52.195 -157.925 52.525 -157.595 ;
        RECT 52.195 -159.285 52.525 -158.955 ;
        RECT 52.195 -160.645 52.525 -160.315 ;
        RECT 52.195 -162.005 52.525 -161.675 ;
        RECT 52.195 -163.365 52.525 -163.035 ;
        RECT 52.195 -164.725 52.525 -164.395 ;
        RECT 52.195 -166.085 52.525 -165.755 ;
        RECT 52.195 -167.445 52.525 -167.115 ;
        RECT 52.195 -168.805 52.525 -168.475 ;
        RECT 52.195 -170.165 52.525 -169.835 ;
        RECT 52.195 -171.525 52.525 -171.195 ;
        RECT 52.195 -172.885 52.525 -172.555 ;
        RECT 52.195 -174.245 52.525 -173.915 ;
        RECT 52.195 -175.605 52.525 -175.275 ;
        RECT 52.195 -176.965 52.525 -176.635 ;
        RECT 52.195 -178.325 52.525 -177.995 ;
        RECT 52.195 -179.685 52.525 -179.355 ;
        RECT 52.195 -181.93 52.525 -180.8 ;
        RECT 52.2 -182.045 52.52 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 241.32 53.885 242.45 ;
        RECT 53.555 239.195 53.885 239.525 ;
        RECT 53.555 237.835 53.885 238.165 ;
        RECT 53.56 237.16 53.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 -1.525 53.885 -1.195 ;
        RECT 53.555 -2.885 53.885 -2.555 ;
        RECT 53.56 -3.56 53.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 53.555 -95.365 53.885 -95.035 ;
        RECT 53.555 -96.725 53.885 -96.395 ;
        RECT 53.555 -98.085 53.885 -97.755 ;
        RECT 53.555 -99.445 53.885 -99.115 ;
        RECT 53.555 -100.805 53.885 -100.475 ;
        RECT 53.555 -102.165 53.885 -101.835 ;
        RECT 53.555 -103.525 53.885 -103.195 ;
        RECT 53.555 -104.885 53.885 -104.555 ;
        RECT 53.555 -106.245 53.885 -105.915 ;
        RECT 53.555 -107.605 53.885 -107.275 ;
        RECT 53.555 -108.965 53.885 -108.635 ;
        RECT 53.555 -110.325 53.885 -109.995 ;
        RECT 53.555 -111.685 53.885 -111.355 ;
        RECT 53.555 -113.045 53.885 -112.715 ;
        RECT 53.555 -114.405 53.885 -114.075 ;
        RECT 53.555 -115.765 53.885 -115.435 ;
        RECT 53.555 -117.125 53.885 -116.795 ;
        RECT 53.555 -118.485 53.885 -118.155 ;
        RECT 53.555 -119.845 53.885 -119.515 ;
        RECT 53.555 -121.205 53.885 -120.875 ;
        RECT 53.555 -122.565 53.885 -122.235 ;
        RECT 53.555 -123.925 53.885 -123.595 ;
        RECT 53.555 -125.285 53.885 -124.955 ;
        RECT 53.555 -126.645 53.885 -126.315 ;
        RECT 53.555 -128.005 53.885 -127.675 ;
        RECT 53.555 -129.365 53.885 -129.035 ;
        RECT 53.555 -130.725 53.885 -130.395 ;
        RECT 53.555 -132.085 53.885 -131.755 ;
        RECT 53.555 -133.445 53.885 -133.115 ;
        RECT 53.555 -134.805 53.885 -134.475 ;
        RECT 53.555 -136.165 53.885 -135.835 ;
        RECT 53.555 -137.525 53.885 -137.195 ;
        RECT 53.555 -138.885 53.885 -138.555 ;
        RECT 53.555 -140.245 53.885 -139.915 ;
        RECT 53.555 -141.605 53.885 -141.275 ;
        RECT 53.555 -142.965 53.885 -142.635 ;
        RECT 53.555 -144.325 53.885 -143.995 ;
        RECT 53.555 -145.685 53.885 -145.355 ;
        RECT 53.555 -147.045 53.885 -146.715 ;
        RECT 53.555 -148.405 53.885 -148.075 ;
        RECT 53.555 -149.765 53.885 -149.435 ;
        RECT 53.555 -151.125 53.885 -150.795 ;
        RECT 53.555 -152.485 53.885 -152.155 ;
        RECT 53.555 -153.845 53.885 -153.515 ;
        RECT 53.555 -155.205 53.885 -154.875 ;
        RECT 53.555 -156.565 53.885 -156.235 ;
        RECT 53.555 -157.925 53.885 -157.595 ;
        RECT 53.555 -159.285 53.885 -158.955 ;
        RECT 53.555 -160.645 53.885 -160.315 ;
        RECT 53.555 -162.005 53.885 -161.675 ;
        RECT 53.555 -163.365 53.885 -163.035 ;
        RECT 53.555 -164.725 53.885 -164.395 ;
        RECT 53.555 -166.085 53.885 -165.755 ;
        RECT 53.555 -167.445 53.885 -167.115 ;
        RECT 53.555 -168.805 53.885 -168.475 ;
        RECT 53.555 -170.165 53.885 -169.835 ;
        RECT 53.555 -171.525 53.885 -171.195 ;
        RECT 53.555 -172.885 53.885 -172.555 ;
        RECT 53.555 -174.245 53.885 -173.915 ;
        RECT 53.555 -175.605 53.885 -175.275 ;
        RECT 53.555 -176.965 53.885 -176.635 ;
        RECT 53.555 -178.325 53.885 -177.995 ;
        RECT 53.555 -179.685 53.885 -179.355 ;
        RECT 53.555 -181.93 53.885 -180.8 ;
        RECT 53.56 -182.045 53.88 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 241.32 55.245 242.45 ;
        RECT 54.915 239.195 55.245 239.525 ;
        RECT 54.915 237.835 55.245 238.165 ;
        RECT 54.92 237.16 55.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 -1.525 55.245 -1.195 ;
        RECT 54.915 -2.885 55.245 -2.555 ;
        RECT 54.92 -3.56 55.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 54.915 -95.365 55.245 -95.035 ;
        RECT 54.915 -96.725 55.245 -96.395 ;
        RECT 54.915 -98.085 55.245 -97.755 ;
        RECT 54.915 -99.445 55.245 -99.115 ;
        RECT 54.915 -100.805 55.245 -100.475 ;
        RECT 54.915 -102.165 55.245 -101.835 ;
        RECT 54.915 -103.525 55.245 -103.195 ;
        RECT 54.915 -104.885 55.245 -104.555 ;
        RECT 54.915 -106.245 55.245 -105.915 ;
        RECT 54.915 -107.605 55.245 -107.275 ;
        RECT 54.915 -108.965 55.245 -108.635 ;
        RECT 54.915 -110.325 55.245 -109.995 ;
        RECT 54.915 -111.685 55.245 -111.355 ;
        RECT 54.915 -113.045 55.245 -112.715 ;
        RECT 54.915 -114.405 55.245 -114.075 ;
        RECT 54.915 -115.765 55.245 -115.435 ;
        RECT 54.915 -117.125 55.245 -116.795 ;
        RECT 54.915 -118.485 55.245 -118.155 ;
        RECT 54.915 -119.845 55.245 -119.515 ;
        RECT 54.915 -121.205 55.245 -120.875 ;
        RECT 54.915 -122.565 55.245 -122.235 ;
        RECT 54.915 -123.925 55.245 -123.595 ;
        RECT 54.915 -125.285 55.245 -124.955 ;
        RECT 54.915 -126.645 55.245 -126.315 ;
        RECT 54.915 -128.005 55.245 -127.675 ;
        RECT 54.915 -129.365 55.245 -129.035 ;
        RECT 54.915 -130.725 55.245 -130.395 ;
        RECT 54.915 -132.085 55.245 -131.755 ;
        RECT 54.915 -133.445 55.245 -133.115 ;
        RECT 54.915 -134.805 55.245 -134.475 ;
        RECT 54.915 -136.165 55.245 -135.835 ;
        RECT 54.915 -137.525 55.245 -137.195 ;
        RECT 54.915 -138.885 55.245 -138.555 ;
        RECT 54.915 -140.245 55.245 -139.915 ;
        RECT 54.915 -141.605 55.245 -141.275 ;
        RECT 54.915 -142.965 55.245 -142.635 ;
        RECT 54.915 -144.325 55.245 -143.995 ;
        RECT 54.915 -145.685 55.245 -145.355 ;
        RECT 54.915 -147.045 55.245 -146.715 ;
        RECT 54.915 -148.405 55.245 -148.075 ;
        RECT 54.915 -149.765 55.245 -149.435 ;
        RECT 54.915 -151.125 55.245 -150.795 ;
        RECT 54.915 -152.485 55.245 -152.155 ;
        RECT 54.915 -153.845 55.245 -153.515 ;
        RECT 54.915 -155.205 55.245 -154.875 ;
        RECT 54.915 -156.565 55.245 -156.235 ;
        RECT 54.915 -157.925 55.245 -157.595 ;
        RECT 54.915 -159.285 55.245 -158.955 ;
        RECT 54.915 -160.645 55.245 -160.315 ;
        RECT 54.915 -162.005 55.245 -161.675 ;
        RECT 54.915 -163.365 55.245 -163.035 ;
        RECT 54.915 -164.725 55.245 -164.395 ;
        RECT 54.915 -166.085 55.245 -165.755 ;
        RECT 54.915 -167.445 55.245 -167.115 ;
        RECT 54.915 -168.805 55.245 -168.475 ;
        RECT 54.915 -170.165 55.245 -169.835 ;
        RECT 54.915 -171.525 55.245 -171.195 ;
        RECT 54.915 -172.885 55.245 -172.555 ;
        RECT 54.915 -174.245 55.245 -173.915 ;
        RECT 54.915 -175.605 55.245 -175.275 ;
        RECT 54.915 -176.965 55.245 -176.635 ;
        RECT 54.915 -178.325 55.245 -177.995 ;
        RECT 54.915 -179.685 55.245 -179.355 ;
        RECT 54.915 -181.93 55.245 -180.8 ;
        RECT 54.92 -182.045 55.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 241.32 56.605 242.45 ;
        RECT 56.275 239.195 56.605 239.525 ;
        RECT 56.275 237.835 56.605 238.165 ;
        RECT 56.28 237.16 56.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 -1.525 56.605 -1.195 ;
        RECT 56.275 -2.885 56.605 -2.555 ;
        RECT 56.28 -3.56 56.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 56.275 -95.365 56.605 -95.035 ;
        RECT 56.275 -96.725 56.605 -96.395 ;
        RECT 56.275 -98.085 56.605 -97.755 ;
        RECT 56.275 -99.445 56.605 -99.115 ;
        RECT 56.275 -100.805 56.605 -100.475 ;
        RECT 56.275 -102.165 56.605 -101.835 ;
        RECT 56.275 -103.525 56.605 -103.195 ;
        RECT 56.275 -104.885 56.605 -104.555 ;
        RECT 56.275 -106.245 56.605 -105.915 ;
        RECT 56.275 -107.605 56.605 -107.275 ;
        RECT 56.275 -108.965 56.605 -108.635 ;
        RECT 56.275 -110.325 56.605 -109.995 ;
        RECT 56.275 -111.685 56.605 -111.355 ;
        RECT 56.275 -113.045 56.605 -112.715 ;
        RECT 56.275 -114.405 56.605 -114.075 ;
        RECT 56.275 -115.765 56.605 -115.435 ;
        RECT 56.275 -117.125 56.605 -116.795 ;
        RECT 56.275 -118.485 56.605 -118.155 ;
        RECT 56.275 -119.845 56.605 -119.515 ;
        RECT 56.275 -121.205 56.605 -120.875 ;
        RECT 56.275 -122.565 56.605 -122.235 ;
        RECT 56.275 -123.925 56.605 -123.595 ;
        RECT 56.275 -125.285 56.605 -124.955 ;
        RECT 56.275 -126.645 56.605 -126.315 ;
        RECT 56.275 -128.005 56.605 -127.675 ;
        RECT 56.275 -129.365 56.605 -129.035 ;
        RECT 56.275 -130.725 56.605 -130.395 ;
        RECT 56.275 -132.085 56.605 -131.755 ;
        RECT 56.275 -133.445 56.605 -133.115 ;
        RECT 56.275 -134.805 56.605 -134.475 ;
        RECT 56.275 -136.165 56.605 -135.835 ;
        RECT 56.275 -137.525 56.605 -137.195 ;
        RECT 56.275 -138.885 56.605 -138.555 ;
        RECT 56.275 -140.245 56.605 -139.915 ;
        RECT 56.275 -141.605 56.605 -141.275 ;
        RECT 56.275 -142.965 56.605 -142.635 ;
        RECT 56.275 -144.325 56.605 -143.995 ;
        RECT 56.275 -145.685 56.605 -145.355 ;
        RECT 56.275 -147.045 56.605 -146.715 ;
        RECT 56.275 -148.405 56.605 -148.075 ;
        RECT 56.275 -149.765 56.605 -149.435 ;
        RECT 56.275 -151.125 56.605 -150.795 ;
        RECT 56.275 -152.485 56.605 -152.155 ;
        RECT 56.275 -153.845 56.605 -153.515 ;
        RECT 56.275 -155.205 56.605 -154.875 ;
        RECT 56.275 -156.565 56.605 -156.235 ;
        RECT 56.275 -157.925 56.605 -157.595 ;
        RECT 56.275 -159.285 56.605 -158.955 ;
        RECT 56.275 -160.645 56.605 -160.315 ;
        RECT 56.275 -162.005 56.605 -161.675 ;
        RECT 56.275 -163.365 56.605 -163.035 ;
        RECT 56.275 -164.725 56.605 -164.395 ;
        RECT 56.275 -166.085 56.605 -165.755 ;
        RECT 56.275 -167.445 56.605 -167.115 ;
        RECT 56.275 -168.805 56.605 -168.475 ;
        RECT 56.275 -170.165 56.605 -169.835 ;
        RECT 56.275 -171.525 56.605 -171.195 ;
        RECT 56.275 -172.885 56.605 -172.555 ;
        RECT 56.275 -174.245 56.605 -173.915 ;
        RECT 56.275 -175.605 56.605 -175.275 ;
        RECT 56.275 -176.965 56.605 -176.635 ;
        RECT 56.275 -178.325 56.605 -177.995 ;
        RECT 56.275 -179.685 56.605 -179.355 ;
        RECT 56.275 -181.93 56.605 -180.8 ;
        RECT 56.28 -182.045 56.6 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 241.32 57.965 242.45 ;
        RECT 57.635 239.195 57.965 239.525 ;
        RECT 57.635 237.835 57.965 238.165 ;
        RECT 57.64 237.16 57.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.635 -99.445 57.965 -99.115 ;
        RECT 57.635 -100.805 57.965 -100.475 ;
        RECT 57.635 -102.165 57.965 -101.835 ;
        RECT 57.635 -103.525 57.965 -103.195 ;
        RECT 57.635 -104.885 57.965 -104.555 ;
        RECT 57.635 -106.245 57.965 -105.915 ;
        RECT 57.635 -107.605 57.965 -107.275 ;
        RECT 57.635 -108.965 57.965 -108.635 ;
        RECT 57.635 -110.325 57.965 -109.995 ;
        RECT 57.635 -111.685 57.965 -111.355 ;
        RECT 57.635 -113.045 57.965 -112.715 ;
        RECT 57.635 -114.405 57.965 -114.075 ;
        RECT 57.635 -115.765 57.965 -115.435 ;
        RECT 57.635 -117.125 57.965 -116.795 ;
        RECT 57.635 -118.485 57.965 -118.155 ;
        RECT 57.635 -119.845 57.965 -119.515 ;
        RECT 57.635 -121.205 57.965 -120.875 ;
        RECT 57.635 -122.565 57.965 -122.235 ;
        RECT 57.635 -123.925 57.965 -123.595 ;
        RECT 57.635 -125.285 57.965 -124.955 ;
        RECT 57.635 -126.645 57.965 -126.315 ;
        RECT 57.635 -128.005 57.965 -127.675 ;
        RECT 57.635 -129.365 57.965 -129.035 ;
        RECT 57.635 -130.725 57.965 -130.395 ;
        RECT 57.635 -132.085 57.965 -131.755 ;
        RECT 57.635 -133.445 57.965 -133.115 ;
        RECT 57.635 -134.805 57.965 -134.475 ;
        RECT 57.635 -136.165 57.965 -135.835 ;
        RECT 57.635 -137.525 57.965 -137.195 ;
        RECT 57.635 -138.885 57.965 -138.555 ;
        RECT 57.635 -140.245 57.965 -139.915 ;
        RECT 57.635 -141.605 57.965 -141.275 ;
        RECT 57.635 -142.965 57.965 -142.635 ;
        RECT 57.635 -144.325 57.965 -143.995 ;
        RECT 57.635 -145.685 57.965 -145.355 ;
        RECT 57.635 -147.045 57.965 -146.715 ;
        RECT 57.635 -148.405 57.965 -148.075 ;
        RECT 57.635 -149.765 57.965 -149.435 ;
        RECT 57.635 -151.125 57.965 -150.795 ;
        RECT 57.635 -152.485 57.965 -152.155 ;
        RECT 57.635 -153.845 57.965 -153.515 ;
        RECT 57.635 -155.205 57.965 -154.875 ;
        RECT 57.635 -156.565 57.965 -156.235 ;
        RECT 57.635 -157.925 57.965 -157.595 ;
        RECT 57.635 -159.285 57.965 -158.955 ;
        RECT 57.635 -160.645 57.965 -160.315 ;
        RECT 57.635 -162.005 57.965 -161.675 ;
        RECT 57.635 -163.365 57.965 -163.035 ;
        RECT 57.635 -164.725 57.965 -164.395 ;
        RECT 57.635 -166.085 57.965 -165.755 ;
        RECT 57.635 -167.445 57.965 -167.115 ;
        RECT 57.635 -168.805 57.965 -168.475 ;
        RECT 57.635 -170.165 57.965 -169.835 ;
        RECT 57.635 -171.525 57.965 -171.195 ;
        RECT 57.635 -172.885 57.965 -172.555 ;
        RECT 57.635 -174.245 57.965 -173.915 ;
        RECT 57.635 -175.605 57.965 -175.275 ;
        RECT 57.635 -176.965 57.965 -176.635 ;
        RECT 57.635 -178.325 57.965 -177.995 ;
        RECT 57.635 -179.685 57.965 -179.355 ;
        RECT 57.635 -181.93 57.965 -180.8 ;
        RECT 57.64 -182.045 57.96 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 57.81 -98.075 58.14 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 241.32 59.325 242.45 ;
        RECT 58.995 239.195 59.325 239.525 ;
        RECT 58.995 237.835 59.325 238.165 ;
        RECT 59 237.16 59.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 58.995 -1.525 59.325 -1.195 ;
        RECT 58.995 -2.885 59.325 -2.555 ;
        RECT 59 -3.56 59.32 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 241.32 60.685 242.45 ;
        RECT 60.355 239.195 60.685 239.525 ;
        RECT 60.355 237.835 60.685 238.165 ;
        RECT 60.36 237.16 60.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 60.355 -1.525 60.685 -1.195 ;
        RECT 60.355 -2.885 60.685 -2.555 ;
        RECT 60.36 -3.56 60.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 241.32 62.045 242.45 ;
        RECT 61.715 239.195 62.045 239.525 ;
        RECT 61.715 237.835 62.045 238.165 ;
        RECT 61.72 237.16 62.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 -1.525 62.045 -1.195 ;
        RECT 61.715 -2.885 62.045 -2.555 ;
        RECT 61.72 -3.56 62.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 61.715 -95.365 62.045 -95.035 ;
        RECT 61.715 -96.725 62.045 -96.395 ;
        RECT 61.715 -98.085 62.045 -97.755 ;
        RECT 61.715 -99.445 62.045 -99.115 ;
        RECT 61.715 -100.805 62.045 -100.475 ;
        RECT 61.715 -102.165 62.045 -101.835 ;
        RECT 61.715 -103.525 62.045 -103.195 ;
        RECT 61.715 -104.885 62.045 -104.555 ;
        RECT 61.715 -106.245 62.045 -105.915 ;
        RECT 61.715 -107.605 62.045 -107.275 ;
        RECT 61.715 -108.965 62.045 -108.635 ;
        RECT 61.715 -110.325 62.045 -109.995 ;
        RECT 61.715 -111.685 62.045 -111.355 ;
        RECT 61.715 -113.045 62.045 -112.715 ;
        RECT 61.715 -114.405 62.045 -114.075 ;
        RECT 61.715 -115.765 62.045 -115.435 ;
        RECT 61.715 -117.125 62.045 -116.795 ;
        RECT 61.715 -118.485 62.045 -118.155 ;
        RECT 61.715 -119.845 62.045 -119.515 ;
        RECT 61.715 -121.205 62.045 -120.875 ;
        RECT 61.715 -122.565 62.045 -122.235 ;
        RECT 61.715 -123.925 62.045 -123.595 ;
        RECT 61.715 -125.285 62.045 -124.955 ;
        RECT 61.715 -126.645 62.045 -126.315 ;
        RECT 61.715 -128.005 62.045 -127.675 ;
        RECT 61.715 -129.365 62.045 -129.035 ;
        RECT 61.715 -130.725 62.045 -130.395 ;
        RECT 61.715 -132.085 62.045 -131.755 ;
        RECT 61.715 -133.445 62.045 -133.115 ;
        RECT 61.715 -134.805 62.045 -134.475 ;
        RECT 61.715 -136.165 62.045 -135.835 ;
        RECT 61.715 -137.525 62.045 -137.195 ;
        RECT 61.715 -138.885 62.045 -138.555 ;
        RECT 61.715 -140.245 62.045 -139.915 ;
        RECT 61.715 -141.605 62.045 -141.275 ;
        RECT 61.715 -142.965 62.045 -142.635 ;
        RECT 61.715 -144.325 62.045 -143.995 ;
        RECT 61.715 -145.685 62.045 -145.355 ;
        RECT 61.715 -147.045 62.045 -146.715 ;
        RECT 61.715 -148.405 62.045 -148.075 ;
        RECT 61.715 -149.765 62.045 -149.435 ;
        RECT 61.715 -151.125 62.045 -150.795 ;
        RECT 61.715 -152.485 62.045 -152.155 ;
        RECT 61.715 -153.845 62.045 -153.515 ;
        RECT 61.715 -155.205 62.045 -154.875 ;
        RECT 61.715 -156.565 62.045 -156.235 ;
        RECT 61.715 -157.925 62.045 -157.595 ;
        RECT 61.715 -159.285 62.045 -158.955 ;
        RECT 61.715 -160.645 62.045 -160.315 ;
        RECT 61.715 -162.005 62.045 -161.675 ;
        RECT 61.715 -163.365 62.045 -163.035 ;
        RECT 61.715 -164.725 62.045 -164.395 ;
        RECT 61.715 -166.085 62.045 -165.755 ;
        RECT 61.715 -167.445 62.045 -167.115 ;
        RECT 61.715 -168.805 62.045 -168.475 ;
        RECT 61.715 -170.165 62.045 -169.835 ;
        RECT 61.715 -171.525 62.045 -171.195 ;
        RECT 61.715 -172.885 62.045 -172.555 ;
        RECT 61.715 -174.245 62.045 -173.915 ;
        RECT 61.715 -175.605 62.045 -175.275 ;
        RECT 61.715 -176.965 62.045 -176.635 ;
        RECT 61.715 -178.325 62.045 -177.995 ;
        RECT 61.715 -179.685 62.045 -179.355 ;
        RECT 61.715 -181.93 62.045 -180.8 ;
        RECT 61.72 -182.045 62.04 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 241.32 63.405 242.45 ;
        RECT 63.075 239.195 63.405 239.525 ;
        RECT 63.075 237.835 63.405 238.165 ;
        RECT 63.08 237.16 63.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 -1.525 63.405 -1.195 ;
        RECT 63.075 -2.885 63.405 -2.555 ;
        RECT 63.08 -3.56 63.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 63.075 -95.365 63.405 -95.035 ;
        RECT 63.075 -96.725 63.405 -96.395 ;
        RECT 63.075 -98.085 63.405 -97.755 ;
        RECT 63.075 -99.445 63.405 -99.115 ;
        RECT 63.075 -100.805 63.405 -100.475 ;
        RECT 63.075 -102.165 63.405 -101.835 ;
        RECT 63.075 -103.525 63.405 -103.195 ;
        RECT 63.075 -104.885 63.405 -104.555 ;
        RECT 63.075 -106.245 63.405 -105.915 ;
        RECT 63.075 -107.605 63.405 -107.275 ;
        RECT 63.075 -108.965 63.405 -108.635 ;
        RECT 63.075 -110.325 63.405 -109.995 ;
        RECT 63.075 -111.685 63.405 -111.355 ;
        RECT 63.075 -113.045 63.405 -112.715 ;
        RECT 63.075 -114.405 63.405 -114.075 ;
        RECT 63.075 -115.765 63.405 -115.435 ;
        RECT 63.075 -117.125 63.405 -116.795 ;
        RECT 63.075 -118.485 63.405 -118.155 ;
        RECT 63.075 -119.845 63.405 -119.515 ;
        RECT 63.075 -121.205 63.405 -120.875 ;
        RECT 63.075 -122.565 63.405 -122.235 ;
        RECT 63.075 -123.925 63.405 -123.595 ;
        RECT 63.075 -125.285 63.405 -124.955 ;
        RECT 63.075 -126.645 63.405 -126.315 ;
        RECT 63.075 -128.005 63.405 -127.675 ;
        RECT 63.075 -129.365 63.405 -129.035 ;
        RECT 63.075 -130.725 63.405 -130.395 ;
        RECT 63.075 -132.085 63.405 -131.755 ;
        RECT 63.075 -133.445 63.405 -133.115 ;
        RECT 63.075 -134.805 63.405 -134.475 ;
        RECT 63.075 -136.165 63.405 -135.835 ;
        RECT 63.075 -137.525 63.405 -137.195 ;
        RECT 63.075 -138.885 63.405 -138.555 ;
        RECT 63.075 -140.245 63.405 -139.915 ;
        RECT 63.075 -141.605 63.405 -141.275 ;
        RECT 63.075 -142.965 63.405 -142.635 ;
        RECT 63.075 -144.325 63.405 -143.995 ;
        RECT 63.075 -145.685 63.405 -145.355 ;
        RECT 63.075 -147.045 63.405 -146.715 ;
        RECT 63.075 -148.405 63.405 -148.075 ;
        RECT 63.075 -149.765 63.405 -149.435 ;
        RECT 63.075 -151.125 63.405 -150.795 ;
        RECT 63.075 -152.485 63.405 -152.155 ;
        RECT 63.075 -153.845 63.405 -153.515 ;
        RECT 63.075 -155.205 63.405 -154.875 ;
        RECT 63.075 -156.565 63.405 -156.235 ;
        RECT 63.075 -157.925 63.405 -157.595 ;
        RECT 63.075 -159.285 63.405 -158.955 ;
        RECT 63.075 -160.645 63.405 -160.315 ;
        RECT 63.075 -162.005 63.405 -161.675 ;
        RECT 63.075 -163.365 63.405 -163.035 ;
        RECT 63.075 -164.725 63.405 -164.395 ;
        RECT 63.075 -166.085 63.405 -165.755 ;
        RECT 63.075 -167.445 63.405 -167.115 ;
        RECT 63.075 -168.805 63.405 -168.475 ;
        RECT 63.075 -170.165 63.405 -169.835 ;
        RECT 63.075 -171.525 63.405 -171.195 ;
        RECT 63.075 -172.885 63.405 -172.555 ;
        RECT 63.075 -174.245 63.405 -173.915 ;
        RECT 63.075 -175.605 63.405 -175.275 ;
        RECT 63.075 -176.965 63.405 -176.635 ;
        RECT 63.075 -178.325 63.405 -177.995 ;
        RECT 63.075 -179.685 63.405 -179.355 ;
        RECT 63.075 -181.93 63.405 -180.8 ;
        RECT 63.08 -182.045 63.4 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.435 241.32 64.765 242.45 ;
        RECT 64.435 239.195 64.765 239.525 ;
        RECT 64.435 237.835 64.765 238.165 ;
        RECT 64.44 237.16 64.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.435 -1.525 64.765 -1.195 ;
        RECT 64.435 -2.885 64.765 -2.555 ;
        RECT 64.44 -3.56 64.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 64.435 -95.365 64.765 -95.035 ;
        RECT 64.435 -96.725 64.765 -96.395 ;
        RECT 64.435 -98.085 64.765 -97.755 ;
        RECT 64.435 -99.445 64.765 -99.115 ;
        RECT 64.435 -100.805 64.765 -100.475 ;
        RECT 64.435 -102.165 64.765 -101.835 ;
        RECT 64.435 -103.525 64.765 -103.195 ;
        RECT 64.435 -104.885 64.765 -104.555 ;
        RECT 64.435 -106.245 64.765 -105.915 ;
        RECT 64.435 -107.605 64.765 -107.275 ;
        RECT 64.435 -108.965 64.765 -108.635 ;
        RECT 64.435 -110.325 64.765 -109.995 ;
        RECT 64.435 -111.685 64.765 -111.355 ;
        RECT 64.435 -113.045 64.765 -112.715 ;
        RECT 64.435 -114.405 64.765 -114.075 ;
        RECT 64.435 -115.765 64.765 -115.435 ;
        RECT 64.435 -117.125 64.765 -116.795 ;
        RECT 64.435 -118.485 64.765 -118.155 ;
        RECT 64.435 -119.845 64.765 -119.515 ;
        RECT 64.435 -121.205 64.765 -120.875 ;
        RECT 64.435 -122.565 64.765 -122.235 ;
        RECT 64.435 -123.925 64.765 -123.595 ;
        RECT 64.435 -125.285 64.765 -124.955 ;
        RECT 64.435 -126.645 64.765 -126.315 ;
        RECT 64.435 -128.005 64.765 -127.675 ;
        RECT 64.435 -129.365 64.765 -129.035 ;
        RECT 64.435 -130.725 64.765 -130.395 ;
        RECT 64.435 -132.085 64.765 -131.755 ;
        RECT 64.435 -133.445 64.765 -133.115 ;
        RECT 64.435 -134.805 64.765 -134.475 ;
        RECT 64.435 -136.165 64.765 -135.835 ;
        RECT 64.435 -137.525 64.765 -137.195 ;
        RECT 64.435 -138.885 64.765 -138.555 ;
        RECT 64.435 -140.245 64.765 -139.915 ;
        RECT 64.435 -141.605 64.765 -141.275 ;
        RECT 64.435 -142.965 64.765 -142.635 ;
        RECT 64.435 -144.325 64.765 -143.995 ;
        RECT 64.435 -145.685 64.765 -145.355 ;
        RECT 64.435 -147.045 64.765 -146.715 ;
        RECT 64.435 -148.405 64.765 -148.075 ;
        RECT 64.435 -149.765 64.765 -149.435 ;
        RECT 64.435 -151.125 64.765 -150.795 ;
        RECT 64.435 -152.485 64.765 -152.155 ;
        RECT 64.435 -153.845 64.765 -153.515 ;
        RECT 64.435 -155.205 64.765 -154.875 ;
        RECT 64.435 -156.565 64.765 -156.235 ;
        RECT 64.435 -157.925 64.765 -157.595 ;
        RECT 64.435 -159.285 64.765 -158.955 ;
        RECT 64.435 -160.645 64.765 -160.315 ;
        RECT 64.435 -162.005 64.765 -161.675 ;
        RECT 64.435 -163.365 64.765 -163.035 ;
        RECT 64.435 -164.725 64.765 -164.395 ;
        RECT 64.435 -166.085 64.765 -165.755 ;
        RECT 64.435 -167.445 64.765 -167.115 ;
        RECT 64.435 -168.805 64.765 -168.475 ;
        RECT 64.435 -170.165 64.765 -169.835 ;
        RECT 64.435 -171.525 64.765 -171.195 ;
        RECT 64.435 -172.885 64.765 -172.555 ;
        RECT 64.435 -174.245 64.765 -173.915 ;
        RECT 64.435 -175.605 64.765 -175.275 ;
        RECT 64.435 -176.965 64.765 -176.635 ;
        RECT 64.435 -178.325 64.765 -177.995 ;
        RECT 64.435 -179.685 64.765 -179.355 ;
        RECT 64.435 -181.93 64.765 -180.8 ;
        RECT 64.44 -182.045 64.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 241.32 66.125 242.45 ;
        RECT 65.795 239.195 66.125 239.525 ;
        RECT 65.795 237.835 66.125 238.165 ;
        RECT 65.8 237.16 66.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 -1.525 66.125 -1.195 ;
        RECT 65.795 -2.885 66.125 -2.555 ;
        RECT 65.8 -3.56 66.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 65.795 -95.365 66.125 -95.035 ;
        RECT 65.795 -96.725 66.125 -96.395 ;
        RECT 65.795 -98.085 66.125 -97.755 ;
        RECT 65.795 -99.445 66.125 -99.115 ;
        RECT 65.795 -100.805 66.125 -100.475 ;
        RECT 65.795 -102.165 66.125 -101.835 ;
        RECT 65.795 -103.525 66.125 -103.195 ;
        RECT 65.795 -104.885 66.125 -104.555 ;
        RECT 65.795 -106.245 66.125 -105.915 ;
        RECT 65.795 -107.605 66.125 -107.275 ;
        RECT 65.795 -108.965 66.125 -108.635 ;
        RECT 65.795 -110.325 66.125 -109.995 ;
        RECT 65.795 -111.685 66.125 -111.355 ;
        RECT 65.795 -113.045 66.125 -112.715 ;
        RECT 65.795 -114.405 66.125 -114.075 ;
        RECT 65.795 -115.765 66.125 -115.435 ;
        RECT 65.795 -117.125 66.125 -116.795 ;
        RECT 65.795 -118.485 66.125 -118.155 ;
        RECT 65.795 -119.845 66.125 -119.515 ;
        RECT 65.795 -121.205 66.125 -120.875 ;
        RECT 65.795 -122.565 66.125 -122.235 ;
        RECT 65.795 -123.925 66.125 -123.595 ;
        RECT 65.795 -125.285 66.125 -124.955 ;
        RECT 65.795 -126.645 66.125 -126.315 ;
        RECT 65.795 -128.005 66.125 -127.675 ;
        RECT 65.795 -129.365 66.125 -129.035 ;
        RECT 65.795 -130.725 66.125 -130.395 ;
        RECT 65.795 -132.085 66.125 -131.755 ;
        RECT 65.795 -133.445 66.125 -133.115 ;
        RECT 65.795 -134.805 66.125 -134.475 ;
        RECT 65.795 -136.165 66.125 -135.835 ;
        RECT 65.795 -137.525 66.125 -137.195 ;
        RECT 65.795 -138.885 66.125 -138.555 ;
        RECT 65.795 -140.245 66.125 -139.915 ;
        RECT 65.795 -141.605 66.125 -141.275 ;
        RECT 65.795 -142.965 66.125 -142.635 ;
        RECT 65.795 -144.325 66.125 -143.995 ;
        RECT 65.795 -145.685 66.125 -145.355 ;
        RECT 65.795 -147.045 66.125 -146.715 ;
        RECT 65.795 -148.405 66.125 -148.075 ;
        RECT 65.795 -149.765 66.125 -149.435 ;
        RECT 65.795 -151.125 66.125 -150.795 ;
        RECT 65.795 -152.485 66.125 -152.155 ;
        RECT 65.795 -153.845 66.125 -153.515 ;
        RECT 65.795 -155.205 66.125 -154.875 ;
        RECT 65.795 -156.565 66.125 -156.235 ;
        RECT 65.795 -157.925 66.125 -157.595 ;
        RECT 65.795 -159.285 66.125 -158.955 ;
        RECT 65.795 -160.645 66.125 -160.315 ;
        RECT 65.795 -162.005 66.125 -161.675 ;
        RECT 65.795 -163.365 66.125 -163.035 ;
        RECT 65.795 -164.725 66.125 -164.395 ;
        RECT 65.795 -166.085 66.125 -165.755 ;
        RECT 65.795 -167.445 66.125 -167.115 ;
        RECT 65.795 -168.805 66.125 -168.475 ;
        RECT 65.795 -170.165 66.125 -169.835 ;
        RECT 65.795 -171.525 66.125 -171.195 ;
        RECT 65.795 -172.885 66.125 -172.555 ;
        RECT 65.795 -174.245 66.125 -173.915 ;
        RECT 65.795 -175.605 66.125 -175.275 ;
        RECT 65.795 -176.965 66.125 -176.635 ;
        RECT 65.795 -178.325 66.125 -177.995 ;
        RECT 65.795 -179.685 66.125 -179.355 ;
        RECT 65.795 -181.93 66.125 -180.8 ;
        RECT 65.8 -182.045 66.12 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 241.32 67.485 242.45 ;
        RECT 67.155 239.195 67.485 239.525 ;
        RECT 67.155 237.835 67.485 238.165 ;
        RECT 67.16 237.16 67.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 -1.525 67.485 -1.195 ;
        RECT 67.155 -2.885 67.485 -2.555 ;
        RECT 67.16 -3.56 67.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 67.155 -164.725 67.485 -164.395 ;
        RECT 67.155 -166.085 67.485 -165.755 ;
        RECT 67.155 -167.445 67.485 -167.115 ;
        RECT 67.155 -168.805 67.485 -168.475 ;
        RECT 67.155 -170.165 67.485 -169.835 ;
        RECT 67.155 -171.525 67.485 -171.195 ;
        RECT 67.155 -172.885 67.485 -172.555 ;
        RECT 67.155 -174.245 67.485 -173.915 ;
        RECT 67.155 -175.605 67.485 -175.275 ;
        RECT 67.155 -176.965 67.485 -176.635 ;
        RECT 67.155 -178.325 67.485 -177.995 ;
        RECT 67.155 -179.685 67.485 -179.355 ;
        RECT 67.155 -181.93 67.485 -180.8 ;
        RECT 67.16 -182.045 67.48 -95.035 ;
        RECT 67.155 -95.365 67.485 -95.035 ;
        RECT 67.155 -96.725 67.485 -96.395 ;
        RECT 67.155 -98.085 67.485 -97.755 ;
        RECT 67.155 -99.445 67.485 -99.115 ;
        RECT 67.155 -100.805 67.485 -100.475 ;
        RECT 67.155 -102.165 67.485 -101.835 ;
        RECT 67.155 -103.525 67.485 -103.195 ;
        RECT 67.155 -104.885 67.485 -104.555 ;
        RECT 67.155 -106.245 67.485 -105.915 ;
        RECT 67.155 -107.605 67.485 -107.275 ;
        RECT 67.155 -108.965 67.485 -108.635 ;
        RECT 67.155 -110.325 67.485 -109.995 ;
        RECT 67.155 -111.685 67.485 -111.355 ;
        RECT 67.155 -113.045 67.485 -112.715 ;
        RECT 67.155 -114.405 67.485 -114.075 ;
        RECT 67.155 -115.765 67.485 -115.435 ;
        RECT 67.155 -117.125 67.485 -116.795 ;
        RECT 67.155 -118.485 67.485 -118.155 ;
        RECT 67.155 -119.845 67.485 -119.515 ;
        RECT 67.155 -121.205 67.485 -120.875 ;
        RECT 67.155 -122.565 67.485 -122.235 ;
        RECT 67.155 -123.925 67.485 -123.595 ;
        RECT 67.155 -125.285 67.485 -124.955 ;
        RECT 67.155 -126.645 67.485 -126.315 ;
        RECT 67.155 -128.005 67.485 -127.675 ;
        RECT 67.155 -129.365 67.485 -129.035 ;
        RECT 67.155 -130.725 67.485 -130.395 ;
        RECT 67.155 -132.085 67.485 -131.755 ;
        RECT 67.155 -133.445 67.485 -133.115 ;
        RECT 67.155 -134.805 67.485 -134.475 ;
        RECT 67.155 -136.165 67.485 -135.835 ;
        RECT 67.155 -137.525 67.485 -137.195 ;
        RECT 67.155 -138.885 67.485 -138.555 ;
        RECT 67.155 -140.245 67.485 -139.915 ;
        RECT 67.155 -141.605 67.485 -141.275 ;
        RECT 67.155 -142.965 67.485 -142.635 ;
        RECT 67.155 -144.325 67.485 -143.995 ;
        RECT 67.155 -145.685 67.485 -145.355 ;
        RECT 67.155 -147.045 67.485 -146.715 ;
        RECT 67.155 -148.405 67.485 -148.075 ;
        RECT 67.155 -149.765 67.485 -149.435 ;
        RECT 67.155 -151.125 67.485 -150.795 ;
        RECT 67.155 -152.485 67.485 -152.155 ;
        RECT 67.155 -153.845 67.485 -153.515 ;
        RECT 67.155 -155.205 67.485 -154.875 ;
        RECT 67.155 -156.565 67.485 -156.235 ;
        RECT 67.155 -157.925 67.485 -157.595 ;
        RECT 67.155 -159.285 67.485 -158.955 ;
        RECT 67.155 -160.645 67.485 -160.315 ;
        RECT 67.155 -162.005 67.485 -161.675 ;
        RECT 67.155 -163.365 67.485 -163.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 -1.525 19.885 -1.195 ;
        RECT 19.555 -2.885 19.885 -2.555 ;
        RECT 19.56 -3.56 19.88 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.555 -95.365 19.885 -95.035 ;
        RECT 19.555 -96.725 19.885 -96.395 ;
        RECT 19.555 -98.085 19.885 -97.755 ;
        RECT 19.555 -99.445 19.885 -99.115 ;
        RECT 19.555 -100.805 19.885 -100.475 ;
        RECT 19.555 -102.165 19.885 -101.835 ;
        RECT 19.555 -103.525 19.885 -103.195 ;
        RECT 19.555 -104.885 19.885 -104.555 ;
        RECT 19.555 -106.245 19.885 -105.915 ;
        RECT 19.555 -107.605 19.885 -107.275 ;
        RECT 19.555 -108.965 19.885 -108.635 ;
        RECT 19.555 -110.325 19.885 -109.995 ;
        RECT 19.555 -111.685 19.885 -111.355 ;
        RECT 19.555 -113.045 19.885 -112.715 ;
        RECT 19.555 -114.405 19.885 -114.075 ;
        RECT 19.555 -115.765 19.885 -115.435 ;
        RECT 19.555 -117.125 19.885 -116.795 ;
        RECT 19.555 -118.485 19.885 -118.155 ;
        RECT 19.555 -119.845 19.885 -119.515 ;
        RECT 19.555 -121.205 19.885 -120.875 ;
        RECT 19.555 -122.565 19.885 -122.235 ;
        RECT 19.555 -123.925 19.885 -123.595 ;
        RECT 19.555 -125.285 19.885 -124.955 ;
        RECT 19.555 -126.645 19.885 -126.315 ;
        RECT 19.555 -128.005 19.885 -127.675 ;
        RECT 19.555 -129.365 19.885 -129.035 ;
        RECT 19.555 -130.725 19.885 -130.395 ;
        RECT 19.555 -132.085 19.885 -131.755 ;
        RECT 19.555 -133.445 19.885 -133.115 ;
        RECT 19.555 -134.805 19.885 -134.475 ;
        RECT 19.555 -136.165 19.885 -135.835 ;
        RECT 19.555 -137.525 19.885 -137.195 ;
        RECT 19.555 -138.885 19.885 -138.555 ;
        RECT 19.555 -140.245 19.885 -139.915 ;
        RECT 19.555 -141.605 19.885 -141.275 ;
        RECT 19.555 -142.965 19.885 -142.635 ;
        RECT 19.555 -144.325 19.885 -143.995 ;
        RECT 19.555 -145.685 19.885 -145.355 ;
        RECT 19.555 -147.045 19.885 -146.715 ;
        RECT 19.555 -148.405 19.885 -148.075 ;
        RECT 19.555 -149.765 19.885 -149.435 ;
        RECT 19.555 -151.125 19.885 -150.795 ;
        RECT 19.555 -152.485 19.885 -152.155 ;
        RECT 19.555 -153.845 19.885 -153.515 ;
        RECT 19.555 -155.205 19.885 -154.875 ;
        RECT 19.555 -156.565 19.885 -156.235 ;
        RECT 19.555 -157.925 19.885 -157.595 ;
        RECT 19.555 -159.285 19.885 -158.955 ;
        RECT 19.555 -160.645 19.885 -160.315 ;
        RECT 19.555 -162.005 19.885 -161.675 ;
        RECT 19.555 -163.365 19.885 -163.035 ;
        RECT 19.555 -164.725 19.885 -164.395 ;
        RECT 19.555 -166.085 19.885 -165.755 ;
        RECT 19.555 -167.445 19.885 -167.115 ;
        RECT 19.555 -168.805 19.885 -168.475 ;
        RECT 19.555 -170.165 19.885 -169.835 ;
        RECT 19.555 -171.525 19.885 -171.195 ;
        RECT 19.555 -172.885 19.885 -172.555 ;
        RECT 19.555 -174.245 19.885 -173.915 ;
        RECT 19.555 -175.605 19.885 -175.275 ;
        RECT 19.555 -176.965 19.885 -176.635 ;
        RECT 19.555 -178.325 19.885 -177.995 ;
        RECT 19.555 -179.685 19.885 -179.355 ;
        RECT 19.555 -181.93 19.885 -180.8 ;
        RECT 19.56 -182.045 19.88 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 241.32 21.245 242.45 ;
        RECT 20.915 239.195 21.245 239.525 ;
        RECT 20.915 237.835 21.245 238.165 ;
        RECT 20.92 237.16 21.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 -1.525 21.245 -1.195 ;
        RECT 20.915 -2.885 21.245 -2.555 ;
        RECT 20.92 -3.56 21.24 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 20.915 -95.365 21.245 -95.035 ;
        RECT 20.915 -96.725 21.245 -96.395 ;
        RECT 20.915 -98.085 21.245 -97.755 ;
        RECT 20.915 -99.445 21.245 -99.115 ;
        RECT 20.915 -100.805 21.245 -100.475 ;
        RECT 20.915 -102.165 21.245 -101.835 ;
        RECT 20.915 -103.525 21.245 -103.195 ;
        RECT 20.915 -104.885 21.245 -104.555 ;
        RECT 20.915 -106.245 21.245 -105.915 ;
        RECT 20.915 -107.605 21.245 -107.275 ;
        RECT 20.915 -108.965 21.245 -108.635 ;
        RECT 20.915 -110.325 21.245 -109.995 ;
        RECT 20.915 -111.685 21.245 -111.355 ;
        RECT 20.915 -113.045 21.245 -112.715 ;
        RECT 20.915 -114.405 21.245 -114.075 ;
        RECT 20.915 -115.765 21.245 -115.435 ;
        RECT 20.915 -117.125 21.245 -116.795 ;
        RECT 20.915 -118.485 21.245 -118.155 ;
        RECT 20.915 -119.845 21.245 -119.515 ;
        RECT 20.915 -121.205 21.245 -120.875 ;
        RECT 20.915 -122.565 21.245 -122.235 ;
        RECT 20.915 -123.925 21.245 -123.595 ;
        RECT 20.915 -125.285 21.245 -124.955 ;
        RECT 20.915 -126.645 21.245 -126.315 ;
        RECT 20.915 -128.005 21.245 -127.675 ;
        RECT 20.915 -129.365 21.245 -129.035 ;
        RECT 20.915 -130.725 21.245 -130.395 ;
        RECT 20.915 -132.085 21.245 -131.755 ;
        RECT 20.915 -133.445 21.245 -133.115 ;
        RECT 20.915 -134.805 21.245 -134.475 ;
        RECT 20.915 -136.165 21.245 -135.835 ;
        RECT 20.915 -137.525 21.245 -137.195 ;
        RECT 20.915 -138.885 21.245 -138.555 ;
        RECT 20.915 -140.245 21.245 -139.915 ;
        RECT 20.915 -141.605 21.245 -141.275 ;
        RECT 20.915 -142.965 21.245 -142.635 ;
        RECT 20.915 -144.325 21.245 -143.995 ;
        RECT 20.915 -145.685 21.245 -145.355 ;
        RECT 20.915 -147.045 21.245 -146.715 ;
        RECT 20.915 -148.405 21.245 -148.075 ;
        RECT 20.915 -149.765 21.245 -149.435 ;
        RECT 20.915 -151.125 21.245 -150.795 ;
        RECT 20.915 -152.485 21.245 -152.155 ;
        RECT 20.915 -153.845 21.245 -153.515 ;
        RECT 20.915 -155.205 21.245 -154.875 ;
        RECT 20.915 -156.565 21.245 -156.235 ;
        RECT 20.915 -157.925 21.245 -157.595 ;
        RECT 20.915 -159.285 21.245 -158.955 ;
        RECT 20.915 -160.645 21.245 -160.315 ;
        RECT 20.915 -162.005 21.245 -161.675 ;
        RECT 20.915 -163.365 21.245 -163.035 ;
        RECT 20.915 -164.725 21.245 -164.395 ;
        RECT 20.915 -166.085 21.245 -165.755 ;
        RECT 20.915 -167.445 21.245 -167.115 ;
        RECT 20.915 -168.805 21.245 -168.475 ;
        RECT 20.915 -170.165 21.245 -169.835 ;
        RECT 20.915 -171.525 21.245 -171.195 ;
        RECT 20.915 -172.885 21.245 -172.555 ;
        RECT 20.915 -174.245 21.245 -173.915 ;
        RECT 20.915 -175.605 21.245 -175.275 ;
        RECT 20.915 -176.965 21.245 -176.635 ;
        RECT 20.915 -178.325 21.245 -177.995 ;
        RECT 20.915 -179.685 21.245 -179.355 ;
        RECT 20.915 -181.93 21.245 -180.8 ;
        RECT 20.92 -182.045 21.24 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 241.32 22.605 242.45 ;
        RECT 22.275 239.195 22.605 239.525 ;
        RECT 22.275 237.835 22.605 238.165 ;
        RECT 22.28 237.16 22.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 -1.525 22.605 -1.195 ;
        RECT 22.275 -2.885 22.605 -2.555 ;
        RECT 22.28 -3.56 22.6 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 22.275 -95.365 22.605 -95.035 ;
        RECT 22.275 -96.725 22.605 -96.395 ;
        RECT 22.275 -98.085 22.605 -97.755 ;
        RECT 22.275 -99.445 22.605 -99.115 ;
        RECT 22.275 -100.805 22.605 -100.475 ;
        RECT 22.275 -102.165 22.605 -101.835 ;
        RECT 22.275 -103.525 22.605 -103.195 ;
        RECT 22.275 -104.885 22.605 -104.555 ;
        RECT 22.275 -106.245 22.605 -105.915 ;
        RECT 22.275 -107.605 22.605 -107.275 ;
        RECT 22.275 -108.965 22.605 -108.635 ;
        RECT 22.275 -110.325 22.605 -109.995 ;
        RECT 22.275 -111.685 22.605 -111.355 ;
        RECT 22.275 -113.045 22.605 -112.715 ;
        RECT 22.275 -114.405 22.605 -114.075 ;
        RECT 22.275 -115.765 22.605 -115.435 ;
        RECT 22.275 -117.125 22.605 -116.795 ;
        RECT 22.275 -118.485 22.605 -118.155 ;
        RECT 22.275 -119.845 22.605 -119.515 ;
        RECT 22.275 -121.205 22.605 -120.875 ;
        RECT 22.275 -122.565 22.605 -122.235 ;
        RECT 22.275 -123.925 22.605 -123.595 ;
        RECT 22.275 -125.285 22.605 -124.955 ;
        RECT 22.275 -126.645 22.605 -126.315 ;
        RECT 22.275 -128.005 22.605 -127.675 ;
        RECT 22.275 -129.365 22.605 -129.035 ;
        RECT 22.275 -130.725 22.605 -130.395 ;
        RECT 22.275 -132.085 22.605 -131.755 ;
        RECT 22.275 -133.445 22.605 -133.115 ;
        RECT 22.275 -134.805 22.605 -134.475 ;
        RECT 22.275 -136.165 22.605 -135.835 ;
        RECT 22.275 -137.525 22.605 -137.195 ;
        RECT 22.275 -138.885 22.605 -138.555 ;
        RECT 22.275 -140.245 22.605 -139.915 ;
        RECT 22.275 -141.605 22.605 -141.275 ;
        RECT 22.275 -142.965 22.605 -142.635 ;
        RECT 22.275 -144.325 22.605 -143.995 ;
        RECT 22.275 -145.685 22.605 -145.355 ;
        RECT 22.275 -147.045 22.605 -146.715 ;
        RECT 22.275 -148.405 22.605 -148.075 ;
        RECT 22.275 -149.765 22.605 -149.435 ;
        RECT 22.275 -151.125 22.605 -150.795 ;
        RECT 22.275 -152.485 22.605 -152.155 ;
        RECT 22.275 -153.845 22.605 -153.515 ;
        RECT 22.275 -155.205 22.605 -154.875 ;
        RECT 22.275 -156.565 22.605 -156.235 ;
        RECT 22.275 -157.925 22.605 -157.595 ;
        RECT 22.275 -159.285 22.605 -158.955 ;
        RECT 22.275 -160.645 22.605 -160.315 ;
        RECT 22.275 -162.005 22.605 -161.675 ;
        RECT 22.275 -163.365 22.605 -163.035 ;
        RECT 22.275 -164.725 22.605 -164.395 ;
        RECT 22.275 -166.085 22.605 -165.755 ;
        RECT 22.275 -167.445 22.605 -167.115 ;
        RECT 22.275 -168.805 22.605 -168.475 ;
        RECT 22.275 -170.165 22.605 -169.835 ;
        RECT 22.275 -171.525 22.605 -171.195 ;
        RECT 22.275 -172.885 22.605 -172.555 ;
        RECT 22.275 -174.245 22.605 -173.915 ;
        RECT 22.275 -175.605 22.605 -175.275 ;
        RECT 22.275 -176.965 22.605 -176.635 ;
        RECT 22.275 -178.325 22.605 -177.995 ;
        RECT 22.275 -179.685 22.605 -179.355 ;
        RECT 22.275 -181.93 22.605 -180.8 ;
        RECT 22.28 -182.045 22.6 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 241.32 23.965 242.45 ;
        RECT 23.635 239.195 23.965 239.525 ;
        RECT 23.635 237.835 23.965 238.165 ;
        RECT 23.64 237.16 23.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 -1.525 23.965 -1.195 ;
        RECT 23.635 -2.885 23.965 -2.555 ;
        RECT 23.64 -3.56 23.96 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 23.635 -95.365 23.965 -95.035 ;
        RECT 23.635 -96.725 23.965 -96.395 ;
        RECT 23.635 -98.085 23.965 -97.755 ;
        RECT 23.635 -99.445 23.965 -99.115 ;
        RECT 23.635 -100.805 23.965 -100.475 ;
        RECT 23.635 -102.165 23.965 -101.835 ;
        RECT 23.635 -103.525 23.965 -103.195 ;
        RECT 23.635 -104.885 23.965 -104.555 ;
        RECT 23.635 -106.245 23.965 -105.915 ;
        RECT 23.635 -107.605 23.965 -107.275 ;
        RECT 23.635 -108.965 23.965 -108.635 ;
        RECT 23.635 -110.325 23.965 -109.995 ;
        RECT 23.635 -111.685 23.965 -111.355 ;
        RECT 23.635 -113.045 23.965 -112.715 ;
        RECT 23.635 -114.405 23.965 -114.075 ;
        RECT 23.635 -115.765 23.965 -115.435 ;
        RECT 23.635 -117.125 23.965 -116.795 ;
        RECT 23.635 -118.485 23.965 -118.155 ;
        RECT 23.635 -119.845 23.965 -119.515 ;
        RECT 23.635 -121.205 23.965 -120.875 ;
        RECT 23.635 -122.565 23.965 -122.235 ;
        RECT 23.635 -123.925 23.965 -123.595 ;
        RECT 23.635 -125.285 23.965 -124.955 ;
        RECT 23.635 -126.645 23.965 -126.315 ;
        RECT 23.635 -128.005 23.965 -127.675 ;
        RECT 23.635 -129.365 23.965 -129.035 ;
        RECT 23.635 -130.725 23.965 -130.395 ;
        RECT 23.635 -132.085 23.965 -131.755 ;
        RECT 23.635 -133.445 23.965 -133.115 ;
        RECT 23.635 -134.805 23.965 -134.475 ;
        RECT 23.635 -136.165 23.965 -135.835 ;
        RECT 23.635 -137.525 23.965 -137.195 ;
        RECT 23.635 -138.885 23.965 -138.555 ;
        RECT 23.635 -140.245 23.965 -139.915 ;
        RECT 23.635 -141.605 23.965 -141.275 ;
        RECT 23.635 -142.965 23.965 -142.635 ;
        RECT 23.635 -144.325 23.965 -143.995 ;
        RECT 23.635 -145.685 23.965 -145.355 ;
        RECT 23.635 -147.045 23.965 -146.715 ;
        RECT 23.635 -148.405 23.965 -148.075 ;
        RECT 23.635 -149.765 23.965 -149.435 ;
        RECT 23.635 -151.125 23.965 -150.795 ;
        RECT 23.635 -152.485 23.965 -152.155 ;
        RECT 23.635 -153.845 23.965 -153.515 ;
        RECT 23.635 -155.205 23.965 -154.875 ;
        RECT 23.635 -156.565 23.965 -156.235 ;
        RECT 23.635 -157.925 23.965 -157.595 ;
        RECT 23.635 -159.285 23.965 -158.955 ;
        RECT 23.635 -160.645 23.965 -160.315 ;
        RECT 23.635 -162.005 23.965 -161.675 ;
        RECT 23.635 -163.365 23.965 -163.035 ;
        RECT 23.635 -164.725 23.965 -164.395 ;
        RECT 23.635 -166.085 23.965 -165.755 ;
        RECT 23.635 -167.445 23.965 -167.115 ;
        RECT 23.635 -168.805 23.965 -168.475 ;
        RECT 23.635 -170.165 23.965 -169.835 ;
        RECT 23.635 -171.525 23.965 -171.195 ;
        RECT 23.635 -172.885 23.965 -172.555 ;
        RECT 23.635 -174.245 23.965 -173.915 ;
        RECT 23.635 -175.605 23.965 -175.275 ;
        RECT 23.635 -176.965 23.965 -176.635 ;
        RECT 23.635 -178.325 23.965 -177.995 ;
        RECT 23.635 -179.685 23.965 -179.355 ;
        RECT 23.635 -181.93 23.965 -180.8 ;
        RECT 23.64 -182.045 23.96 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 241.32 25.325 242.45 ;
        RECT 24.995 239.195 25.325 239.525 ;
        RECT 24.995 237.835 25.325 238.165 ;
        RECT 25 237.16 25.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 24.995 -99.445 25.325 -99.115 ;
        RECT 24.995 -100.805 25.325 -100.475 ;
        RECT 24.995 -102.165 25.325 -101.835 ;
        RECT 24.995 -103.525 25.325 -103.195 ;
        RECT 24.995 -104.885 25.325 -104.555 ;
        RECT 24.995 -106.245 25.325 -105.915 ;
        RECT 24.995 -107.605 25.325 -107.275 ;
        RECT 24.995 -108.965 25.325 -108.635 ;
        RECT 24.995 -110.325 25.325 -109.995 ;
        RECT 24.995 -111.685 25.325 -111.355 ;
        RECT 24.995 -113.045 25.325 -112.715 ;
        RECT 24.995 -114.405 25.325 -114.075 ;
        RECT 24.995 -115.765 25.325 -115.435 ;
        RECT 24.995 -117.125 25.325 -116.795 ;
        RECT 24.995 -118.485 25.325 -118.155 ;
        RECT 24.995 -119.845 25.325 -119.515 ;
        RECT 24.995 -121.205 25.325 -120.875 ;
        RECT 24.995 -122.565 25.325 -122.235 ;
        RECT 24.995 -123.925 25.325 -123.595 ;
        RECT 24.995 -125.285 25.325 -124.955 ;
        RECT 24.995 -126.645 25.325 -126.315 ;
        RECT 24.995 -128.005 25.325 -127.675 ;
        RECT 24.995 -129.365 25.325 -129.035 ;
        RECT 24.995 -130.725 25.325 -130.395 ;
        RECT 24.995 -132.085 25.325 -131.755 ;
        RECT 24.995 -133.445 25.325 -133.115 ;
        RECT 24.995 -134.805 25.325 -134.475 ;
        RECT 24.995 -136.165 25.325 -135.835 ;
        RECT 24.995 -137.525 25.325 -137.195 ;
        RECT 24.995 -138.885 25.325 -138.555 ;
        RECT 24.995 -140.245 25.325 -139.915 ;
        RECT 24.995 -141.605 25.325 -141.275 ;
        RECT 24.995 -142.965 25.325 -142.635 ;
        RECT 24.995 -144.325 25.325 -143.995 ;
        RECT 24.995 -145.685 25.325 -145.355 ;
        RECT 24.995 -147.045 25.325 -146.715 ;
        RECT 24.995 -148.405 25.325 -148.075 ;
        RECT 24.995 -149.765 25.325 -149.435 ;
        RECT 24.995 -151.125 25.325 -150.795 ;
        RECT 24.995 -152.485 25.325 -152.155 ;
        RECT 24.995 -153.845 25.325 -153.515 ;
        RECT 24.995 -155.205 25.325 -154.875 ;
        RECT 24.995 -156.565 25.325 -156.235 ;
        RECT 24.995 -157.925 25.325 -157.595 ;
        RECT 24.995 -159.285 25.325 -158.955 ;
        RECT 24.995 -160.645 25.325 -160.315 ;
        RECT 24.995 -162.005 25.325 -161.675 ;
        RECT 24.995 -163.365 25.325 -163.035 ;
        RECT 24.995 -164.725 25.325 -164.395 ;
        RECT 24.995 -166.085 25.325 -165.755 ;
        RECT 24.995 -167.445 25.325 -167.115 ;
        RECT 24.995 -168.805 25.325 -168.475 ;
        RECT 24.995 -170.165 25.325 -169.835 ;
        RECT 24.995 -171.525 25.325 -171.195 ;
        RECT 24.995 -172.885 25.325 -172.555 ;
        RECT 24.995 -174.245 25.325 -173.915 ;
        RECT 24.995 -175.605 25.325 -175.275 ;
        RECT 24.995 -176.965 25.325 -176.635 ;
        RECT 24.995 -178.325 25.325 -177.995 ;
        RECT 24.995 -179.685 25.325 -179.355 ;
        RECT 24.995 -181.93 25.325 -180.8 ;
        RECT 25 -182.045 25.32 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 25.11 -98.075 25.44 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 241.32 26.685 242.45 ;
        RECT 26.355 239.195 26.685 239.525 ;
        RECT 26.355 237.835 26.685 238.165 ;
        RECT 26.36 237.16 26.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 26.355 -1.525 26.685 -1.195 ;
        RECT 26.355 -2.885 26.685 -2.555 ;
        RECT 26.36 -3.56 26.68 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 241.32 28.045 242.45 ;
        RECT 27.715 239.195 28.045 239.525 ;
        RECT 27.715 237.835 28.045 238.165 ;
        RECT 27.72 237.16 28.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 27.715 -1.525 28.045 -1.195 ;
        RECT 27.715 -2.885 28.045 -2.555 ;
        RECT 27.72 -3.56 28.04 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 241.32 29.405 242.45 ;
        RECT 29.075 239.195 29.405 239.525 ;
        RECT 29.075 237.835 29.405 238.165 ;
        RECT 29.08 237.16 29.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 -1.525 29.405 -1.195 ;
        RECT 29.075 -2.885 29.405 -2.555 ;
        RECT 29.08 -3.56 29.4 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 29.075 -95.365 29.405 -95.035 ;
        RECT 29.075 -96.725 29.405 -96.395 ;
        RECT 29.075 -98.085 29.405 -97.755 ;
        RECT 29.075 -99.445 29.405 -99.115 ;
        RECT 29.075 -100.805 29.405 -100.475 ;
        RECT 29.075 -102.165 29.405 -101.835 ;
        RECT 29.075 -103.525 29.405 -103.195 ;
        RECT 29.075 -104.885 29.405 -104.555 ;
        RECT 29.075 -106.245 29.405 -105.915 ;
        RECT 29.075 -107.605 29.405 -107.275 ;
        RECT 29.075 -108.965 29.405 -108.635 ;
        RECT 29.075 -110.325 29.405 -109.995 ;
        RECT 29.075 -111.685 29.405 -111.355 ;
        RECT 29.075 -113.045 29.405 -112.715 ;
        RECT 29.075 -114.405 29.405 -114.075 ;
        RECT 29.075 -115.765 29.405 -115.435 ;
        RECT 29.075 -117.125 29.405 -116.795 ;
        RECT 29.075 -118.485 29.405 -118.155 ;
        RECT 29.075 -119.845 29.405 -119.515 ;
        RECT 29.075 -121.205 29.405 -120.875 ;
        RECT 29.075 -122.565 29.405 -122.235 ;
        RECT 29.075 -123.925 29.405 -123.595 ;
        RECT 29.075 -125.285 29.405 -124.955 ;
        RECT 29.075 -126.645 29.405 -126.315 ;
        RECT 29.075 -128.005 29.405 -127.675 ;
        RECT 29.075 -129.365 29.405 -129.035 ;
        RECT 29.075 -130.725 29.405 -130.395 ;
        RECT 29.075 -132.085 29.405 -131.755 ;
        RECT 29.075 -133.445 29.405 -133.115 ;
        RECT 29.075 -134.805 29.405 -134.475 ;
        RECT 29.075 -136.165 29.405 -135.835 ;
        RECT 29.075 -137.525 29.405 -137.195 ;
        RECT 29.075 -138.885 29.405 -138.555 ;
        RECT 29.075 -140.245 29.405 -139.915 ;
        RECT 29.075 -141.605 29.405 -141.275 ;
        RECT 29.075 -142.965 29.405 -142.635 ;
        RECT 29.075 -144.325 29.405 -143.995 ;
        RECT 29.075 -145.685 29.405 -145.355 ;
        RECT 29.075 -147.045 29.405 -146.715 ;
        RECT 29.075 -148.405 29.405 -148.075 ;
        RECT 29.075 -149.765 29.405 -149.435 ;
        RECT 29.075 -151.125 29.405 -150.795 ;
        RECT 29.075 -152.485 29.405 -152.155 ;
        RECT 29.075 -153.845 29.405 -153.515 ;
        RECT 29.075 -155.205 29.405 -154.875 ;
        RECT 29.075 -156.565 29.405 -156.235 ;
        RECT 29.075 -157.925 29.405 -157.595 ;
        RECT 29.075 -159.285 29.405 -158.955 ;
        RECT 29.075 -160.645 29.405 -160.315 ;
        RECT 29.075 -162.005 29.405 -161.675 ;
        RECT 29.075 -163.365 29.405 -163.035 ;
        RECT 29.075 -164.725 29.405 -164.395 ;
        RECT 29.075 -166.085 29.405 -165.755 ;
        RECT 29.075 -167.445 29.405 -167.115 ;
        RECT 29.075 -168.805 29.405 -168.475 ;
        RECT 29.075 -170.165 29.405 -169.835 ;
        RECT 29.075 -171.525 29.405 -171.195 ;
        RECT 29.075 -172.885 29.405 -172.555 ;
        RECT 29.075 -174.245 29.405 -173.915 ;
        RECT 29.075 -175.605 29.405 -175.275 ;
        RECT 29.075 -176.965 29.405 -176.635 ;
        RECT 29.075 -178.325 29.405 -177.995 ;
        RECT 29.075 -179.685 29.405 -179.355 ;
        RECT 29.075 -181.93 29.405 -180.8 ;
        RECT 29.08 -182.045 29.4 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 241.32 30.765 242.45 ;
        RECT 30.435 239.195 30.765 239.525 ;
        RECT 30.435 237.835 30.765 238.165 ;
        RECT 30.44 237.16 30.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 -1.525 30.765 -1.195 ;
        RECT 30.435 -2.885 30.765 -2.555 ;
        RECT 30.44 -3.56 30.76 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 30.435 -95.365 30.765 -95.035 ;
        RECT 30.435 -96.725 30.765 -96.395 ;
        RECT 30.435 -98.085 30.765 -97.755 ;
        RECT 30.435 -99.445 30.765 -99.115 ;
        RECT 30.435 -100.805 30.765 -100.475 ;
        RECT 30.435 -102.165 30.765 -101.835 ;
        RECT 30.435 -103.525 30.765 -103.195 ;
        RECT 30.435 -104.885 30.765 -104.555 ;
        RECT 30.435 -106.245 30.765 -105.915 ;
        RECT 30.435 -107.605 30.765 -107.275 ;
        RECT 30.435 -108.965 30.765 -108.635 ;
        RECT 30.435 -110.325 30.765 -109.995 ;
        RECT 30.435 -111.685 30.765 -111.355 ;
        RECT 30.435 -113.045 30.765 -112.715 ;
        RECT 30.435 -114.405 30.765 -114.075 ;
        RECT 30.435 -115.765 30.765 -115.435 ;
        RECT 30.435 -117.125 30.765 -116.795 ;
        RECT 30.435 -118.485 30.765 -118.155 ;
        RECT 30.435 -119.845 30.765 -119.515 ;
        RECT 30.435 -121.205 30.765 -120.875 ;
        RECT 30.435 -122.565 30.765 -122.235 ;
        RECT 30.435 -123.925 30.765 -123.595 ;
        RECT 30.435 -125.285 30.765 -124.955 ;
        RECT 30.435 -126.645 30.765 -126.315 ;
        RECT 30.435 -128.005 30.765 -127.675 ;
        RECT 30.435 -129.365 30.765 -129.035 ;
        RECT 30.435 -130.725 30.765 -130.395 ;
        RECT 30.435 -132.085 30.765 -131.755 ;
        RECT 30.435 -133.445 30.765 -133.115 ;
        RECT 30.435 -134.805 30.765 -134.475 ;
        RECT 30.435 -136.165 30.765 -135.835 ;
        RECT 30.435 -137.525 30.765 -137.195 ;
        RECT 30.435 -138.885 30.765 -138.555 ;
        RECT 30.435 -140.245 30.765 -139.915 ;
        RECT 30.435 -141.605 30.765 -141.275 ;
        RECT 30.435 -142.965 30.765 -142.635 ;
        RECT 30.435 -144.325 30.765 -143.995 ;
        RECT 30.435 -145.685 30.765 -145.355 ;
        RECT 30.435 -147.045 30.765 -146.715 ;
        RECT 30.435 -148.405 30.765 -148.075 ;
        RECT 30.435 -149.765 30.765 -149.435 ;
        RECT 30.435 -151.125 30.765 -150.795 ;
        RECT 30.435 -152.485 30.765 -152.155 ;
        RECT 30.435 -153.845 30.765 -153.515 ;
        RECT 30.435 -155.205 30.765 -154.875 ;
        RECT 30.435 -156.565 30.765 -156.235 ;
        RECT 30.435 -157.925 30.765 -157.595 ;
        RECT 30.435 -159.285 30.765 -158.955 ;
        RECT 30.435 -160.645 30.765 -160.315 ;
        RECT 30.435 -162.005 30.765 -161.675 ;
        RECT 30.435 -163.365 30.765 -163.035 ;
        RECT 30.435 -164.725 30.765 -164.395 ;
        RECT 30.435 -166.085 30.765 -165.755 ;
        RECT 30.435 -167.445 30.765 -167.115 ;
        RECT 30.435 -168.805 30.765 -168.475 ;
        RECT 30.435 -170.165 30.765 -169.835 ;
        RECT 30.435 -171.525 30.765 -171.195 ;
        RECT 30.435 -172.885 30.765 -172.555 ;
        RECT 30.435 -174.245 30.765 -173.915 ;
        RECT 30.435 -175.605 30.765 -175.275 ;
        RECT 30.435 -176.965 30.765 -176.635 ;
        RECT 30.435 -178.325 30.765 -177.995 ;
        RECT 30.435 -179.685 30.765 -179.355 ;
        RECT 30.435 -181.93 30.765 -180.8 ;
        RECT 30.44 -182.045 30.76 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 241.32 32.125 242.45 ;
        RECT 31.795 239.195 32.125 239.525 ;
        RECT 31.795 237.835 32.125 238.165 ;
        RECT 31.8 237.16 32.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 -1.525 32.125 -1.195 ;
        RECT 31.795 -2.885 32.125 -2.555 ;
        RECT 31.8 -3.56 32.12 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 31.795 -95.365 32.125 -95.035 ;
        RECT 31.795 -96.725 32.125 -96.395 ;
        RECT 31.795 -98.085 32.125 -97.755 ;
        RECT 31.795 -99.445 32.125 -99.115 ;
        RECT 31.795 -100.805 32.125 -100.475 ;
        RECT 31.795 -102.165 32.125 -101.835 ;
        RECT 31.795 -103.525 32.125 -103.195 ;
        RECT 31.795 -104.885 32.125 -104.555 ;
        RECT 31.795 -106.245 32.125 -105.915 ;
        RECT 31.795 -107.605 32.125 -107.275 ;
        RECT 31.795 -108.965 32.125 -108.635 ;
        RECT 31.795 -110.325 32.125 -109.995 ;
        RECT 31.795 -111.685 32.125 -111.355 ;
        RECT 31.795 -113.045 32.125 -112.715 ;
        RECT 31.795 -114.405 32.125 -114.075 ;
        RECT 31.795 -115.765 32.125 -115.435 ;
        RECT 31.795 -117.125 32.125 -116.795 ;
        RECT 31.795 -118.485 32.125 -118.155 ;
        RECT 31.795 -119.845 32.125 -119.515 ;
        RECT 31.795 -121.205 32.125 -120.875 ;
        RECT 31.795 -122.565 32.125 -122.235 ;
        RECT 31.795 -123.925 32.125 -123.595 ;
        RECT 31.795 -125.285 32.125 -124.955 ;
        RECT 31.795 -126.645 32.125 -126.315 ;
        RECT 31.795 -128.005 32.125 -127.675 ;
        RECT 31.795 -129.365 32.125 -129.035 ;
        RECT 31.795 -130.725 32.125 -130.395 ;
        RECT 31.795 -132.085 32.125 -131.755 ;
        RECT 31.795 -133.445 32.125 -133.115 ;
        RECT 31.795 -134.805 32.125 -134.475 ;
        RECT 31.795 -136.165 32.125 -135.835 ;
        RECT 31.795 -137.525 32.125 -137.195 ;
        RECT 31.795 -138.885 32.125 -138.555 ;
        RECT 31.795 -140.245 32.125 -139.915 ;
        RECT 31.795 -141.605 32.125 -141.275 ;
        RECT 31.795 -142.965 32.125 -142.635 ;
        RECT 31.795 -144.325 32.125 -143.995 ;
        RECT 31.795 -145.685 32.125 -145.355 ;
        RECT 31.795 -147.045 32.125 -146.715 ;
        RECT 31.795 -148.405 32.125 -148.075 ;
        RECT 31.795 -149.765 32.125 -149.435 ;
        RECT 31.795 -151.125 32.125 -150.795 ;
        RECT 31.795 -152.485 32.125 -152.155 ;
        RECT 31.795 -153.845 32.125 -153.515 ;
        RECT 31.795 -155.205 32.125 -154.875 ;
        RECT 31.795 -156.565 32.125 -156.235 ;
        RECT 31.795 -157.925 32.125 -157.595 ;
        RECT 31.795 -159.285 32.125 -158.955 ;
        RECT 31.795 -160.645 32.125 -160.315 ;
        RECT 31.795 -162.005 32.125 -161.675 ;
        RECT 31.795 -163.365 32.125 -163.035 ;
        RECT 31.795 -164.725 32.125 -164.395 ;
        RECT 31.795 -166.085 32.125 -165.755 ;
        RECT 31.795 -167.445 32.125 -167.115 ;
        RECT 31.795 -168.805 32.125 -168.475 ;
        RECT 31.795 -170.165 32.125 -169.835 ;
        RECT 31.795 -171.525 32.125 -171.195 ;
        RECT 31.795 -172.885 32.125 -172.555 ;
        RECT 31.795 -174.245 32.125 -173.915 ;
        RECT 31.795 -175.605 32.125 -175.275 ;
        RECT 31.795 -176.965 32.125 -176.635 ;
        RECT 31.795 -178.325 32.125 -177.995 ;
        RECT 31.795 -179.685 32.125 -179.355 ;
        RECT 31.795 -181.93 32.125 -180.8 ;
        RECT 31.8 -182.045 32.12 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 241.32 33.485 242.45 ;
        RECT 33.155 239.195 33.485 239.525 ;
        RECT 33.155 237.835 33.485 238.165 ;
        RECT 33.16 237.16 33.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 -1.525 33.485 -1.195 ;
        RECT 33.155 -2.885 33.485 -2.555 ;
        RECT 33.16 -3.56 33.48 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 33.155 -95.365 33.485 -95.035 ;
        RECT 33.155 -96.725 33.485 -96.395 ;
        RECT 33.155 -98.085 33.485 -97.755 ;
        RECT 33.155 -99.445 33.485 -99.115 ;
        RECT 33.155 -100.805 33.485 -100.475 ;
        RECT 33.155 -102.165 33.485 -101.835 ;
        RECT 33.155 -103.525 33.485 -103.195 ;
        RECT 33.155 -104.885 33.485 -104.555 ;
        RECT 33.155 -106.245 33.485 -105.915 ;
        RECT 33.155 -107.605 33.485 -107.275 ;
        RECT 33.155 -108.965 33.485 -108.635 ;
        RECT 33.155 -110.325 33.485 -109.995 ;
        RECT 33.155 -111.685 33.485 -111.355 ;
        RECT 33.155 -113.045 33.485 -112.715 ;
        RECT 33.155 -114.405 33.485 -114.075 ;
        RECT 33.155 -115.765 33.485 -115.435 ;
        RECT 33.155 -117.125 33.485 -116.795 ;
        RECT 33.155 -118.485 33.485 -118.155 ;
        RECT 33.155 -119.845 33.485 -119.515 ;
        RECT 33.155 -121.205 33.485 -120.875 ;
        RECT 33.155 -122.565 33.485 -122.235 ;
        RECT 33.155 -123.925 33.485 -123.595 ;
        RECT 33.155 -125.285 33.485 -124.955 ;
        RECT 33.155 -126.645 33.485 -126.315 ;
        RECT 33.155 -128.005 33.485 -127.675 ;
        RECT 33.155 -129.365 33.485 -129.035 ;
        RECT 33.155 -130.725 33.485 -130.395 ;
        RECT 33.155 -132.085 33.485 -131.755 ;
        RECT 33.155 -133.445 33.485 -133.115 ;
        RECT 33.155 -134.805 33.485 -134.475 ;
        RECT 33.155 -136.165 33.485 -135.835 ;
        RECT 33.155 -137.525 33.485 -137.195 ;
        RECT 33.155 -138.885 33.485 -138.555 ;
        RECT 33.155 -140.245 33.485 -139.915 ;
        RECT 33.155 -141.605 33.485 -141.275 ;
        RECT 33.155 -142.965 33.485 -142.635 ;
        RECT 33.155 -144.325 33.485 -143.995 ;
        RECT 33.155 -145.685 33.485 -145.355 ;
        RECT 33.155 -147.045 33.485 -146.715 ;
        RECT 33.155 -148.405 33.485 -148.075 ;
        RECT 33.155 -149.765 33.485 -149.435 ;
        RECT 33.155 -151.125 33.485 -150.795 ;
        RECT 33.155 -152.485 33.485 -152.155 ;
        RECT 33.155 -153.845 33.485 -153.515 ;
        RECT 33.155 -155.205 33.485 -154.875 ;
        RECT 33.155 -156.565 33.485 -156.235 ;
        RECT 33.155 -157.925 33.485 -157.595 ;
        RECT 33.155 -159.285 33.485 -158.955 ;
        RECT 33.155 -160.645 33.485 -160.315 ;
        RECT 33.155 -162.005 33.485 -161.675 ;
        RECT 33.155 -163.365 33.485 -163.035 ;
        RECT 33.155 -164.725 33.485 -164.395 ;
        RECT 33.155 -166.085 33.485 -165.755 ;
        RECT 33.155 -167.445 33.485 -167.115 ;
        RECT 33.155 -168.805 33.485 -168.475 ;
        RECT 33.155 -170.165 33.485 -169.835 ;
        RECT 33.155 -171.525 33.485 -171.195 ;
        RECT 33.155 -172.885 33.485 -172.555 ;
        RECT 33.155 -174.245 33.485 -173.915 ;
        RECT 33.155 -175.605 33.485 -175.275 ;
        RECT 33.155 -176.965 33.485 -176.635 ;
        RECT 33.155 -178.325 33.485 -177.995 ;
        RECT 33.155 -179.685 33.485 -179.355 ;
        RECT 33.155 -181.93 33.485 -180.8 ;
        RECT 33.16 -182.045 33.48 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 241.32 34.845 242.45 ;
        RECT 34.515 239.195 34.845 239.525 ;
        RECT 34.515 237.835 34.845 238.165 ;
        RECT 34.52 237.16 34.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 -1.525 34.845 -1.195 ;
        RECT 34.515 -2.885 34.845 -2.555 ;
        RECT 34.52 -3.56 34.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 34.515 -95.365 34.845 -95.035 ;
        RECT 34.515 -96.725 34.845 -96.395 ;
        RECT 34.515 -98.085 34.845 -97.755 ;
        RECT 34.515 -99.445 34.845 -99.115 ;
        RECT 34.515 -100.805 34.845 -100.475 ;
        RECT 34.515 -102.165 34.845 -101.835 ;
        RECT 34.515 -103.525 34.845 -103.195 ;
        RECT 34.515 -104.885 34.845 -104.555 ;
        RECT 34.515 -106.245 34.845 -105.915 ;
        RECT 34.515 -107.605 34.845 -107.275 ;
        RECT 34.515 -108.965 34.845 -108.635 ;
        RECT 34.515 -110.325 34.845 -109.995 ;
        RECT 34.515 -111.685 34.845 -111.355 ;
        RECT 34.515 -113.045 34.845 -112.715 ;
        RECT 34.515 -114.405 34.845 -114.075 ;
        RECT 34.515 -115.765 34.845 -115.435 ;
        RECT 34.515 -117.125 34.845 -116.795 ;
        RECT 34.515 -118.485 34.845 -118.155 ;
        RECT 34.515 -119.845 34.845 -119.515 ;
        RECT 34.515 -121.205 34.845 -120.875 ;
        RECT 34.515 -122.565 34.845 -122.235 ;
        RECT 34.515 -123.925 34.845 -123.595 ;
        RECT 34.515 -125.285 34.845 -124.955 ;
        RECT 34.515 -126.645 34.845 -126.315 ;
        RECT 34.515 -128.005 34.845 -127.675 ;
        RECT 34.515 -129.365 34.845 -129.035 ;
        RECT 34.515 -130.725 34.845 -130.395 ;
        RECT 34.515 -132.085 34.845 -131.755 ;
        RECT 34.515 -133.445 34.845 -133.115 ;
        RECT 34.515 -134.805 34.845 -134.475 ;
        RECT 34.515 -136.165 34.845 -135.835 ;
        RECT 34.515 -137.525 34.845 -137.195 ;
        RECT 34.515 -138.885 34.845 -138.555 ;
        RECT 34.515 -140.245 34.845 -139.915 ;
        RECT 34.515 -141.605 34.845 -141.275 ;
        RECT 34.515 -142.965 34.845 -142.635 ;
        RECT 34.515 -144.325 34.845 -143.995 ;
        RECT 34.515 -145.685 34.845 -145.355 ;
        RECT 34.515 -147.045 34.845 -146.715 ;
        RECT 34.515 -148.405 34.845 -148.075 ;
        RECT 34.515 -149.765 34.845 -149.435 ;
        RECT 34.515 -151.125 34.845 -150.795 ;
        RECT 34.515 -152.485 34.845 -152.155 ;
        RECT 34.515 -153.845 34.845 -153.515 ;
        RECT 34.515 -155.205 34.845 -154.875 ;
        RECT 34.515 -156.565 34.845 -156.235 ;
        RECT 34.515 -157.925 34.845 -157.595 ;
        RECT 34.515 -159.285 34.845 -158.955 ;
        RECT 34.515 -160.645 34.845 -160.315 ;
        RECT 34.515 -162.005 34.845 -161.675 ;
        RECT 34.515 -163.365 34.845 -163.035 ;
        RECT 34.515 -164.725 34.845 -164.395 ;
        RECT 34.515 -166.085 34.845 -165.755 ;
        RECT 34.515 -167.445 34.845 -167.115 ;
        RECT 34.515 -168.805 34.845 -168.475 ;
        RECT 34.515 -170.165 34.845 -169.835 ;
        RECT 34.515 -171.525 34.845 -171.195 ;
        RECT 34.515 -172.885 34.845 -172.555 ;
        RECT 34.515 -174.245 34.845 -173.915 ;
        RECT 34.515 -175.605 34.845 -175.275 ;
        RECT 34.515 -176.965 34.845 -176.635 ;
        RECT 34.515 -178.325 34.845 -177.995 ;
        RECT 34.515 -179.685 34.845 -179.355 ;
        RECT 34.515 -181.93 34.845 -180.8 ;
        RECT 34.52 -182.045 34.84 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 241.32 36.205 242.45 ;
        RECT 35.875 239.195 36.205 239.525 ;
        RECT 35.875 237.835 36.205 238.165 ;
        RECT 35.88 237.16 36.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 35.875 -99.445 36.205 -99.115 ;
        RECT 35.875 -100.805 36.205 -100.475 ;
        RECT 35.875 -102.165 36.205 -101.835 ;
        RECT 35.875 -103.525 36.205 -103.195 ;
        RECT 35.875 -104.885 36.205 -104.555 ;
        RECT 35.875 -106.245 36.205 -105.915 ;
        RECT 35.875 -107.605 36.205 -107.275 ;
        RECT 35.875 -108.965 36.205 -108.635 ;
        RECT 35.875 -110.325 36.205 -109.995 ;
        RECT 35.875 -111.685 36.205 -111.355 ;
        RECT 35.875 -113.045 36.205 -112.715 ;
        RECT 35.875 -114.405 36.205 -114.075 ;
        RECT 35.875 -115.765 36.205 -115.435 ;
        RECT 35.875 -117.125 36.205 -116.795 ;
        RECT 35.875 -118.485 36.205 -118.155 ;
        RECT 35.875 -119.845 36.205 -119.515 ;
        RECT 35.875 -121.205 36.205 -120.875 ;
        RECT 35.875 -122.565 36.205 -122.235 ;
        RECT 35.875 -123.925 36.205 -123.595 ;
        RECT 35.875 -125.285 36.205 -124.955 ;
        RECT 35.875 -126.645 36.205 -126.315 ;
        RECT 35.875 -128.005 36.205 -127.675 ;
        RECT 35.875 -129.365 36.205 -129.035 ;
        RECT 35.875 -130.725 36.205 -130.395 ;
        RECT 35.875 -132.085 36.205 -131.755 ;
        RECT 35.875 -133.445 36.205 -133.115 ;
        RECT 35.875 -134.805 36.205 -134.475 ;
        RECT 35.875 -136.165 36.205 -135.835 ;
        RECT 35.875 -137.525 36.205 -137.195 ;
        RECT 35.875 -138.885 36.205 -138.555 ;
        RECT 35.875 -140.245 36.205 -139.915 ;
        RECT 35.875 -141.605 36.205 -141.275 ;
        RECT 35.875 -142.965 36.205 -142.635 ;
        RECT 35.875 -144.325 36.205 -143.995 ;
        RECT 35.875 -145.685 36.205 -145.355 ;
        RECT 35.875 -147.045 36.205 -146.715 ;
        RECT 35.875 -148.405 36.205 -148.075 ;
        RECT 35.875 -149.765 36.205 -149.435 ;
        RECT 35.875 -151.125 36.205 -150.795 ;
        RECT 35.875 -152.485 36.205 -152.155 ;
        RECT 35.875 -153.845 36.205 -153.515 ;
        RECT 35.875 -155.205 36.205 -154.875 ;
        RECT 35.875 -156.565 36.205 -156.235 ;
        RECT 35.875 -157.925 36.205 -157.595 ;
        RECT 35.875 -159.285 36.205 -158.955 ;
        RECT 35.875 -160.645 36.205 -160.315 ;
        RECT 35.875 -162.005 36.205 -161.675 ;
        RECT 35.875 -163.365 36.205 -163.035 ;
        RECT 35.875 -164.725 36.205 -164.395 ;
        RECT 35.875 -166.085 36.205 -165.755 ;
        RECT 35.875 -167.445 36.205 -167.115 ;
        RECT 35.875 -168.805 36.205 -168.475 ;
        RECT 35.875 -170.165 36.205 -169.835 ;
        RECT 35.875 -171.525 36.205 -171.195 ;
        RECT 35.875 -172.885 36.205 -172.555 ;
        RECT 35.875 -174.245 36.205 -173.915 ;
        RECT 35.875 -175.605 36.205 -175.275 ;
        RECT 35.875 -176.965 36.205 -176.635 ;
        RECT 35.875 -178.325 36.205 -177.995 ;
        RECT 35.875 -179.685 36.205 -179.355 ;
        RECT 35.875 -181.93 36.205 -180.8 ;
        RECT 35.88 -182.045 36.2 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 36.01 -98.075 36.34 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 241.32 37.565 242.45 ;
        RECT 37.235 239.195 37.565 239.525 ;
        RECT 37.235 237.835 37.565 238.165 ;
        RECT 37.24 237.16 37.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 37.235 -1.525 37.565 -1.195 ;
        RECT 37.235 -2.885 37.565 -2.555 ;
        RECT 37.24 -3.56 37.56 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 241.32 38.925 242.45 ;
        RECT 38.595 239.195 38.925 239.525 ;
        RECT 38.595 237.835 38.925 238.165 ;
        RECT 38.6 237.16 38.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 38.595 -1.525 38.925 -1.195 ;
        RECT 38.595 -2.885 38.925 -2.555 ;
        RECT 38.6 -3.56 38.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.955 241.32 40.285 242.45 ;
        RECT 39.955 239.195 40.285 239.525 ;
        RECT 39.955 237.835 40.285 238.165 ;
        RECT 39.96 237.16 40.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.955 -1.525 40.285 -1.195 ;
        RECT 39.955 -2.885 40.285 -2.555 ;
        RECT 39.96 -3.56 40.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 39.955 -95.365 40.285 -95.035 ;
        RECT 39.955 -96.725 40.285 -96.395 ;
        RECT 39.955 -98.085 40.285 -97.755 ;
        RECT 39.955 -99.445 40.285 -99.115 ;
        RECT 39.955 -100.805 40.285 -100.475 ;
        RECT 39.955 -102.165 40.285 -101.835 ;
        RECT 39.955 -103.525 40.285 -103.195 ;
        RECT 39.955 -104.885 40.285 -104.555 ;
        RECT 39.955 -106.245 40.285 -105.915 ;
        RECT 39.955 -107.605 40.285 -107.275 ;
        RECT 39.955 -108.965 40.285 -108.635 ;
        RECT 39.955 -110.325 40.285 -109.995 ;
        RECT 39.955 -111.685 40.285 -111.355 ;
        RECT 39.955 -113.045 40.285 -112.715 ;
        RECT 39.955 -114.405 40.285 -114.075 ;
        RECT 39.955 -115.765 40.285 -115.435 ;
        RECT 39.955 -117.125 40.285 -116.795 ;
        RECT 39.955 -118.485 40.285 -118.155 ;
        RECT 39.955 -119.845 40.285 -119.515 ;
        RECT 39.955 -121.205 40.285 -120.875 ;
        RECT 39.955 -122.565 40.285 -122.235 ;
        RECT 39.955 -123.925 40.285 -123.595 ;
        RECT 39.955 -125.285 40.285 -124.955 ;
        RECT 39.955 -126.645 40.285 -126.315 ;
        RECT 39.955 -128.005 40.285 -127.675 ;
        RECT 39.955 -129.365 40.285 -129.035 ;
        RECT 39.955 -130.725 40.285 -130.395 ;
        RECT 39.955 -132.085 40.285 -131.755 ;
        RECT 39.955 -133.445 40.285 -133.115 ;
        RECT 39.955 -134.805 40.285 -134.475 ;
        RECT 39.955 -136.165 40.285 -135.835 ;
        RECT 39.955 -137.525 40.285 -137.195 ;
        RECT 39.955 -138.885 40.285 -138.555 ;
        RECT 39.955 -140.245 40.285 -139.915 ;
        RECT 39.955 -141.605 40.285 -141.275 ;
        RECT 39.955 -142.965 40.285 -142.635 ;
        RECT 39.955 -144.325 40.285 -143.995 ;
        RECT 39.955 -145.685 40.285 -145.355 ;
        RECT 39.955 -147.045 40.285 -146.715 ;
        RECT 39.955 -148.405 40.285 -148.075 ;
        RECT 39.955 -149.765 40.285 -149.435 ;
        RECT 39.955 -151.125 40.285 -150.795 ;
        RECT 39.955 -152.485 40.285 -152.155 ;
        RECT 39.955 -153.845 40.285 -153.515 ;
        RECT 39.955 -155.205 40.285 -154.875 ;
        RECT 39.955 -156.565 40.285 -156.235 ;
        RECT 39.955 -157.925 40.285 -157.595 ;
        RECT 39.955 -159.285 40.285 -158.955 ;
        RECT 39.955 -160.645 40.285 -160.315 ;
        RECT 39.955 -162.005 40.285 -161.675 ;
        RECT 39.955 -163.365 40.285 -163.035 ;
        RECT 39.955 -164.725 40.285 -164.395 ;
        RECT 39.955 -166.085 40.285 -165.755 ;
        RECT 39.955 -167.445 40.285 -167.115 ;
        RECT 39.955 -168.805 40.285 -168.475 ;
        RECT 39.955 -170.165 40.285 -169.835 ;
        RECT 39.955 -171.525 40.285 -171.195 ;
        RECT 39.955 -172.885 40.285 -172.555 ;
        RECT 39.955 -174.245 40.285 -173.915 ;
        RECT 39.955 -175.605 40.285 -175.275 ;
        RECT 39.955 -176.965 40.285 -176.635 ;
        RECT 39.955 -178.325 40.285 -177.995 ;
        RECT 39.955 -179.685 40.285 -179.355 ;
        RECT 39.955 -181.93 40.285 -180.8 ;
        RECT 39.96 -182.045 40.28 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 241.32 41.645 242.45 ;
        RECT 41.315 239.195 41.645 239.525 ;
        RECT 41.315 237.835 41.645 238.165 ;
        RECT 41.32 237.16 41.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 -1.525 41.645 -1.195 ;
        RECT 41.315 -2.885 41.645 -2.555 ;
        RECT 41.32 -3.56 41.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 41.315 -95.365 41.645 -95.035 ;
        RECT 41.315 -96.725 41.645 -96.395 ;
        RECT 41.315 -98.085 41.645 -97.755 ;
        RECT 41.315 -99.445 41.645 -99.115 ;
        RECT 41.315 -100.805 41.645 -100.475 ;
        RECT 41.315 -102.165 41.645 -101.835 ;
        RECT 41.315 -103.525 41.645 -103.195 ;
        RECT 41.315 -104.885 41.645 -104.555 ;
        RECT 41.315 -106.245 41.645 -105.915 ;
        RECT 41.315 -107.605 41.645 -107.275 ;
        RECT 41.315 -108.965 41.645 -108.635 ;
        RECT 41.315 -110.325 41.645 -109.995 ;
        RECT 41.315 -111.685 41.645 -111.355 ;
        RECT 41.315 -113.045 41.645 -112.715 ;
        RECT 41.315 -114.405 41.645 -114.075 ;
        RECT 41.315 -115.765 41.645 -115.435 ;
        RECT 41.315 -117.125 41.645 -116.795 ;
        RECT 41.315 -118.485 41.645 -118.155 ;
        RECT 41.315 -119.845 41.645 -119.515 ;
        RECT 41.315 -121.205 41.645 -120.875 ;
        RECT 41.315 -122.565 41.645 -122.235 ;
        RECT 41.315 -123.925 41.645 -123.595 ;
        RECT 41.315 -125.285 41.645 -124.955 ;
        RECT 41.315 -126.645 41.645 -126.315 ;
        RECT 41.315 -128.005 41.645 -127.675 ;
        RECT 41.315 -129.365 41.645 -129.035 ;
        RECT 41.315 -130.725 41.645 -130.395 ;
        RECT 41.315 -132.085 41.645 -131.755 ;
        RECT 41.315 -133.445 41.645 -133.115 ;
        RECT 41.315 -134.805 41.645 -134.475 ;
        RECT 41.315 -136.165 41.645 -135.835 ;
        RECT 41.315 -137.525 41.645 -137.195 ;
        RECT 41.315 -138.885 41.645 -138.555 ;
        RECT 41.315 -140.245 41.645 -139.915 ;
        RECT 41.315 -141.605 41.645 -141.275 ;
        RECT 41.315 -142.965 41.645 -142.635 ;
        RECT 41.315 -144.325 41.645 -143.995 ;
        RECT 41.315 -145.685 41.645 -145.355 ;
        RECT 41.315 -147.045 41.645 -146.715 ;
        RECT 41.315 -148.405 41.645 -148.075 ;
        RECT 41.315 -149.765 41.645 -149.435 ;
        RECT 41.315 -151.125 41.645 -150.795 ;
        RECT 41.315 -152.485 41.645 -152.155 ;
        RECT 41.315 -153.845 41.645 -153.515 ;
        RECT 41.315 -155.205 41.645 -154.875 ;
        RECT 41.315 -156.565 41.645 -156.235 ;
        RECT 41.315 -157.925 41.645 -157.595 ;
        RECT 41.315 -159.285 41.645 -158.955 ;
        RECT 41.315 -160.645 41.645 -160.315 ;
        RECT 41.315 -162.005 41.645 -161.675 ;
        RECT 41.315 -163.365 41.645 -163.035 ;
        RECT 41.315 -164.725 41.645 -164.395 ;
        RECT 41.315 -166.085 41.645 -165.755 ;
        RECT 41.315 -167.445 41.645 -167.115 ;
        RECT 41.315 -168.805 41.645 -168.475 ;
        RECT 41.315 -170.165 41.645 -169.835 ;
        RECT 41.315 -171.525 41.645 -171.195 ;
        RECT 41.315 -172.885 41.645 -172.555 ;
        RECT 41.315 -174.245 41.645 -173.915 ;
        RECT 41.315 -175.605 41.645 -175.275 ;
        RECT 41.315 -176.965 41.645 -176.635 ;
        RECT 41.315 -178.325 41.645 -177.995 ;
        RECT 41.315 -179.685 41.645 -179.355 ;
        RECT 41.315 -181.93 41.645 -180.8 ;
        RECT 41.32 -182.045 41.64 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 241.32 43.005 242.45 ;
        RECT 42.675 239.195 43.005 239.525 ;
        RECT 42.675 237.835 43.005 238.165 ;
        RECT 42.68 237.16 43 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 -1.525 43.005 -1.195 ;
        RECT 42.675 -2.885 43.005 -2.555 ;
        RECT 42.68 -3.56 43 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 42.675 -129.365 43.005 -129.035 ;
        RECT 42.675 -130.725 43.005 -130.395 ;
        RECT 42.675 -132.085 43.005 -131.755 ;
        RECT 42.675 -133.445 43.005 -133.115 ;
        RECT 42.675 -134.805 43.005 -134.475 ;
        RECT 42.675 -136.165 43.005 -135.835 ;
        RECT 42.675 -137.525 43.005 -137.195 ;
        RECT 42.675 -138.885 43.005 -138.555 ;
        RECT 42.675 -140.245 43.005 -139.915 ;
        RECT 42.675 -141.605 43.005 -141.275 ;
        RECT 42.675 -142.965 43.005 -142.635 ;
        RECT 42.675 -144.325 43.005 -143.995 ;
        RECT 42.675 -145.685 43.005 -145.355 ;
        RECT 42.675 -147.045 43.005 -146.715 ;
        RECT 42.675 -148.405 43.005 -148.075 ;
        RECT 42.675 -149.765 43.005 -149.435 ;
        RECT 42.675 -151.125 43.005 -150.795 ;
        RECT 42.675 -152.485 43.005 -152.155 ;
        RECT 42.675 -153.845 43.005 -153.515 ;
        RECT 42.675 -155.205 43.005 -154.875 ;
        RECT 42.675 -156.565 43.005 -156.235 ;
        RECT 42.675 -157.925 43.005 -157.595 ;
        RECT 42.675 -159.285 43.005 -158.955 ;
        RECT 42.675 -160.645 43.005 -160.315 ;
        RECT 42.675 -162.005 43.005 -161.675 ;
        RECT 42.675 -163.365 43.005 -163.035 ;
        RECT 42.675 -164.725 43.005 -164.395 ;
        RECT 42.675 -166.085 43.005 -165.755 ;
        RECT 42.675 -167.445 43.005 -167.115 ;
        RECT 42.675 -168.805 43.005 -168.475 ;
        RECT 42.675 -170.165 43.005 -169.835 ;
        RECT 42.675 -171.525 43.005 -171.195 ;
        RECT 42.675 -172.885 43.005 -172.555 ;
        RECT 42.675 -174.245 43.005 -173.915 ;
        RECT 42.675 -175.605 43.005 -175.275 ;
        RECT 42.675 -176.965 43.005 -176.635 ;
        RECT 42.675 -178.325 43.005 -177.995 ;
        RECT 42.675 -179.685 43.005 -179.355 ;
        RECT 42.675 -181.93 43.005 -180.8 ;
        RECT 42.68 -182.045 43 -95.035 ;
        RECT 42.675 -95.365 43.005 -95.035 ;
        RECT 42.675 -96.725 43.005 -96.395 ;
        RECT 42.675 -98.085 43.005 -97.755 ;
        RECT 42.675 -99.445 43.005 -99.115 ;
        RECT 42.675 -100.805 43.005 -100.475 ;
        RECT 42.675 -102.165 43.005 -101.835 ;
        RECT 42.675 -103.525 43.005 -103.195 ;
        RECT 42.675 -104.885 43.005 -104.555 ;
        RECT 42.675 -106.245 43.005 -105.915 ;
        RECT 42.675 -107.605 43.005 -107.275 ;
        RECT 42.675 -108.965 43.005 -108.635 ;
        RECT 42.675 -110.325 43.005 -109.995 ;
        RECT 42.675 -111.685 43.005 -111.355 ;
        RECT 42.675 -113.045 43.005 -112.715 ;
        RECT 42.675 -114.405 43.005 -114.075 ;
        RECT 42.675 -115.765 43.005 -115.435 ;
        RECT 42.675 -117.125 43.005 -116.795 ;
        RECT 42.675 -118.485 43.005 -118.155 ;
        RECT 42.675 -119.845 43.005 -119.515 ;
        RECT 42.675 -121.205 43.005 -120.875 ;
        RECT 42.675 -122.565 43.005 -122.235 ;
        RECT 42.675 -123.925 43.005 -123.595 ;
        RECT 42.675 -125.285 43.005 -124.955 ;
        RECT 42.675 -126.645 43.005 -126.315 ;
        RECT 42.675 -128.005 43.005 -127.675 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.845 -51.845 -0.515 -51.515 ;
        RECT -0.845 -53.205 -0.515 -52.875 ;
        RECT -0.845 -54.565 -0.515 -54.235 ;
        RECT -0.845 -55.925 -0.515 -55.595 ;
        RECT -0.845 -57.285 -0.515 -56.955 ;
        RECT -0.845 -58.645 -0.515 -58.315 ;
        RECT -0.845 -60.005 -0.515 -59.675 ;
        RECT -0.845 -61.365 -0.515 -61.035 ;
        RECT -0.845 -62.725 -0.515 -62.395 ;
        RECT -0.845 -64.085 -0.515 -63.755 ;
        RECT -0.845 -65.445 -0.515 -65.115 ;
        RECT -0.845 -68.165 -0.515 -67.835 ;
        RECT -0.845 -69.525 -0.515 -69.195 ;
        RECT -0.845 -70.885 -0.515 -70.555 ;
        RECT -0.845 -72.245 -0.515 -71.915 ;
        RECT -0.845 -73.605 -0.515 -73.275 ;
        RECT -0.845 -74.965 -0.515 -74.635 ;
        RECT -0.845 -76.325 -0.515 -75.995 ;
        RECT -0.845 -77.685 -0.515 -77.355 ;
        RECT -0.845 -79.045 -0.515 -78.715 ;
        RECT -0.845 -80.405 -0.515 -80.075 ;
        RECT -0.845 -81.765 -0.515 -81.435 ;
        RECT -0.845 -83.125 -0.515 -82.795 ;
        RECT -0.845 -84.485 -0.515 -84.155 ;
        RECT -0.845 -85.845 -0.515 -85.515 ;
        RECT -0.845 -87.205 -0.515 -86.875 ;
        RECT -0.845 -88.565 -0.515 -88.235 ;
        RECT -0.845 -91.285 -0.515 -90.955 ;
        RECT -0.845 -92.645 -0.515 -92.315 ;
        RECT -0.845 -94.005 -0.515 -93.675 ;
        RECT -0.845 -95.365 -0.515 -95.035 ;
        RECT -0.845 -96.725 -0.515 -96.395 ;
        RECT -0.845 -98.085 -0.515 -97.755 ;
        RECT -0.845 -99.445 -0.515 -99.115 ;
        RECT -0.845 -100.805 -0.515 -100.475 ;
        RECT -0.845 -102.165 -0.515 -101.835 ;
        RECT -0.845 -103.525 -0.515 -103.195 ;
        RECT -0.845 -104.885 -0.515 -104.555 ;
        RECT -0.845 -106.245 -0.515 -105.915 ;
        RECT -0.845 -107.605 -0.515 -107.275 ;
        RECT -0.845 -108.965 -0.515 -108.635 ;
        RECT -0.845 -110.325 -0.515 -109.995 ;
        RECT -0.845 -111.685 -0.515 -111.355 ;
        RECT -0.845 -113.045 -0.515 -112.715 ;
        RECT -0.845 -114.405 -0.515 -114.075 ;
        RECT -0.845 -115.765 -0.515 -115.435 ;
        RECT -0.845 -117.125 -0.515 -116.795 ;
        RECT -0.845 -118.485 -0.515 -118.155 ;
        RECT -0.845 -119.845 -0.515 -119.515 ;
        RECT -0.845 -121.205 -0.515 -120.875 ;
        RECT -0.845 -122.565 -0.515 -122.235 ;
        RECT -0.845 -123.925 -0.515 -123.595 ;
        RECT -0.845 -125.285 -0.515 -124.955 ;
        RECT -0.845 -126.645 -0.515 -126.315 ;
        RECT -0.845 -128.005 -0.515 -127.675 ;
        RECT -0.845 -129.365 -0.515 -129.035 ;
        RECT -0.845 -130.725 -0.515 -130.395 ;
        RECT -0.845 -132.085 -0.515 -131.755 ;
        RECT -0.845 -133.445 -0.515 -133.115 ;
        RECT -0.845 -134.805 -0.515 -134.475 ;
        RECT -0.845 -136.165 -0.515 -135.835 ;
        RECT -0.845 -137.525 -0.515 -137.195 ;
        RECT -0.845 -138.885 -0.515 -138.555 ;
        RECT -0.845 -140.245 -0.515 -139.915 ;
        RECT -0.845 -141.605 -0.515 -141.275 ;
        RECT -0.845 -142.965 -0.515 -142.635 ;
        RECT -0.845 -144.325 -0.515 -143.995 ;
        RECT -0.845 -145.685 -0.515 -145.355 ;
        RECT -0.845 -147.045 -0.515 -146.715 ;
        RECT -0.845 -148.405 -0.515 -148.075 ;
        RECT -0.845 -149.765 -0.515 -149.435 ;
        RECT -0.845 -151.125 -0.515 -150.795 ;
        RECT -0.845 -152.485 -0.515 -152.155 ;
        RECT -0.845 -153.845 -0.515 -153.515 ;
        RECT -0.845 -155.205 -0.515 -154.875 ;
        RECT -0.845 -156.565 -0.515 -156.235 ;
        RECT -0.845 -157.925 -0.515 -157.595 ;
        RECT -0.845 -159.285 -0.515 -158.955 ;
        RECT -0.845 -160.645 -0.515 -160.315 ;
        RECT -0.845 -162.005 -0.515 -161.675 ;
        RECT -0.845 -163.365 -0.515 -163.035 ;
        RECT -0.845 -164.725 -0.515 -164.395 ;
        RECT -0.845 -166.085 -0.515 -165.755 ;
        RECT -0.845 -167.445 -0.515 -167.115 ;
        RECT -0.845 -168.805 -0.515 -168.475 ;
        RECT -0.845 -170.165 -0.515 -169.835 ;
        RECT -0.845 -171.525 -0.515 -171.195 ;
        RECT -0.845 -172.885 -0.515 -172.555 ;
        RECT -0.845 -174.245 -0.515 -173.915 ;
        RECT -0.845 -175.605 -0.515 -175.275 ;
        RECT -0.845 -176.965 -0.515 -176.635 ;
        RECT -0.845 -178.325 -0.515 -177.995 ;
        RECT -0.845 -179.685 -0.515 -179.355 ;
        RECT -0.845 -181.93 -0.515 -180.8 ;
        RECT -0.84 -182.045 -0.52 -50.84 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 241.32 0.845 242.45 ;
        RECT 0.515 239.195 0.845 239.525 ;
        RECT 0.515 237.835 0.845 238.165 ;
        RECT 0.52 237.16 0.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 -1.525 0.845 -1.195 ;
        RECT 0.515 -2.885 0.845 -2.555 ;
        RECT 0.52 -3.56 0.84 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 0.515 -95.365 0.845 -95.035 ;
        RECT 0.515 -96.725 0.845 -96.395 ;
        RECT 0.515 -98.085 0.845 -97.755 ;
        RECT 0.515 -99.445 0.845 -99.115 ;
        RECT 0.515 -100.805 0.845 -100.475 ;
        RECT 0.515 -102.165 0.845 -101.835 ;
        RECT 0.515 -103.525 0.845 -103.195 ;
        RECT 0.515 -104.885 0.845 -104.555 ;
        RECT 0.515 -106.245 0.845 -105.915 ;
        RECT 0.515 -107.605 0.845 -107.275 ;
        RECT 0.515 -108.965 0.845 -108.635 ;
        RECT 0.515 -110.325 0.845 -109.995 ;
        RECT 0.515 -111.685 0.845 -111.355 ;
        RECT 0.515 -113.045 0.845 -112.715 ;
        RECT 0.515 -114.405 0.845 -114.075 ;
        RECT 0.515 -115.765 0.845 -115.435 ;
        RECT 0.515 -117.125 0.845 -116.795 ;
        RECT 0.515 -118.485 0.845 -118.155 ;
        RECT 0.515 -119.845 0.845 -119.515 ;
        RECT 0.515 -121.205 0.845 -120.875 ;
        RECT 0.515 -122.565 0.845 -122.235 ;
        RECT 0.515 -123.925 0.845 -123.595 ;
        RECT 0.515 -125.285 0.845 -124.955 ;
        RECT 0.515 -126.645 0.845 -126.315 ;
        RECT 0.515 -128.005 0.845 -127.675 ;
        RECT 0.515 -129.365 0.845 -129.035 ;
        RECT 0.515 -130.725 0.845 -130.395 ;
        RECT 0.515 -132.085 0.845 -131.755 ;
        RECT 0.515 -133.445 0.845 -133.115 ;
        RECT 0.515 -134.805 0.845 -134.475 ;
        RECT 0.515 -136.165 0.845 -135.835 ;
        RECT 0.515 -137.525 0.845 -137.195 ;
        RECT 0.515 -138.885 0.845 -138.555 ;
        RECT 0.515 -140.245 0.845 -139.915 ;
        RECT 0.515 -141.605 0.845 -141.275 ;
        RECT 0.515 -142.965 0.845 -142.635 ;
        RECT 0.515 -144.325 0.845 -143.995 ;
        RECT 0.515 -145.685 0.845 -145.355 ;
        RECT 0.515 -147.045 0.845 -146.715 ;
        RECT 0.515 -148.405 0.845 -148.075 ;
        RECT 0.515 -149.765 0.845 -149.435 ;
        RECT 0.515 -151.125 0.845 -150.795 ;
        RECT 0.515 -152.485 0.845 -152.155 ;
        RECT 0.515 -153.845 0.845 -153.515 ;
        RECT 0.515 -155.205 0.845 -154.875 ;
        RECT 0.515 -156.565 0.845 -156.235 ;
        RECT 0.515 -157.925 0.845 -157.595 ;
        RECT 0.515 -159.285 0.845 -158.955 ;
        RECT 0.515 -160.645 0.845 -160.315 ;
        RECT 0.515 -162.005 0.845 -161.675 ;
        RECT 0.515 -163.365 0.845 -163.035 ;
        RECT 0.515 -164.725 0.845 -164.395 ;
        RECT 0.515 -166.085 0.845 -165.755 ;
        RECT 0.515 -167.445 0.845 -167.115 ;
        RECT 0.515 -168.805 0.845 -168.475 ;
        RECT 0.515 -170.165 0.845 -169.835 ;
        RECT 0.515 -171.525 0.845 -171.195 ;
        RECT 0.515 -172.885 0.845 -172.555 ;
        RECT 0.515 -174.245 0.845 -173.915 ;
        RECT 0.515 -175.605 0.845 -175.275 ;
        RECT 0.515 -176.965 0.845 -176.635 ;
        RECT 0.515 -178.325 0.845 -177.995 ;
        RECT 0.515 -179.685 0.845 -179.355 ;
        RECT 0.515 -181.93 0.845 -180.8 ;
        RECT 0.52 -182.045 0.84 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 241.32 2.205 242.45 ;
        RECT 1.875 239.195 2.205 239.525 ;
        RECT 1.875 237.835 2.205 238.165 ;
        RECT 1.88 237.16 2.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 -1.525 2.205 -1.195 ;
        RECT 1.875 -2.885 2.205 -2.555 ;
        RECT 1.88 -3.56 2.2 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.875 -95.365 2.205 -95.035 ;
        RECT 1.875 -96.725 2.205 -96.395 ;
        RECT 1.875 -98.085 2.205 -97.755 ;
        RECT 1.875 -99.445 2.205 -99.115 ;
        RECT 1.875 -100.805 2.205 -100.475 ;
        RECT 1.875 -102.165 2.205 -101.835 ;
        RECT 1.875 -103.525 2.205 -103.195 ;
        RECT 1.875 -104.885 2.205 -104.555 ;
        RECT 1.875 -106.245 2.205 -105.915 ;
        RECT 1.875 -107.605 2.205 -107.275 ;
        RECT 1.875 -108.965 2.205 -108.635 ;
        RECT 1.875 -110.325 2.205 -109.995 ;
        RECT 1.875 -111.685 2.205 -111.355 ;
        RECT 1.875 -113.045 2.205 -112.715 ;
        RECT 1.875 -114.405 2.205 -114.075 ;
        RECT 1.875 -115.765 2.205 -115.435 ;
        RECT 1.875 -117.125 2.205 -116.795 ;
        RECT 1.875 -118.485 2.205 -118.155 ;
        RECT 1.875 -119.845 2.205 -119.515 ;
        RECT 1.875 -121.205 2.205 -120.875 ;
        RECT 1.875 -122.565 2.205 -122.235 ;
        RECT 1.875 -123.925 2.205 -123.595 ;
        RECT 1.875 -125.285 2.205 -124.955 ;
        RECT 1.875 -126.645 2.205 -126.315 ;
        RECT 1.875 -128.005 2.205 -127.675 ;
        RECT 1.875 -129.365 2.205 -129.035 ;
        RECT 1.875 -130.725 2.205 -130.395 ;
        RECT 1.875 -132.085 2.205 -131.755 ;
        RECT 1.875 -133.445 2.205 -133.115 ;
        RECT 1.875 -134.805 2.205 -134.475 ;
        RECT 1.875 -136.165 2.205 -135.835 ;
        RECT 1.875 -137.525 2.205 -137.195 ;
        RECT 1.875 -138.885 2.205 -138.555 ;
        RECT 1.875 -140.245 2.205 -139.915 ;
        RECT 1.875 -141.605 2.205 -141.275 ;
        RECT 1.875 -142.965 2.205 -142.635 ;
        RECT 1.875 -144.325 2.205 -143.995 ;
        RECT 1.875 -145.685 2.205 -145.355 ;
        RECT 1.875 -147.045 2.205 -146.715 ;
        RECT 1.875 -148.405 2.205 -148.075 ;
        RECT 1.875 -149.765 2.205 -149.435 ;
        RECT 1.875 -151.125 2.205 -150.795 ;
        RECT 1.875 -152.485 2.205 -152.155 ;
        RECT 1.875 -153.845 2.205 -153.515 ;
        RECT 1.875 -155.205 2.205 -154.875 ;
        RECT 1.875 -156.565 2.205 -156.235 ;
        RECT 1.875 -157.925 2.205 -157.595 ;
        RECT 1.875 -159.285 2.205 -158.955 ;
        RECT 1.875 -160.645 2.205 -160.315 ;
        RECT 1.875 -162.005 2.205 -161.675 ;
        RECT 1.875 -163.365 2.205 -163.035 ;
        RECT 1.875 -164.725 2.205 -164.395 ;
        RECT 1.875 -166.085 2.205 -165.755 ;
        RECT 1.875 -167.445 2.205 -167.115 ;
        RECT 1.875 -168.805 2.205 -168.475 ;
        RECT 1.875 -170.165 2.205 -169.835 ;
        RECT 1.875 -171.525 2.205 -171.195 ;
        RECT 1.875 -172.885 2.205 -172.555 ;
        RECT 1.875 -174.245 2.205 -173.915 ;
        RECT 1.875 -175.605 2.205 -175.275 ;
        RECT 1.875 -176.965 2.205 -176.635 ;
        RECT 1.875 -178.325 2.205 -177.995 ;
        RECT 1.875 -179.685 2.205 -179.355 ;
        RECT 1.875 -181.93 2.205 -180.8 ;
        RECT 1.88 -182.045 2.2 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 241.32 3.565 242.45 ;
        RECT 3.235 239.195 3.565 239.525 ;
        RECT 3.235 237.835 3.565 238.165 ;
        RECT 3.24 237.16 3.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.235 -99.445 3.565 -99.115 ;
        RECT 3.235 -100.805 3.565 -100.475 ;
        RECT 3.235 -102.165 3.565 -101.835 ;
        RECT 3.235 -103.525 3.565 -103.195 ;
        RECT 3.235 -104.885 3.565 -104.555 ;
        RECT 3.235 -106.245 3.565 -105.915 ;
        RECT 3.235 -107.605 3.565 -107.275 ;
        RECT 3.235 -108.965 3.565 -108.635 ;
        RECT 3.235 -110.325 3.565 -109.995 ;
        RECT 3.235 -111.685 3.565 -111.355 ;
        RECT 3.235 -113.045 3.565 -112.715 ;
        RECT 3.235 -114.405 3.565 -114.075 ;
        RECT 3.235 -115.765 3.565 -115.435 ;
        RECT 3.235 -117.125 3.565 -116.795 ;
        RECT 3.235 -118.485 3.565 -118.155 ;
        RECT 3.235 -119.845 3.565 -119.515 ;
        RECT 3.235 -121.205 3.565 -120.875 ;
        RECT 3.235 -122.565 3.565 -122.235 ;
        RECT 3.235 -123.925 3.565 -123.595 ;
        RECT 3.235 -125.285 3.565 -124.955 ;
        RECT 3.235 -126.645 3.565 -126.315 ;
        RECT 3.235 -128.005 3.565 -127.675 ;
        RECT 3.235 -129.365 3.565 -129.035 ;
        RECT 3.235 -130.725 3.565 -130.395 ;
        RECT 3.235 -132.085 3.565 -131.755 ;
        RECT 3.235 -133.445 3.565 -133.115 ;
        RECT 3.235 -134.805 3.565 -134.475 ;
        RECT 3.235 -136.165 3.565 -135.835 ;
        RECT 3.235 -137.525 3.565 -137.195 ;
        RECT 3.235 -138.885 3.565 -138.555 ;
        RECT 3.235 -140.245 3.565 -139.915 ;
        RECT 3.235 -141.605 3.565 -141.275 ;
        RECT 3.235 -142.965 3.565 -142.635 ;
        RECT 3.235 -144.325 3.565 -143.995 ;
        RECT 3.235 -145.685 3.565 -145.355 ;
        RECT 3.235 -147.045 3.565 -146.715 ;
        RECT 3.235 -148.405 3.565 -148.075 ;
        RECT 3.235 -149.765 3.565 -149.435 ;
        RECT 3.235 -151.125 3.565 -150.795 ;
        RECT 3.235 -152.485 3.565 -152.155 ;
        RECT 3.235 -153.845 3.565 -153.515 ;
        RECT 3.235 -155.205 3.565 -154.875 ;
        RECT 3.235 -156.565 3.565 -156.235 ;
        RECT 3.235 -157.925 3.565 -157.595 ;
        RECT 3.235 -159.285 3.565 -158.955 ;
        RECT 3.235 -160.645 3.565 -160.315 ;
        RECT 3.235 -162.005 3.565 -161.675 ;
        RECT 3.235 -163.365 3.565 -163.035 ;
        RECT 3.235 -164.725 3.565 -164.395 ;
        RECT 3.235 -166.085 3.565 -165.755 ;
        RECT 3.235 -167.445 3.565 -167.115 ;
        RECT 3.235 -168.805 3.565 -168.475 ;
        RECT 3.235 -170.165 3.565 -169.835 ;
        RECT 3.235 -171.525 3.565 -171.195 ;
        RECT 3.235 -172.885 3.565 -172.555 ;
        RECT 3.235 -174.245 3.565 -173.915 ;
        RECT 3.235 -175.605 3.565 -175.275 ;
        RECT 3.235 -176.965 3.565 -176.635 ;
        RECT 3.235 -178.325 3.565 -177.995 ;
        RECT 3.235 -179.685 3.565 -179.355 ;
        RECT 3.235 -181.93 3.565 -180.8 ;
        RECT 3.24 -182.045 3.56 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 3.31 -98.075 3.64 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 241.32 4.925 242.45 ;
        RECT 4.595 239.195 4.925 239.525 ;
        RECT 4.595 237.835 4.925 238.165 ;
        RECT 4.6 237.16 4.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 4.595 -1.525 4.925 -1.195 ;
        RECT 4.595 -2.885 4.925 -2.555 ;
        RECT 4.6 -3.56 4.92 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 241.32 6.285 242.45 ;
        RECT 5.955 239.195 6.285 239.525 ;
        RECT 5.955 237.835 6.285 238.165 ;
        RECT 5.96 237.16 6.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.955 -1.525 6.285 -1.195 ;
        RECT 5.955 -2.885 6.285 -2.555 ;
        RECT 5.96 -3.56 6.28 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 241.32 7.645 242.45 ;
        RECT 7.315 239.195 7.645 239.525 ;
        RECT 7.315 237.835 7.645 238.165 ;
        RECT 7.32 237.16 7.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 -1.525 7.645 -1.195 ;
        RECT 7.315 -2.885 7.645 -2.555 ;
        RECT 7.32 -3.56 7.64 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 7.315 -95.365 7.645 -95.035 ;
        RECT 7.315 -96.725 7.645 -96.395 ;
        RECT 7.315 -98.085 7.645 -97.755 ;
        RECT 7.315 -99.445 7.645 -99.115 ;
        RECT 7.315 -100.805 7.645 -100.475 ;
        RECT 7.315 -102.165 7.645 -101.835 ;
        RECT 7.315 -103.525 7.645 -103.195 ;
        RECT 7.315 -104.885 7.645 -104.555 ;
        RECT 7.315 -106.245 7.645 -105.915 ;
        RECT 7.315 -107.605 7.645 -107.275 ;
        RECT 7.315 -108.965 7.645 -108.635 ;
        RECT 7.315 -110.325 7.645 -109.995 ;
        RECT 7.315 -111.685 7.645 -111.355 ;
        RECT 7.315 -113.045 7.645 -112.715 ;
        RECT 7.315 -114.405 7.645 -114.075 ;
        RECT 7.315 -115.765 7.645 -115.435 ;
        RECT 7.315 -117.125 7.645 -116.795 ;
        RECT 7.315 -118.485 7.645 -118.155 ;
        RECT 7.315 -119.845 7.645 -119.515 ;
        RECT 7.315 -121.205 7.645 -120.875 ;
        RECT 7.315 -122.565 7.645 -122.235 ;
        RECT 7.315 -123.925 7.645 -123.595 ;
        RECT 7.315 -125.285 7.645 -124.955 ;
        RECT 7.315 -126.645 7.645 -126.315 ;
        RECT 7.315 -128.005 7.645 -127.675 ;
        RECT 7.315 -129.365 7.645 -129.035 ;
        RECT 7.315 -130.725 7.645 -130.395 ;
        RECT 7.315 -132.085 7.645 -131.755 ;
        RECT 7.315 -133.445 7.645 -133.115 ;
        RECT 7.315 -134.805 7.645 -134.475 ;
        RECT 7.315 -136.165 7.645 -135.835 ;
        RECT 7.315 -137.525 7.645 -137.195 ;
        RECT 7.315 -138.885 7.645 -138.555 ;
        RECT 7.315 -140.245 7.645 -139.915 ;
        RECT 7.315 -141.605 7.645 -141.275 ;
        RECT 7.315 -142.965 7.645 -142.635 ;
        RECT 7.315 -144.325 7.645 -143.995 ;
        RECT 7.315 -145.685 7.645 -145.355 ;
        RECT 7.315 -147.045 7.645 -146.715 ;
        RECT 7.315 -148.405 7.645 -148.075 ;
        RECT 7.315 -149.765 7.645 -149.435 ;
        RECT 7.315 -151.125 7.645 -150.795 ;
        RECT 7.315 -152.485 7.645 -152.155 ;
        RECT 7.315 -153.845 7.645 -153.515 ;
        RECT 7.315 -155.205 7.645 -154.875 ;
        RECT 7.315 -156.565 7.645 -156.235 ;
        RECT 7.315 -157.925 7.645 -157.595 ;
        RECT 7.315 -159.285 7.645 -158.955 ;
        RECT 7.315 -160.645 7.645 -160.315 ;
        RECT 7.315 -162.005 7.645 -161.675 ;
        RECT 7.315 -163.365 7.645 -163.035 ;
        RECT 7.315 -164.725 7.645 -164.395 ;
        RECT 7.315 -166.085 7.645 -165.755 ;
        RECT 7.315 -167.445 7.645 -167.115 ;
        RECT 7.315 -168.805 7.645 -168.475 ;
        RECT 7.315 -170.165 7.645 -169.835 ;
        RECT 7.315 -171.525 7.645 -171.195 ;
        RECT 7.315 -172.885 7.645 -172.555 ;
        RECT 7.315 -174.245 7.645 -173.915 ;
        RECT 7.315 -175.605 7.645 -175.275 ;
        RECT 7.315 -176.965 7.645 -176.635 ;
        RECT 7.315 -178.325 7.645 -177.995 ;
        RECT 7.315 -179.685 7.645 -179.355 ;
        RECT 7.315 -181.93 7.645 -180.8 ;
        RECT 7.32 -182.045 7.64 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 241.32 9.005 242.45 ;
        RECT 8.675 239.195 9.005 239.525 ;
        RECT 8.675 237.835 9.005 238.165 ;
        RECT 8.68 237.16 9 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 -1.525 9.005 -1.195 ;
        RECT 8.675 -2.885 9.005 -2.555 ;
        RECT 8.68 -3.56 9 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 8.675 -95.365 9.005 -95.035 ;
        RECT 8.675 -96.725 9.005 -96.395 ;
        RECT 8.675 -98.085 9.005 -97.755 ;
        RECT 8.675 -99.445 9.005 -99.115 ;
        RECT 8.675 -100.805 9.005 -100.475 ;
        RECT 8.675 -102.165 9.005 -101.835 ;
        RECT 8.675 -103.525 9.005 -103.195 ;
        RECT 8.675 -104.885 9.005 -104.555 ;
        RECT 8.675 -106.245 9.005 -105.915 ;
        RECT 8.675 -107.605 9.005 -107.275 ;
        RECT 8.675 -108.965 9.005 -108.635 ;
        RECT 8.675 -110.325 9.005 -109.995 ;
        RECT 8.675 -111.685 9.005 -111.355 ;
        RECT 8.675 -113.045 9.005 -112.715 ;
        RECT 8.675 -114.405 9.005 -114.075 ;
        RECT 8.675 -115.765 9.005 -115.435 ;
        RECT 8.675 -117.125 9.005 -116.795 ;
        RECT 8.675 -118.485 9.005 -118.155 ;
        RECT 8.675 -119.845 9.005 -119.515 ;
        RECT 8.675 -121.205 9.005 -120.875 ;
        RECT 8.675 -122.565 9.005 -122.235 ;
        RECT 8.675 -123.925 9.005 -123.595 ;
        RECT 8.675 -125.285 9.005 -124.955 ;
        RECT 8.675 -126.645 9.005 -126.315 ;
        RECT 8.675 -128.005 9.005 -127.675 ;
        RECT 8.675 -129.365 9.005 -129.035 ;
        RECT 8.675 -130.725 9.005 -130.395 ;
        RECT 8.675 -132.085 9.005 -131.755 ;
        RECT 8.675 -133.445 9.005 -133.115 ;
        RECT 8.675 -134.805 9.005 -134.475 ;
        RECT 8.675 -136.165 9.005 -135.835 ;
        RECT 8.675 -137.525 9.005 -137.195 ;
        RECT 8.675 -138.885 9.005 -138.555 ;
        RECT 8.675 -140.245 9.005 -139.915 ;
        RECT 8.675 -141.605 9.005 -141.275 ;
        RECT 8.675 -142.965 9.005 -142.635 ;
        RECT 8.675 -144.325 9.005 -143.995 ;
        RECT 8.675 -145.685 9.005 -145.355 ;
        RECT 8.675 -147.045 9.005 -146.715 ;
        RECT 8.675 -148.405 9.005 -148.075 ;
        RECT 8.675 -149.765 9.005 -149.435 ;
        RECT 8.675 -151.125 9.005 -150.795 ;
        RECT 8.675 -152.485 9.005 -152.155 ;
        RECT 8.675 -153.845 9.005 -153.515 ;
        RECT 8.675 -155.205 9.005 -154.875 ;
        RECT 8.675 -156.565 9.005 -156.235 ;
        RECT 8.675 -157.925 9.005 -157.595 ;
        RECT 8.675 -159.285 9.005 -158.955 ;
        RECT 8.675 -160.645 9.005 -160.315 ;
        RECT 8.675 -162.005 9.005 -161.675 ;
        RECT 8.675 -163.365 9.005 -163.035 ;
        RECT 8.675 -164.725 9.005 -164.395 ;
        RECT 8.675 -166.085 9.005 -165.755 ;
        RECT 8.675 -167.445 9.005 -167.115 ;
        RECT 8.675 -168.805 9.005 -168.475 ;
        RECT 8.675 -170.165 9.005 -169.835 ;
        RECT 8.675 -171.525 9.005 -171.195 ;
        RECT 8.675 -172.885 9.005 -172.555 ;
        RECT 8.675 -174.245 9.005 -173.915 ;
        RECT 8.675 -175.605 9.005 -175.275 ;
        RECT 8.675 -176.965 9.005 -176.635 ;
        RECT 8.675 -178.325 9.005 -177.995 ;
        RECT 8.675 -179.685 9.005 -179.355 ;
        RECT 8.675 -181.93 9.005 -180.8 ;
        RECT 8.68 -182.045 9 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 241.32 10.365 242.45 ;
        RECT 10.035 239.195 10.365 239.525 ;
        RECT 10.035 237.835 10.365 238.165 ;
        RECT 10.04 237.16 10.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 -1.525 10.365 -1.195 ;
        RECT 10.035 -2.885 10.365 -2.555 ;
        RECT 10.04 -3.56 10.36 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 10.035 -95.365 10.365 -95.035 ;
        RECT 10.035 -96.725 10.365 -96.395 ;
        RECT 10.035 -98.085 10.365 -97.755 ;
        RECT 10.035 -99.445 10.365 -99.115 ;
        RECT 10.035 -100.805 10.365 -100.475 ;
        RECT 10.035 -102.165 10.365 -101.835 ;
        RECT 10.035 -103.525 10.365 -103.195 ;
        RECT 10.035 -104.885 10.365 -104.555 ;
        RECT 10.035 -106.245 10.365 -105.915 ;
        RECT 10.035 -107.605 10.365 -107.275 ;
        RECT 10.035 -108.965 10.365 -108.635 ;
        RECT 10.035 -110.325 10.365 -109.995 ;
        RECT 10.035 -111.685 10.365 -111.355 ;
        RECT 10.035 -113.045 10.365 -112.715 ;
        RECT 10.035 -114.405 10.365 -114.075 ;
        RECT 10.035 -115.765 10.365 -115.435 ;
        RECT 10.035 -117.125 10.365 -116.795 ;
        RECT 10.035 -118.485 10.365 -118.155 ;
        RECT 10.035 -119.845 10.365 -119.515 ;
        RECT 10.035 -121.205 10.365 -120.875 ;
        RECT 10.035 -122.565 10.365 -122.235 ;
        RECT 10.035 -123.925 10.365 -123.595 ;
        RECT 10.035 -125.285 10.365 -124.955 ;
        RECT 10.035 -126.645 10.365 -126.315 ;
        RECT 10.035 -128.005 10.365 -127.675 ;
        RECT 10.035 -129.365 10.365 -129.035 ;
        RECT 10.035 -130.725 10.365 -130.395 ;
        RECT 10.035 -132.085 10.365 -131.755 ;
        RECT 10.035 -133.445 10.365 -133.115 ;
        RECT 10.035 -134.805 10.365 -134.475 ;
        RECT 10.035 -136.165 10.365 -135.835 ;
        RECT 10.035 -137.525 10.365 -137.195 ;
        RECT 10.035 -138.885 10.365 -138.555 ;
        RECT 10.035 -140.245 10.365 -139.915 ;
        RECT 10.035 -141.605 10.365 -141.275 ;
        RECT 10.035 -142.965 10.365 -142.635 ;
        RECT 10.035 -144.325 10.365 -143.995 ;
        RECT 10.035 -145.685 10.365 -145.355 ;
        RECT 10.035 -147.045 10.365 -146.715 ;
        RECT 10.035 -148.405 10.365 -148.075 ;
        RECT 10.035 -149.765 10.365 -149.435 ;
        RECT 10.035 -151.125 10.365 -150.795 ;
        RECT 10.035 -152.485 10.365 -152.155 ;
        RECT 10.035 -153.845 10.365 -153.515 ;
        RECT 10.035 -155.205 10.365 -154.875 ;
        RECT 10.035 -156.565 10.365 -156.235 ;
        RECT 10.035 -157.925 10.365 -157.595 ;
        RECT 10.035 -159.285 10.365 -158.955 ;
        RECT 10.035 -160.645 10.365 -160.315 ;
        RECT 10.035 -162.005 10.365 -161.675 ;
        RECT 10.035 -163.365 10.365 -163.035 ;
        RECT 10.035 -164.725 10.365 -164.395 ;
        RECT 10.035 -166.085 10.365 -165.755 ;
        RECT 10.035 -167.445 10.365 -167.115 ;
        RECT 10.035 -168.805 10.365 -168.475 ;
        RECT 10.035 -170.165 10.365 -169.835 ;
        RECT 10.035 -171.525 10.365 -171.195 ;
        RECT 10.035 -172.885 10.365 -172.555 ;
        RECT 10.035 -174.245 10.365 -173.915 ;
        RECT 10.035 -175.605 10.365 -175.275 ;
        RECT 10.035 -176.965 10.365 -176.635 ;
        RECT 10.035 -178.325 10.365 -177.995 ;
        RECT 10.035 -179.685 10.365 -179.355 ;
        RECT 10.035 -181.93 10.365 -180.8 ;
        RECT 10.04 -182.045 10.36 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 241.32 11.725 242.45 ;
        RECT 11.395 239.195 11.725 239.525 ;
        RECT 11.395 237.835 11.725 238.165 ;
        RECT 11.4 237.16 11.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 -1.525 11.725 -1.195 ;
        RECT 11.395 -2.885 11.725 -2.555 ;
        RECT 11.4 -3.56 11.72 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 11.395 -95.365 11.725 -95.035 ;
        RECT 11.395 -96.725 11.725 -96.395 ;
        RECT 11.395 -98.085 11.725 -97.755 ;
        RECT 11.395 -99.445 11.725 -99.115 ;
        RECT 11.395 -100.805 11.725 -100.475 ;
        RECT 11.395 -102.165 11.725 -101.835 ;
        RECT 11.395 -103.525 11.725 -103.195 ;
        RECT 11.395 -104.885 11.725 -104.555 ;
        RECT 11.395 -106.245 11.725 -105.915 ;
        RECT 11.395 -107.605 11.725 -107.275 ;
        RECT 11.395 -108.965 11.725 -108.635 ;
        RECT 11.395 -110.325 11.725 -109.995 ;
        RECT 11.395 -111.685 11.725 -111.355 ;
        RECT 11.395 -113.045 11.725 -112.715 ;
        RECT 11.395 -114.405 11.725 -114.075 ;
        RECT 11.395 -115.765 11.725 -115.435 ;
        RECT 11.395 -117.125 11.725 -116.795 ;
        RECT 11.395 -118.485 11.725 -118.155 ;
        RECT 11.395 -119.845 11.725 -119.515 ;
        RECT 11.395 -121.205 11.725 -120.875 ;
        RECT 11.395 -122.565 11.725 -122.235 ;
        RECT 11.395 -123.925 11.725 -123.595 ;
        RECT 11.395 -125.285 11.725 -124.955 ;
        RECT 11.395 -126.645 11.725 -126.315 ;
        RECT 11.395 -128.005 11.725 -127.675 ;
        RECT 11.395 -129.365 11.725 -129.035 ;
        RECT 11.395 -130.725 11.725 -130.395 ;
        RECT 11.395 -132.085 11.725 -131.755 ;
        RECT 11.395 -133.445 11.725 -133.115 ;
        RECT 11.395 -134.805 11.725 -134.475 ;
        RECT 11.395 -136.165 11.725 -135.835 ;
        RECT 11.395 -137.525 11.725 -137.195 ;
        RECT 11.395 -138.885 11.725 -138.555 ;
        RECT 11.395 -140.245 11.725 -139.915 ;
        RECT 11.395 -141.605 11.725 -141.275 ;
        RECT 11.395 -142.965 11.725 -142.635 ;
        RECT 11.395 -144.325 11.725 -143.995 ;
        RECT 11.395 -145.685 11.725 -145.355 ;
        RECT 11.395 -147.045 11.725 -146.715 ;
        RECT 11.395 -148.405 11.725 -148.075 ;
        RECT 11.395 -149.765 11.725 -149.435 ;
        RECT 11.395 -151.125 11.725 -150.795 ;
        RECT 11.395 -152.485 11.725 -152.155 ;
        RECT 11.395 -153.845 11.725 -153.515 ;
        RECT 11.395 -155.205 11.725 -154.875 ;
        RECT 11.395 -156.565 11.725 -156.235 ;
        RECT 11.395 -157.925 11.725 -157.595 ;
        RECT 11.395 -159.285 11.725 -158.955 ;
        RECT 11.395 -160.645 11.725 -160.315 ;
        RECT 11.395 -162.005 11.725 -161.675 ;
        RECT 11.395 -163.365 11.725 -163.035 ;
        RECT 11.395 -164.725 11.725 -164.395 ;
        RECT 11.395 -166.085 11.725 -165.755 ;
        RECT 11.395 -167.445 11.725 -167.115 ;
        RECT 11.395 -168.805 11.725 -168.475 ;
        RECT 11.395 -170.165 11.725 -169.835 ;
        RECT 11.395 -171.525 11.725 -171.195 ;
        RECT 11.395 -172.885 11.725 -172.555 ;
        RECT 11.395 -174.245 11.725 -173.915 ;
        RECT 11.395 -175.605 11.725 -175.275 ;
        RECT 11.395 -176.965 11.725 -176.635 ;
        RECT 11.395 -178.325 11.725 -177.995 ;
        RECT 11.395 -179.685 11.725 -179.355 ;
        RECT 11.395 -181.93 11.725 -180.8 ;
        RECT 11.4 -182.045 11.72 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 241.32 13.085 242.45 ;
        RECT 12.755 239.195 13.085 239.525 ;
        RECT 12.755 237.835 13.085 238.165 ;
        RECT 12.76 237.16 13.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 -1.525 13.085 -1.195 ;
        RECT 12.755 -2.885 13.085 -2.555 ;
        RECT 12.76 -3.56 13.08 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 12.755 -95.365 13.085 -95.035 ;
        RECT 12.755 -96.725 13.085 -96.395 ;
        RECT 12.755 -98.085 13.085 -97.755 ;
        RECT 12.755 -99.445 13.085 -99.115 ;
        RECT 12.755 -100.805 13.085 -100.475 ;
        RECT 12.755 -102.165 13.085 -101.835 ;
        RECT 12.755 -103.525 13.085 -103.195 ;
        RECT 12.755 -104.885 13.085 -104.555 ;
        RECT 12.755 -106.245 13.085 -105.915 ;
        RECT 12.755 -107.605 13.085 -107.275 ;
        RECT 12.755 -108.965 13.085 -108.635 ;
        RECT 12.755 -110.325 13.085 -109.995 ;
        RECT 12.755 -111.685 13.085 -111.355 ;
        RECT 12.755 -113.045 13.085 -112.715 ;
        RECT 12.755 -114.405 13.085 -114.075 ;
        RECT 12.755 -115.765 13.085 -115.435 ;
        RECT 12.755 -117.125 13.085 -116.795 ;
        RECT 12.755 -118.485 13.085 -118.155 ;
        RECT 12.755 -119.845 13.085 -119.515 ;
        RECT 12.755 -121.205 13.085 -120.875 ;
        RECT 12.755 -122.565 13.085 -122.235 ;
        RECT 12.755 -123.925 13.085 -123.595 ;
        RECT 12.755 -125.285 13.085 -124.955 ;
        RECT 12.755 -126.645 13.085 -126.315 ;
        RECT 12.755 -128.005 13.085 -127.675 ;
        RECT 12.755 -129.365 13.085 -129.035 ;
        RECT 12.755 -130.725 13.085 -130.395 ;
        RECT 12.755 -132.085 13.085 -131.755 ;
        RECT 12.755 -133.445 13.085 -133.115 ;
        RECT 12.755 -134.805 13.085 -134.475 ;
        RECT 12.755 -136.165 13.085 -135.835 ;
        RECT 12.755 -137.525 13.085 -137.195 ;
        RECT 12.755 -138.885 13.085 -138.555 ;
        RECT 12.755 -140.245 13.085 -139.915 ;
        RECT 12.755 -141.605 13.085 -141.275 ;
        RECT 12.755 -142.965 13.085 -142.635 ;
        RECT 12.755 -144.325 13.085 -143.995 ;
        RECT 12.755 -145.685 13.085 -145.355 ;
        RECT 12.755 -147.045 13.085 -146.715 ;
        RECT 12.755 -148.405 13.085 -148.075 ;
        RECT 12.755 -149.765 13.085 -149.435 ;
        RECT 12.755 -151.125 13.085 -150.795 ;
        RECT 12.755 -152.485 13.085 -152.155 ;
        RECT 12.755 -153.845 13.085 -153.515 ;
        RECT 12.755 -155.205 13.085 -154.875 ;
        RECT 12.755 -156.565 13.085 -156.235 ;
        RECT 12.755 -157.925 13.085 -157.595 ;
        RECT 12.755 -159.285 13.085 -158.955 ;
        RECT 12.755 -160.645 13.085 -160.315 ;
        RECT 12.755 -162.005 13.085 -161.675 ;
        RECT 12.755 -163.365 13.085 -163.035 ;
        RECT 12.755 -164.725 13.085 -164.395 ;
        RECT 12.755 -166.085 13.085 -165.755 ;
        RECT 12.755 -167.445 13.085 -167.115 ;
        RECT 12.755 -168.805 13.085 -168.475 ;
        RECT 12.755 -170.165 13.085 -169.835 ;
        RECT 12.755 -171.525 13.085 -171.195 ;
        RECT 12.755 -172.885 13.085 -172.555 ;
        RECT 12.755 -174.245 13.085 -173.915 ;
        RECT 12.755 -175.605 13.085 -175.275 ;
        RECT 12.755 -176.965 13.085 -176.635 ;
        RECT 12.755 -178.325 13.085 -177.995 ;
        RECT 12.755 -179.685 13.085 -179.355 ;
        RECT 12.755 -181.93 13.085 -180.8 ;
        RECT 12.76 -182.045 13.08 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 241.32 14.445 242.45 ;
        RECT 14.115 239.195 14.445 239.525 ;
        RECT 14.115 237.835 14.445 238.165 ;
        RECT 14.12 237.16 14.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.115 -99.445 14.445 -99.115 ;
        RECT 14.115 -100.805 14.445 -100.475 ;
        RECT 14.115 -102.165 14.445 -101.835 ;
        RECT 14.115 -103.525 14.445 -103.195 ;
        RECT 14.115 -104.885 14.445 -104.555 ;
        RECT 14.115 -106.245 14.445 -105.915 ;
        RECT 14.115 -107.605 14.445 -107.275 ;
        RECT 14.115 -108.965 14.445 -108.635 ;
        RECT 14.115 -110.325 14.445 -109.995 ;
        RECT 14.115 -111.685 14.445 -111.355 ;
        RECT 14.115 -113.045 14.445 -112.715 ;
        RECT 14.115 -114.405 14.445 -114.075 ;
        RECT 14.115 -115.765 14.445 -115.435 ;
        RECT 14.115 -117.125 14.445 -116.795 ;
        RECT 14.115 -118.485 14.445 -118.155 ;
        RECT 14.115 -119.845 14.445 -119.515 ;
        RECT 14.115 -121.205 14.445 -120.875 ;
        RECT 14.115 -122.565 14.445 -122.235 ;
        RECT 14.115 -123.925 14.445 -123.595 ;
        RECT 14.115 -125.285 14.445 -124.955 ;
        RECT 14.115 -126.645 14.445 -126.315 ;
        RECT 14.115 -128.005 14.445 -127.675 ;
        RECT 14.115 -129.365 14.445 -129.035 ;
        RECT 14.115 -130.725 14.445 -130.395 ;
        RECT 14.115 -132.085 14.445 -131.755 ;
        RECT 14.115 -133.445 14.445 -133.115 ;
        RECT 14.115 -134.805 14.445 -134.475 ;
        RECT 14.115 -136.165 14.445 -135.835 ;
        RECT 14.115 -137.525 14.445 -137.195 ;
        RECT 14.115 -138.885 14.445 -138.555 ;
        RECT 14.115 -140.245 14.445 -139.915 ;
        RECT 14.115 -141.605 14.445 -141.275 ;
        RECT 14.115 -142.965 14.445 -142.635 ;
        RECT 14.115 -144.325 14.445 -143.995 ;
        RECT 14.115 -145.685 14.445 -145.355 ;
        RECT 14.115 -147.045 14.445 -146.715 ;
        RECT 14.115 -148.405 14.445 -148.075 ;
        RECT 14.115 -149.765 14.445 -149.435 ;
        RECT 14.115 -151.125 14.445 -150.795 ;
        RECT 14.115 -152.485 14.445 -152.155 ;
        RECT 14.115 -153.845 14.445 -153.515 ;
        RECT 14.115 -155.205 14.445 -154.875 ;
        RECT 14.115 -156.565 14.445 -156.235 ;
        RECT 14.115 -157.925 14.445 -157.595 ;
        RECT 14.115 -159.285 14.445 -158.955 ;
        RECT 14.115 -160.645 14.445 -160.315 ;
        RECT 14.115 -162.005 14.445 -161.675 ;
        RECT 14.115 -163.365 14.445 -163.035 ;
        RECT 14.115 -164.725 14.445 -164.395 ;
        RECT 14.115 -166.085 14.445 -165.755 ;
        RECT 14.115 -167.445 14.445 -167.115 ;
        RECT 14.115 -168.805 14.445 -168.475 ;
        RECT 14.115 -170.165 14.445 -169.835 ;
        RECT 14.115 -171.525 14.445 -171.195 ;
        RECT 14.115 -172.885 14.445 -172.555 ;
        RECT 14.115 -174.245 14.445 -173.915 ;
        RECT 14.115 -175.605 14.445 -175.275 ;
        RECT 14.115 -176.965 14.445 -176.635 ;
        RECT 14.115 -178.325 14.445 -177.995 ;
        RECT 14.115 -179.685 14.445 -179.355 ;
        RECT 14.115 -181.93 14.445 -180.8 ;
        RECT 14.12 -182.045 14.44 -98.44 ;
    END
    PORT
      LAYER met3 ;
        RECT 14.21 -98.075 14.54 -0.51 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 241.32 15.805 242.45 ;
        RECT 15.475 239.195 15.805 239.525 ;
        RECT 15.475 237.835 15.805 238.165 ;
        RECT 15.48 237.16 15.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 15.475 -1.525 15.805 -1.195 ;
        RECT 15.475 -2.885 15.805 -2.555 ;
        RECT 15.48 -3.56 15.8 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 241.32 17.165 242.45 ;
        RECT 16.835 239.195 17.165 239.525 ;
        RECT 16.835 237.835 17.165 238.165 ;
        RECT 16.84 237.16 17.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 16.835 -1.525 17.165 -1.195 ;
        RECT 16.835 -2.885 17.165 -2.555 ;
        RECT 16.84 -3.56 17.16 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 241.32 18.525 242.45 ;
        RECT 18.195 239.195 18.525 239.525 ;
        RECT 18.195 237.835 18.525 238.165 ;
        RECT 18.2 237.16 18.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 -1.525 18.525 -1.195 ;
        RECT 18.195 -2.885 18.525 -2.555 ;
        RECT 18.2 -3.56 18.52 -0.52 ;
    END
    PORT
      LAYER met3 ;
        RECT 18.195 -95.365 18.525 -95.035 ;
        RECT 18.195 -96.725 18.525 -96.395 ;
        RECT 18.195 -98.085 18.525 -97.755 ;
        RECT 18.195 -99.445 18.525 -99.115 ;
        RECT 18.195 -100.805 18.525 -100.475 ;
        RECT 18.195 -102.165 18.525 -101.835 ;
        RECT 18.195 -103.525 18.525 -103.195 ;
        RECT 18.195 -104.885 18.525 -104.555 ;
        RECT 18.195 -106.245 18.525 -105.915 ;
        RECT 18.195 -107.605 18.525 -107.275 ;
        RECT 18.195 -108.965 18.525 -108.635 ;
        RECT 18.195 -110.325 18.525 -109.995 ;
        RECT 18.195 -111.685 18.525 -111.355 ;
        RECT 18.195 -113.045 18.525 -112.715 ;
        RECT 18.195 -114.405 18.525 -114.075 ;
        RECT 18.195 -115.765 18.525 -115.435 ;
        RECT 18.195 -117.125 18.525 -116.795 ;
        RECT 18.195 -118.485 18.525 -118.155 ;
        RECT 18.195 -119.845 18.525 -119.515 ;
        RECT 18.195 -121.205 18.525 -120.875 ;
        RECT 18.195 -122.565 18.525 -122.235 ;
        RECT 18.195 -123.925 18.525 -123.595 ;
        RECT 18.195 -125.285 18.525 -124.955 ;
        RECT 18.195 -126.645 18.525 -126.315 ;
        RECT 18.195 -128.005 18.525 -127.675 ;
        RECT 18.195 -129.365 18.525 -129.035 ;
        RECT 18.195 -130.725 18.525 -130.395 ;
        RECT 18.195 -132.085 18.525 -131.755 ;
        RECT 18.195 -133.445 18.525 -133.115 ;
        RECT 18.195 -134.805 18.525 -134.475 ;
        RECT 18.195 -136.165 18.525 -135.835 ;
        RECT 18.195 -137.525 18.525 -137.195 ;
        RECT 18.195 -138.885 18.525 -138.555 ;
        RECT 18.195 -140.245 18.525 -139.915 ;
        RECT 18.195 -141.605 18.525 -141.275 ;
        RECT 18.195 -142.965 18.525 -142.635 ;
        RECT 18.195 -144.325 18.525 -143.995 ;
        RECT 18.195 -145.685 18.525 -145.355 ;
        RECT 18.195 -147.045 18.525 -146.715 ;
        RECT 18.195 -148.405 18.525 -148.075 ;
        RECT 18.195 -149.765 18.525 -149.435 ;
        RECT 18.195 -151.125 18.525 -150.795 ;
        RECT 18.195 -152.485 18.525 -152.155 ;
        RECT 18.195 -153.845 18.525 -153.515 ;
        RECT 18.195 -155.205 18.525 -154.875 ;
        RECT 18.195 -156.565 18.525 -156.235 ;
        RECT 18.195 -157.925 18.525 -157.595 ;
        RECT 18.195 -159.285 18.525 -158.955 ;
        RECT 18.195 -160.645 18.525 -160.315 ;
        RECT 18.195 -162.005 18.525 -161.675 ;
        RECT 18.195 -163.365 18.525 -163.035 ;
        RECT 18.195 -164.725 18.525 -164.395 ;
        RECT 18.195 -166.085 18.525 -165.755 ;
        RECT 18.195 -167.445 18.525 -167.115 ;
        RECT 18.195 -168.805 18.525 -168.475 ;
        RECT 18.195 -170.165 18.525 -169.835 ;
        RECT 18.195 -171.525 18.525 -171.195 ;
        RECT 18.195 -172.885 18.525 -172.555 ;
        RECT 18.195 -174.245 18.525 -173.915 ;
        RECT 18.195 -175.605 18.525 -175.275 ;
        RECT 18.195 -176.965 18.525 -176.635 ;
        RECT 18.195 -178.325 18.525 -177.995 ;
        RECT 18.195 -179.685 18.525 -179.355 ;
        RECT 18.195 -181.93 18.525 -180.8 ;
        RECT 18.2 -182.045 18.52 -95.035 ;
    END
    PORT
      LAYER met3 ;
        RECT 19.56 237.16 19.88 242.565 ;
        RECT 19.555 241.32 19.885 242.45 ;
        RECT 19.555 239.195 19.885 239.525 ;
        RECT 19.555 237.835 19.885 238.165 ;
    END
    PORT
      LAYER met3 ;
        RECT -6.285 241.32 -5.955 242.45 ;
        RECT -6.285 239.195 -5.955 239.525 ;
        RECT -6.285 237.835 -5.955 238.165 ;
        RECT -6.285 -1.525 -5.955 -1.195 ;
        RECT -6.285 -2.885 -5.955 -2.555 ;
        RECT -6.285 -4.245 -5.955 -3.915 ;
        RECT -6.285 -5.605 -5.955 -5.275 ;
        RECT -6.285 -6.965 -5.955 -6.635 ;
        RECT -6.285 -8.325 -5.955 -7.995 ;
        RECT -6.285 -9.685 -5.955 -9.355 ;
        RECT -6.285 -12.405 -5.955 -12.075 ;
        RECT -6.285 -13.765 -5.955 -13.435 ;
        RECT -6.285 -15.125 -5.955 -14.795 ;
        RECT -6.285 -16.485 -5.955 -16.155 ;
        RECT -6.285 -17.845 -5.955 -17.515 ;
        RECT -6.285 -24.645 -5.955 -24.315 ;
        RECT -6.285 -26.005 -5.955 -25.675 ;
        RECT -6.285 -27.365 -5.955 -27.035 ;
        RECT -6.285 -28.725 -5.955 -28.395 ;
        RECT -6.285 -30.085 -5.955 -29.755 ;
        RECT -6.285 -31.445 -5.955 -31.115 ;
        RECT -6.285 -32.805 -5.955 -32.475 ;
        RECT -6.285 -34.165 -5.955 -33.835 ;
        RECT -6.285 -35.525 -5.955 -35.195 ;
        RECT -6.285 -36.885 -5.955 -36.555 ;
        RECT -6.285 -38.245 -5.955 -37.915 ;
        RECT -6.285 -39.605 -5.955 -39.275 ;
        RECT -6.285 -42.325 -5.955 -41.995 ;
        RECT -6.285 -45.045 -5.955 -44.715 ;
        RECT -6.285 -46.405 -5.955 -46.075 ;
        RECT -6.285 -47.765 -5.955 -47.435 ;
        RECT -6.285 -49.125 -5.955 -48.795 ;
        RECT -6.285 -51.845 -5.955 -51.515 ;
        RECT -6.285 -53.205 -5.955 -52.875 ;
        RECT -6.285 -54.565 -5.955 -54.235 ;
        RECT -6.285 -55.925 -5.955 -55.595 ;
        RECT -6.285 -57.285 -5.955 -56.955 ;
        RECT -6.285 -58.645 -5.955 -58.315 ;
        RECT -6.285 -60.005 -5.955 -59.675 ;
        RECT -6.285 -61.365 -5.955 -61.035 ;
        RECT -6.285 -62.725 -5.955 -62.395 ;
        RECT -6.285 -64.085 -5.955 -63.755 ;
        RECT -6.285 -65.445 -5.955 -65.115 ;
        RECT -6.285 -68.165 -5.955 -67.835 ;
        RECT -6.285 -69.525 -5.955 -69.195 ;
        RECT -6.285 -70.885 -5.955 -70.555 ;
        RECT -6.285 -72.245 -5.955 -71.915 ;
        RECT -6.285 -73.605 -5.955 -73.275 ;
        RECT -6.285 -74.965 -5.955 -74.635 ;
        RECT -6.285 -76.325 -5.955 -75.995 ;
        RECT -6.285 -77.685 -5.955 -77.355 ;
        RECT -6.285 -79.045 -5.955 -78.715 ;
        RECT -6.285 -80.405 -5.955 -80.075 ;
        RECT -6.285 -81.765 -5.955 -81.435 ;
        RECT -6.285 -83.125 -5.955 -82.795 ;
        RECT -6.285 -84.485 -5.955 -84.155 ;
        RECT -6.285 -85.845 -5.955 -85.515 ;
        RECT -6.285 -87.205 -5.955 -86.875 ;
        RECT -6.285 -88.565 -5.955 -88.235 ;
        RECT -6.285 -91.285 -5.955 -90.955 ;
        RECT -6.285 -92.645 -5.955 -92.315 ;
        RECT -6.285 -94.005 -5.955 -93.675 ;
        RECT -6.285 -95.365 -5.955 -95.035 ;
        RECT -6.285 -96.725 -5.955 -96.395 ;
        RECT -6.285 -98.085 -5.955 -97.755 ;
        RECT -6.285 -99.445 -5.955 -99.115 ;
        RECT -6.285 -100.805 -5.955 -100.475 ;
        RECT -6.285 -102.165 -5.955 -101.835 ;
        RECT -6.285 -103.525 -5.955 -103.195 ;
        RECT -6.285 -104.885 -5.955 -104.555 ;
        RECT -6.285 -106.245 -5.955 -105.915 ;
        RECT -6.285 -107.605 -5.955 -107.275 ;
        RECT -6.285 -108.965 -5.955 -108.635 ;
        RECT -6.285 -110.325 -5.955 -109.995 ;
        RECT -6.285 -111.685 -5.955 -111.355 ;
        RECT -6.285 -113.045 -5.955 -112.715 ;
        RECT -6.285 -114.405 -5.955 -114.075 ;
        RECT -6.285 -115.765 -5.955 -115.435 ;
        RECT -6.285 -117.125 -5.955 -116.795 ;
        RECT -6.285 -118.485 -5.955 -118.155 ;
        RECT -6.285 -119.845 -5.955 -119.515 ;
        RECT -6.285 -121.205 -5.955 -120.875 ;
        RECT -6.285 -122.565 -5.955 -122.235 ;
        RECT -6.285 -123.925 -5.955 -123.595 ;
        RECT -6.285 -125.285 -5.955 -124.955 ;
        RECT -6.285 -126.645 -5.955 -126.315 ;
        RECT -6.285 -128.005 -5.955 -127.675 ;
        RECT -6.285 -129.365 -5.955 -129.035 ;
        RECT -6.285 -130.725 -5.955 -130.395 ;
        RECT -6.285 -132.085 -5.955 -131.755 ;
        RECT -6.285 -133.445 -5.955 -133.115 ;
        RECT -6.285 -134.805 -5.955 -134.475 ;
        RECT -6.285 -136.165 -5.955 -135.835 ;
        RECT -6.285 -137.525 -5.955 -137.195 ;
        RECT -6.285 -138.885 -5.955 -138.555 ;
        RECT -6.285 -140.245 -5.955 -139.915 ;
        RECT -6.285 -141.605 -5.955 -141.275 ;
        RECT -6.285 -142.965 -5.955 -142.635 ;
        RECT -6.285 -144.325 -5.955 -143.995 ;
        RECT -6.285 -145.685 -5.955 -145.355 ;
        RECT -6.285 -147.045 -5.955 -146.715 ;
        RECT -6.285 -148.405 -5.955 -148.075 ;
        RECT -6.285 -149.765 -5.955 -149.435 ;
        RECT -6.285 -151.125 -5.955 -150.795 ;
        RECT -6.285 -152.485 -5.955 -152.155 ;
        RECT -6.285 -153.845 -5.955 -153.515 ;
        RECT -6.285 -155.205 -5.955 -154.875 ;
        RECT -6.285 -156.565 -5.955 -156.235 ;
        RECT -6.285 -157.925 -5.955 -157.595 ;
        RECT -6.285 -159.285 -5.955 -158.955 ;
        RECT -6.285 -160.645 -5.955 -160.315 ;
        RECT -6.285 -162.005 -5.955 -161.675 ;
        RECT -6.285 -163.365 -5.955 -163.035 ;
        RECT -6.285 -164.725 -5.955 -164.395 ;
        RECT -6.285 -166.085 -5.955 -165.755 ;
        RECT -6.285 -167.445 -5.955 -167.115 ;
        RECT -6.285 -168.805 -5.955 -168.475 ;
        RECT -6.285 -170.165 -5.955 -169.835 ;
        RECT -6.285 -171.525 -5.955 -171.195 ;
        RECT -6.285 -172.885 -5.955 -172.555 ;
        RECT -6.285 -174.245 -5.955 -173.915 ;
        RECT -6.285 -175.605 -5.955 -175.275 ;
        RECT -6.285 -176.965 -5.955 -176.635 ;
        RECT -6.285 -178.325 -5.955 -177.995 ;
        RECT -6.285 -179.685 -5.955 -179.355 ;
        RECT -6.285 -181.93 -5.955 -180.8 ;
        RECT -6.28 -182.045 -5.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -4.925 241.32 -4.595 242.45 ;
        RECT -4.925 239.195 -4.595 239.525 ;
        RECT -4.925 237.835 -4.595 238.165 ;
        RECT -4.925 235.975 -4.595 236.305 ;
        RECT -4.925 233.925 -4.595 234.255 ;
        RECT -4.925 231.995 -4.595 232.325 ;
        RECT -4.925 230.155 -4.595 230.485 ;
        RECT -4.925 228.665 -4.595 228.995 ;
        RECT -4.925 226.995 -4.595 227.325 ;
        RECT -4.925 225.505 -4.595 225.835 ;
        RECT -4.925 223.835 -4.595 224.165 ;
        RECT -4.925 222.345 -4.595 222.675 ;
        RECT -4.925 220.675 -4.595 221.005 ;
        RECT -4.925 219.185 -4.595 219.515 ;
        RECT -4.925 217.775 -4.595 218.105 ;
        RECT -4.925 215.935 -4.595 216.265 ;
        RECT -4.925 214.445 -4.595 214.775 ;
        RECT -4.925 212.775 -4.595 213.105 ;
        RECT -4.925 211.285 -4.595 211.615 ;
        RECT -4.925 209.615 -4.595 209.945 ;
        RECT -4.925 208.125 -4.595 208.455 ;
        RECT -4.925 206.455 -4.595 206.785 ;
        RECT -4.925 204.965 -4.595 205.295 ;
        RECT -4.925 203.555 -4.595 203.885 ;
        RECT -4.925 201.715 -4.595 202.045 ;
        RECT -4.925 200.225 -4.595 200.555 ;
        RECT -4.925 198.555 -4.595 198.885 ;
        RECT -4.925 197.065 -4.595 197.395 ;
        RECT -4.925 195.395 -4.595 195.725 ;
        RECT -4.925 193.905 -4.595 194.235 ;
        RECT -4.925 192.235 -4.595 192.565 ;
        RECT -4.925 190.745 -4.595 191.075 ;
        RECT -4.925 189.335 -4.595 189.665 ;
        RECT -4.925 187.495 -4.595 187.825 ;
        RECT -4.925 186.005 -4.595 186.335 ;
        RECT -4.925 184.335 -4.595 184.665 ;
        RECT -4.925 182.845 -4.595 183.175 ;
        RECT -4.925 181.175 -4.595 181.505 ;
        RECT -4.925 179.685 -4.595 180.015 ;
        RECT -4.925 178.015 -4.595 178.345 ;
        RECT -4.925 176.525 -4.595 176.855 ;
        RECT -4.925 175.115 -4.595 175.445 ;
        RECT -4.925 173.275 -4.595 173.605 ;
        RECT -4.925 171.785 -4.595 172.115 ;
        RECT -4.925 170.115 -4.595 170.445 ;
        RECT -4.925 168.625 -4.595 168.955 ;
        RECT -4.925 166.955 -4.595 167.285 ;
        RECT -4.925 165.465 -4.595 165.795 ;
        RECT -4.925 163.795 -4.595 164.125 ;
        RECT -4.925 162.305 -4.595 162.635 ;
        RECT -4.925 160.895 -4.595 161.225 ;
        RECT -4.925 159.055 -4.595 159.385 ;
        RECT -4.925 157.565 -4.595 157.895 ;
        RECT -4.925 155.895 -4.595 156.225 ;
        RECT -4.925 154.405 -4.595 154.735 ;
        RECT -4.925 152.735 -4.595 153.065 ;
        RECT -4.925 151.245 -4.595 151.575 ;
        RECT -4.925 149.575 -4.595 149.905 ;
        RECT -4.925 148.085 -4.595 148.415 ;
        RECT -4.925 146.675 -4.595 147.005 ;
        RECT -4.925 144.835 -4.595 145.165 ;
        RECT -4.925 143.345 -4.595 143.675 ;
        RECT -4.925 141.675 -4.595 142.005 ;
        RECT -4.925 140.185 -4.595 140.515 ;
        RECT -4.925 138.515 -4.595 138.845 ;
        RECT -4.925 137.025 -4.595 137.355 ;
        RECT -4.925 135.355 -4.595 135.685 ;
        RECT -4.925 133.865 -4.595 134.195 ;
        RECT -4.925 132.455 -4.595 132.785 ;
        RECT -4.925 130.615 -4.595 130.945 ;
        RECT -4.925 129.125 -4.595 129.455 ;
        RECT -4.925 127.455 -4.595 127.785 ;
        RECT -4.925 125.965 -4.595 126.295 ;
        RECT -4.925 124.295 -4.595 124.625 ;
        RECT -4.925 122.805 -4.595 123.135 ;
        RECT -4.925 121.135 -4.595 121.465 ;
        RECT -4.925 119.645 -4.595 119.975 ;
        RECT -4.925 118.235 -4.595 118.565 ;
        RECT -4.925 116.395 -4.595 116.725 ;
        RECT -4.925 114.905 -4.595 115.235 ;
        RECT -4.925 113.235 -4.595 113.565 ;
        RECT -4.925 111.745 -4.595 112.075 ;
        RECT -4.925 110.075 -4.595 110.405 ;
        RECT -4.925 108.585 -4.595 108.915 ;
        RECT -4.925 106.915 -4.595 107.245 ;
        RECT -4.925 105.425 -4.595 105.755 ;
        RECT -4.925 104.015 -4.595 104.345 ;
        RECT -4.925 102.175 -4.595 102.505 ;
        RECT -4.925 100.685 -4.595 101.015 ;
        RECT -4.925 99.015 -4.595 99.345 ;
        RECT -4.925 97.525 -4.595 97.855 ;
        RECT -4.925 95.855 -4.595 96.185 ;
        RECT -4.925 94.365 -4.595 94.695 ;
        RECT -4.925 92.695 -4.595 93.025 ;
        RECT -4.925 91.205 -4.595 91.535 ;
        RECT -4.925 89.795 -4.595 90.125 ;
        RECT -4.925 87.955 -4.595 88.285 ;
        RECT -4.925 86.465 -4.595 86.795 ;
        RECT -4.925 84.795 -4.595 85.125 ;
        RECT -4.925 83.305 -4.595 83.635 ;
        RECT -4.925 81.635 -4.595 81.965 ;
        RECT -4.925 80.145 -4.595 80.475 ;
        RECT -4.925 78.475 -4.595 78.805 ;
        RECT -4.925 76.985 -4.595 77.315 ;
        RECT -4.925 75.575 -4.595 75.905 ;
        RECT -4.925 73.735 -4.595 74.065 ;
        RECT -4.925 72.245 -4.595 72.575 ;
        RECT -4.925 70.575 -4.595 70.905 ;
        RECT -4.925 69.085 -4.595 69.415 ;
        RECT -4.925 67.415 -4.595 67.745 ;
        RECT -4.925 65.925 -4.595 66.255 ;
        RECT -4.925 64.255 -4.595 64.585 ;
        RECT -4.925 62.765 -4.595 63.095 ;
        RECT -4.925 61.355 -4.595 61.685 ;
        RECT -4.925 59.515 -4.595 59.845 ;
        RECT -4.925 58.025 -4.595 58.355 ;
        RECT -4.925 56.355 -4.595 56.685 ;
        RECT -4.925 54.865 -4.595 55.195 ;
        RECT -4.925 53.195 -4.595 53.525 ;
        RECT -4.925 51.705 -4.595 52.035 ;
        RECT -4.925 50.035 -4.595 50.365 ;
        RECT -4.925 48.545 -4.595 48.875 ;
        RECT -4.925 47.135 -4.595 47.465 ;
        RECT -4.925 45.295 -4.595 45.625 ;
        RECT -4.925 43.805 -4.595 44.135 ;
        RECT -4.925 42.135 -4.595 42.465 ;
        RECT -4.925 40.645 -4.595 40.975 ;
        RECT -4.925 38.975 -4.595 39.305 ;
        RECT -4.925 37.485 -4.595 37.815 ;
        RECT -4.925 35.815 -4.595 36.145 ;
        RECT -4.925 34.325 -4.595 34.655 ;
        RECT -4.925 32.915 -4.595 33.245 ;
        RECT -4.925 31.075 -4.595 31.405 ;
        RECT -4.925 29.585 -4.595 29.915 ;
        RECT -4.925 27.915 -4.595 28.245 ;
        RECT -4.925 26.425 -4.595 26.755 ;
        RECT -4.925 24.755 -4.595 25.085 ;
        RECT -4.925 23.265 -4.595 23.595 ;
        RECT -4.925 21.595 -4.595 21.925 ;
        RECT -4.925 20.105 -4.595 20.435 ;
        RECT -4.925 18.695 -4.595 19.025 ;
        RECT -4.925 16.855 -4.595 17.185 ;
        RECT -4.925 15.365 -4.595 15.695 ;
        RECT -4.925 13.695 -4.595 14.025 ;
        RECT -4.925 12.205 -4.595 12.535 ;
        RECT -4.925 10.535 -4.595 10.865 ;
        RECT -4.925 9.045 -4.595 9.375 ;
        RECT -4.925 7.375 -4.595 7.705 ;
        RECT -4.925 5.885 -4.595 6.215 ;
        RECT -4.925 4.475 -4.595 4.805 ;
        RECT -4.925 2.115 -4.595 2.445 ;
        RECT -4.925 0.06 -4.595 0.39 ;
        RECT -4.925 -1.525 -4.595 -1.195 ;
        RECT -4.925 -2.885 -4.595 -2.555 ;
        RECT -4.925 -4.245 -4.595 -3.915 ;
        RECT -4.925 -5.605 -4.595 -5.275 ;
        RECT -4.925 -6.965 -4.595 -6.635 ;
        RECT -4.925 -8.325 -4.595 -7.995 ;
        RECT -4.925 -9.685 -4.595 -9.355 ;
        RECT -4.925 -12.405 -4.595 -12.075 ;
        RECT -4.925 -13.765 -4.595 -13.435 ;
        RECT -4.925 -15.125 -4.595 -14.795 ;
        RECT -4.925 -16.485 -4.595 -16.155 ;
        RECT -4.925 -17.845 -4.595 -17.515 ;
        RECT -4.925 -24.645 -4.595 -24.315 ;
        RECT -4.925 -26.005 -4.595 -25.675 ;
        RECT -4.925 -27.365 -4.595 -27.035 ;
        RECT -4.925 -28.725 -4.595 -28.395 ;
        RECT -4.925 -30.085 -4.595 -29.755 ;
        RECT -4.925 -31.445 -4.595 -31.115 ;
        RECT -4.925 -32.805 -4.595 -32.475 ;
        RECT -4.925 -34.165 -4.595 -33.835 ;
        RECT -4.925 -35.525 -4.595 -35.195 ;
        RECT -4.925 -36.885 -4.595 -36.555 ;
        RECT -4.925 -38.245 -4.595 -37.915 ;
        RECT -4.925 -39.605 -4.595 -39.275 ;
        RECT -4.925 -42.325 -4.595 -41.995 ;
        RECT -4.925 -45.045 -4.595 -44.715 ;
        RECT -4.925 -46.405 -4.595 -46.075 ;
        RECT -4.925 -47.765 -4.595 -47.435 ;
        RECT -4.925 -49.125 -4.595 -48.795 ;
        RECT -4.925 -51.845 -4.595 -51.515 ;
        RECT -4.925 -53.205 -4.595 -52.875 ;
        RECT -4.925 -54.565 -4.595 -54.235 ;
        RECT -4.925 -55.925 -4.595 -55.595 ;
        RECT -4.925 -57.285 -4.595 -56.955 ;
        RECT -4.925 -58.645 -4.595 -58.315 ;
        RECT -4.925 -60.005 -4.595 -59.675 ;
        RECT -4.925 -61.365 -4.595 -61.035 ;
        RECT -4.925 -62.725 -4.595 -62.395 ;
        RECT -4.925 -64.085 -4.595 -63.755 ;
        RECT -4.925 -65.445 -4.595 -65.115 ;
        RECT -4.925 -68.165 -4.595 -67.835 ;
        RECT -4.925 -69.525 -4.595 -69.195 ;
        RECT -4.925 -70.885 -4.595 -70.555 ;
        RECT -4.925 -72.245 -4.595 -71.915 ;
        RECT -4.925 -73.605 -4.595 -73.275 ;
        RECT -4.925 -74.965 -4.595 -74.635 ;
        RECT -4.925 -76.325 -4.595 -75.995 ;
        RECT -4.925 -77.685 -4.595 -77.355 ;
        RECT -4.925 -79.045 -4.595 -78.715 ;
        RECT -4.925 -80.405 -4.595 -80.075 ;
        RECT -4.925 -81.765 -4.595 -81.435 ;
        RECT -4.925 -83.125 -4.595 -82.795 ;
        RECT -4.925 -84.485 -4.595 -84.155 ;
        RECT -4.925 -85.845 -4.595 -85.515 ;
        RECT -4.925 -87.205 -4.595 -86.875 ;
        RECT -4.925 -88.565 -4.595 -88.235 ;
        RECT -4.925 -91.285 -4.595 -90.955 ;
        RECT -4.925 -92.645 -4.595 -92.315 ;
        RECT -4.925 -94.005 -4.595 -93.675 ;
        RECT -4.925 -95.365 -4.595 -95.035 ;
        RECT -4.925 -96.725 -4.595 -96.395 ;
        RECT -4.925 -98.085 -4.595 -97.755 ;
        RECT -4.925 -99.445 -4.595 -99.115 ;
        RECT -4.925 -100.805 -4.595 -100.475 ;
        RECT -4.925 -102.165 -4.595 -101.835 ;
        RECT -4.925 -103.525 -4.595 -103.195 ;
        RECT -4.925 -104.885 -4.595 -104.555 ;
        RECT -4.925 -106.245 -4.595 -105.915 ;
        RECT -4.925 -107.605 -4.595 -107.275 ;
        RECT -4.925 -108.965 -4.595 -108.635 ;
        RECT -4.925 -110.325 -4.595 -109.995 ;
        RECT -4.925 -111.685 -4.595 -111.355 ;
        RECT -4.925 -113.045 -4.595 -112.715 ;
        RECT -4.925 -114.405 -4.595 -114.075 ;
        RECT -4.925 -115.765 -4.595 -115.435 ;
        RECT -4.925 -117.125 -4.595 -116.795 ;
        RECT -4.925 -118.485 -4.595 -118.155 ;
        RECT -4.925 -119.845 -4.595 -119.515 ;
        RECT -4.925 -121.205 -4.595 -120.875 ;
        RECT -4.925 -122.565 -4.595 -122.235 ;
        RECT -4.925 -123.925 -4.595 -123.595 ;
        RECT -4.925 -125.285 -4.595 -124.955 ;
        RECT -4.925 -126.645 -4.595 -126.315 ;
        RECT -4.925 -128.005 -4.595 -127.675 ;
        RECT -4.925 -129.365 -4.595 -129.035 ;
        RECT -4.925 -130.725 -4.595 -130.395 ;
        RECT -4.925 -132.085 -4.595 -131.755 ;
        RECT -4.925 -133.445 -4.595 -133.115 ;
        RECT -4.925 -134.805 -4.595 -134.475 ;
        RECT -4.925 -136.165 -4.595 -135.835 ;
        RECT -4.925 -137.525 -4.595 -137.195 ;
        RECT -4.925 -138.885 -4.595 -138.555 ;
        RECT -4.925 -140.245 -4.595 -139.915 ;
        RECT -4.925 -141.605 -4.595 -141.275 ;
        RECT -4.925 -142.965 -4.595 -142.635 ;
        RECT -4.925 -144.325 -4.595 -143.995 ;
        RECT -4.925 -145.685 -4.595 -145.355 ;
        RECT -4.925 -147.045 -4.595 -146.715 ;
        RECT -4.925 -148.405 -4.595 -148.075 ;
        RECT -4.925 -149.765 -4.595 -149.435 ;
        RECT -4.925 -151.125 -4.595 -150.795 ;
        RECT -4.925 -152.485 -4.595 -152.155 ;
        RECT -4.925 -153.845 -4.595 -153.515 ;
        RECT -4.925 -155.205 -4.595 -154.875 ;
        RECT -4.925 -156.565 -4.595 -156.235 ;
        RECT -4.925 -157.925 -4.595 -157.595 ;
        RECT -4.925 -159.285 -4.595 -158.955 ;
        RECT -4.925 -160.645 -4.595 -160.315 ;
        RECT -4.925 -162.005 -4.595 -161.675 ;
        RECT -4.925 -163.365 -4.595 -163.035 ;
        RECT -4.925 -164.725 -4.595 -164.395 ;
        RECT -4.925 -166.085 -4.595 -165.755 ;
        RECT -4.925 -167.445 -4.595 -167.115 ;
        RECT -4.925 -168.805 -4.595 -168.475 ;
        RECT -4.925 -170.165 -4.595 -169.835 ;
        RECT -4.925 -171.525 -4.595 -171.195 ;
        RECT -4.925 -172.885 -4.595 -172.555 ;
        RECT -4.925 -174.245 -4.595 -173.915 ;
        RECT -4.925 -175.605 -4.595 -175.275 ;
        RECT -4.925 -176.965 -4.595 -176.635 ;
        RECT -4.925 -178.325 -4.595 -177.995 ;
        RECT -4.925 -179.685 -4.595 -179.355 ;
        RECT -4.925 -181.93 -4.595 -180.8 ;
        RECT -4.92 -182.045 -4.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -3.565 241.32 -3.235 242.45 ;
        RECT -3.565 239.195 -3.235 239.525 ;
        RECT -3.565 237.835 -3.235 238.165 ;
        RECT -3.565 235.975 -3.235 236.305 ;
        RECT -3.565 233.925 -3.235 234.255 ;
        RECT -3.565 231.995 -3.235 232.325 ;
        RECT -3.565 230.155 -3.235 230.485 ;
        RECT -3.565 228.665 -3.235 228.995 ;
        RECT -3.565 226.995 -3.235 227.325 ;
        RECT -3.565 225.505 -3.235 225.835 ;
        RECT -3.565 223.835 -3.235 224.165 ;
        RECT -3.565 222.345 -3.235 222.675 ;
        RECT -3.565 220.675 -3.235 221.005 ;
        RECT -3.565 219.185 -3.235 219.515 ;
        RECT -3.565 217.775 -3.235 218.105 ;
        RECT -3.565 215.935 -3.235 216.265 ;
        RECT -3.565 214.445 -3.235 214.775 ;
        RECT -3.565 212.775 -3.235 213.105 ;
        RECT -3.565 211.285 -3.235 211.615 ;
        RECT -3.565 209.615 -3.235 209.945 ;
        RECT -3.565 208.125 -3.235 208.455 ;
        RECT -3.565 206.455 -3.235 206.785 ;
        RECT -3.565 204.965 -3.235 205.295 ;
        RECT -3.565 203.555 -3.235 203.885 ;
        RECT -3.565 201.715 -3.235 202.045 ;
        RECT -3.565 200.225 -3.235 200.555 ;
        RECT -3.565 198.555 -3.235 198.885 ;
        RECT -3.565 197.065 -3.235 197.395 ;
        RECT -3.565 195.395 -3.235 195.725 ;
        RECT -3.565 193.905 -3.235 194.235 ;
        RECT -3.565 192.235 -3.235 192.565 ;
        RECT -3.565 190.745 -3.235 191.075 ;
        RECT -3.565 189.335 -3.235 189.665 ;
        RECT -3.565 187.495 -3.235 187.825 ;
        RECT -3.565 186.005 -3.235 186.335 ;
        RECT -3.565 184.335 -3.235 184.665 ;
        RECT -3.565 182.845 -3.235 183.175 ;
        RECT -3.565 181.175 -3.235 181.505 ;
        RECT -3.565 179.685 -3.235 180.015 ;
        RECT -3.565 178.015 -3.235 178.345 ;
        RECT -3.565 176.525 -3.235 176.855 ;
        RECT -3.565 175.115 -3.235 175.445 ;
        RECT -3.565 173.275 -3.235 173.605 ;
        RECT -3.565 171.785 -3.235 172.115 ;
        RECT -3.565 170.115 -3.235 170.445 ;
        RECT -3.565 168.625 -3.235 168.955 ;
        RECT -3.565 166.955 -3.235 167.285 ;
        RECT -3.565 165.465 -3.235 165.795 ;
        RECT -3.565 163.795 -3.235 164.125 ;
        RECT -3.565 162.305 -3.235 162.635 ;
        RECT -3.565 160.895 -3.235 161.225 ;
        RECT -3.565 159.055 -3.235 159.385 ;
        RECT -3.565 157.565 -3.235 157.895 ;
        RECT -3.565 155.895 -3.235 156.225 ;
        RECT -3.565 154.405 -3.235 154.735 ;
        RECT -3.565 152.735 -3.235 153.065 ;
        RECT -3.565 151.245 -3.235 151.575 ;
        RECT -3.565 149.575 -3.235 149.905 ;
        RECT -3.565 148.085 -3.235 148.415 ;
        RECT -3.565 146.675 -3.235 147.005 ;
        RECT -3.565 144.835 -3.235 145.165 ;
        RECT -3.565 143.345 -3.235 143.675 ;
        RECT -3.565 141.675 -3.235 142.005 ;
        RECT -3.565 140.185 -3.235 140.515 ;
        RECT -3.565 138.515 -3.235 138.845 ;
        RECT -3.565 137.025 -3.235 137.355 ;
        RECT -3.565 135.355 -3.235 135.685 ;
        RECT -3.565 133.865 -3.235 134.195 ;
        RECT -3.565 132.455 -3.235 132.785 ;
        RECT -3.565 130.615 -3.235 130.945 ;
        RECT -3.565 129.125 -3.235 129.455 ;
        RECT -3.565 127.455 -3.235 127.785 ;
        RECT -3.565 125.965 -3.235 126.295 ;
        RECT -3.565 124.295 -3.235 124.625 ;
        RECT -3.565 122.805 -3.235 123.135 ;
        RECT -3.565 121.135 -3.235 121.465 ;
        RECT -3.565 119.645 -3.235 119.975 ;
        RECT -3.565 118.235 -3.235 118.565 ;
        RECT -3.565 116.395 -3.235 116.725 ;
        RECT -3.565 114.905 -3.235 115.235 ;
        RECT -3.565 113.235 -3.235 113.565 ;
        RECT -3.565 111.745 -3.235 112.075 ;
        RECT -3.565 110.075 -3.235 110.405 ;
        RECT -3.565 108.585 -3.235 108.915 ;
        RECT -3.565 106.915 -3.235 107.245 ;
        RECT -3.565 105.425 -3.235 105.755 ;
        RECT -3.565 104.015 -3.235 104.345 ;
        RECT -3.565 102.175 -3.235 102.505 ;
        RECT -3.565 100.685 -3.235 101.015 ;
        RECT -3.565 99.015 -3.235 99.345 ;
        RECT -3.565 97.525 -3.235 97.855 ;
        RECT -3.565 95.855 -3.235 96.185 ;
        RECT -3.565 94.365 -3.235 94.695 ;
        RECT -3.565 92.695 -3.235 93.025 ;
        RECT -3.565 91.205 -3.235 91.535 ;
        RECT -3.565 89.795 -3.235 90.125 ;
        RECT -3.565 87.955 -3.235 88.285 ;
        RECT -3.565 86.465 -3.235 86.795 ;
        RECT -3.565 84.795 -3.235 85.125 ;
        RECT -3.565 83.305 -3.235 83.635 ;
        RECT -3.565 81.635 -3.235 81.965 ;
        RECT -3.565 80.145 -3.235 80.475 ;
        RECT -3.565 78.475 -3.235 78.805 ;
        RECT -3.565 76.985 -3.235 77.315 ;
        RECT -3.565 75.575 -3.235 75.905 ;
        RECT -3.565 73.735 -3.235 74.065 ;
        RECT -3.565 72.245 -3.235 72.575 ;
        RECT -3.565 70.575 -3.235 70.905 ;
        RECT -3.565 69.085 -3.235 69.415 ;
        RECT -3.565 67.415 -3.235 67.745 ;
        RECT -3.565 65.925 -3.235 66.255 ;
        RECT -3.565 64.255 -3.235 64.585 ;
        RECT -3.565 62.765 -3.235 63.095 ;
        RECT -3.565 61.355 -3.235 61.685 ;
        RECT -3.565 59.515 -3.235 59.845 ;
        RECT -3.565 58.025 -3.235 58.355 ;
        RECT -3.565 56.355 -3.235 56.685 ;
        RECT -3.565 54.865 -3.235 55.195 ;
        RECT -3.565 53.195 -3.235 53.525 ;
        RECT -3.565 51.705 -3.235 52.035 ;
        RECT -3.565 50.035 -3.235 50.365 ;
        RECT -3.565 48.545 -3.235 48.875 ;
        RECT -3.565 47.135 -3.235 47.465 ;
        RECT -3.565 45.295 -3.235 45.625 ;
        RECT -3.565 43.805 -3.235 44.135 ;
        RECT -3.565 42.135 -3.235 42.465 ;
        RECT -3.565 40.645 -3.235 40.975 ;
        RECT -3.565 38.975 -3.235 39.305 ;
        RECT -3.565 37.485 -3.235 37.815 ;
        RECT -3.565 35.815 -3.235 36.145 ;
        RECT -3.565 34.325 -3.235 34.655 ;
        RECT -3.565 32.915 -3.235 33.245 ;
        RECT -3.565 31.075 -3.235 31.405 ;
        RECT -3.565 29.585 -3.235 29.915 ;
        RECT -3.565 27.915 -3.235 28.245 ;
        RECT -3.565 26.425 -3.235 26.755 ;
        RECT -3.565 24.755 -3.235 25.085 ;
        RECT -3.565 23.265 -3.235 23.595 ;
        RECT -3.565 21.595 -3.235 21.925 ;
        RECT -3.565 20.105 -3.235 20.435 ;
        RECT -3.565 18.695 -3.235 19.025 ;
        RECT -3.565 16.855 -3.235 17.185 ;
        RECT -3.565 15.365 -3.235 15.695 ;
        RECT -3.565 13.695 -3.235 14.025 ;
        RECT -3.565 12.205 -3.235 12.535 ;
        RECT -3.565 10.535 -3.235 10.865 ;
        RECT -3.565 9.045 -3.235 9.375 ;
        RECT -3.565 7.375 -3.235 7.705 ;
        RECT -3.565 5.885 -3.235 6.215 ;
        RECT -3.565 4.475 -3.235 4.805 ;
        RECT -3.565 2.115 -3.235 2.445 ;
        RECT -3.565 0.06 -3.235 0.39 ;
        RECT -3.565 -1.525 -3.235 -1.195 ;
        RECT -3.565 -2.885 -3.235 -2.555 ;
        RECT -3.565 -4.245 -3.235 -3.915 ;
        RECT -3.565 -5.605 -3.235 -5.275 ;
        RECT -3.565 -6.965 -3.235 -6.635 ;
        RECT -3.565 -8.325 -3.235 -7.995 ;
        RECT -3.565 -9.685 -3.235 -9.355 ;
        RECT -3.565 -12.405 -3.235 -12.075 ;
        RECT -3.565 -13.765 -3.235 -13.435 ;
        RECT -3.565 -15.125 -3.235 -14.795 ;
        RECT -3.565 -16.485 -3.235 -16.155 ;
        RECT -3.565 -17.845 -3.235 -17.515 ;
        RECT -3.565 -24.645 -3.235 -24.315 ;
        RECT -3.565 -26.005 -3.235 -25.675 ;
        RECT -3.565 -27.365 -3.235 -27.035 ;
        RECT -3.565 -28.725 -3.235 -28.395 ;
        RECT -3.565 -30.085 -3.235 -29.755 ;
        RECT -3.565 -31.445 -3.235 -31.115 ;
        RECT -3.565 -32.805 -3.235 -32.475 ;
        RECT -3.565 -34.165 -3.235 -33.835 ;
        RECT -3.565 -35.525 -3.235 -35.195 ;
        RECT -3.565 -36.885 -3.235 -36.555 ;
        RECT -3.565 -38.245 -3.235 -37.915 ;
        RECT -3.565 -39.605 -3.235 -39.275 ;
        RECT -3.565 -42.325 -3.235 -41.995 ;
        RECT -3.565 -45.045 -3.235 -44.715 ;
        RECT -3.565 -46.405 -3.235 -46.075 ;
        RECT -3.565 -47.765 -3.235 -47.435 ;
        RECT -3.565 -49.125 -3.235 -48.795 ;
        RECT -3.565 -51.845 -3.235 -51.515 ;
        RECT -3.565 -53.205 -3.235 -52.875 ;
        RECT -3.565 -54.565 -3.235 -54.235 ;
        RECT -3.565 -55.925 -3.235 -55.595 ;
        RECT -3.565 -57.285 -3.235 -56.955 ;
        RECT -3.565 -58.645 -3.235 -58.315 ;
        RECT -3.565 -60.005 -3.235 -59.675 ;
        RECT -3.565 -61.365 -3.235 -61.035 ;
        RECT -3.565 -62.725 -3.235 -62.395 ;
        RECT -3.565 -64.085 -3.235 -63.755 ;
        RECT -3.565 -65.445 -3.235 -65.115 ;
        RECT -3.565 -68.165 -3.235 -67.835 ;
        RECT -3.565 -69.525 -3.235 -69.195 ;
        RECT -3.565 -70.885 -3.235 -70.555 ;
        RECT -3.565 -72.245 -3.235 -71.915 ;
        RECT -3.565 -73.605 -3.235 -73.275 ;
        RECT -3.565 -74.965 -3.235 -74.635 ;
        RECT -3.565 -76.325 -3.235 -75.995 ;
        RECT -3.565 -77.685 -3.235 -77.355 ;
        RECT -3.565 -79.045 -3.235 -78.715 ;
        RECT -3.565 -80.405 -3.235 -80.075 ;
        RECT -3.565 -81.765 -3.235 -81.435 ;
        RECT -3.565 -83.125 -3.235 -82.795 ;
        RECT -3.565 -84.485 -3.235 -84.155 ;
        RECT -3.565 -85.845 -3.235 -85.515 ;
        RECT -3.565 -87.205 -3.235 -86.875 ;
        RECT -3.565 -88.565 -3.235 -88.235 ;
        RECT -3.565 -91.285 -3.235 -90.955 ;
        RECT -3.565 -92.645 -3.235 -92.315 ;
        RECT -3.565 -94.005 -3.235 -93.675 ;
        RECT -3.565 -95.365 -3.235 -95.035 ;
        RECT -3.565 -96.725 -3.235 -96.395 ;
        RECT -3.565 -98.085 -3.235 -97.755 ;
        RECT -3.565 -99.445 -3.235 -99.115 ;
        RECT -3.565 -100.805 -3.235 -100.475 ;
        RECT -3.565 -102.165 -3.235 -101.835 ;
        RECT -3.565 -103.525 -3.235 -103.195 ;
        RECT -3.565 -104.885 -3.235 -104.555 ;
        RECT -3.565 -106.245 -3.235 -105.915 ;
        RECT -3.565 -107.605 -3.235 -107.275 ;
        RECT -3.565 -108.965 -3.235 -108.635 ;
        RECT -3.565 -110.325 -3.235 -109.995 ;
        RECT -3.565 -111.685 -3.235 -111.355 ;
        RECT -3.565 -113.045 -3.235 -112.715 ;
        RECT -3.565 -114.405 -3.235 -114.075 ;
        RECT -3.565 -115.765 -3.235 -115.435 ;
        RECT -3.565 -117.125 -3.235 -116.795 ;
        RECT -3.565 -118.485 -3.235 -118.155 ;
        RECT -3.565 -119.845 -3.235 -119.515 ;
        RECT -3.565 -121.205 -3.235 -120.875 ;
        RECT -3.565 -122.565 -3.235 -122.235 ;
        RECT -3.565 -123.925 -3.235 -123.595 ;
        RECT -3.565 -125.285 -3.235 -124.955 ;
        RECT -3.565 -126.645 -3.235 -126.315 ;
        RECT -3.565 -128.005 -3.235 -127.675 ;
        RECT -3.565 -129.365 -3.235 -129.035 ;
        RECT -3.565 -130.725 -3.235 -130.395 ;
        RECT -3.565 -132.085 -3.235 -131.755 ;
        RECT -3.565 -133.445 -3.235 -133.115 ;
        RECT -3.565 -134.805 -3.235 -134.475 ;
        RECT -3.565 -136.165 -3.235 -135.835 ;
        RECT -3.565 -137.525 -3.235 -137.195 ;
        RECT -3.565 -138.885 -3.235 -138.555 ;
        RECT -3.565 -140.245 -3.235 -139.915 ;
        RECT -3.565 -141.605 -3.235 -141.275 ;
        RECT -3.565 -142.965 -3.235 -142.635 ;
        RECT -3.565 -144.325 -3.235 -143.995 ;
        RECT -3.565 -145.685 -3.235 -145.355 ;
        RECT -3.565 -147.045 -3.235 -146.715 ;
        RECT -3.565 -148.405 -3.235 -148.075 ;
        RECT -3.565 -149.765 -3.235 -149.435 ;
        RECT -3.565 -151.125 -3.235 -150.795 ;
        RECT -3.565 -152.485 -3.235 -152.155 ;
        RECT -3.565 -153.845 -3.235 -153.515 ;
        RECT -3.565 -155.205 -3.235 -154.875 ;
        RECT -3.565 -156.565 -3.235 -156.235 ;
        RECT -3.565 -157.925 -3.235 -157.595 ;
        RECT -3.565 -159.285 -3.235 -158.955 ;
        RECT -3.565 -160.645 -3.235 -160.315 ;
        RECT -3.565 -162.005 -3.235 -161.675 ;
        RECT -3.565 -163.365 -3.235 -163.035 ;
        RECT -3.565 -164.725 -3.235 -164.395 ;
        RECT -3.565 -166.085 -3.235 -165.755 ;
        RECT -3.565 -167.445 -3.235 -167.115 ;
        RECT -3.565 -168.805 -3.235 -168.475 ;
        RECT -3.565 -170.165 -3.235 -169.835 ;
        RECT -3.565 -171.525 -3.235 -171.195 ;
        RECT -3.565 -172.885 -3.235 -172.555 ;
        RECT -3.565 -174.245 -3.235 -173.915 ;
        RECT -3.565 -175.605 -3.235 -175.275 ;
        RECT -3.565 -176.965 -3.235 -176.635 ;
        RECT -3.565 -178.325 -3.235 -177.995 ;
        RECT -3.565 -179.685 -3.235 -179.355 ;
        RECT -3.565 -181.93 -3.235 -180.8 ;
        RECT -3.56 -182.045 -3.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.205 241.32 -1.875 242.45 ;
        RECT -2.205 239.195 -1.875 239.525 ;
        RECT -2.205 237.835 -1.875 238.165 ;
        RECT -2.205 235.975 -1.875 236.305 ;
        RECT -2.205 233.925 -1.875 234.255 ;
        RECT -2.205 231.995 -1.875 232.325 ;
        RECT -2.205 230.155 -1.875 230.485 ;
        RECT -2.205 228.665 -1.875 228.995 ;
        RECT -2.205 226.995 -1.875 227.325 ;
        RECT -2.205 225.505 -1.875 225.835 ;
        RECT -2.205 223.835 -1.875 224.165 ;
        RECT -2.205 222.345 -1.875 222.675 ;
        RECT -2.205 220.675 -1.875 221.005 ;
        RECT -2.205 219.185 -1.875 219.515 ;
        RECT -2.205 217.775 -1.875 218.105 ;
        RECT -2.205 215.935 -1.875 216.265 ;
        RECT -2.205 214.445 -1.875 214.775 ;
        RECT -2.205 212.775 -1.875 213.105 ;
        RECT -2.205 211.285 -1.875 211.615 ;
        RECT -2.205 209.615 -1.875 209.945 ;
        RECT -2.205 208.125 -1.875 208.455 ;
        RECT -2.205 206.455 -1.875 206.785 ;
        RECT -2.205 204.965 -1.875 205.295 ;
        RECT -2.205 203.555 -1.875 203.885 ;
        RECT -2.205 201.715 -1.875 202.045 ;
        RECT -2.205 200.225 -1.875 200.555 ;
        RECT -2.205 198.555 -1.875 198.885 ;
        RECT -2.205 197.065 -1.875 197.395 ;
        RECT -2.205 195.395 -1.875 195.725 ;
        RECT -2.205 193.905 -1.875 194.235 ;
        RECT -2.205 192.235 -1.875 192.565 ;
        RECT -2.205 190.745 -1.875 191.075 ;
        RECT -2.205 189.335 -1.875 189.665 ;
        RECT -2.205 187.495 -1.875 187.825 ;
        RECT -2.205 186.005 -1.875 186.335 ;
        RECT -2.205 184.335 -1.875 184.665 ;
        RECT -2.205 182.845 -1.875 183.175 ;
        RECT -2.205 181.175 -1.875 181.505 ;
        RECT -2.205 179.685 -1.875 180.015 ;
        RECT -2.205 178.015 -1.875 178.345 ;
        RECT -2.205 176.525 -1.875 176.855 ;
        RECT -2.205 175.115 -1.875 175.445 ;
        RECT -2.205 173.275 -1.875 173.605 ;
        RECT -2.205 171.785 -1.875 172.115 ;
        RECT -2.205 170.115 -1.875 170.445 ;
        RECT -2.205 168.625 -1.875 168.955 ;
        RECT -2.205 166.955 -1.875 167.285 ;
        RECT -2.205 165.465 -1.875 165.795 ;
        RECT -2.205 163.795 -1.875 164.125 ;
        RECT -2.205 162.305 -1.875 162.635 ;
        RECT -2.205 160.895 -1.875 161.225 ;
        RECT -2.205 159.055 -1.875 159.385 ;
        RECT -2.205 157.565 -1.875 157.895 ;
        RECT -2.205 155.895 -1.875 156.225 ;
        RECT -2.205 154.405 -1.875 154.735 ;
        RECT -2.205 152.735 -1.875 153.065 ;
        RECT -2.205 151.245 -1.875 151.575 ;
        RECT -2.205 149.575 -1.875 149.905 ;
        RECT -2.205 148.085 -1.875 148.415 ;
        RECT -2.205 146.675 -1.875 147.005 ;
        RECT -2.205 144.835 -1.875 145.165 ;
        RECT -2.205 143.345 -1.875 143.675 ;
        RECT -2.205 141.675 -1.875 142.005 ;
        RECT -2.205 140.185 -1.875 140.515 ;
        RECT -2.205 138.515 -1.875 138.845 ;
        RECT -2.205 137.025 -1.875 137.355 ;
        RECT -2.205 135.355 -1.875 135.685 ;
        RECT -2.205 133.865 -1.875 134.195 ;
        RECT -2.205 132.455 -1.875 132.785 ;
        RECT -2.205 130.615 -1.875 130.945 ;
        RECT -2.205 129.125 -1.875 129.455 ;
        RECT -2.205 127.455 -1.875 127.785 ;
        RECT -2.205 125.965 -1.875 126.295 ;
        RECT -2.205 124.295 -1.875 124.625 ;
        RECT -2.205 122.805 -1.875 123.135 ;
        RECT -2.205 121.135 -1.875 121.465 ;
        RECT -2.205 119.645 -1.875 119.975 ;
        RECT -2.205 118.235 -1.875 118.565 ;
        RECT -2.205 116.395 -1.875 116.725 ;
        RECT -2.205 114.905 -1.875 115.235 ;
        RECT -2.205 113.235 -1.875 113.565 ;
        RECT -2.205 111.745 -1.875 112.075 ;
        RECT -2.205 110.075 -1.875 110.405 ;
        RECT -2.205 108.585 -1.875 108.915 ;
        RECT -2.205 106.915 -1.875 107.245 ;
        RECT -2.205 105.425 -1.875 105.755 ;
        RECT -2.205 104.015 -1.875 104.345 ;
        RECT -2.205 102.175 -1.875 102.505 ;
        RECT -2.205 100.685 -1.875 101.015 ;
        RECT -2.205 99.015 -1.875 99.345 ;
        RECT -2.205 97.525 -1.875 97.855 ;
        RECT -2.205 95.855 -1.875 96.185 ;
        RECT -2.205 94.365 -1.875 94.695 ;
        RECT -2.205 92.695 -1.875 93.025 ;
        RECT -2.205 91.205 -1.875 91.535 ;
        RECT -2.205 89.795 -1.875 90.125 ;
        RECT -2.205 87.955 -1.875 88.285 ;
        RECT -2.205 86.465 -1.875 86.795 ;
        RECT -2.205 84.795 -1.875 85.125 ;
        RECT -2.205 83.305 -1.875 83.635 ;
        RECT -2.205 81.635 -1.875 81.965 ;
        RECT -2.205 80.145 -1.875 80.475 ;
        RECT -2.205 78.475 -1.875 78.805 ;
        RECT -2.205 76.985 -1.875 77.315 ;
        RECT -2.205 75.575 -1.875 75.905 ;
        RECT -2.205 73.735 -1.875 74.065 ;
        RECT -2.205 72.245 -1.875 72.575 ;
        RECT -2.205 70.575 -1.875 70.905 ;
        RECT -2.205 69.085 -1.875 69.415 ;
        RECT -2.205 67.415 -1.875 67.745 ;
        RECT -2.205 65.925 -1.875 66.255 ;
        RECT -2.205 64.255 -1.875 64.585 ;
        RECT -2.205 62.765 -1.875 63.095 ;
        RECT -2.205 61.355 -1.875 61.685 ;
        RECT -2.205 59.515 -1.875 59.845 ;
        RECT -2.205 58.025 -1.875 58.355 ;
        RECT -2.205 56.355 -1.875 56.685 ;
        RECT -2.205 54.865 -1.875 55.195 ;
        RECT -2.205 53.195 -1.875 53.525 ;
        RECT -2.205 51.705 -1.875 52.035 ;
        RECT -2.205 50.035 -1.875 50.365 ;
        RECT -2.205 48.545 -1.875 48.875 ;
        RECT -2.205 47.135 -1.875 47.465 ;
        RECT -2.205 45.295 -1.875 45.625 ;
        RECT -2.205 43.805 -1.875 44.135 ;
        RECT -2.205 42.135 -1.875 42.465 ;
        RECT -2.205 40.645 -1.875 40.975 ;
        RECT -2.205 38.975 -1.875 39.305 ;
        RECT -2.205 37.485 -1.875 37.815 ;
        RECT -2.205 35.815 -1.875 36.145 ;
        RECT -2.205 34.325 -1.875 34.655 ;
        RECT -2.205 32.915 -1.875 33.245 ;
        RECT -2.205 31.075 -1.875 31.405 ;
        RECT -2.205 29.585 -1.875 29.915 ;
        RECT -2.205 27.915 -1.875 28.245 ;
        RECT -2.205 26.425 -1.875 26.755 ;
        RECT -2.205 24.755 -1.875 25.085 ;
        RECT -2.205 23.265 -1.875 23.595 ;
        RECT -2.205 21.595 -1.875 21.925 ;
        RECT -2.205 20.105 -1.875 20.435 ;
        RECT -2.205 18.695 -1.875 19.025 ;
        RECT -2.205 16.855 -1.875 17.185 ;
        RECT -2.205 15.365 -1.875 15.695 ;
        RECT -2.205 13.695 -1.875 14.025 ;
        RECT -2.205 12.205 -1.875 12.535 ;
        RECT -2.205 10.535 -1.875 10.865 ;
        RECT -2.205 9.045 -1.875 9.375 ;
        RECT -2.205 7.375 -1.875 7.705 ;
        RECT -2.205 5.885 -1.875 6.215 ;
        RECT -2.205 4.475 -1.875 4.805 ;
        RECT -2.205 2.115 -1.875 2.445 ;
        RECT -2.205 0.06 -1.875 0.39 ;
        RECT -2.205 -1.525 -1.875 -1.195 ;
        RECT -2.205 -2.885 -1.875 -2.555 ;
        RECT -2.205 -4.245 -1.875 -3.915 ;
        RECT -2.205 -5.605 -1.875 -5.275 ;
        RECT -2.205 -6.965 -1.875 -6.635 ;
        RECT -2.205 -8.325 -1.875 -7.995 ;
        RECT -2.205 -9.685 -1.875 -9.355 ;
        RECT -2.205 -12.405 -1.875 -12.075 ;
        RECT -2.205 -13.765 -1.875 -13.435 ;
        RECT -2.205 -15.125 -1.875 -14.795 ;
        RECT -2.205 -16.485 -1.875 -16.155 ;
        RECT -2.205 -17.845 -1.875 -17.515 ;
        RECT -2.205 -24.645 -1.875 -24.315 ;
        RECT -2.205 -26.005 -1.875 -25.675 ;
        RECT -2.205 -27.365 -1.875 -27.035 ;
        RECT -2.205 -28.725 -1.875 -28.395 ;
        RECT -2.205 -30.085 -1.875 -29.755 ;
        RECT -2.205 -31.445 -1.875 -31.115 ;
        RECT -2.205 -32.805 -1.875 -32.475 ;
        RECT -2.205 -34.165 -1.875 -33.835 ;
        RECT -2.205 -35.525 -1.875 -35.195 ;
        RECT -2.205 -36.885 -1.875 -36.555 ;
        RECT -2.205 -38.245 -1.875 -37.915 ;
        RECT -2.205 -39.605 -1.875 -39.275 ;
        RECT -2.205 -42.325 -1.875 -41.995 ;
        RECT -2.205 -45.045 -1.875 -44.715 ;
        RECT -2.205 -46.405 -1.875 -46.075 ;
        RECT -2.205 -47.765 -1.875 -47.435 ;
        RECT -2.205 -49.125 -1.875 -48.795 ;
        RECT -2.205 -51.845 -1.875 -51.515 ;
        RECT -2.205 -53.205 -1.875 -52.875 ;
        RECT -2.205 -54.565 -1.875 -54.235 ;
        RECT -2.205 -55.925 -1.875 -55.595 ;
        RECT -2.205 -57.285 -1.875 -56.955 ;
        RECT -2.205 -58.645 -1.875 -58.315 ;
        RECT -2.205 -60.005 -1.875 -59.675 ;
        RECT -2.205 -61.365 -1.875 -61.035 ;
        RECT -2.205 -62.725 -1.875 -62.395 ;
        RECT -2.205 -64.085 -1.875 -63.755 ;
        RECT -2.205 -65.445 -1.875 -65.115 ;
        RECT -2.205 -68.165 -1.875 -67.835 ;
        RECT -2.205 -69.525 -1.875 -69.195 ;
        RECT -2.205 -70.885 -1.875 -70.555 ;
        RECT -2.205 -72.245 -1.875 -71.915 ;
        RECT -2.205 -73.605 -1.875 -73.275 ;
        RECT -2.205 -74.965 -1.875 -74.635 ;
        RECT -2.205 -76.325 -1.875 -75.995 ;
        RECT -2.205 -77.685 -1.875 -77.355 ;
        RECT -2.205 -79.045 -1.875 -78.715 ;
        RECT -2.205 -80.405 -1.875 -80.075 ;
        RECT -2.205 -81.765 -1.875 -81.435 ;
        RECT -2.205 -83.125 -1.875 -82.795 ;
        RECT -2.205 -84.485 -1.875 -84.155 ;
        RECT -2.205 -85.845 -1.875 -85.515 ;
        RECT -2.205 -87.205 -1.875 -86.875 ;
        RECT -2.205 -88.565 -1.875 -88.235 ;
        RECT -2.205 -91.285 -1.875 -90.955 ;
        RECT -2.205 -92.645 -1.875 -92.315 ;
        RECT -2.205 -94.005 -1.875 -93.675 ;
        RECT -2.205 -95.365 -1.875 -95.035 ;
        RECT -2.205 -96.725 -1.875 -96.395 ;
        RECT -2.205 -98.085 -1.875 -97.755 ;
        RECT -2.205 -99.445 -1.875 -99.115 ;
        RECT -2.205 -100.805 -1.875 -100.475 ;
        RECT -2.205 -102.165 -1.875 -101.835 ;
        RECT -2.205 -103.525 -1.875 -103.195 ;
        RECT -2.205 -104.885 -1.875 -104.555 ;
        RECT -2.205 -106.245 -1.875 -105.915 ;
        RECT -2.205 -107.605 -1.875 -107.275 ;
        RECT -2.205 -108.965 -1.875 -108.635 ;
        RECT -2.205 -110.325 -1.875 -109.995 ;
        RECT -2.205 -111.685 -1.875 -111.355 ;
        RECT -2.205 -113.045 -1.875 -112.715 ;
        RECT -2.205 -114.405 -1.875 -114.075 ;
        RECT -2.205 -115.765 -1.875 -115.435 ;
        RECT -2.205 -117.125 -1.875 -116.795 ;
        RECT -2.205 -118.485 -1.875 -118.155 ;
        RECT -2.205 -119.845 -1.875 -119.515 ;
        RECT -2.205 -121.205 -1.875 -120.875 ;
        RECT -2.205 -122.565 -1.875 -122.235 ;
        RECT -2.205 -123.925 -1.875 -123.595 ;
        RECT -2.205 -125.285 -1.875 -124.955 ;
        RECT -2.205 -126.645 -1.875 -126.315 ;
        RECT -2.205 -128.005 -1.875 -127.675 ;
        RECT -2.205 -129.365 -1.875 -129.035 ;
        RECT -2.205 -130.725 -1.875 -130.395 ;
        RECT -2.205 -132.085 -1.875 -131.755 ;
        RECT -2.205 -133.445 -1.875 -133.115 ;
        RECT -2.205 -134.805 -1.875 -134.475 ;
        RECT -2.205 -136.165 -1.875 -135.835 ;
        RECT -2.205 -137.525 -1.875 -137.195 ;
        RECT -2.205 -138.885 -1.875 -138.555 ;
        RECT -2.205 -140.245 -1.875 -139.915 ;
        RECT -2.205 -141.605 -1.875 -141.275 ;
        RECT -2.205 -142.965 -1.875 -142.635 ;
        RECT -2.205 -144.325 -1.875 -143.995 ;
        RECT -2.205 -145.685 -1.875 -145.355 ;
        RECT -2.205 -147.045 -1.875 -146.715 ;
        RECT -2.205 -148.405 -1.875 -148.075 ;
        RECT -2.205 -149.765 -1.875 -149.435 ;
        RECT -2.205 -151.125 -1.875 -150.795 ;
        RECT -2.205 -152.485 -1.875 -152.155 ;
        RECT -2.205 -153.845 -1.875 -153.515 ;
        RECT -2.205 -155.205 -1.875 -154.875 ;
        RECT -2.205 -156.565 -1.875 -156.235 ;
        RECT -2.205 -157.925 -1.875 -157.595 ;
        RECT -2.205 -159.285 -1.875 -158.955 ;
        RECT -2.205 -160.645 -1.875 -160.315 ;
        RECT -2.205 -162.005 -1.875 -161.675 ;
        RECT -2.205 -163.365 -1.875 -163.035 ;
        RECT -2.205 -164.725 -1.875 -164.395 ;
        RECT -2.205 -166.085 -1.875 -165.755 ;
        RECT -2.205 -167.445 -1.875 -167.115 ;
        RECT -2.205 -168.805 -1.875 -168.475 ;
        RECT -2.205 -170.165 -1.875 -169.835 ;
        RECT -2.205 -171.525 -1.875 -171.195 ;
        RECT -2.205 -172.885 -1.875 -172.555 ;
        RECT -2.205 -174.245 -1.875 -173.915 ;
        RECT -2.205 -175.605 -1.875 -175.275 ;
        RECT -2.205 -176.965 -1.875 -176.635 ;
        RECT -2.205 -178.325 -1.875 -177.995 ;
        RECT -2.205 -179.685 -1.875 -179.355 ;
        RECT -2.205 -181.93 -1.875 -180.8 ;
        RECT -2.2 -182.045 -1.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -0.845 -28.725 -0.515 -28.395 ;
        RECT -0.845 -30.085 -0.515 -29.755 ;
        RECT -0.845 -31.445 -0.515 -31.115 ;
        RECT -0.845 -32.805 -0.515 -32.475 ;
        RECT -0.845 -34.165 -0.515 -33.835 ;
        RECT -0.84 -36.2 -0.52 242.565 ;
        RECT -0.845 241.32 -0.515 242.45 ;
        RECT -0.845 239.195 -0.515 239.525 ;
        RECT -0.845 237.835 -0.515 238.165 ;
        RECT -0.845 235.975 -0.515 236.305 ;
        RECT -0.845 233.925 -0.515 234.255 ;
        RECT -0.845 231.995 -0.515 232.325 ;
        RECT -0.845 230.155 -0.515 230.485 ;
        RECT -0.845 228.665 -0.515 228.995 ;
        RECT -0.845 226.995 -0.515 227.325 ;
        RECT -0.845 225.505 -0.515 225.835 ;
        RECT -0.845 223.835 -0.515 224.165 ;
        RECT -0.845 222.345 -0.515 222.675 ;
        RECT -0.845 220.675 -0.515 221.005 ;
        RECT -0.845 219.185 -0.515 219.515 ;
        RECT -0.845 217.775 -0.515 218.105 ;
        RECT -0.845 215.935 -0.515 216.265 ;
        RECT -0.845 214.445 -0.515 214.775 ;
        RECT -0.845 212.775 -0.515 213.105 ;
        RECT -0.845 211.285 -0.515 211.615 ;
        RECT -0.845 209.615 -0.515 209.945 ;
        RECT -0.845 208.125 -0.515 208.455 ;
        RECT -0.845 206.455 -0.515 206.785 ;
        RECT -0.845 204.965 -0.515 205.295 ;
        RECT -0.845 203.555 -0.515 203.885 ;
        RECT -0.845 201.715 -0.515 202.045 ;
        RECT -0.845 200.225 -0.515 200.555 ;
        RECT -0.845 198.555 -0.515 198.885 ;
        RECT -0.845 197.065 -0.515 197.395 ;
        RECT -0.845 195.395 -0.515 195.725 ;
        RECT -0.845 193.905 -0.515 194.235 ;
        RECT -0.845 192.235 -0.515 192.565 ;
        RECT -0.845 190.745 -0.515 191.075 ;
        RECT -0.845 189.335 -0.515 189.665 ;
        RECT -0.845 187.495 -0.515 187.825 ;
        RECT -0.845 186.005 -0.515 186.335 ;
        RECT -0.845 184.335 -0.515 184.665 ;
        RECT -0.845 182.845 -0.515 183.175 ;
        RECT -0.845 181.175 -0.515 181.505 ;
        RECT -0.845 179.685 -0.515 180.015 ;
        RECT -0.845 178.015 -0.515 178.345 ;
        RECT -0.845 176.525 -0.515 176.855 ;
        RECT -0.845 175.115 -0.515 175.445 ;
        RECT -0.845 173.275 -0.515 173.605 ;
        RECT -0.845 171.785 -0.515 172.115 ;
        RECT -0.845 170.115 -0.515 170.445 ;
        RECT -0.845 168.625 -0.515 168.955 ;
        RECT -0.845 166.955 -0.515 167.285 ;
        RECT -0.845 165.465 -0.515 165.795 ;
        RECT -0.845 163.795 -0.515 164.125 ;
        RECT -0.845 162.305 -0.515 162.635 ;
        RECT -0.845 160.895 -0.515 161.225 ;
        RECT -0.845 159.055 -0.515 159.385 ;
        RECT -0.845 157.565 -0.515 157.895 ;
        RECT -0.845 155.895 -0.515 156.225 ;
        RECT -0.845 154.405 -0.515 154.735 ;
        RECT -0.845 152.735 -0.515 153.065 ;
        RECT -0.845 151.245 -0.515 151.575 ;
        RECT -0.845 149.575 -0.515 149.905 ;
        RECT -0.845 148.085 -0.515 148.415 ;
        RECT -0.845 146.675 -0.515 147.005 ;
        RECT -0.845 144.835 -0.515 145.165 ;
        RECT -0.845 143.345 -0.515 143.675 ;
        RECT -0.845 141.675 -0.515 142.005 ;
        RECT -0.845 140.185 -0.515 140.515 ;
        RECT -0.845 138.515 -0.515 138.845 ;
        RECT -0.845 137.025 -0.515 137.355 ;
        RECT -0.845 135.355 -0.515 135.685 ;
        RECT -0.845 133.865 -0.515 134.195 ;
        RECT -0.845 132.455 -0.515 132.785 ;
        RECT -0.845 130.615 -0.515 130.945 ;
        RECT -0.845 129.125 -0.515 129.455 ;
        RECT -0.845 127.455 -0.515 127.785 ;
        RECT -0.845 125.965 -0.515 126.295 ;
        RECT -0.845 124.295 -0.515 124.625 ;
        RECT -0.845 122.805 -0.515 123.135 ;
        RECT -0.845 121.135 -0.515 121.465 ;
        RECT -0.845 119.645 -0.515 119.975 ;
        RECT -0.845 118.235 -0.515 118.565 ;
        RECT -0.845 116.395 -0.515 116.725 ;
        RECT -0.845 114.905 -0.515 115.235 ;
        RECT -0.845 113.235 -0.515 113.565 ;
        RECT -0.845 111.745 -0.515 112.075 ;
        RECT -0.845 110.075 -0.515 110.405 ;
        RECT -0.845 108.585 -0.515 108.915 ;
        RECT -0.845 106.915 -0.515 107.245 ;
        RECT -0.845 105.425 -0.515 105.755 ;
        RECT -0.845 104.015 -0.515 104.345 ;
        RECT -0.845 102.175 -0.515 102.505 ;
        RECT -0.845 100.685 -0.515 101.015 ;
        RECT -0.845 99.015 -0.515 99.345 ;
        RECT -0.845 97.525 -0.515 97.855 ;
        RECT -0.845 95.855 -0.515 96.185 ;
        RECT -0.845 94.365 -0.515 94.695 ;
        RECT -0.845 92.695 -0.515 93.025 ;
        RECT -0.845 91.205 -0.515 91.535 ;
        RECT -0.845 89.795 -0.515 90.125 ;
        RECT -0.845 87.955 -0.515 88.285 ;
        RECT -0.845 86.465 -0.515 86.795 ;
        RECT -0.845 84.795 -0.515 85.125 ;
        RECT -0.845 83.305 -0.515 83.635 ;
        RECT -0.845 81.635 -0.515 81.965 ;
        RECT -0.845 80.145 -0.515 80.475 ;
        RECT -0.845 78.475 -0.515 78.805 ;
        RECT -0.845 76.985 -0.515 77.315 ;
        RECT -0.845 75.575 -0.515 75.905 ;
        RECT -0.845 73.735 -0.515 74.065 ;
        RECT -0.845 72.245 -0.515 72.575 ;
        RECT -0.845 70.575 -0.515 70.905 ;
        RECT -0.845 69.085 -0.515 69.415 ;
        RECT -0.845 67.415 -0.515 67.745 ;
        RECT -0.845 65.925 -0.515 66.255 ;
        RECT -0.845 64.255 -0.515 64.585 ;
        RECT -0.845 62.765 -0.515 63.095 ;
        RECT -0.845 61.355 -0.515 61.685 ;
        RECT -0.845 59.515 -0.515 59.845 ;
        RECT -0.845 58.025 -0.515 58.355 ;
        RECT -0.845 56.355 -0.515 56.685 ;
        RECT -0.845 54.865 -0.515 55.195 ;
        RECT -0.845 53.195 -0.515 53.525 ;
        RECT -0.845 51.705 -0.515 52.035 ;
        RECT -0.845 50.035 -0.515 50.365 ;
        RECT -0.845 48.545 -0.515 48.875 ;
        RECT -0.845 47.135 -0.515 47.465 ;
        RECT -0.845 45.295 -0.515 45.625 ;
        RECT -0.845 43.805 -0.515 44.135 ;
        RECT -0.845 42.135 -0.515 42.465 ;
        RECT -0.845 40.645 -0.515 40.975 ;
        RECT -0.845 38.975 -0.515 39.305 ;
        RECT -0.845 37.485 -0.515 37.815 ;
        RECT -0.845 35.815 -0.515 36.145 ;
        RECT -0.845 34.325 -0.515 34.655 ;
        RECT -0.845 32.915 -0.515 33.245 ;
        RECT -0.845 31.075 -0.515 31.405 ;
        RECT -0.845 29.585 -0.515 29.915 ;
        RECT -0.845 27.915 -0.515 28.245 ;
        RECT -0.845 26.425 -0.515 26.755 ;
        RECT -0.845 24.755 -0.515 25.085 ;
        RECT -0.845 23.265 -0.515 23.595 ;
        RECT -0.845 21.595 -0.515 21.925 ;
        RECT -0.845 20.105 -0.515 20.435 ;
        RECT -0.845 18.695 -0.515 19.025 ;
        RECT -0.845 16.855 -0.515 17.185 ;
        RECT -0.845 15.365 -0.515 15.695 ;
        RECT -0.845 13.695 -0.515 14.025 ;
        RECT -0.845 12.205 -0.515 12.535 ;
        RECT -0.845 10.535 -0.515 10.865 ;
        RECT -0.845 9.045 -0.515 9.375 ;
        RECT -0.845 7.375 -0.515 7.705 ;
        RECT -0.845 5.885 -0.515 6.215 ;
        RECT -0.845 4.475 -0.515 4.805 ;
        RECT -0.845 2.115 -0.515 2.445 ;
        RECT -0.845 0.06 -0.515 0.39 ;
        RECT -0.845 -1.525 -0.515 -1.195 ;
        RECT -0.845 -2.885 -0.515 -2.555 ;
        RECT -0.845 -4.245 -0.515 -3.915 ;
        RECT -0.845 -5.605 -0.515 -5.275 ;
        RECT -0.845 -6.965 -0.515 -6.635 ;
        RECT -0.845 -8.325 -0.515 -7.995 ;
        RECT -0.845 -9.685 -0.515 -9.355 ;
        RECT -0.845 -12.405 -0.515 -12.075 ;
        RECT -0.845 -13.765 -0.515 -13.435 ;
        RECT -0.845 -15.125 -0.515 -14.795 ;
        RECT -0.845 -16.485 -0.515 -16.155 ;
        RECT -0.845 -24.645 -0.515 -24.315 ;
        RECT -0.845 -26.005 -0.515 -25.675 ;
        RECT -0.845 -27.365 -0.515 -27.035 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 -160.645 -14.115 -160.315 ;
        RECT -14.445 -162.005 -14.115 -161.675 ;
        RECT -14.445 -163.365 -14.115 -163.035 ;
        RECT -14.445 -164.725 -14.115 -164.395 ;
        RECT -14.445 -166.085 -14.115 -165.755 ;
        RECT -14.445 -167.445 -14.115 -167.115 ;
        RECT -14.44 -167.445 -14.12 -159.64 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 -174.245 -14.115 -173.915 ;
        RECT -14.445 -175.605 -14.115 -175.275 ;
        RECT -14.445 -176.685 -14.115 -176.355 ;
        RECT -14.445 -178.325 -14.115 -177.995 ;
        RECT -14.445 -179.685 -14.115 -179.355 ;
        RECT -14.445 -181.93 -14.115 -180.8 ;
        RECT -14.44 -182.045 -14.12 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -13.085 241.32 -12.755 242.45 ;
        RECT -13.085 239.195 -12.755 239.525 ;
        RECT -13.085 237.835 -12.755 238.165 ;
        RECT -13.085 236.475 -12.755 236.805 ;
        RECT -13.085 235.115 -12.755 235.445 ;
        RECT -13.085 233.755 -12.755 234.085 ;
        RECT -13.085 232.395 -12.755 232.725 ;
        RECT -13.085 231.035 -12.755 231.365 ;
        RECT -13.085 229.675 -12.755 230.005 ;
        RECT -13.085 228.315 -12.755 228.645 ;
        RECT -13.085 226.955 -12.755 227.285 ;
        RECT -13.085 225.595 -12.755 225.925 ;
        RECT -13.085 224.235 -12.755 224.565 ;
        RECT -13.085 222.875 -12.755 223.205 ;
        RECT -13.085 221.515 -12.755 221.845 ;
        RECT -13.085 220.155 -12.755 220.485 ;
        RECT -13.085 218.795 -12.755 219.125 ;
        RECT -13.085 217.435 -12.755 217.765 ;
        RECT -13.085 216.075 -12.755 216.405 ;
        RECT -13.085 214.715 -12.755 215.045 ;
        RECT -13.085 213.355 -12.755 213.685 ;
        RECT -13.085 211.995 -12.755 212.325 ;
        RECT -13.085 210.635 -12.755 210.965 ;
        RECT -13.085 209.275 -12.755 209.605 ;
        RECT -13.085 207.915 -12.755 208.245 ;
        RECT -13.085 206.555 -12.755 206.885 ;
        RECT -13.085 205.195 -12.755 205.525 ;
        RECT -13.085 203.835 -12.755 204.165 ;
        RECT -13.085 202.475 -12.755 202.805 ;
        RECT -13.085 201.115 -12.755 201.445 ;
        RECT -13.085 199.755 -12.755 200.085 ;
        RECT -13.085 198.395 -12.755 198.725 ;
        RECT -13.085 197.035 -12.755 197.365 ;
        RECT -13.085 195.675 -12.755 196.005 ;
        RECT -13.085 194.315 -12.755 194.645 ;
        RECT -13.085 192.955 -12.755 193.285 ;
        RECT -13.085 191.595 -12.755 191.925 ;
        RECT -13.085 190.235 -12.755 190.565 ;
        RECT -13.085 188.875 -12.755 189.205 ;
        RECT -13.085 187.515 -12.755 187.845 ;
        RECT -13.085 186.155 -12.755 186.485 ;
        RECT -13.085 184.795 -12.755 185.125 ;
        RECT -13.085 183.435 -12.755 183.765 ;
        RECT -13.085 182.075 -12.755 182.405 ;
        RECT -13.085 180.715 -12.755 181.045 ;
        RECT -13.085 179.355 -12.755 179.685 ;
        RECT -13.085 177.995 -12.755 178.325 ;
        RECT -13.085 176.635 -12.755 176.965 ;
        RECT -13.085 175.275 -12.755 175.605 ;
        RECT -13.085 173.915 -12.755 174.245 ;
        RECT -13.085 172.555 -12.755 172.885 ;
        RECT -13.085 171.195 -12.755 171.525 ;
        RECT -13.085 169.835 -12.755 170.165 ;
        RECT -13.085 168.475 -12.755 168.805 ;
        RECT -13.085 167.115 -12.755 167.445 ;
        RECT -13.085 165.755 -12.755 166.085 ;
        RECT -13.085 164.395 -12.755 164.725 ;
        RECT -13.085 163.035 -12.755 163.365 ;
        RECT -13.085 161.675 -12.755 162.005 ;
        RECT -13.085 160.315 -12.755 160.645 ;
        RECT -13.085 158.955 -12.755 159.285 ;
        RECT -13.085 157.595 -12.755 157.925 ;
        RECT -13.085 156.235 -12.755 156.565 ;
        RECT -13.085 154.875 -12.755 155.205 ;
        RECT -13.085 153.515 -12.755 153.845 ;
        RECT -13.085 152.155 -12.755 152.485 ;
        RECT -13.085 150.795 -12.755 151.125 ;
        RECT -13.085 149.435 -12.755 149.765 ;
        RECT -13.085 148.075 -12.755 148.405 ;
        RECT -13.085 146.715 -12.755 147.045 ;
        RECT -13.085 145.355 -12.755 145.685 ;
        RECT -13.085 143.995 -12.755 144.325 ;
        RECT -13.085 142.635 -12.755 142.965 ;
        RECT -13.085 141.275 -12.755 141.605 ;
        RECT -13.085 139.915 -12.755 140.245 ;
        RECT -13.085 138.555 -12.755 138.885 ;
        RECT -13.085 137.195 -12.755 137.525 ;
        RECT -13.085 135.835 -12.755 136.165 ;
        RECT -13.085 134.475 -12.755 134.805 ;
        RECT -13.085 133.115 -12.755 133.445 ;
        RECT -13.085 131.755 -12.755 132.085 ;
        RECT -13.085 130.395 -12.755 130.725 ;
        RECT -13.085 129.035 -12.755 129.365 ;
        RECT -13.085 127.675 -12.755 128.005 ;
        RECT -13.085 126.315 -12.755 126.645 ;
        RECT -13.085 124.955 -12.755 125.285 ;
        RECT -13.085 123.595 -12.755 123.925 ;
        RECT -13.085 122.235 -12.755 122.565 ;
        RECT -13.085 120.875 -12.755 121.205 ;
        RECT -13.085 119.515 -12.755 119.845 ;
        RECT -13.085 118.155 -12.755 118.485 ;
        RECT -13.085 116.795 -12.755 117.125 ;
        RECT -13.085 115.435 -12.755 115.765 ;
        RECT -13.085 114.075 -12.755 114.405 ;
        RECT -13.085 112.715 -12.755 113.045 ;
        RECT -13.085 111.355 -12.755 111.685 ;
        RECT -13.085 109.995 -12.755 110.325 ;
        RECT -13.085 108.635 -12.755 108.965 ;
        RECT -13.085 107.275 -12.755 107.605 ;
        RECT -13.085 105.915 -12.755 106.245 ;
        RECT -13.085 104.555 -12.755 104.885 ;
        RECT -13.085 103.195 -12.755 103.525 ;
        RECT -13.085 101.835 -12.755 102.165 ;
        RECT -13.085 100.475 -12.755 100.805 ;
        RECT -13.085 99.115 -12.755 99.445 ;
        RECT -13.085 97.755 -12.755 98.085 ;
        RECT -13.085 96.395 -12.755 96.725 ;
        RECT -13.085 95.035 -12.755 95.365 ;
        RECT -13.085 93.675 -12.755 94.005 ;
        RECT -13.085 92.315 -12.755 92.645 ;
        RECT -13.085 90.955 -12.755 91.285 ;
        RECT -13.085 89.595 -12.755 89.925 ;
        RECT -13.085 88.235 -12.755 88.565 ;
        RECT -13.085 86.875 -12.755 87.205 ;
        RECT -13.085 85.515 -12.755 85.845 ;
        RECT -13.085 84.155 -12.755 84.485 ;
        RECT -13.085 82.795 -12.755 83.125 ;
        RECT -13.085 81.435 -12.755 81.765 ;
        RECT -13.085 80.075 -12.755 80.405 ;
        RECT -13.085 78.715 -12.755 79.045 ;
        RECT -13.085 77.355 -12.755 77.685 ;
        RECT -13.085 75.995 -12.755 76.325 ;
        RECT -13.085 74.635 -12.755 74.965 ;
        RECT -13.085 73.275 -12.755 73.605 ;
        RECT -13.085 71.915 -12.755 72.245 ;
        RECT -13.085 70.555 -12.755 70.885 ;
        RECT -13.085 69.195 -12.755 69.525 ;
        RECT -13.085 67.835 -12.755 68.165 ;
        RECT -13.085 66.475 -12.755 66.805 ;
        RECT -13.085 65.115 -12.755 65.445 ;
        RECT -13.085 63.755 -12.755 64.085 ;
        RECT -13.085 62.395 -12.755 62.725 ;
        RECT -13.085 61.035 -12.755 61.365 ;
        RECT -13.085 59.675 -12.755 60.005 ;
        RECT -13.085 58.315 -12.755 58.645 ;
        RECT -13.085 56.955 -12.755 57.285 ;
        RECT -13.085 55.595 -12.755 55.925 ;
        RECT -13.085 54.235 -12.755 54.565 ;
        RECT -13.085 52.875 -12.755 53.205 ;
        RECT -13.085 51.515 -12.755 51.845 ;
        RECT -13.085 50.155 -12.755 50.485 ;
        RECT -13.085 48.795 -12.755 49.125 ;
        RECT -13.085 47.435 -12.755 47.765 ;
        RECT -13.085 46.075 -12.755 46.405 ;
        RECT -13.085 44.715 -12.755 45.045 ;
        RECT -13.085 43.355 -12.755 43.685 ;
        RECT -13.085 41.995 -12.755 42.325 ;
        RECT -13.085 40.635 -12.755 40.965 ;
        RECT -13.085 39.275 -12.755 39.605 ;
        RECT -13.085 37.915 -12.755 38.245 ;
        RECT -13.085 36.555 -12.755 36.885 ;
        RECT -13.085 35.195 -12.755 35.525 ;
        RECT -13.085 33.835 -12.755 34.165 ;
        RECT -13.085 32.475 -12.755 32.805 ;
        RECT -13.085 31.115 -12.755 31.445 ;
        RECT -13.085 29.755 -12.755 30.085 ;
        RECT -13.085 28.395 -12.755 28.725 ;
        RECT -13.085 27.035 -12.755 27.365 ;
        RECT -13.085 25.675 -12.755 26.005 ;
        RECT -13.085 24.315 -12.755 24.645 ;
        RECT -13.085 22.955 -12.755 23.285 ;
        RECT -13.085 21.595 -12.755 21.925 ;
        RECT -13.085 20.235 -12.755 20.565 ;
        RECT -13.085 18.875 -12.755 19.205 ;
        RECT -13.085 17.515 -12.755 17.845 ;
        RECT -13.085 16.155 -12.755 16.485 ;
        RECT -13.085 14.795 -12.755 15.125 ;
        RECT -13.085 13.435 -12.755 13.765 ;
        RECT -13.085 12.075 -12.755 12.405 ;
        RECT -13.085 10.715 -12.755 11.045 ;
        RECT -13.085 9.355 -12.755 9.685 ;
        RECT -13.085 7.995 -12.755 8.325 ;
        RECT -13.085 6.635 -12.755 6.965 ;
        RECT -13.085 5.275 -12.755 5.605 ;
        RECT -13.085 3.915 -12.755 4.245 ;
        RECT -13.085 2.555 -12.755 2.885 ;
        RECT -13.085 1.195 -12.755 1.525 ;
        RECT -13.085 -0.165 -12.755 0.165 ;
        RECT -13.085 -2.885 -12.755 -2.555 ;
        RECT -13.085 -4.245 -12.755 -3.915 ;
        RECT -13.085 -5.605 -12.755 -5.275 ;
        RECT -13.085 -8.325 -12.755 -7.995 ;
        RECT -13.085 -9.685 -12.755 -9.355 ;
        RECT -13.085 -12.405 -12.755 -12.075 ;
        RECT -13.085 -13.765 -12.755 -13.435 ;
        RECT -13.085 -14.95 -12.755 -14.62 ;
        RECT -13.085 -17.845 -12.755 -17.515 ;
        RECT -13.085 -19.79 -12.755 -19.46 ;
        RECT -13.085 -27.365 -12.755 -27.035 ;
        RECT -13.085 -28.725 -12.755 -28.395 ;
        RECT -13.085 -30.085 -12.755 -29.755 ;
        RECT -13.085 -31.445 -12.755 -31.115 ;
        RECT -13.085 -32.805 -12.755 -32.475 ;
        RECT -13.085 -35.525 -12.755 -35.195 ;
        RECT -13.085 -36.885 -12.755 -36.555 ;
        RECT -13.085 -37.93 -12.755 -37.6 ;
        RECT -13.085 -42.77 -12.755 -42.44 ;
        RECT -13.085 -51.845 -12.755 -51.515 ;
        RECT -13.085 -53.205 -12.755 -52.875 ;
        RECT -13.085 -54.565 -12.755 -54.235 ;
        RECT -13.085 -55.925 -12.755 -55.595 ;
        RECT -13.085 -57.285 -12.755 -56.955 ;
        RECT -13.085 -58.645 -12.755 -58.315 ;
        RECT -13.085 -60.005 -12.755 -59.675 ;
        RECT -13.085 -61.365 -12.755 -61.035 ;
        RECT -13.085 -62.725 -12.755 -62.395 ;
        RECT -13.085 -64.085 -12.755 -63.755 ;
        RECT -13.085 -65.445 -12.755 -65.115 ;
        RECT -13.085 -68.165 -12.755 -67.835 ;
        RECT -13.085 -69.525 -12.755 -69.195 ;
        RECT -13.085 -70.885 -12.755 -70.555 ;
        RECT -13.085 -72.245 -12.755 -71.915 ;
        RECT -13.085 -74.965 -12.755 -74.635 ;
        RECT -13.085 -76.71 -12.755 -76.38 ;
        RECT -13.085 -77.685 -12.755 -77.355 ;
        RECT -13.085 -79.045 -12.755 -78.715 ;
        RECT -13.085 -81.765 -12.755 -81.435 ;
        RECT -13.085 -83.125 -12.755 -82.795 ;
        RECT -13.085 -84.485 -12.755 -84.155 ;
        RECT -13.085 -85.25 -12.755 -84.92 ;
        RECT -13.085 -87.205 -12.755 -86.875 ;
        RECT -13.085 -91.285 -12.755 -90.955 ;
        RECT -13.085 -92.645 -12.755 -92.315 ;
        RECT -13.085 -94.005 -12.755 -93.675 ;
        RECT -13.085 -96.725 -12.755 -96.395 ;
        RECT -13.085 -98.085 -12.755 -97.755 ;
        RECT -13.085 -98.89 -12.755 -98.56 ;
        RECT -13.085 -100.805 -12.755 -100.475 ;
        RECT -13.085 -102.165 -12.755 -101.835 ;
        RECT -13.085 -104.885 -12.755 -104.555 ;
        RECT -13.085 -107.43 -12.755 -107.1 ;
        RECT -13.085 -114.405 -12.755 -114.075 ;
        RECT -13.085 -115.765 -12.755 -115.435 ;
        RECT -13.085 -117.125 -12.755 -116.795 ;
        RECT -13.085 -118.485 -12.755 -118.155 ;
        RECT -13.085 -119.845 -12.755 -119.515 ;
        RECT -13.085 -121.205 -12.755 -120.875 ;
        RECT -13.085 -132.085 -12.755 -131.755 ;
        RECT -13.085 -134.805 -12.755 -134.475 ;
        RECT -13.085 -136.165 -12.755 -135.835 ;
        RECT -13.085 -137.525 -12.755 -137.195 ;
        RECT -13.085 -141.605 -12.755 -141.275 ;
        RECT -13.085 -144.325 -12.755 -143.995 ;
        RECT -13.085 -147.045 -12.755 -146.715 ;
        RECT -13.085 -148.405 -12.755 -148.075 ;
        RECT -13.085 -151.125 -12.755 -150.795 ;
        RECT -13.085 -152.485 -12.755 -152.155 ;
        RECT -13.085 -156.565 -12.755 -156.235 ;
        RECT -13.085 -159.285 -12.755 -158.955 ;
        RECT -13.085 -160.645 -12.755 -160.315 ;
        RECT -13.085 -162.005 -12.755 -161.675 ;
        RECT -13.085 -163.365 -12.755 -163.035 ;
        RECT -13.085 -164.725 -12.755 -164.395 ;
        RECT -13.085 -166.085 -12.755 -165.755 ;
        RECT -13.085 -171.525 -12.755 -171.195 ;
        RECT -13.085 -172.885 -12.755 -172.555 ;
        RECT -13.085 -174.245 -12.755 -173.915 ;
        RECT -13.085 -175.605 -12.755 -175.275 ;
        RECT -13.085 -176.685 -12.755 -176.355 ;
        RECT -13.085 -178.325 -12.755 -177.995 ;
        RECT -13.085 -179.685 -12.755 -179.355 ;
        RECT -13.085 -181.93 -12.755 -180.8 ;
        RECT -13.08 -182.045 -12.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.725 241.32 -11.395 242.45 ;
        RECT -11.725 239.195 -11.395 239.525 ;
        RECT -11.725 237.835 -11.395 238.165 ;
        RECT -11.725 236.475 -11.395 236.805 ;
        RECT -11.725 235.115 -11.395 235.445 ;
        RECT -11.725 233.755 -11.395 234.085 ;
        RECT -11.725 232.395 -11.395 232.725 ;
        RECT -11.725 231.035 -11.395 231.365 ;
        RECT -11.725 229.675 -11.395 230.005 ;
        RECT -11.725 228.315 -11.395 228.645 ;
        RECT -11.725 226.955 -11.395 227.285 ;
        RECT -11.725 225.595 -11.395 225.925 ;
        RECT -11.725 224.235 -11.395 224.565 ;
        RECT -11.725 222.875 -11.395 223.205 ;
        RECT -11.725 221.515 -11.395 221.845 ;
        RECT -11.725 220.155 -11.395 220.485 ;
        RECT -11.725 218.795 -11.395 219.125 ;
        RECT -11.725 217.435 -11.395 217.765 ;
        RECT -11.725 216.075 -11.395 216.405 ;
        RECT -11.725 214.715 -11.395 215.045 ;
        RECT -11.725 213.355 -11.395 213.685 ;
        RECT -11.725 211.995 -11.395 212.325 ;
        RECT -11.725 210.635 -11.395 210.965 ;
        RECT -11.725 209.275 -11.395 209.605 ;
        RECT -11.725 207.915 -11.395 208.245 ;
        RECT -11.725 206.555 -11.395 206.885 ;
        RECT -11.725 205.195 -11.395 205.525 ;
        RECT -11.725 203.835 -11.395 204.165 ;
        RECT -11.725 202.475 -11.395 202.805 ;
        RECT -11.725 201.115 -11.395 201.445 ;
        RECT -11.725 199.755 -11.395 200.085 ;
        RECT -11.725 198.395 -11.395 198.725 ;
        RECT -11.725 197.035 -11.395 197.365 ;
        RECT -11.725 195.675 -11.395 196.005 ;
        RECT -11.725 194.315 -11.395 194.645 ;
        RECT -11.725 192.955 -11.395 193.285 ;
        RECT -11.725 191.595 -11.395 191.925 ;
        RECT -11.725 190.235 -11.395 190.565 ;
        RECT -11.725 188.875 -11.395 189.205 ;
        RECT -11.725 187.515 -11.395 187.845 ;
        RECT -11.725 186.155 -11.395 186.485 ;
        RECT -11.725 184.795 -11.395 185.125 ;
        RECT -11.725 183.435 -11.395 183.765 ;
        RECT -11.725 182.075 -11.395 182.405 ;
        RECT -11.725 180.715 -11.395 181.045 ;
        RECT -11.725 179.355 -11.395 179.685 ;
        RECT -11.725 177.995 -11.395 178.325 ;
        RECT -11.725 176.635 -11.395 176.965 ;
        RECT -11.725 175.275 -11.395 175.605 ;
        RECT -11.725 173.915 -11.395 174.245 ;
        RECT -11.725 172.555 -11.395 172.885 ;
        RECT -11.725 171.195 -11.395 171.525 ;
        RECT -11.725 169.835 -11.395 170.165 ;
        RECT -11.725 168.475 -11.395 168.805 ;
        RECT -11.725 167.115 -11.395 167.445 ;
        RECT -11.725 165.755 -11.395 166.085 ;
        RECT -11.725 164.395 -11.395 164.725 ;
        RECT -11.725 163.035 -11.395 163.365 ;
        RECT -11.725 161.675 -11.395 162.005 ;
        RECT -11.725 160.315 -11.395 160.645 ;
        RECT -11.725 158.955 -11.395 159.285 ;
        RECT -11.725 157.595 -11.395 157.925 ;
        RECT -11.725 156.235 -11.395 156.565 ;
        RECT -11.725 154.875 -11.395 155.205 ;
        RECT -11.725 153.515 -11.395 153.845 ;
        RECT -11.725 152.155 -11.395 152.485 ;
        RECT -11.725 150.795 -11.395 151.125 ;
        RECT -11.725 149.435 -11.395 149.765 ;
        RECT -11.725 148.075 -11.395 148.405 ;
        RECT -11.725 146.715 -11.395 147.045 ;
        RECT -11.725 145.355 -11.395 145.685 ;
        RECT -11.725 143.995 -11.395 144.325 ;
        RECT -11.725 142.635 -11.395 142.965 ;
        RECT -11.725 141.275 -11.395 141.605 ;
        RECT -11.725 139.915 -11.395 140.245 ;
        RECT -11.725 138.555 -11.395 138.885 ;
        RECT -11.725 137.195 -11.395 137.525 ;
        RECT -11.725 135.835 -11.395 136.165 ;
        RECT -11.725 134.475 -11.395 134.805 ;
        RECT -11.725 133.115 -11.395 133.445 ;
        RECT -11.725 131.755 -11.395 132.085 ;
        RECT -11.725 130.395 -11.395 130.725 ;
        RECT -11.725 129.035 -11.395 129.365 ;
        RECT -11.725 127.675 -11.395 128.005 ;
        RECT -11.725 126.315 -11.395 126.645 ;
        RECT -11.725 124.955 -11.395 125.285 ;
        RECT -11.725 123.595 -11.395 123.925 ;
        RECT -11.725 122.235 -11.395 122.565 ;
        RECT -11.725 120.875 -11.395 121.205 ;
        RECT -11.725 119.515 -11.395 119.845 ;
        RECT -11.725 118.155 -11.395 118.485 ;
        RECT -11.725 116.795 -11.395 117.125 ;
        RECT -11.725 115.435 -11.395 115.765 ;
        RECT -11.725 114.075 -11.395 114.405 ;
        RECT -11.725 112.715 -11.395 113.045 ;
        RECT -11.725 111.355 -11.395 111.685 ;
        RECT -11.725 109.995 -11.395 110.325 ;
        RECT -11.725 108.635 -11.395 108.965 ;
        RECT -11.725 107.275 -11.395 107.605 ;
        RECT -11.725 105.915 -11.395 106.245 ;
        RECT -11.725 104.555 -11.395 104.885 ;
        RECT -11.725 103.195 -11.395 103.525 ;
        RECT -11.725 101.835 -11.395 102.165 ;
        RECT -11.725 100.475 -11.395 100.805 ;
        RECT -11.725 99.115 -11.395 99.445 ;
        RECT -11.725 97.755 -11.395 98.085 ;
        RECT -11.725 96.395 -11.395 96.725 ;
        RECT -11.725 95.035 -11.395 95.365 ;
        RECT -11.725 93.675 -11.395 94.005 ;
        RECT -11.725 92.315 -11.395 92.645 ;
        RECT -11.725 90.955 -11.395 91.285 ;
        RECT -11.725 89.595 -11.395 89.925 ;
        RECT -11.725 88.235 -11.395 88.565 ;
        RECT -11.725 86.875 -11.395 87.205 ;
        RECT -11.725 85.515 -11.395 85.845 ;
        RECT -11.725 84.155 -11.395 84.485 ;
        RECT -11.725 82.795 -11.395 83.125 ;
        RECT -11.725 81.435 -11.395 81.765 ;
        RECT -11.725 80.075 -11.395 80.405 ;
        RECT -11.725 78.715 -11.395 79.045 ;
        RECT -11.725 77.355 -11.395 77.685 ;
        RECT -11.725 75.995 -11.395 76.325 ;
        RECT -11.725 74.635 -11.395 74.965 ;
        RECT -11.725 73.275 -11.395 73.605 ;
        RECT -11.725 71.915 -11.395 72.245 ;
        RECT -11.725 70.555 -11.395 70.885 ;
        RECT -11.725 69.195 -11.395 69.525 ;
        RECT -11.725 67.835 -11.395 68.165 ;
        RECT -11.725 66.475 -11.395 66.805 ;
        RECT -11.725 65.115 -11.395 65.445 ;
        RECT -11.725 63.755 -11.395 64.085 ;
        RECT -11.725 62.395 -11.395 62.725 ;
        RECT -11.725 61.035 -11.395 61.365 ;
        RECT -11.725 59.675 -11.395 60.005 ;
        RECT -11.725 58.315 -11.395 58.645 ;
        RECT -11.725 56.955 -11.395 57.285 ;
        RECT -11.725 55.595 -11.395 55.925 ;
        RECT -11.725 54.235 -11.395 54.565 ;
        RECT -11.725 52.875 -11.395 53.205 ;
        RECT -11.725 51.515 -11.395 51.845 ;
        RECT -11.725 50.155 -11.395 50.485 ;
        RECT -11.725 48.795 -11.395 49.125 ;
        RECT -11.725 47.435 -11.395 47.765 ;
        RECT -11.725 46.075 -11.395 46.405 ;
        RECT -11.725 44.715 -11.395 45.045 ;
        RECT -11.725 43.355 -11.395 43.685 ;
        RECT -11.725 41.995 -11.395 42.325 ;
        RECT -11.725 40.635 -11.395 40.965 ;
        RECT -11.725 39.275 -11.395 39.605 ;
        RECT -11.725 37.915 -11.395 38.245 ;
        RECT -11.725 36.555 -11.395 36.885 ;
        RECT -11.725 35.195 -11.395 35.525 ;
        RECT -11.725 33.835 -11.395 34.165 ;
        RECT -11.725 32.475 -11.395 32.805 ;
        RECT -11.725 31.115 -11.395 31.445 ;
        RECT -11.725 29.755 -11.395 30.085 ;
        RECT -11.725 28.395 -11.395 28.725 ;
        RECT -11.725 27.035 -11.395 27.365 ;
        RECT -11.725 25.675 -11.395 26.005 ;
        RECT -11.725 24.315 -11.395 24.645 ;
        RECT -11.725 22.955 -11.395 23.285 ;
        RECT -11.725 21.595 -11.395 21.925 ;
        RECT -11.725 20.235 -11.395 20.565 ;
        RECT -11.725 18.875 -11.395 19.205 ;
        RECT -11.725 17.515 -11.395 17.845 ;
        RECT -11.725 16.155 -11.395 16.485 ;
        RECT -11.725 14.795 -11.395 15.125 ;
        RECT -11.725 13.435 -11.395 13.765 ;
        RECT -11.725 12.075 -11.395 12.405 ;
        RECT -11.725 10.715 -11.395 11.045 ;
        RECT -11.725 9.355 -11.395 9.685 ;
        RECT -11.725 7.995 -11.395 8.325 ;
        RECT -11.725 6.635 -11.395 6.965 ;
        RECT -11.725 5.275 -11.395 5.605 ;
        RECT -11.725 3.915 -11.395 4.245 ;
        RECT -11.725 2.555 -11.395 2.885 ;
        RECT -11.725 1.195 -11.395 1.525 ;
        RECT -11.725 -0.165 -11.395 0.165 ;
        RECT -11.725 -2.885 -11.395 -2.555 ;
        RECT -11.725 -4.245 -11.395 -3.915 ;
        RECT -11.725 -5.605 -11.395 -5.275 ;
        RECT -11.725 -6.965 -11.395 -6.635 ;
        RECT -11.725 -8.325 -11.395 -7.995 ;
        RECT -11.725 -9.685 -11.395 -9.355 ;
        RECT -11.725 -12.405 -11.395 -12.075 ;
        RECT -11.725 -13.765 -11.395 -13.435 ;
        RECT -11.725 -14.95 -11.395 -14.62 ;
        RECT -11.725 -17.845 -11.395 -17.515 ;
        RECT -11.72 -17.845 -11.4 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -11.725 -107.43 -11.395 -107.1 ;
        RECT -11.725 -114.405 -11.395 -114.075 ;
        RECT -11.725 -115.765 -11.395 -115.435 ;
        RECT -11.725 -117.125 -11.395 -116.795 ;
        RECT -11.725 -118.485 -11.395 -118.155 ;
        RECT -11.725 -119.845 -11.395 -119.515 ;
        RECT -11.725 -121.205 -11.395 -120.875 ;
        RECT -11.725 -128.005 -11.395 -127.675 ;
        RECT -11.725 -130.725 -11.395 -130.395 ;
        RECT -11.725 -132.085 -11.395 -131.755 ;
        RECT -11.725 -134.805 -11.395 -134.475 ;
        RECT -11.725 -136.165 -11.395 -135.835 ;
        RECT -11.725 -137.525 -11.395 -137.195 ;
        RECT -11.725 -138.885 -11.395 -138.555 ;
        RECT -11.725 -140.245 -11.395 -139.915 ;
        RECT -11.725 -141.605 -11.395 -141.275 ;
        RECT -11.725 -142.965 -11.395 -142.635 ;
        RECT -11.725 -144.325 -11.395 -143.995 ;
        RECT -11.725 -147.045 -11.395 -146.715 ;
        RECT -11.725 -148.405 -11.395 -148.075 ;
        RECT -11.725 -151.125 -11.395 -150.795 ;
        RECT -11.725 -152.485 -11.395 -152.155 ;
        RECT -11.725 -155.205 -11.395 -154.875 ;
        RECT -11.725 -156.565 -11.395 -156.235 ;
        RECT -11.725 -159.285 -11.395 -158.955 ;
        RECT -11.725 -160.645 -11.395 -160.315 ;
        RECT -11.725 -162.005 -11.395 -161.675 ;
        RECT -11.725 -163.365 -11.395 -163.035 ;
        RECT -11.725 -164.725 -11.395 -164.395 ;
        RECT -11.725 -166.085 -11.395 -165.755 ;
        RECT -11.725 -171.525 -11.395 -171.195 ;
        RECT -11.725 -172.885 -11.395 -172.555 ;
        RECT -11.725 -174.245 -11.395 -173.915 ;
        RECT -11.725 -175.605 -11.395 -175.275 ;
        RECT -11.725 -176.685 -11.395 -176.355 ;
        RECT -11.725 -178.325 -11.395 -177.995 ;
        RECT -11.725 -179.685 -11.395 -179.355 ;
        RECT -11.725 -181.93 -11.395 -180.8 ;
        RECT -11.72 -182.045 -11.4 -105.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.365 241.32 -10.035 242.45 ;
        RECT -10.365 239.195 -10.035 239.525 ;
        RECT -10.365 237.835 -10.035 238.165 ;
        RECT -10.365 236.475 -10.035 236.805 ;
        RECT -10.365 235.115 -10.035 235.445 ;
        RECT -10.365 233.755 -10.035 234.085 ;
        RECT -10.365 232.395 -10.035 232.725 ;
        RECT -10.365 231.035 -10.035 231.365 ;
        RECT -10.365 221.515 -10.035 221.845 ;
        RECT -10.365 217.435 -10.035 217.765 ;
        RECT -10.365 213.355 -10.035 213.685 ;
        RECT -10.365 210.635 -10.035 210.965 ;
        RECT -10.365 203.835 -10.035 204.165 ;
        RECT -10.365 202.475 -10.035 202.805 ;
        RECT -10.365 199.755 -10.035 200.085 ;
        RECT -10.365 192.955 -10.035 193.285 ;
        RECT -10.365 190.235 -10.035 190.565 ;
        RECT -10.365 188.875 -10.035 189.205 ;
        RECT -10.365 184.795 -10.035 185.125 ;
        RECT -10.365 182.075 -10.035 182.405 ;
        RECT -10.365 175.275 -10.035 175.605 ;
        RECT -10.365 173.915 -10.035 174.245 ;
        RECT -10.365 171.195 -10.035 171.525 ;
        RECT -10.365 164.395 -10.035 164.725 ;
        RECT -10.365 161.675 -10.035 162.005 ;
        RECT -10.365 160.315 -10.035 160.645 ;
        RECT -10.365 153.515 -10.035 153.845 ;
        RECT -10.365 150.795 -10.035 151.125 ;
        RECT -10.365 146.715 -10.035 147.045 ;
        RECT -10.365 145.355 -10.035 145.685 ;
        RECT -10.365 142.635 -10.035 142.965 ;
        RECT -10.365 135.835 -10.035 136.165 ;
        RECT -10.365 133.115 -10.035 133.445 ;
        RECT -10.365 131.755 -10.035 132.085 ;
        RECT -10.365 124.955 -10.035 125.285 ;
        RECT -10.365 122.235 -10.035 122.565 ;
        RECT -10.365 118.155 -10.035 118.485 ;
        RECT -10.365 114.075 -10.035 114.405 ;
        RECT -10.365 104.555 -10.035 104.885 ;
        RECT -10.365 103.195 -10.035 103.525 ;
        RECT -10.365 96.395 -10.035 96.725 ;
        RECT -10.365 93.675 -10.035 94.005 ;
        RECT -10.365 89.595 -10.035 89.925 ;
        RECT -10.365 85.515 -10.035 85.845 ;
        RECT -10.365 82.795 -10.035 83.125 ;
        RECT -10.365 75.995 -10.035 76.325 ;
        RECT -10.365 74.635 -10.035 74.965 ;
        RECT -10.365 65.115 -10.035 65.445 ;
        RECT -10.365 61.035 -10.035 61.365 ;
        RECT -10.365 56.955 -10.035 57.285 ;
        RECT -10.365 54.235 -10.035 54.565 ;
        RECT -10.365 47.435 -10.035 47.765 ;
        RECT -10.365 46.075 -10.035 46.405 ;
        RECT -10.365 43.355 -10.035 43.685 ;
        RECT -10.365 36.555 -10.035 36.885 ;
        RECT -10.365 33.835 -10.035 34.165 ;
        RECT -10.365 32.475 -10.035 32.805 ;
        RECT -10.365 28.395 -10.035 28.725 ;
        RECT -10.365 25.675 -10.035 26.005 ;
        RECT -10.365 18.875 -10.035 19.205 ;
        RECT -10.365 17.515 -10.035 17.845 ;
        RECT -10.365 14.795 -10.035 15.125 ;
        RECT -10.365 7.995 -10.035 8.325 ;
        RECT -10.365 5.275 -10.035 5.605 ;
        RECT -10.365 3.915 -10.035 4.245 ;
        RECT -10.365 2.555 -10.035 2.885 ;
        RECT -10.365 1.195 -10.035 1.525 ;
        RECT -10.365 -0.165 -10.035 0.165 ;
        RECT -10.365 -2.885 -10.035 -2.555 ;
        RECT -10.365 -4.245 -10.035 -3.915 ;
        RECT -10.365 -5.605 -10.035 -5.275 ;
        RECT -10.365 -6.965 -10.035 -6.635 ;
        RECT -10.365 -8.325 -10.035 -7.995 ;
        RECT -10.365 -9.685 -10.035 -9.355 ;
        RECT -10.365 -12.405 -10.035 -12.075 ;
        RECT -10.365 -13.765 -10.035 -13.435 ;
        RECT -10.365 -14.95 -10.035 -14.62 ;
        RECT -10.365 -17.845 -10.035 -17.515 ;
        RECT -10.365 -19.79 -10.035 -19.46 ;
        RECT -10.365 -26.005 -10.035 -25.675 ;
        RECT -10.365 -27.365 -10.035 -27.035 ;
        RECT -10.365 -28.725 -10.035 -28.395 ;
        RECT -10.365 -30.085 -10.035 -29.755 ;
        RECT -10.365 -31.445 -10.035 -31.115 ;
        RECT -10.365 -32.805 -10.035 -32.475 ;
        RECT -10.365 -35.525 -10.035 -35.195 ;
        RECT -10.365 -36.885 -10.035 -36.555 ;
        RECT -10.365 -37.93 -10.035 -37.6 ;
        RECT -10.365 -42.77 -10.035 -42.44 ;
        RECT -10.365 -51.845 -10.035 -51.515 ;
        RECT -10.365 -53.205 -10.035 -52.875 ;
        RECT -10.365 -54.565 -10.035 -54.235 ;
        RECT -10.365 -55.925 -10.035 -55.595 ;
        RECT -10.365 -57.285 -10.035 -56.955 ;
        RECT -10.365 -58.645 -10.035 -58.315 ;
        RECT -10.365 -60.005 -10.035 -59.675 ;
        RECT -10.365 -61.365 -10.035 -61.035 ;
        RECT -10.365 -62.725 -10.035 -62.395 ;
        RECT -10.365 -64.085 -10.035 -63.755 ;
        RECT -10.365 -65.445 -10.035 -65.115 ;
        RECT -10.365 -68.165 -10.035 -67.835 ;
        RECT -10.365 -69.525 -10.035 -69.195 ;
        RECT -10.365 -70.885 -10.035 -70.555 ;
        RECT -10.365 -72.245 -10.035 -71.915 ;
        RECT -10.365 -74.965 -10.035 -74.635 ;
        RECT -10.365 -76.71 -10.035 -76.38 ;
        RECT -10.365 -77.685 -10.035 -77.355 ;
        RECT -10.365 -79.045 -10.035 -78.715 ;
        RECT -10.365 -81.765 -10.035 -81.435 ;
        RECT -10.365 -83.125 -10.035 -82.795 ;
        RECT -10.365 -84.485 -10.035 -84.155 ;
        RECT -10.365 -85.25 -10.035 -84.92 ;
        RECT -10.365 -87.205 -10.035 -86.875 ;
        RECT -10.365 -91.285 -10.035 -90.955 ;
        RECT -10.365 -92.645 -10.035 -92.315 ;
        RECT -10.365 -94.005 -10.035 -93.675 ;
        RECT -10.365 -96.725 -10.035 -96.395 ;
        RECT -10.365 -98.085 -10.035 -97.755 ;
        RECT -10.365 -98.89 -10.035 -98.56 ;
        RECT -10.365 -100.805 -10.035 -100.475 ;
        RECT -10.365 -102.165 -10.035 -101.835 ;
        RECT -10.365 -104.885 -10.035 -104.555 ;
        RECT -10.365 -107.43 -10.035 -107.1 ;
        RECT -10.365 -114.405 -10.035 -114.075 ;
        RECT -10.365 -115.765 -10.035 -115.435 ;
        RECT -10.365 -117.125 -10.035 -116.795 ;
        RECT -10.365 -118.485 -10.035 -118.155 ;
        RECT -10.365 -119.845 -10.035 -119.515 ;
        RECT -10.365 -121.205 -10.035 -120.875 ;
        RECT -10.365 -125.285 -10.035 -124.955 ;
        RECT -10.365 -128.005 -10.035 -127.675 ;
        RECT -10.365 -129.365 -10.035 -129.035 ;
        RECT -10.365 -130.725 -10.035 -130.395 ;
        RECT -10.365 -132.085 -10.035 -131.755 ;
        RECT -10.365 -134.805 -10.035 -134.475 ;
        RECT -10.365 -136.165 -10.035 -135.835 ;
        RECT -10.365 -137.525 -10.035 -137.195 ;
        RECT -10.365 -138.885 -10.035 -138.555 ;
        RECT -10.365 -140.245 -10.035 -139.915 ;
        RECT -10.365 -141.605 -10.035 -141.275 ;
        RECT -10.365 -142.965 -10.035 -142.635 ;
        RECT -10.365 -144.325 -10.035 -143.995 ;
        RECT -10.365 -147.045 -10.035 -146.715 ;
        RECT -10.365 -148.405 -10.035 -148.075 ;
        RECT -10.365 -149.765 -10.035 -149.435 ;
        RECT -10.365 -151.125 -10.035 -150.795 ;
        RECT -10.365 -152.485 -10.035 -152.155 ;
        RECT -10.365 -153.845 -10.035 -153.515 ;
        RECT -10.365 -155.205 -10.035 -154.875 ;
        RECT -10.365 -156.565 -10.035 -156.235 ;
        RECT -10.365 -157.925 -10.035 -157.595 ;
        RECT -10.365 -159.285 -10.035 -158.955 ;
        RECT -10.365 -160.645 -10.035 -160.315 ;
        RECT -10.365 -162.005 -10.035 -161.675 ;
        RECT -10.365 -163.365 -10.035 -163.035 ;
        RECT -10.365 -164.725 -10.035 -164.395 ;
        RECT -10.365 -166.085 -10.035 -165.755 ;
        RECT -10.36 -168.12 -10.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -10.365 -175.605 -10.035 -175.275 ;
        RECT -10.365 -178.325 -10.035 -177.995 ;
        RECT -10.365 -179.685 -10.035 -179.355 ;
        RECT -10.365 -181.93 -10.035 -180.8 ;
        RECT -10.36 -182.045 -10.04 -173.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.005 241.32 -8.675 242.45 ;
        RECT -9.005 239.195 -8.675 239.525 ;
        RECT -9.005 237.835 -8.675 238.165 ;
        RECT -9.005 236.475 -8.675 236.805 ;
        RECT -9.005 235.115 -8.675 235.445 ;
        RECT -9.005 233.755 -8.675 234.085 ;
        RECT -9.005 232.395 -8.675 232.725 ;
        RECT -9.005 231.035 -8.675 231.365 ;
        RECT -9.005 221.515 -8.675 221.845 ;
        RECT -9.005 217.435 -8.675 217.765 ;
        RECT -9.005 213.355 -8.675 213.685 ;
        RECT -9.005 210.635 -8.675 210.965 ;
        RECT -9.005 203.835 -8.675 204.165 ;
        RECT -9.005 202.475 -8.675 202.805 ;
        RECT -9.005 199.755 -8.675 200.085 ;
        RECT -9.005 192.955 -8.675 193.285 ;
        RECT -9.005 190.235 -8.675 190.565 ;
        RECT -9.005 188.875 -8.675 189.205 ;
        RECT -9.005 184.795 -8.675 185.125 ;
        RECT -9.005 182.075 -8.675 182.405 ;
        RECT -9.005 175.275 -8.675 175.605 ;
        RECT -9.005 173.915 -8.675 174.245 ;
        RECT -9.005 171.195 -8.675 171.525 ;
        RECT -9.005 164.395 -8.675 164.725 ;
        RECT -9.005 161.675 -8.675 162.005 ;
        RECT -9.005 160.315 -8.675 160.645 ;
        RECT -9.005 153.515 -8.675 153.845 ;
        RECT -9.005 150.795 -8.675 151.125 ;
        RECT -9.005 146.715 -8.675 147.045 ;
        RECT -9.005 145.355 -8.675 145.685 ;
        RECT -9.005 142.635 -8.675 142.965 ;
        RECT -9.005 135.835 -8.675 136.165 ;
        RECT -9.005 133.115 -8.675 133.445 ;
        RECT -9.005 131.755 -8.675 132.085 ;
        RECT -9.005 124.955 -8.675 125.285 ;
        RECT -9.005 122.235 -8.675 122.565 ;
        RECT -9.005 118.155 -8.675 118.485 ;
        RECT -9.005 114.075 -8.675 114.405 ;
        RECT -9.005 104.555 -8.675 104.885 ;
        RECT -9.005 103.195 -8.675 103.525 ;
        RECT -9.005 96.395 -8.675 96.725 ;
        RECT -9.005 93.675 -8.675 94.005 ;
        RECT -9.005 89.595 -8.675 89.925 ;
        RECT -9.005 85.515 -8.675 85.845 ;
        RECT -9.005 82.795 -8.675 83.125 ;
        RECT -9.005 75.995 -8.675 76.325 ;
        RECT -9.005 74.635 -8.675 74.965 ;
        RECT -9.005 65.115 -8.675 65.445 ;
        RECT -9.005 61.035 -8.675 61.365 ;
        RECT -9.005 56.955 -8.675 57.285 ;
        RECT -9.005 54.235 -8.675 54.565 ;
        RECT -9.005 47.435 -8.675 47.765 ;
        RECT -9.005 46.075 -8.675 46.405 ;
        RECT -9.005 43.355 -8.675 43.685 ;
        RECT -9.005 36.555 -8.675 36.885 ;
        RECT -9.005 33.835 -8.675 34.165 ;
        RECT -9.005 32.475 -8.675 32.805 ;
        RECT -9.005 28.395 -8.675 28.725 ;
        RECT -9.005 25.675 -8.675 26.005 ;
        RECT -9.005 18.875 -8.675 19.205 ;
        RECT -9.005 17.515 -8.675 17.845 ;
        RECT -9.005 14.795 -8.675 15.125 ;
        RECT -9.005 7.995 -8.675 8.325 ;
        RECT -9.005 5.275 -8.675 5.605 ;
        RECT -9.005 3.915 -8.675 4.245 ;
        RECT -9.005 2.555 -8.675 2.885 ;
        RECT -9.005 1.195 -8.675 1.525 ;
        RECT -9.005 -0.165 -8.675 0.165 ;
        RECT -9.005 -2.885 -8.675 -2.555 ;
        RECT -9.005 -4.245 -8.675 -3.915 ;
        RECT -9.005 -5.605 -8.675 -5.275 ;
        RECT -9.005 -6.965 -8.675 -6.635 ;
        RECT -9.005 -8.325 -8.675 -7.995 ;
        RECT -9.005 -9.685 -8.675 -9.355 ;
        RECT -9.005 -11.045 -8.675 -10.715 ;
        RECT -9.005 -12.405 -8.675 -12.075 ;
        RECT -9.005 -13.765 -8.675 -13.435 ;
        RECT -9.005 -15.125 -8.675 -14.795 ;
        RECT -9.005 -16.485 -8.675 -16.155 ;
        RECT -9.005 -17.845 -8.675 -17.515 ;
        RECT -9.005 -19.205 -8.675 -18.875 ;
        RECT -9 -22.6 -8.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -9.005 -110.325 -8.675 -109.995 ;
        RECT -9.005 -111.685 -8.675 -111.355 ;
        RECT -9.005 -113.045 -8.675 -112.715 ;
        RECT -9.005 -114.405 -8.675 -114.075 ;
        RECT -9.005 -115.765 -8.675 -115.435 ;
        RECT -9.005 -117.125 -8.675 -116.795 ;
        RECT -9.005 -118.485 -8.675 -118.155 ;
        RECT -9.005 -119.845 -8.675 -119.515 ;
        RECT -9.005 -121.205 -8.675 -120.875 ;
        RECT -9.005 -123.925 -8.675 -123.595 ;
        RECT -9.005 -125.285 -8.675 -124.955 ;
        RECT -9.005 -126.645 -8.675 -126.315 ;
        RECT -9.005 -128.005 -8.675 -127.675 ;
        RECT -9.005 -129.365 -8.675 -129.035 ;
        RECT -9.005 -130.725 -8.675 -130.395 ;
        RECT -9.005 -132.085 -8.675 -131.755 ;
        RECT -9.005 -133.445 -8.675 -133.115 ;
        RECT -9.005 -134.805 -8.675 -134.475 ;
        RECT -9.005 -136.165 -8.675 -135.835 ;
        RECT -9.005 -137.525 -8.675 -137.195 ;
        RECT -9.005 -138.885 -8.675 -138.555 ;
        RECT -9.005 -140.245 -8.675 -139.915 ;
        RECT -9.005 -141.605 -8.675 -141.275 ;
        RECT -9.005 -142.965 -8.675 -142.635 ;
        RECT -9.005 -144.325 -8.675 -143.995 ;
        RECT -9.005 -145.685 -8.675 -145.355 ;
        RECT -9.005 -147.045 -8.675 -146.715 ;
        RECT -9.005 -148.405 -8.675 -148.075 ;
        RECT -9.005 -149.765 -8.675 -149.435 ;
        RECT -9.005 -151.125 -8.675 -150.795 ;
        RECT -9.005 -152.485 -8.675 -152.155 ;
        RECT -9.005 -153.845 -8.675 -153.515 ;
        RECT -9.005 -155.205 -8.675 -154.875 ;
        RECT -9.005 -156.565 -8.675 -156.235 ;
        RECT -9.005 -157.925 -8.675 -157.595 ;
        RECT -9.005 -159.285 -8.675 -158.955 ;
        RECT -9.005 -160.645 -8.675 -160.315 ;
        RECT -9.005 -162.005 -8.675 -161.675 ;
        RECT -9.005 -163.365 -8.675 -163.035 ;
        RECT -9.005 -164.725 -8.675 -164.395 ;
        RECT -9.005 -166.085 -8.675 -165.755 ;
        RECT -9 -166.76 -8.68 -109.32 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.645 241.32 -7.315 242.45 ;
        RECT -7.645 239.195 -7.315 239.525 ;
        RECT -7.645 237.835 -7.315 238.165 ;
        RECT -7.645 236.475 -7.315 236.805 ;
        RECT -7.645 235.115 -7.315 235.445 ;
        RECT -7.645 233.755 -7.315 234.085 ;
        RECT -7.645 232.395 -7.315 232.725 ;
        RECT -7.645 231.035 -7.315 231.365 ;
        RECT -7.645 221.515 -7.315 221.845 ;
        RECT -7.645 217.435 -7.315 217.765 ;
        RECT -7.645 213.355 -7.315 213.685 ;
        RECT -7.645 210.635 -7.315 210.965 ;
        RECT -7.645 203.835 -7.315 204.165 ;
        RECT -7.645 202.475 -7.315 202.805 ;
        RECT -7.645 199.755 -7.315 200.085 ;
        RECT -7.645 192.955 -7.315 193.285 ;
        RECT -7.645 190.235 -7.315 190.565 ;
        RECT -7.645 188.875 -7.315 189.205 ;
        RECT -7.645 184.795 -7.315 185.125 ;
        RECT -7.645 182.075 -7.315 182.405 ;
        RECT -7.645 175.275 -7.315 175.605 ;
        RECT -7.645 173.915 -7.315 174.245 ;
        RECT -7.645 171.195 -7.315 171.525 ;
        RECT -7.645 164.395 -7.315 164.725 ;
        RECT -7.645 161.675 -7.315 162.005 ;
        RECT -7.645 160.315 -7.315 160.645 ;
        RECT -7.645 153.515 -7.315 153.845 ;
        RECT -7.645 150.795 -7.315 151.125 ;
        RECT -7.645 146.715 -7.315 147.045 ;
        RECT -7.645 145.355 -7.315 145.685 ;
        RECT -7.645 142.635 -7.315 142.965 ;
        RECT -7.645 135.835 -7.315 136.165 ;
        RECT -7.645 133.115 -7.315 133.445 ;
        RECT -7.645 131.755 -7.315 132.085 ;
        RECT -7.645 124.955 -7.315 125.285 ;
        RECT -7.645 122.235 -7.315 122.565 ;
        RECT -7.645 118.155 -7.315 118.485 ;
        RECT -7.645 114.075 -7.315 114.405 ;
        RECT -7.645 104.555 -7.315 104.885 ;
        RECT -7.645 103.195 -7.315 103.525 ;
        RECT -7.645 96.395 -7.315 96.725 ;
        RECT -7.645 93.675 -7.315 94.005 ;
        RECT -7.645 89.595 -7.315 89.925 ;
        RECT -7.645 85.515 -7.315 85.845 ;
        RECT -7.645 82.795 -7.315 83.125 ;
        RECT -7.645 75.995 -7.315 76.325 ;
        RECT -7.645 74.635 -7.315 74.965 ;
        RECT -7.645 65.115 -7.315 65.445 ;
        RECT -7.645 61.035 -7.315 61.365 ;
        RECT -7.645 56.955 -7.315 57.285 ;
        RECT -7.645 54.235 -7.315 54.565 ;
        RECT -7.645 47.435 -7.315 47.765 ;
        RECT -7.645 46.075 -7.315 46.405 ;
        RECT -7.645 43.355 -7.315 43.685 ;
        RECT -7.645 36.555 -7.315 36.885 ;
        RECT -7.645 33.835 -7.315 34.165 ;
        RECT -7.645 32.475 -7.315 32.805 ;
        RECT -7.645 28.395 -7.315 28.725 ;
        RECT -7.645 25.675 -7.315 26.005 ;
        RECT -7.645 18.875 -7.315 19.205 ;
        RECT -7.645 17.515 -7.315 17.845 ;
        RECT -7.645 14.795 -7.315 15.125 ;
        RECT -7.645 7.995 -7.315 8.325 ;
        RECT -7.645 5.275 -7.315 5.605 ;
        RECT -7.645 3.915 -7.315 4.245 ;
        RECT -7.645 2.555 -7.315 2.885 ;
        RECT -7.645 1.195 -7.315 1.525 ;
        RECT -7.645 -0.165 -7.315 0.165 ;
        RECT -7.645 -2.885 -7.315 -2.555 ;
        RECT -7.645 -4.245 -7.315 -3.915 ;
        RECT -7.645 -5.605 -7.315 -5.275 ;
        RECT -7.645 -6.965 -7.315 -6.635 ;
        RECT -7.645 -8.325 -7.315 -7.995 ;
        RECT -7.645 -9.685 -7.315 -9.355 ;
        RECT -7.645 -12.405 -7.315 -12.075 ;
        RECT -7.645 -13.765 -7.315 -13.435 ;
        RECT -7.645 -15.125 -7.315 -14.795 ;
        RECT -7.645 -16.485 -7.315 -16.155 ;
        RECT -7.645 -17.845 -7.315 -17.515 ;
        RECT -7.64 -18.52 -7.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -7.645 -160.645 -7.315 -160.315 ;
        RECT -7.645 -162.005 -7.315 -161.675 ;
        RECT -7.645 -163.365 -7.315 -163.035 ;
        RECT -7.645 -164.725 -7.315 -164.395 ;
        RECT -7.645 -166.085 -7.315 -165.755 ;
        RECT -7.645 -167.445 -7.315 -167.115 ;
        RECT -7.645 -168.805 -7.315 -168.475 ;
        RECT -7.645 -170.165 -7.315 -169.835 ;
        RECT -7.645 -171.525 -7.315 -171.195 ;
        RECT -7.645 -172.885 -7.315 -172.555 ;
        RECT -7.645 -174.245 -7.315 -173.915 ;
        RECT -7.645 -175.605 -7.315 -175.275 ;
        RECT -7.645 -176.965 -7.315 -176.635 ;
        RECT -7.645 -178.325 -7.315 -177.995 ;
        RECT -7.645 -179.685 -7.315 -179.355 ;
        RECT -7.645 -181.93 -7.315 -180.8 ;
        RECT -7.64 -182.045 -7.32 -105.915 ;
        RECT -7.645 -106.245 -7.315 -105.915 ;
        RECT -7.645 -107.605 -7.315 -107.275 ;
        RECT -7.645 -108.965 -7.315 -108.635 ;
        RECT -7.645 -110.325 -7.315 -109.995 ;
        RECT -7.645 -111.685 -7.315 -111.355 ;
        RECT -7.645 -113.045 -7.315 -112.715 ;
        RECT -7.645 -114.405 -7.315 -114.075 ;
        RECT -7.645 -115.765 -7.315 -115.435 ;
        RECT -7.645 -117.125 -7.315 -116.795 ;
        RECT -7.645 -118.485 -7.315 -118.155 ;
        RECT -7.645 -119.845 -7.315 -119.515 ;
        RECT -7.645 -121.205 -7.315 -120.875 ;
        RECT -7.645 -123.925 -7.315 -123.595 ;
        RECT -7.645 -125.285 -7.315 -124.955 ;
        RECT -7.645 -126.645 -7.315 -126.315 ;
        RECT -7.645 -128.005 -7.315 -127.675 ;
        RECT -7.645 -129.365 -7.315 -129.035 ;
        RECT -7.645 -130.725 -7.315 -130.395 ;
        RECT -7.645 -132.085 -7.315 -131.755 ;
        RECT -7.645 -133.445 -7.315 -133.115 ;
        RECT -7.645 -134.805 -7.315 -134.475 ;
        RECT -7.645 -136.165 -7.315 -135.835 ;
        RECT -7.645 -137.525 -7.315 -137.195 ;
        RECT -7.645 -138.885 -7.315 -138.555 ;
        RECT -7.645 -140.245 -7.315 -139.915 ;
        RECT -7.645 -141.605 -7.315 -141.275 ;
        RECT -7.645 -142.965 -7.315 -142.635 ;
        RECT -7.645 -144.325 -7.315 -143.995 ;
        RECT -7.645 -145.685 -7.315 -145.355 ;
        RECT -7.645 -147.045 -7.315 -146.715 ;
        RECT -7.645 -148.405 -7.315 -148.075 ;
        RECT -7.645 -149.765 -7.315 -149.435 ;
        RECT -7.645 -151.125 -7.315 -150.795 ;
        RECT -7.645 -152.485 -7.315 -152.155 ;
        RECT -7.645 -153.845 -7.315 -153.515 ;
        RECT -7.645 -155.205 -7.315 -154.875 ;
        RECT -7.645 -156.565 -7.315 -156.235 ;
        RECT -7.645 -157.925 -7.315 -157.595 ;
        RECT -7.645 -159.285 -7.315 -158.955 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 -28.725 -19.555 -28.395 ;
        RECT -19.885 -30.085 -19.555 -29.755 ;
        RECT -19.885 -31.445 -19.555 -31.115 ;
        RECT -19.885 -32.805 -19.555 -32.475 ;
        RECT -19.885 -35.525 -19.555 -35.195 ;
        RECT -19.885 -36.885 -19.555 -36.555 ;
        RECT -19.885 -37.93 -19.555 -37.6 ;
        RECT -19.885 -40.965 -19.555 -40.635 ;
        RECT -19.885 -42.77 -19.555 -42.44 ;
        RECT -19.885 -43.685 -19.555 -43.355 ;
        RECT -19.885 -50.485 -19.555 -50.155 ;
        RECT -19.885 -51.845 -19.555 -51.515 ;
        RECT -19.885 -53.205 -19.555 -52.875 ;
        RECT -19.885 -54.565 -19.555 -54.235 ;
        RECT -19.885 -55.925 -19.555 -55.595 ;
        RECT -19.885 -57.285 -19.555 -56.955 ;
        RECT -19.885 -58.645 -19.555 -58.315 ;
        RECT -19.885 -60.005 -19.555 -59.675 ;
        RECT -19.885 -61.365 -19.555 -61.035 ;
        RECT -19.885 -62.725 -19.555 -62.395 ;
        RECT -19.885 -64.085 -19.555 -63.755 ;
        RECT -19.885 -65.445 -19.555 -65.115 ;
        RECT -19.885 -68.165 -19.555 -67.835 ;
        RECT -19.885 -69.525 -19.555 -69.195 ;
        RECT -19.885 -70.885 -19.555 -70.555 ;
        RECT -19.885 -72.245 -19.555 -71.915 ;
        RECT -19.885 -74.965 -19.555 -74.635 ;
        RECT -19.885 -76.71 -19.555 -76.38 ;
        RECT -19.885 -77.685 -19.555 -77.355 ;
        RECT -19.885 -79.045 -19.555 -78.715 ;
        RECT -19.885 -81.765 -19.555 -81.435 ;
        RECT -19.885 -83.125 -19.555 -82.795 ;
        RECT -19.885 -84.485 -19.555 -84.155 ;
        RECT -19.885 -85.25 -19.555 -84.92 ;
        RECT -19.885 -87.205 -19.555 -86.875 ;
        RECT -19.885 -89.925 -19.555 -89.595 ;
        RECT -19.885 -91.285 -19.555 -90.955 ;
        RECT -19.885 -92.645 -19.555 -92.315 ;
        RECT -19.885 -94.005 -19.555 -93.675 ;
        RECT -19.885 -96.725 -19.555 -96.395 ;
        RECT -19.885 -98.085 -19.555 -97.755 ;
        RECT -19.885 -98.89 -19.555 -98.56 ;
        RECT -19.885 -100.805 -19.555 -100.475 ;
        RECT -19.885 -102.165 -19.555 -101.835 ;
        RECT -19.885 -104.885 -19.555 -104.555 ;
        RECT -19.885 -107.43 -19.555 -107.1 ;
        RECT -19.88 -110.32 -19.56 -27.72 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 -117.125 -19.555 -116.795 ;
        RECT -19.885 -118.485 -19.555 -118.155 ;
        RECT -19.885 -125.285 -19.555 -124.955 ;
        RECT -19.885 -126.645 -19.555 -126.315 ;
        RECT -19.885 -128.005 -19.555 -127.675 ;
        RECT -19.885 -130.725 -19.555 -130.395 ;
        RECT -19.885 -141.605 -19.555 -141.275 ;
        RECT -19.885 -144.325 -19.555 -143.995 ;
        RECT -19.885 -145.685 -19.555 -145.355 ;
        RECT -19.885 -147.045 -19.555 -146.715 ;
        RECT -19.885 -148.405 -19.555 -148.075 ;
        RECT -19.885 -149.765 -19.555 -149.435 ;
        RECT -19.885 -153.845 -19.555 -153.515 ;
        RECT -19.885 -159.285 -19.555 -158.955 ;
        RECT -19.885 -160.645 -19.555 -160.315 ;
        RECT -19.885 -162.005 -19.555 -161.675 ;
        RECT -19.885 -163.365 -19.555 -163.035 ;
        RECT -19.885 -164.725 -19.555 -164.395 ;
        RECT -19.885 -166.085 -19.555 -165.755 ;
        RECT -19.885 -167.445 -19.555 -167.115 ;
        RECT -19.88 -167.445 -19.56 -115.44 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 -174.245 -19.555 -173.915 ;
        RECT -19.885 -175.605 -19.555 -175.275 ;
        RECT -19.885 -176.685 -19.555 -176.355 ;
        RECT -19.885 -178.325 -19.555 -177.995 ;
        RECT -19.885 -179.685 -19.555 -179.355 ;
        RECT -19.885 -181.93 -19.555 -180.8 ;
        RECT -19.88 -182.045 -19.56 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 241.32 -18.195 242.45 ;
        RECT -18.525 239.195 -18.195 239.525 ;
        RECT -18.525 237.835 -18.195 238.165 ;
        RECT -18.525 236.475 -18.195 236.805 ;
        RECT -18.525 235.115 -18.195 235.445 ;
        RECT -18.525 233.755 -18.195 234.085 ;
        RECT -18.525 232.395 -18.195 232.725 ;
        RECT -18.525 231.035 -18.195 231.365 ;
        RECT -18.525 229.675 -18.195 230.005 ;
        RECT -18.525 228.315 -18.195 228.645 ;
        RECT -18.525 226.955 -18.195 227.285 ;
        RECT -18.525 225.595 -18.195 225.925 ;
        RECT -18.525 224.235 -18.195 224.565 ;
        RECT -18.525 222.875 -18.195 223.205 ;
        RECT -18.525 221.515 -18.195 221.845 ;
        RECT -18.525 220.155 -18.195 220.485 ;
        RECT -18.525 218.795 -18.195 219.125 ;
        RECT -18.525 217.435 -18.195 217.765 ;
        RECT -18.525 216.075 -18.195 216.405 ;
        RECT -18.525 214.715 -18.195 215.045 ;
        RECT -18.525 213.355 -18.195 213.685 ;
        RECT -18.525 211.995 -18.195 212.325 ;
        RECT -18.525 210.635 -18.195 210.965 ;
        RECT -18.525 209.275 -18.195 209.605 ;
        RECT -18.525 207.915 -18.195 208.245 ;
        RECT -18.525 206.555 -18.195 206.885 ;
        RECT -18.525 205.195 -18.195 205.525 ;
        RECT -18.525 203.835 -18.195 204.165 ;
        RECT -18.525 202.475 -18.195 202.805 ;
        RECT -18.525 201.115 -18.195 201.445 ;
        RECT -18.525 199.755 -18.195 200.085 ;
        RECT -18.525 198.395 -18.195 198.725 ;
        RECT -18.525 197.035 -18.195 197.365 ;
        RECT -18.525 195.675 -18.195 196.005 ;
        RECT -18.525 194.315 -18.195 194.645 ;
        RECT -18.525 192.955 -18.195 193.285 ;
        RECT -18.525 191.595 -18.195 191.925 ;
        RECT -18.525 190.235 -18.195 190.565 ;
        RECT -18.525 188.875 -18.195 189.205 ;
        RECT -18.525 187.515 -18.195 187.845 ;
        RECT -18.525 186.155 -18.195 186.485 ;
        RECT -18.525 184.795 -18.195 185.125 ;
        RECT -18.525 183.435 -18.195 183.765 ;
        RECT -18.525 182.075 -18.195 182.405 ;
        RECT -18.525 180.715 -18.195 181.045 ;
        RECT -18.525 179.355 -18.195 179.685 ;
        RECT -18.525 177.995 -18.195 178.325 ;
        RECT -18.525 176.635 -18.195 176.965 ;
        RECT -18.525 175.275 -18.195 175.605 ;
        RECT -18.525 173.915 -18.195 174.245 ;
        RECT -18.525 172.555 -18.195 172.885 ;
        RECT -18.525 171.195 -18.195 171.525 ;
        RECT -18.525 169.835 -18.195 170.165 ;
        RECT -18.525 168.475 -18.195 168.805 ;
        RECT -18.525 167.115 -18.195 167.445 ;
        RECT -18.525 165.755 -18.195 166.085 ;
        RECT -18.525 164.395 -18.195 164.725 ;
        RECT -18.525 163.035 -18.195 163.365 ;
        RECT -18.525 161.675 -18.195 162.005 ;
        RECT -18.525 160.315 -18.195 160.645 ;
        RECT -18.525 158.955 -18.195 159.285 ;
        RECT -18.525 157.595 -18.195 157.925 ;
        RECT -18.525 156.235 -18.195 156.565 ;
        RECT -18.525 154.875 -18.195 155.205 ;
        RECT -18.525 153.515 -18.195 153.845 ;
        RECT -18.525 152.155 -18.195 152.485 ;
        RECT -18.525 150.795 -18.195 151.125 ;
        RECT -18.525 149.435 -18.195 149.765 ;
        RECT -18.525 148.075 -18.195 148.405 ;
        RECT -18.525 146.715 -18.195 147.045 ;
        RECT -18.525 145.355 -18.195 145.685 ;
        RECT -18.525 143.995 -18.195 144.325 ;
        RECT -18.525 142.635 -18.195 142.965 ;
        RECT -18.525 141.275 -18.195 141.605 ;
        RECT -18.525 139.915 -18.195 140.245 ;
        RECT -18.525 138.555 -18.195 138.885 ;
        RECT -18.525 137.195 -18.195 137.525 ;
        RECT -18.525 135.835 -18.195 136.165 ;
        RECT -18.525 134.475 -18.195 134.805 ;
        RECT -18.525 133.115 -18.195 133.445 ;
        RECT -18.525 131.755 -18.195 132.085 ;
        RECT -18.525 130.395 -18.195 130.725 ;
        RECT -18.525 129.035 -18.195 129.365 ;
        RECT -18.525 127.675 -18.195 128.005 ;
        RECT -18.525 126.315 -18.195 126.645 ;
        RECT -18.525 124.955 -18.195 125.285 ;
        RECT -18.525 123.595 -18.195 123.925 ;
        RECT -18.525 122.235 -18.195 122.565 ;
        RECT -18.525 120.875 -18.195 121.205 ;
        RECT -18.525 119.515 -18.195 119.845 ;
        RECT -18.525 118.155 -18.195 118.485 ;
        RECT -18.525 116.795 -18.195 117.125 ;
        RECT -18.525 115.435 -18.195 115.765 ;
        RECT -18.525 114.075 -18.195 114.405 ;
        RECT -18.525 112.715 -18.195 113.045 ;
        RECT -18.525 111.355 -18.195 111.685 ;
        RECT -18.525 109.995 -18.195 110.325 ;
        RECT -18.525 108.635 -18.195 108.965 ;
        RECT -18.525 107.275 -18.195 107.605 ;
        RECT -18.525 105.915 -18.195 106.245 ;
        RECT -18.525 104.555 -18.195 104.885 ;
        RECT -18.525 103.195 -18.195 103.525 ;
        RECT -18.525 101.835 -18.195 102.165 ;
        RECT -18.525 100.475 -18.195 100.805 ;
        RECT -18.525 99.115 -18.195 99.445 ;
        RECT -18.525 97.755 -18.195 98.085 ;
        RECT -18.525 96.395 -18.195 96.725 ;
        RECT -18.525 95.035 -18.195 95.365 ;
        RECT -18.525 93.675 -18.195 94.005 ;
        RECT -18.525 92.315 -18.195 92.645 ;
        RECT -18.525 90.955 -18.195 91.285 ;
        RECT -18.525 89.595 -18.195 89.925 ;
        RECT -18.525 88.235 -18.195 88.565 ;
        RECT -18.525 86.875 -18.195 87.205 ;
        RECT -18.525 85.515 -18.195 85.845 ;
        RECT -18.525 84.155 -18.195 84.485 ;
        RECT -18.525 82.795 -18.195 83.125 ;
        RECT -18.525 81.435 -18.195 81.765 ;
        RECT -18.525 80.075 -18.195 80.405 ;
        RECT -18.525 78.715 -18.195 79.045 ;
        RECT -18.525 77.355 -18.195 77.685 ;
        RECT -18.525 75.995 -18.195 76.325 ;
        RECT -18.525 74.635 -18.195 74.965 ;
        RECT -18.525 73.275 -18.195 73.605 ;
        RECT -18.525 71.915 -18.195 72.245 ;
        RECT -18.525 70.555 -18.195 70.885 ;
        RECT -18.525 69.195 -18.195 69.525 ;
        RECT -18.525 67.835 -18.195 68.165 ;
        RECT -18.525 66.475 -18.195 66.805 ;
        RECT -18.525 65.115 -18.195 65.445 ;
        RECT -18.525 63.755 -18.195 64.085 ;
        RECT -18.525 62.395 -18.195 62.725 ;
        RECT -18.525 61.035 -18.195 61.365 ;
        RECT -18.525 59.675 -18.195 60.005 ;
        RECT -18.525 58.315 -18.195 58.645 ;
        RECT -18.525 56.955 -18.195 57.285 ;
        RECT -18.525 55.595 -18.195 55.925 ;
        RECT -18.525 54.235 -18.195 54.565 ;
        RECT -18.525 52.875 -18.195 53.205 ;
        RECT -18.525 51.515 -18.195 51.845 ;
        RECT -18.525 50.155 -18.195 50.485 ;
        RECT -18.525 48.795 -18.195 49.125 ;
        RECT -18.525 47.435 -18.195 47.765 ;
        RECT -18.525 46.075 -18.195 46.405 ;
        RECT -18.525 44.715 -18.195 45.045 ;
        RECT -18.525 43.355 -18.195 43.685 ;
        RECT -18.525 41.995 -18.195 42.325 ;
        RECT -18.525 40.635 -18.195 40.965 ;
        RECT -18.525 39.275 -18.195 39.605 ;
        RECT -18.525 37.915 -18.195 38.245 ;
        RECT -18.525 36.555 -18.195 36.885 ;
        RECT -18.525 35.195 -18.195 35.525 ;
        RECT -18.525 33.835 -18.195 34.165 ;
        RECT -18.525 32.475 -18.195 32.805 ;
        RECT -18.525 31.115 -18.195 31.445 ;
        RECT -18.525 29.755 -18.195 30.085 ;
        RECT -18.525 28.395 -18.195 28.725 ;
        RECT -18.525 27.035 -18.195 27.365 ;
        RECT -18.525 25.675 -18.195 26.005 ;
        RECT -18.525 24.315 -18.195 24.645 ;
        RECT -18.525 22.955 -18.195 23.285 ;
        RECT -18.525 21.595 -18.195 21.925 ;
        RECT -18.525 20.235 -18.195 20.565 ;
        RECT -18.525 18.875 -18.195 19.205 ;
        RECT -18.525 17.515 -18.195 17.845 ;
        RECT -18.525 16.155 -18.195 16.485 ;
        RECT -18.525 14.795 -18.195 15.125 ;
        RECT -18.525 13.435 -18.195 13.765 ;
        RECT -18.525 12.075 -18.195 12.405 ;
        RECT -18.525 10.715 -18.195 11.045 ;
        RECT -18.525 9.355 -18.195 9.685 ;
        RECT -18.525 7.995 -18.195 8.325 ;
        RECT -18.525 6.635 -18.195 6.965 ;
        RECT -18.525 5.275 -18.195 5.605 ;
        RECT -18.525 3.915 -18.195 4.245 ;
        RECT -18.525 2.555 -18.195 2.885 ;
        RECT -18.525 1.195 -18.195 1.525 ;
        RECT -18.525 -0.165 -18.195 0.165 ;
        RECT -18.525 -2.885 -18.195 -2.555 ;
        RECT -18.525 -4.245 -18.195 -3.915 ;
        RECT -18.525 -8.325 -18.195 -7.995 ;
        RECT -18.525 -9.685 -18.195 -9.355 ;
        RECT -18.525 -14.95 -18.195 -14.62 ;
        RECT -18.525 -17.845 -18.195 -17.515 ;
        RECT -18.525 -19.79 -18.195 -19.46 ;
        RECT -18.525 -20.565 -18.195 -20.235 ;
        RECT -18.52 -21.24 -18.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 -27.365 -18.195 -27.035 ;
        RECT -18.525 -28.725 -18.195 -28.395 ;
        RECT -18.525 -30.085 -18.195 -29.755 ;
        RECT -18.525 -31.445 -18.195 -31.115 ;
        RECT -18.525 -32.805 -18.195 -32.475 ;
        RECT -18.525 -35.525 -18.195 -35.195 ;
        RECT -18.525 -36.885 -18.195 -36.555 ;
        RECT -18.525 -37.93 -18.195 -37.6 ;
        RECT -18.525 -40.965 -18.195 -40.635 ;
        RECT -18.525 -42.77 -18.195 -42.44 ;
        RECT -18.525 -43.685 -18.195 -43.355 ;
        RECT -18.525 -50.485 -18.195 -50.155 ;
        RECT -18.525 -51.845 -18.195 -51.515 ;
        RECT -18.525 -53.205 -18.195 -52.875 ;
        RECT -18.525 -54.565 -18.195 -54.235 ;
        RECT -18.525 -55.925 -18.195 -55.595 ;
        RECT -18.525 -57.285 -18.195 -56.955 ;
        RECT -18.525 -58.645 -18.195 -58.315 ;
        RECT -18.525 -60.005 -18.195 -59.675 ;
        RECT -18.525 -61.365 -18.195 -61.035 ;
        RECT -18.525 -62.725 -18.195 -62.395 ;
        RECT -18.525 -64.085 -18.195 -63.755 ;
        RECT -18.525 -65.445 -18.195 -65.115 ;
        RECT -18.525 -68.165 -18.195 -67.835 ;
        RECT -18.525 -69.525 -18.195 -69.195 ;
        RECT -18.525 -70.885 -18.195 -70.555 ;
        RECT -18.525 -72.245 -18.195 -71.915 ;
        RECT -18.525 -74.965 -18.195 -74.635 ;
        RECT -18.525 -76.71 -18.195 -76.38 ;
        RECT -18.525 -77.685 -18.195 -77.355 ;
        RECT -18.525 -79.045 -18.195 -78.715 ;
        RECT -18.525 -81.765 -18.195 -81.435 ;
        RECT -18.525 -83.125 -18.195 -82.795 ;
        RECT -18.525 -84.485 -18.195 -84.155 ;
        RECT -18.525 -85.25 -18.195 -84.92 ;
        RECT -18.525 -87.205 -18.195 -86.875 ;
        RECT -18.525 -89.925 -18.195 -89.595 ;
        RECT -18.525 -91.285 -18.195 -90.955 ;
        RECT -18.525 -92.645 -18.195 -92.315 ;
        RECT -18.525 -94.005 -18.195 -93.675 ;
        RECT -18.525 -96.725 -18.195 -96.395 ;
        RECT -18.525 -98.085 -18.195 -97.755 ;
        RECT -18.525 -98.89 -18.195 -98.56 ;
        RECT -18.525 -100.805 -18.195 -100.475 ;
        RECT -18.525 -102.165 -18.195 -101.835 ;
        RECT -18.525 -107.43 -18.195 -107.1 ;
        RECT -18.52 -108.96 -18.2 -26.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -18.525 -114.405 -18.195 -114.075 ;
        RECT -18.525 -115.765 -18.195 -115.435 ;
        RECT -18.525 -117.125 -18.195 -116.795 ;
        RECT -18.525 -118.485 -18.195 -118.155 ;
        RECT -18.525 -126.645 -18.195 -126.315 ;
        RECT -18.525 -128.005 -18.195 -127.675 ;
        RECT -18.525 -141.605 -18.195 -141.275 ;
        RECT -18.525 -144.325 -18.195 -143.995 ;
        RECT -18.525 -148.405 -18.195 -148.075 ;
        RECT -18.525 -153.845 -18.195 -153.515 ;
        RECT -18.525 -159.285 -18.195 -158.955 ;
        RECT -18.525 -160.645 -18.195 -160.315 ;
        RECT -18.525 -162.005 -18.195 -161.675 ;
        RECT -18.525 -163.365 -18.195 -163.035 ;
        RECT -18.525 -164.725 -18.195 -164.395 ;
        RECT -18.525 -166.085 -18.195 -165.755 ;
        RECT -18.525 -167.445 -18.195 -167.115 ;
        RECT -18.525 -168.805 -18.195 -168.475 ;
        RECT -18.525 -171.525 -18.195 -171.195 ;
        RECT -18.525 -174.245 -18.195 -173.915 ;
        RECT -18.525 -175.605 -18.195 -175.275 ;
        RECT -18.525 -176.685 -18.195 -176.355 ;
        RECT -18.525 -178.325 -18.195 -177.995 ;
        RECT -18.525 -179.685 -18.195 -179.355 ;
        RECT -18.525 -181.93 -18.195 -180.8 ;
        RECT -18.52 -182.045 -18.2 -114.075 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 241.32 -16.835 242.45 ;
        RECT -17.165 239.195 -16.835 239.525 ;
        RECT -17.165 237.835 -16.835 238.165 ;
        RECT -17.165 236.475 -16.835 236.805 ;
        RECT -17.165 235.115 -16.835 235.445 ;
        RECT -17.165 233.755 -16.835 234.085 ;
        RECT -17.165 232.395 -16.835 232.725 ;
        RECT -17.165 231.035 -16.835 231.365 ;
        RECT -17.165 229.675 -16.835 230.005 ;
        RECT -17.165 228.315 -16.835 228.645 ;
        RECT -17.165 226.955 -16.835 227.285 ;
        RECT -17.165 225.595 -16.835 225.925 ;
        RECT -17.165 224.235 -16.835 224.565 ;
        RECT -17.165 222.875 -16.835 223.205 ;
        RECT -17.165 221.515 -16.835 221.845 ;
        RECT -17.165 220.155 -16.835 220.485 ;
        RECT -17.165 218.795 -16.835 219.125 ;
        RECT -17.165 217.435 -16.835 217.765 ;
        RECT -17.165 216.075 -16.835 216.405 ;
        RECT -17.165 214.715 -16.835 215.045 ;
        RECT -17.165 213.355 -16.835 213.685 ;
        RECT -17.165 211.995 -16.835 212.325 ;
        RECT -17.165 210.635 -16.835 210.965 ;
        RECT -17.165 209.275 -16.835 209.605 ;
        RECT -17.165 207.915 -16.835 208.245 ;
        RECT -17.165 206.555 -16.835 206.885 ;
        RECT -17.165 205.195 -16.835 205.525 ;
        RECT -17.165 203.835 -16.835 204.165 ;
        RECT -17.165 202.475 -16.835 202.805 ;
        RECT -17.165 201.115 -16.835 201.445 ;
        RECT -17.165 199.755 -16.835 200.085 ;
        RECT -17.165 198.395 -16.835 198.725 ;
        RECT -17.165 197.035 -16.835 197.365 ;
        RECT -17.165 195.675 -16.835 196.005 ;
        RECT -17.165 194.315 -16.835 194.645 ;
        RECT -17.165 192.955 -16.835 193.285 ;
        RECT -17.165 191.595 -16.835 191.925 ;
        RECT -17.165 190.235 -16.835 190.565 ;
        RECT -17.165 188.875 -16.835 189.205 ;
        RECT -17.165 187.515 -16.835 187.845 ;
        RECT -17.165 186.155 -16.835 186.485 ;
        RECT -17.165 184.795 -16.835 185.125 ;
        RECT -17.165 183.435 -16.835 183.765 ;
        RECT -17.165 182.075 -16.835 182.405 ;
        RECT -17.165 180.715 -16.835 181.045 ;
        RECT -17.165 179.355 -16.835 179.685 ;
        RECT -17.165 177.995 -16.835 178.325 ;
        RECT -17.165 176.635 -16.835 176.965 ;
        RECT -17.165 175.275 -16.835 175.605 ;
        RECT -17.165 173.915 -16.835 174.245 ;
        RECT -17.165 172.555 -16.835 172.885 ;
        RECT -17.165 171.195 -16.835 171.525 ;
        RECT -17.165 169.835 -16.835 170.165 ;
        RECT -17.165 168.475 -16.835 168.805 ;
        RECT -17.165 167.115 -16.835 167.445 ;
        RECT -17.165 165.755 -16.835 166.085 ;
        RECT -17.165 164.395 -16.835 164.725 ;
        RECT -17.165 163.035 -16.835 163.365 ;
        RECT -17.165 161.675 -16.835 162.005 ;
        RECT -17.165 160.315 -16.835 160.645 ;
        RECT -17.165 158.955 -16.835 159.285 ;
        RECT -17.165 157.595 -16.835 157.925 ;
        RECT -17.165 156.235 -16.835 156.565 ;
        RECT -17.165 154.875 -16.835 155.205 ;
        RECT -17.165 153.515 -16.835 153.845 ;
        RECT -17.165 152.155 -16.835 152.485 ;
        RECT -17.165 150.795 -16.835 151.125 ;
        RECT -17.165 149.435 -16.835 149.765 ;
        RECT -17.165 148.075 -16.835 148.405 ;
        RECT -17.165 146.715 -16.835 147.045 ;
        RECT -17.165 145.355 -16.835 145.685 ;
        RECT -17.165 143.995 -16.835 144.325 ;
        RECT -17.165 142.635 -16.835 142.965 ;
        RECT -17.165 141.275 -16.835 141.605 ;
        RECT -17.165 139.915 -16.835 140.245 ;
        RECT -17.165 138.555 -16.835 138.885 ;
        RECT -17.165 137.195 -16.835 137.525 ;
        RECT -17.165 135.835 -16.835 136.165 ;
        RECT -17.165 134.475 -16.835 134.805 ;
        RECT -17.165 133.115 -16.835 133.445 ;
        RECT -17.165 131.755 -16.835 132.085 ;
        RECT -17.165 130.395 -16.835 130.725 ;
        RECT -17.165 129.035 -16.835 129.365 ;
        RECT -17.165 127.675 -16.835 128.005 ;
        RECT -17.165 126.315 -16.835 126.645 ;
        RECT -17.165 124.955 -16.835 125.285 ;
        RECT -17.165 123.595 -16.835 123.925 ;
        RECT -17.165 122.235 -16.835 122.565 ;
        RECT -17.165 120.875 -16.835 121.205 ;
        RECT -17.165 119.515 -16.835 119.845 ;
        RECT -17.165 118.155 -16.835 118.485 ;
        RECT -17.165 116.795 -16.835 117.125 ;
        RECT -17.165 115.435 -16.835 115.765 ;
        RECT -17.165 114.075 -16.835 114.405 ;
        RECT -17.165 112.715 -16.835 113.045 ;
        RECT -17.165 111.355 -16.835 111.685 ;
        RECT -17.165 109.995 -16.835 110.325 ;
        RECT -17.165 108.635 -16.835 108.965 ;
        RECT -17.165 107.275 -16.835 107.605 ;
        RECT -17.165 105.915 -16.835 106.245 ;
        RECT -17.165 104.555 -16.835 104.885 ;
        RECT -17.165 103.195 -16.835 103.525 ;
        RECT -17.165 101.835 -16.835 102.165 ;
        RECT -17.165 100.475 -16.835 100.805 ;
        RECT -17.165 99.115 -16.835 99.445 ;
        RECT -17.165 97.755 -16.835 98.085 ;
        RECT -17.165 96.395 -16.835 96.725 ;
        RECT -17.165 95.035 -16.835 95.365 ;
        RECT -17.165 93.675 -16.835 94.005 ;
        RECT -17.165 92.315 -16.835 92.645 ;
        RECT -17.165 90.955 -16.835 91.285 ;
        RECT -17.165 89.595 -16.835 89.925 ;
        RECT -17.165 88.235 -16.835 88.565 ;
        RECT -17.165 86.875 -16.835 87.205 ;
        RECT -17.165 85.515 -16.835 85.845 ;
        RECT -17.165 84.155 -16.835 84.485 ;
        RECT -17.165 82.795 -16.835 83.125 ;
        RECT -17.165 81.435 -16.835 81.765 ;
        RECT -17.165 80.075 -16.835 80.405 ;
        RECT -17.165 78.715 -16.835 79.045 ;
        RECT -17.165 77.355 -16.835 77.685 ;
        RECT -17.165 75.995 -16.835 76.325 ;
        RECT -17.165 74.635 -16.835 74.965 ;
        RECT -17.165 73.275 -16.835 73.605 ;
        RECT -17.165 71.915 -16.835 72.245 ;
        RECT -17.165 70.555 -16.835 70.885 ;
        RECT -17.165 69.195 -16.835 69.525 ;
        RECT -17.165 67.835 -16.835 68.165 ;
        RECT -17.165 66.475 -16.835 66.805 ;
        RECT -17.165 65.115 -16.835 65.445 ;
        RECT -17.165 63.755 -16.835 64.085 ;
        RECT -17.165 62.395 -16.835 62.725 ;
        RECT -17.165 61.035 -16.835 61.365 ;
        RECT -17.165 59.675 -16.835 60.005 ;
        RECT -17.165 58.315 -16.835 58.645 ;
        RECT -17.165 56.955 -16.835 57.285 ;
        RECT -17.165 55.595 -16.835 55.925 ;
        RECT -17.165 54.235 -16.835 54.565 ;
        RECT -17.165 52.875 -16.835 53.205 ;
        RECT -17.165 51.515 -16.835 51.845 ;
        RECT -17.165 50.155 -16.835 50.485 ;
        RECT -17.165 48.795 -16.835 49.125 ;
        RECT -17.165 47.435 -16.835 47.765 ;
        RECT -17.165 46.075 -16.835 46.405 ;
        RECT -17.165 44.715 -16.835 45.045 ;
        RECT -17.165 43.355 -16.835 43.685 ;
        RECT -17.165 41.995 -16.835 42.325 ;
        RECT -17.165 40.635 -16.835 40.965 ;
        RECT -17.165 39.275 -16.835 39.605 ;
        RECT -17.165 37.915 -16.835 38.245 ;
        RECT -17.165 36.555 -16.835 36.885 ;
        RECT -17.165 35.195 -16.835 35.525 ;
        RECT -17.165 33.835 -16.835 34.165 ;
        RECT -17.165 32.475 -16.835 32.805 ;
        RECT -17.165 31.115 -16.835 31.445 ;
        RECT -17.165 29.755 -16.835 30.085 ;
        RECT -17.165 28.395 -16.835 28.725 ;
        RECT -17.165 27.035 -16.835 27.365 ;
        RECT -17.165 25.675 -16.835 26.005 ;
        RECT -17.165 24.315 -16.835 24.645 ;
        RECT -17.165 22.955 -16.835 23.285 ;
        RECT -17.165 21.595 -16.835 21.925 ;
        RECT -17.165 20.235 -16.835 20.565 ;
        RECT -17.165 18.875 -16.835 19.205 ;
        RECT -17.165 17.515 -16.835 17.845 ;
        RECT -17.165 16.155 -16.835 16.485 ;
        RECT -17.165 14.795 -16.835 15.125 ;
        RECT -17.165 13.435 -16.835 13.765 ;
        RECT -17.165 12.075 -16.835 12.405 ;
        RECT -17.165 10.715 -16.835 11.045 ;
        RECT -17.165 9.355 -16.835 9.685 ;
        RECT -17.165 7.995 -16.835 8.325 ;
        RECT -17.165 6.635 -16.835 6.965 ;
        RECT -17.165 5.275 -16.835 5.605 ;
        RECT -17.165 3.915 -16.835 4.245 ;
        RECT -17.165 2.555 -16.835 2.885 ;
        RECT -17.165 1.195 -16.835 1.525 ;
        RECT -17.165 -0.165 -16.835 0.165 ;
        RECT -17.165 -2.885 -16.835 -2.555 ;
        RECT -17.165 -4.245 -16.835 -3.915 ;
        RECT -17.165 -8.325 -16.835 -7.995 ;
        RECT -17.165 -9.685 -16.835 -9.355 ;
        RECT -17.165 -12.405 -16.835 -12.075 ;
        RECT -17.16 -12.405 -16.84 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 -27.365 -16.835 -27.035 ;
        RECT -17.165 -28.725 -16.835 -28.395 ;
        RECT -17.165 -30.085 -16.835 -29.755 ;
        RECT -17.165 -31.445 -16.835 -31.115 ;
        RECT -17.165 -32.805 -16.835 -32.475 ;
        RECT -17.165 -35.525 -16.835 -35.195 ;
        RECT -17.165 -36.885 -16.835 -36.555 ;
        RECT -17.165 -37.93 -16.835 -37.6 ;
        RECT -17.165 -42.77 -16.835 -42.44 ;
        RECT -17.165 -43.685 -16.835 -43.355 ;
        RECT -17.165 -51.845 -16.835 -51.515 ;
        RECT -17.165 -53.205 -16.835 -52.875 ;
        RECT -17.165 -54.565 -16.835 -54.235 ;
        RECT -17.165 -55.925 -16.835 -55.595 ;
        RECT -17.165 -57.285 -16.835 -56.955 ;
        RECT -17.165 -58.645 -16.835 -58.315 ;
        RECT -17.165 -60.005 -16.835 -59.675 ;
        RECT -17.165 -61.365 -16.835 -61.035 ;
        RECT -17.165 -62.725 -16.835 -62.395 ;
        RECT -17.165 -64.085 -16.835 -63.755 ;
        RECT -17.165 -65.445 -16.835 -65.115 ;
        RECT -17.165 -68.165 -16.835 -67.835 ;
        RECT -17.165 -69.525 -16.835 -69.195 ;
        RECT -17.165 -70.885 -16.835 -70.555 ;
        RECT -17.165 -72.245 -16.835 -71.915 ;
        RECT -17.165 -74.965 -16.835 -74.635 ;
        RECT -17.165 -76.71 -16.835 -76.38 ;
        RECT -17.165 -77.685 -16.835 -77.355 ;
        RECT -17.165 -79.045 -16.835 -78.715 ;
        RECT -17.165 -81.765 -16.835 -81.435 ;
        RECT -17.165 -83.125 -16.835 -82.795 ;
        RECT -17.165 -84.485 -16.835 -84.155 ;
        RECT -17.165 -85.25 -16.835 -84.92 ;
        RECT -17.165 -87.205 -16.835 -86.875 ;
        RECT -17.165 -89.925 -16.835 -89.595 ;
        RECT -17.165 -91.285 -16.835 -90.955 ;
        RECT -17.165 -92.645 -16.835 -92.315 ;
        RECT -17.165 -94.005 -16.835 -93.675 ;
        RECT -17.165 -96.725 -16.835 -96.395 ;
        RECT -17.165 -98.085 -16.835 -97.755 ;
        RECT -17.165 -98.89 -16.835 -98.56 ;
        RECT -17.165 -100.805 -16.835 -100.475 ;
        RECT -17.165 -102.165 -16.835 -101.835 ;
        RECT -17.165 -107.43 -16.835 -107.1 ;
        RECT -17.165 -114.405 -16.835 -114.075 ;
        RECT -17.165 -115.765 -16.835 -115.435 ;
        RECT -17.16 -115.765 -16.84 -26.36 ;
    END
    PORT
      LAYER met3 ;
        RECT -17.165 -175.605 -16.835 -175.275 ;
        RECT -17.165 -176.685 -16.835 -176.355 ;
        RECT -17.165 -178.325 -16.835 -177.995 ;
        RECT -17.165 -179.685 -16.835 -179.355 ;
        RECT -17.165 -181.93 -16.835 -180.8 ;
        RECT -17.16 -182.045 -16.84 -175.275 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 241.32 -15.475 242.45 ;
        RECT -15.805 239.195 -15.475 239.525 ;
        RECT -15.805 237.835 -15.475 238.165 ;
        RECT -15.805 236.475 -15.475 236.805 ;
        RECT -15.805 235.115 -15.475 235.445 ;
        RECT -15.805 233.755 -15.475 234.085 ;
        RECT -15.805 232.395 -15.475 232.725 ;
        RECT -15.805 231.035 -15.475 231.365 ;
        RECT -15.805 229.675 -15.475 230.005 ;
        RECT -15.805 228.315 -15.475 228.645 ;
        RECT -15.805 226.955 -15.475 227.285 ;
        RECT -15.805 225.595 -15.475 225.925 ;
        RECT -15.805 224.235 -15.475 224.565 ;
        RECT -15.805 222.875 -15.475 223.205 ;
        RECT -15.805 221.515 -15.475 221.845 ;
        RECT -15.805 220.155 -15.475 220.485 ;
        RECT -15.805 218.795 -15.475 219.125 ;
        RECT -15.805 217.435 -15.475 217.765 ;
        RECT -15.805 216.075 -15.475 216.405 ;
        RECT -15.805 214.715 -15.475 215.045 ;
        RECT -15.805 213.355 -15.475 213.685 ;
        RECT -15.805 211.995 -15.475 212.325 ;
        RECT -15.805 210.635 -15.475 210.965 ;
        RECT -15.805 209.275 -15.475 209.605 ;
        RECT -15.805 207.915 -15.475 208.245 ;
        RECT -15.805 206.555 -15.475 206.885 ;
        RECT -15.805 205.195 -15.475 205.525 ;
        RECT -15.805 203.835 -15.475 204.165 ;
        RECT -15.805 202.475 -15.475 202.805 ;
        RECT -15.805 201.115 -15.475 201.445 ;
        RECT -15.805 199.755 -15.475 200.085 ;
        RECT -15.805 198.395 -15.475 198.725 ;
        RECT -15.805 197.035 -15.475 197.365 ;
        RECT -15.805 195.675 -15.475 196.005 ;
        RECT -15.805 194.315 -15.475 194.645 ;
        RECT -15.805 192.955 -15.475 193.285 ;
        RECT -15.805 191.595 -15.475 191.925 ;
        RECT -15.805 190.235 -15.475 190.565 ;
        RECT -15.805 188.875 -15.475 189.205 ;
        RECT -15.805 187.515 -15.475 187.845 ;
        RECT -15.805 186.155 -15.475 186.485 ;
        RECT -15.805 184.795 -15.475 185.125 ;
        RECT -15.805 183.435 -15.475 183.765 ;
        RECT -15.805 182.075 -15.475 182.405 ;
        RECT -15.805 180.715 -15.475 181.045 ;
        RECT -15.805 179.355 -15.475 179.685 ;
        RECT -15.805 177.995 -15.475 178.325 ;
        RECT -15.805 176.635 -15.475 176.965 ;
        RECT -15.805 175.275 -15.475 175.605 ;
        RECT -15.805 173.915 -15.475 174.245 ;
        RECT -15.805 172.555 -15.475 172.885 ;
        RECT -15.805 171.195 -15.475 171.525 ;
        RECT -15.805 169.835 -15.475 170.165 ;
        RECT -15.805 168.475 -15.475 168.805 ;
        RECT -15.805 167.115 -15.475 167.445 ;
        RECT -15.805 165.755 -15.475 166.085 ;
        RECT -15.805 164.395 -15.475 164.725 ;
        RECT -15.805 163.035 -15.475 163.365 ;
        RECT -15.805 161.675 -15.475 162.005 ;
        RECT -15.805 160.315 -15.475 160.645 ;
        RECT -15.805 158.955 -15.475 159.285 ;
        RECT -15.805 157.595 -15.475 157.925 ;
        RECT -15.805 156.235 -15.475 156.565 ;
        RECT -15.805 154.875 -15.475 155.205 ;
        RECT -15.805 153.515 -15.475 153.845 ;
        RECT -15.805 152.155 -15.475 152.485 ;
        RECT -15.805 150.795 -15.475 151.125 ;
        RECT -15.805 149.435 -15.475 149.765 ;
        RECT -15.805 148.075 -15.475 148.405 ;
        RECT -15.805 146.715 -15.475 147.045 ;
        RECT -15.805 145.355 -15.475 145.685 ;
        RECT -15.805 143.995 -15.475 144.325 ;
        RECT -15.805 142.635 -15.475 142.965 ;
        RECT -15.805 141.275 -15.475 141.605 ;
        RECT -15.805 139.915 -15.475 140.245 ;
        RECT -15.805 138.555 -15.475 138.885 ;
        RECT -15.805 137.195 -15.475 137.525 ;
        RECT -15.805 135.835 -15.475 136.165 ;
        RECT -15.805 134.475 -15.475 134.805 ;
        RECT -15.805 133.115 -15.475 133.445 ;
        RECT -15.805 131.755 -15.475 132.085 ;
        RECT -15.805 130.395 -15.475 130.725 ;
        RECT -15.805 129.035 -15.475 129.365 ;
        RECT -15.805 127.675 -15.475 128.005 ;
        RECT -15.805 126.315 -15.475 126.645 ;
        RECT -15.805 124.955 -15.475 125.285 ;
        RECT -15.805 123.595 -15.475 123.925 ;
        RECT -15.805 122.235 -15.475 122.565 ;
        RECT -15.805 120.875 -15.475 121.205 ;
        RECT -15.805 119.515 -15.475 119.845 ;
        RECT -15.805 118.155 -15.475 118.485 ;
        RECT -15.805 116.795 -15.475 117.125 ;
        RECT -15.805 115.435 -15.475 115.765 ;
        RECT -15.805 114.075 -15.475 114.405 ;
        RECT -15.805 112.715 -15.475 113.045 ;
        RECT -15.805 111.355 -15.475 111.685 ;
        RECT -15.805 109.995 -15.475 110.325 ;
        RECT -15.805 108.635 -15.475 108.965 ;
        RECT -15.805 107.275 -15.475 107.605 ;
        RECT -15.805 105.915 -15.475 106.245 ;
        RECT -15.805 104.555 -15.475 104.885 ;
        RECT -15.805 103.195 -15.475 103.525 ;
        RECT -15.805 101.835 -15.475 102.165 ;
        RECT -15.805 100.475 -15.475 100.805 ;
        RECT -15.805 99.115 -15.475 99.445 ;
        RECT -15.805 97.755 -15.475 98.085 ;
        RECT -15.805 96.395 -15.475 96.725 ;
        RECT -15.805 95.035 -15.475 95.365 ;
        RECT -15.805 93.675 -15.475 94.005 ;
        RECT -15.805 92.315 -15.475 92.645 ;
        RECT -15.805 90.955 -15.475 91.285 ;
        RECT -15.805 89.595 -15.475 89.925 ;
        RECT -15.805 88.235 -15.475 88.565 ;
        RECT -15.805 86.875 -15.475 87.205 ;
        RECT -15.805 85.515 -15.475 85.845 ;
        RECT -15.805 84.155 -15.475 84.485 ;
        RECT -15.805 82.795 -15.475 83.125 ;
        RECT -15.805 81.435 -15.475 81.765 ;
        RECT -15.805 80.075 -15.475 80.405 ;
        RECT -15.805 78.715 -15.475 79.045 ;
        RECT -15.805 77.355 -15.475 77.685 ;
        RECT -15.805 75.995 -15.475 76.325 ;
        RECT -15.805 74.635 -15.475 74.965 ;
        RECT -15.805 73.275 -15.475 73.605 ;
        RECT -15.805 71.915 -15.475 72.245 ;
        RECT -15.805 70.555 -15.475 70.885 ;
        RECT -15.805 69.195 -15.475 69.525 ;
        RECT -15.805 67.835 -15.475 68.165 ;
        RECT -15.805 66.475 -15.475 66.805 ;
        RECT -15.805 65.115 -15.475 65.445 ;
        RECT -15.805 63.755 -15.475 64.085 ;
        RECT -15.805 62.395 -15.475 62.725 ;
        RECT -15.805 61.035 -15.475 61.365 ;
        RECT -15.805 59.675 -15.475 60.005 ;
        RECT -15.805 58.315 -15.475 58.645 ;
        RECT -15.805 56.955 -15.475 57.285 ;
        RECT -15.805 55.595 -15.475 55.925 ;
        RECT -15.805 54.235 -15.475 54.565 ;
        RECT -15.805 52.875 -15.475 53.205 ;
        RECT -15.805 51.515 -15.475 51.845 ;
        RECT -15.805 50.155 -15.475 50.485 ;
        RECT -15.805 48.795 -15.475 49.125 ;
        RECT -15.805 47.435 -15.475 47.765 ;
        RECT -15.805 46.075 -15.475 46.405 ;
        RECT -15.805 44.715 -15.475 45.045 ;
        RECT -15.805 43.355 -15.475 43.685 ;
        RECT -15.805 41.995 -15.475 42.325 ;
        RECT -15.805 40.635 -15.475 40.965 ;
        RECT -15.805 39.275 -15.475 39.605 ;
        RECT -15.805 37.915 -15.475 38.245 ;
        RECT -15.805 36.555 -15.475 36.885 ;
        RECT -15.805 35.195 -15.475 35.525 ;
        RECT -15.805 33.835 -15.475 34.165 ;
        RECT -15.805 32.475 -15.475 32.805 ;
        RECT -15.805 31.115 -15.475 31.445 ;
        RECT -15.805 29.755 -15.475 30.085 ;
        RECT -15.805 28.395 -15.475 28.725 ;
        RECT -15.805 27.035 -15.475 27.365 ;
        RECT -15.805 25.675 -15.475 26.005 ;
        RECT -15.805 24.315 -15.475 24.645 ;
        RECT -15.805 22.955 -15.475 23.285 ;
        RECT -15.805 21.595 -15.475 21.925 ;
        RECT -15.805 20.235 -15.475 20.565 ;
        RECT -15.805 18.875 -15.475 19.205 ;
        RECT -15.805 17.515 -15.475 17.845 ;
        RECT -15.805 16.155 -15.475 16.485 ;
        RECT -15.805 14.795 -15.475 15.125 ;
        RECT -15.805 13.435 -15.475 13.765 ;
        RECT -15.805 12.075 -15.475 12.405 ;
        RECT -15.805 10.715 -15.475 11.045 ;
        RECT -15.805 9.355 -15.475 9.685 ;
        RECT -15.805 7.995 -15.475 8.325 ;
        RECT -15.805 6.635 -15.475 6.965 ;
        RECT -15.805 5.275 -15.475 5.605 ;
        RECT -15.805 3.915 -15.475 4.245 ;
        RECT -15.805 2.555 -15.475 2.885 ;
        RECT -15.805 1.195 -15.475 1.525 ;
        RECT -15.805 -0.165 -15.475 0.165 ;
        RECT -15.805 -2.885 -15.475 -2.555 ;
        RECT -15.805 -4.245 -15.475 -3.915 ;
        RECT -15.805 -5.605 -15.475 -5.275 ;
        RECT -15.805 -8.325 -15.475 -7.995 ;
        RECT -15.805 -9.685 -15.475 -9.355 ;
        RECT -15.805 -12.405 -15.475 -12.075 ;
        RECT -15.805 -13.765 -15.475 -13.435 ;
        RECT -15.805 -14.95 -15.475 -14.62 ;
        RECT -15.805 -17.845 -15.475 -17.515 ;
        RECT -15.805 -19.79 -15.475 -19.46 ;
        RECT -15.805 -20.565 -15.475 -20.235 ;
        RECT -15.8 -20.565 -15.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -15.805 -107.43 -15.475 -107.1 ;
        RECT -15.805 -114.405 -15.475 -114.075 ;
        RECT -15.805 -115.765 -15.475 -115.435 ;
        RECT -15.805 -117.125 -15.475 -116.795 ;
        RECT -15.805 -118.485 -15.475 -118.155 ;
        RECT -15.805 -122.565 -15.475 -122.235 ;
        RECT -15.805 -128.005 -15.475 -127.675 ;
        RECT -15.805 -137.525 -15.475 -137.195 ;
        RECT -15.805 -141.605 -15.475 -141.275 ;
        RECT -15.805 -144.325 -15.475 -143.995 ;
        RECT -15.805 -159.285 -15.475 -158.955 ;
        RECT -15.805 -160.645 -15.475 -160.315 ;
        RECT -15.805 -162.005 -15.475 -161.675 ;
        RECT -15.805 -163.365 -15.475 -163.035 ;
        RECT -15.805 -164.725 -15.475 -164.395 ;
        RECT -15.805 -166.085 -15.475 -165.755 ;
        RECT -15.805 -167.445 -15.475 -167.115 ;
        RECT -15.805 -171.525 -15.475 -171.195 ;
        RECT -15.805 -172.885 -15.475 -172.555 ;
        RECT -15.805 -175.605 -15.475 -175.275 ;
        RECT -15.805 -176.685 -15.475 -176.355 ;
        RECT -15.805 -178.325 -15.475 -177.995 ;
        RECT -15.805 -179.685 -15.475 -179.355 ;
        RECT -15.805 -181.93 -15.475 -180.8 ;
        RECT -15.8 -182.045 -15.48 -105.92 ;
    END
    PORT
      LAYER met3 ;
        RECT -14.445 89.595 -14.115 89.925 ;
        RECT -14.445 88.235 -14.115 88.565 ;
        RECT -14.445 86.875 -14.115 87.205 ;
        RECT -14.445 85.515 -14.115 85.845 ;
        RECT -14.445 84.155 -14.115 84.485 ;
        RECT -14.445 82.795 -14.115 83.125 ;
        RECT -14.445 81.435 -14.115 81.765 ;
        RECT -14.445 80.075 -14.115 80.405 ;
        RECT -14.445 78.715 -14.115 79.045 ;
        RECT -14.445 77.355 -14.115 77.685 ;
        RECT -14.445 75.995 -14.115 76.325 ;
        RECT -14.445 74.635 -14.115 74.965 ;
        RECT -14.445 73.275 -14.115 73.605 ;
        RECT -14.445 71.915 -14.115 72.245 ;
        RECT -14.445 70.555 -14.115 70.885 ;
        RECT -14.445 69.195 -14.115 69.525 ;
        RECT -14.445 67.835 -14.115 68.165 ;
        RECT -14.445 66.475 -14.115 66.805 ;
        RECT -14.445 65.115 -14.115 65.445 ;
        RECT -14.445 63.755 -14.115 64.085 ;
        RECT -14.445 62.395 -14.115 62.725 ;
        RECT -14.445 61.035 -14.115 61.365 ;
        RECT -14.445 59.675 -14.115 60.005 ;
        RECT -14.445 58.315 -14.115 58.645 ;
        RECT -14.445 56.955 -14.115 57.285 ;
        RECT -14.445 55.595 -14.115 55.925 ;
        RECT -14.445 54.235 -14.115 54.565 ;
        RECT -14.445 52.875 -14.115 53.205 ;
        RECT -14.445 51.515 -14.115 51.845 ;
        RECT -14.445 50.155 -14.115 50.485 ;
        RECT -14.445 48.795 -14.115 49.125 ;
        RECT -14.445 47.435 -14.115 47.765 ;
        RECT -14.445 46.075 -14.115 46.405 ;
        RECT -14.445 44.715 -14.115 45.045 ;
        RECT -14.445 43.355 -14.115 43.685 ;
        RECT -14.445 41.995 -14.115 42.325 ;
        RECT -14.445 40.635 -14.115 40.965 ;
        RECT -14.445 39.275 -14.115 39.605 ;
        RECT -14.445 37.915 -14.115 38.245 ;
        RECT -14.445 36.555 -14.115 36.885 ;
        RECT -14.445 35.195 -14.115 35.525 ;
        RECT -14.445 33.835 -14.115 34.165 ;
        RECT -14.445 32.475 -14.115 32.805 ;
        RECT -14.445 31.115 -14.115 31.445 ;
        RECT -14.445 29.755 -14.115 30.085 ;
        RECT -14.445 28.395 -14.115 28.725 ;
        RECT -14.445 27.035 -14.115 27.365 ;
        RECT -14.445 25.675 -14.115 26.005 ;
        RECT -14.445 24.315 -14.115 24.645 ;
        RECT -14.445 22.955 -14.115 23.285 ;
        RECT -14.445 21.595 -14.115 21.925 ;
        RECT -14.445 20.235 -14.115 20.565 ;
        RECT -14.445 18.875 -14.115 19.205 ;
        RECT -14.445 17.515 -14.115 17.845 ;
        RECT -14.445 16.155 -14.115 16.485 ;
        RECT -14.445 14.795 -14.115 15.125 ;
        RECT -14.445 13.435 -14.115 13.765 ;
        RECT -14.445 12.075 -14.115 12.405 ;
        RECT -14.445 10.715 -14.115 11.045 ;
        RECT -14.445 9.355 -14.115 9.685 ;
        RECT -14.445 7.995 -14.115 8.325 ;
        RECT -14.445 6.635 -14.115 6.965 ;
        RECT -14.445 5.275 -14.115 5.605 ;
        RECT -14.445 3.915 -14.115 4.245 ;
        RECT -14.445 2.555 -14.115 2.885 ;
        RECT -14.445 1.195 -14.115 1.525 ;
        RECT -14.445 -0.165 -14.115 0.165 ;
        RECT -14.445 -2.885 -14.115 -2.555 ;
        RECT -14.445 -4.245 -14.115 -3.915 ;
        RECT -14.445 -5.605 -14.115 -5.275 ;
        RECT -14.445 -8.325 -14.115 -7.995 ;
        RECT -14.445 -9.685 -14.115 -9.355 ;
        RECT -14.445 -12.405 -14.115 -12.075 ;
        RECT -14.445 -13.765 -14.115 -13.435 ;
        RECT -14.445 -14.95 -14.115 -14.62 ;
        RECT -14.445 -17.845 -14.115 -17.515 ;
        RECT -14.445 -19.79 -14.115 -19.46 ;
        RECT -14.445 -27.365 -14.115 -27.035 ;
        RECT -14.445 -28.725 -14.115 -28.395 ;
        RECT -14.445 -30.085 -14.115 -29.755 ;
        RECT -14.445 -31.445 -14.115 -31.115 ;
        RECT -14.445 -32.805 -14.115 -32.475 ;
        RECT -14.445 -35.525 -14.115 -35.195 ;
        RECT -14.445 -36.885 -14.115 -36.555 ;
        RECT -14.445 -37.93 -14.115 -37.6 ;
        RECT -14.445 -42.77 -14.115 -42.44 ;
        RECT -14.445 -51.845 -14.115 -51.515 ;
        RECT -14.445 -53.205 -14.115 -52.875 ;
        RECT -14.445 -54.565 -14.115 -54.235 ;
        RECT -14.445 -55.925 -14.115 -55.595 ;
        RECT -14.445 -57.285 -14.115 -56.955 ;
        RECT -14.445 -58.645 -14.115 -58.315 ;
        RECT -14.445 -60.005 -14.115 -59.675 ;
        RECT -14.445 -61.365 -14.115 -61.035 ;
        RECT -14.445 -62.725 -14.115 -62.395 ;
        RECT -14.445 -64.085 -14.115 -63.755 ;
        RECT -14.445 -65.445 -14.115 -65.115 ;
        RECT -14.445 -68.165 -14.115 -67.835 ;
        RECT -14.445 -69.525 -14.115 -69.195 ;
        RECT -14.445 -70.885 -14.115 -70.555 ;
        RECT -14.445 -72.245 -14.115 -71.915 ;
        RECT -14.445 -74.965 -14.115 -74.635 ;
        RECT -14.445 -76.71 -14.115 -76.38 ;
        RECT -14.445 -77.685 -14.115 -77.355 ;
        RECT -14.445 -79.045 -14.115 -78.715 ;
        RECT -14.445 -81.765 -14.115 -81.435 ;
        RECT -14.445 -83.125 -14.115 -82.795 ;
        RECT -14.445 -84.485 -14.115 -84.155 ;
        RECT -14.445 -85.25 -14.115 -84.92 ;
        RECT -14.445 -87.205 -14.115 -86.875 ;
        RECT -14.44 -89.24 -14.12 242.565 ;
        RECT -14.445 241.32 -14.115 242.45 ;
        RECT -14.445 239.195 -14.115 239.525 ;
        RECT -14.445 237.835 -14.115 238.165 ;
        RECT -14.445 236.475 -14.115 236.805 ;
        RECT -14.445 235.115 -14.115 235.445 ;
        RECT -14.445 233.755 -14.115 234.085 ;
        RECT -14.445 232.395 -14.115 232.725 ;
        RECT -14.445 231.035 -14.115 231.365 ;
        RECT -14.445 229.675 -14.115 230.005 ;
        RECT -14.445 228.315 -14.115 228.645 ;
        RECT -14.445 226.955 -14.115 227.285 ;
        RECT -14.445 225.595 -14.115 225.925 ;
        RECT -14.445 224.235 -14.115 224.565 ;
        RECT -14.445 222.875 -14.115 223.205 ;
        RECT -14.445 221.515 -14.115 221.845 ;
        RECT -14.445 220.155 -14.115 220.485 ;
        RECT -14.445 218.795 -14.115 219.125 ;
        RECT -14.445 217.435 -14.115 217.765 ;
        RECT -14.445 216.075 -14.115 216.405 ;
        RECT -14.445 214.715 -14.115 215.045 ;
        RECT -14.445 213.355 -14.115 213.685 ;
        RECT -14.445 211.995 -14.115 212.325 ;
        RECT -14.445 210.635 -14.115 210.965 ;
        RECT -14.445 209.275 -14.115 209.605 ;
        RECT -14.445 207.915 -14.115 208.245 ;
        RECT -14.445 206.555 -14.115 206.885 ;
        RECT -14.445 205.195 -14.115 205.525 ;
        RECT -14.445 203.835 -14.115 204.165 ;
        RECT -14.445 202.475 -14.115 202.805 ;
        RECT -14.445 201.115 -14.115 201.445 ;
        RECT -14.445 199.755 -14.115 200.085 ;
        RECT -14.445 198.395 -14.115 198.725 ;
        RECT -14.445 197.035 -14.115 197.365 ;
        RECT -14.445 195.675 -14.115 196.005 ;
        RECT -14.445 194.315 -14.115 194.645 ;
        RECT -14.445 192.955 -14.115 193.285 ;
        RECT -14.445 191.595 -14.115 191.925 ;
        RECT -14.445 190.235 -14.115 190.565 ;
        RECT -14.445 188.875 -14.115 189.205 ;
        RECT -14.445 187.515 -14.115 187.845 ;
        RECT -14.445 186.155 -14.115 186.485 ;
        RECT -14.445 184.795 -14.115 185.125 ;
        RECT -14.445 183.435 -14.115 183.765 ;
        RECT -14.445 182.075 -14.115 182.405 ;
        RECT -14.445 180.715 -14.115 181.045 ;
        RECT -14.445 179.355 -14.115 179.685 ;
        RECT -14.445 177.995 -14.115 178.325 ;
        RECT -14.445 176.635 -14.115 176.965 ;
        RECT -14.445 175.275 -14.115 175.605 ;
        RECT -14.445 173.915 -14.115 174.245 ;
        RECT -14.445 172.555 -14.115 172.885 ;
        RECT -14.445 171.195 -14.115 171.525 ;
        RECT -14.445 169.835 -14.115 170.165 ;
        RECT -14.445 168.475 -14.115 168.805 ;
        RECT -14.445 167.115 -14.115 167.445 ;
        RECT -14.445 165.755 -14.115 166.085 ;
        RECT -14.445 164.395 -14.115 164.725 ;
        RECT -14.445 163.035 -14.115 163.365 ;
        RECT -14.445 161.675 -14.115 162.005 ;
        RECT -14.445 160.315 -14.115 160.645 ;
        RECT -14.445 158.955 -14.115 159.285 ;
        RECT -14.445 157.595 -14.115 157.925 ;
        RECT -14.445 156.235 -14.115 156.565 ;
        RECT -14.445 154.875 -14.115 155.205 ;
        RECT -14.445 153.515 -14.115 153.845 ;
        RECT -14.445 152.155 -14.115 152.485 ;
        RECT -14.445 150.795 -14.115 151.125 ;
        RECT -14.445 149.435 -14.115 149.765 ;
        RECT -14.445 148.075 -14.115 148.405 ;
        RECT -14.445 146.715 -14.115 147.045 ;
        RECT -14.445 145.355 -14.115 145.685 ;
        RECT -14.445 143.995 -14.115 144.325 ;
        RECT -14.445 142.635 -14.115 142.965 ;
        RECT -14.445 141.275 -14.115 141.605 ;
        RECT -14.445 139.915 -14.115 140.245 ;
        RECT -14.445 138.555 -14.115 138.885 ;
        RECT -14.445 137.195 -14.115 137.525 ;
        RECT -14.445 135.835 -14.115 136.165 ;
        RECT -14.445 134.475 -14.115 134.805 ;
        RECT -14.445 133.115 -14.115 133.445 ;
        RECT -14.445 131.755 -14.115 132.085 ;
        RECT -14.445 130.395 -14.115 130.725 ;
        RECT -14.445 129.035 -14.115 129.365 ;
        RECT -14.445 127.675 -14.115 128.005 ;
        RECT -14.445 126.315 -14.115 126.645 ;
        RECT -14.445 124.955 -14.115 125.285 ;
        RECT -14.445 123.595 -14.115 123.925 ;
        RECT -14.445 122.235 -14.115 122.565 ;
        RECT -14.445 120.875 -14.115 121.205 ;
        RECT -14.445 119.515 -14.115 119.845 ;
        RECT -14.445 118.155 -14.115 118.485 ;
        RECT -14.445 116.795 -14.115 117.125 ;
        RECT -14.445 115.435 -14.115 115.765 ;
        RECT -14.445 114.075 -14.115 114.405 ;
        RECT -14.445 112.715 -14.115 113.045 ;
        RECT -14.445 111.355 -14.115 111.685 ;
        RECT -14.445 109.995 -14.115 110.325 ;
        RECT -14.445 108.635 -14.115 108.965 ;
        RECT -14.445 107.275 -14.115 107.605 ;
        RECT -14.445 105.915 -14.115 106.245 ;
        RECT -14.445 104.555 -14.115 104.885 ;
        RECT -14.445 103.195 -14.115 103.525 ;
        RECT -14.445 101.835 -14.115 102.165 ;
        RECT -14.445 100.475 -14.115 100.805 ;
        RECT -14.445 99.115 -14.115 99.445 ;
        RECT -14.445 97.755 -14.115 98.085 ;
        RECT -14.445 96.395 -14.115 96.725 ;
        RECT -14.445 95.035 -14.115 95.365 ;
        RECT -14.445 93.675 -14.115 94.005 ;
        RECT -14.445 92.315 -14.115 92.645 ;
        RECT -14.445 90.955 -14.115 91.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -23.965 241.32 -23.635 242.45 ;
        RECT -23.965 239.195 -23.635 239.525 ;
        RECT -23.965 237.835 -23.635 238.165 ;
        RECT -23.965 236.475 -23.635 236.805 ;
        RECT -23.965 235.115 -23.635 235.445 ;
        RECT -23.965 233.755 -23.635 234.085 ;
        RECT -23.965 232.395 -23.635 232.725 ;
        RECT -23.965 231.035 -23.635 231.365 ;
        RECT -23.965 229.675 -23.635 230.005 ;
        RECT -23.965 228.315 -23.635 228.645 ;
        RECT -23.965 226.955 -23.635 227.285 ;
        RECT -23.965 225.595 -23.635 225.925 ;
        RECT -23.965 224.235 -23.635 224.565 ;
        RECT -23.965 222.875 -23.635 223.205 ;
        RECT -23.965 221.515 -23.635 221.845 ;
        RECT -23.965 220.155 -23.635 220.485 ;
        RECT -23.965 218.795 -23.635 219.125 ;
        RECT -23.965 217.435 -23.635 217.765 ;
        RECT -23.965 216.075 -23.635 216.405 ;
        RECT -23.965 214.715 -23.635 215.045 ;
        RECT -23.965 213.355 -23.635 213.685 ;
        RECT -23.965 211.995 -23.635 212.325 ;
        RECT -23.965 210.635 -23.635 210.965 ;
        RECT -23.965 209.275 -23.635 209.605 ;
        RECT -23.965 207.915 -23.635 208.245 ;
        RECT -23.965 206.555 -23.635 206.885 ;
        RECT -23.965 205.195 -23.635 205.525 ;
        RECT -23.965 203.835 -23.635 204.165 ;
        RECT -23.965 202.475 -23.635 202.805 ;
        RECT -23.965 201.115 -23.635 201.445 ;
        RECT -23.965 199.755 -23.635 200.085 ;
        RECT -23.965 198.395 -23.635 198.725 ;
        RECT -23.965 197.035 -23.635 197.365 ;
        RECT -23.965 195.675 -23.635 196.005 ;
        RECT -23.965 194.315 -23.635 194.645 ;
        RECT -23.965 192.955 -23.635 193.285 ;
        RECT -23.965 191.595 -23.635 191.925 ;
        RECT -23.965 190.235 -23.635 190.565 ;
        RECT -23.965 188.875 -23.635 189.205 ;
        RECT -23.965 187.515 -23.635 187.845 ;
        RECT -23.965 186.155 -23.635 186.485 ;
        RECT -23.965 184.795 -23.635 185.125 ;
        RECT -23.965 183.435 -23.635 183.765 ;
        RECT -23.965 182.075 -23.635 182.405 ;
        RECT -23.965 180.715 -23.635 181.045 ;
        RECT -23.965 179.355 -23.635 179.685 ;
        RECT -23.965 177.995 -23.635 178.325 ;
        RECT -23.965 176.635 -23.635 176.965 ;
        RECT -23.965 175.275 -23.635 175.605 ;
        RECT -23.965 173.915 -23.635 174.245 ;
        RECT -23.965 172.555 -23.635 172.885 ;
        RECT -23.965 171.195 -23.635 171.525 ;
        RECT -23.965 169.835 -23.635 170.165 ;
        RECT -23.965 168.475 -23.635 168.805 ;
        RECT -23.965 167.115 -23.635 167.445 ;
        RECT -23.965 165.755 -23.635 166.085 ;
        RECT -23.965 164.395 -23.635 164.725 ;
        RECT -23.965 163.035 -23.635 163.365 ;
        RECT -23.965 161.675 -23.635 162.005 ;
        RECT -23.965 160.315 -23.635 160.645 ;
        RECT -23.965 158.955 -23.635 159.285 ;
        RECT -23.965 157.595 -23.635 157.925 ;
        RECT -23.965 156.235 -23.635 156.565 ;
        RECT -23.965 154.875 -23.635 155.205 ;
        RECT -23.965 153.515 -23.635 153.845 ;
        RECT -23.965 152.155 -23.635 152.485 ;
        RECT -23.965 150.795 -23.635 151.125 ;
        RECT -23.965 149.435 -23.635 149.765 ;
        RECT -23.965 148.075 -23.635 148.405 ;
        RECT -23.965 146.715 -23.635 147.045 ;
        RECT -23.965 145.355 -23.635 145.685 ;
        RECT -23.965 143.995 -23.635 144.325 ;
        RECT -23.965 142.635 -23.635 142.965 ;
        RECT -23.965 141.275 -23.635 141.605 ;
        RECT -23.965 139.915 -23.635 140.245 ;
        RECT -23.965 138.555 -23.635 138.885 ;
        RECT -23.965 137.195 -23.635 137.525 ;
        RECT -23.965 135.835 -23.635 136.165 ;
        RECT -23.965 134.475 -23.635 134.805 ;
        RECT -23.965 133.115 -23.635 133.445 ;
        RECT -23.965 131.755 -23.635 132.085 ;
        RECT -23.965 130.395 -23.635 130.725 ;
        RECT -23.965 129.035 -23.635 129.365 ;
        RECT -23.965 127.675 -23.635 128.005 ;
        RECT -23.965 126.315 -23.635 126.645 ;
        RECT -23.965 124.955 -23.635 125.285 ;
        RECT -23.965 123.595 -23.635 123.925 ;
        RECT -23.965 122.235 -23.635 122.565 ;
        RECT -23.965 120.875 -23.635 121.205 ;
        RECT -23.965 119.515 -23.635 119.845 ;
        RECT -23.965 118.155 -23.635 118.485 ;
        RECT -23.965 116.795 -23.635 117.125 ;
        RECT -23.965 115.435 -23.635 115.765 ;
        RECT -23.965 114.075 -23.635 114.405 ;
        RECT -23.965 112.715 -23.635 113.045 ;
        RECT -23.965 111.355 -23.635 111.685 ;
        RECT -23.965 109.995 -23.635 110.325 ;
        RECT -23.965 108.635 -23.635 108.965 ;
        RECT -23.965 107.275 -23.635 107.605 ;
        RECT -23.965 105.915 -23.635 106.245 ;
        RECT -23.965 104.555 -23.635 104.885 ;
        RECT -23.965 103.195 -23.635 103.525 ;
        RECT -23.965 101.835 -23.635 102.165 ;
        RECT -23.965 100.475 -23.635 100.805 ;
        RECT -23.965 99.115 -23.635 99.445 ;
        RECT -23.965 97.755 -23.635 98.085 ;
        RECT -23.965 96.395 -23.635 96.725 ;
        RECT -23.965 95.035 -23.635 95.365 ;
        RECT -23.965 93.675 -23.635 94.005 ;
        RECT -23.965 92.315 -23.635 92.645 ;
        RECT -23.965 90.955 -23.635 91.285 ;
        RECT -23.965 89.595 -23.635 89.925 ;
        RECT -23.965 88.235 -23.635 88.565 ;
        RECT -23.965 86.875 -23.635 87.205 ;
        RECT -23.965 85.515 -23.635 85.845 ;
        RECT -23.965 84.155 -23.635 84.485 ;
        RECT -23.965 82.795 -23.635 83.125 ;
        RECT -23.965 81.435 -23.635 81.765 ;
        RECT -23.965 80.075 -23.635 80.405 ;
        RECT -23.965 78.715 -23.635 79.045 ;
        RECT -23.965 77.355 -23.635 77.685 ;
        RECT -23.965 75.995 -23.635 76.325 ;
        RECT -23.965 74.635 -23.635 74.965 ;
        RECT -23.965 73.275 -23.635 73.605 ;
        RECT -23.965 71.915 -23.635 72.245 ;
        RECT -23.965 70.555 -23.635 70.885 ;
        RECT -23.965 69.195 -23.635 69.525 ;
        RECT -23.965 67.835 -23.635 68.165 ;
        RECT -23.965 66.475 -23.635 66.805 ;
        RECT -23.965 65.115 -23.635 65.445 ;
        RECT -23.965 63.755 -23.635 64.085 ;
        RECT -23.965 62.395 -23.635 62.725 ;
        RECT -23.965 61.035 -23.635 61.365 ;
        RECT -23.965 59.675 -23.635 60.005 ;
        RECT -23.965 58.315 -23.635 58.645 ;
        RECT -23.965 56.955 -23.635 57.285 ;
        RECT -23.965 55.595 -23.635 55.925 ;
        RECT -23.965 54.235 -23.635 54.565 ;
        RECT -23.965 52.875 -23.635 53.205 ;
        RECT -23.965 51.515 -23.635 51.845 ;
        RECT -23.965 50.155 -23.635 50.485 ;
        RECT -23.965 48.795 -23.635 49.125 ;
        RECT -23.965 47.435 -23.635 47.765 ;
        RECT -23.965 46.075 -23.635 46.405 ;
        RECT -23.965 44.715 -23.635 45.045 ;
        RECT -23.965 43.355 -23.635 43.685 ;
        RECT -23.965 41.995 -23.635 42.325 ;
        RECT -23.965 40.635 -23.635 40.965 ;
        RECT -23.965 39.275 -23.635 39.605 ;
        RECT -23.965 37.915 -23.635 38.245 ;
        RECT -23.965 36.555 -23.635 36.885 ;
        RECT -23.965 35.195 -23.635 35.525 ;
        RECT -23.965 33.835 -23.635 34.165 ;
        RECT -23.965 32.475 -23.635 32.805 ;
        RECT -23.965 31.115 -23.635 31.445 ;
        RECT -23.965 29.755 -23.635 30.085 ;
        RECT -23.965 28.395 -23.635 28.725 ;
        RECT -23.965 27.035 -23.635 27.365 ;
        RECT -23.965 25.675 -23.635 26.005 ;
        RECT -23.965 24.315 -23.635 24.645 ;
        RECT -23.965 22.955 -23.635 23.285 ;
        RECT -23.965 21.595 -23.635 21.925 ;
        RECT -23.965 20.235 -23.635 20.565 ;
        RECT -23.965 18.875 -23.635 19.205 ;
        RECT -23.965 17.515 -23.635 17.845 ;
        RECT -23.965 16.155 -23.635 16.485 ;
        RECT -23.965 14.795 -23.635 15.125 ;
        RECT -23.965 13.435 -23.635 13.765 ;
        RECT -23.965 12.075 -23.635 12.405 ;
        RECT -23.965 10.715 -23.635 11.045 ;
        RECT -23.965 9.355 -23.635 9.685 ;
        RECT -23.965 7.995 -23.635 8.325 ;
        RECT -23.965 6.635 -23.635 6.965 ;
        RECT -23.965 5.275 -23.635 5.605 ;
        RECT -23.965 3.915 -23.635 4.245 ;
        RECT -23.965 2.555 -23.635 2.885 ;
        RECT -23.965 1.195 -23.635 1.525 ;
        RECT -23.965 -0.165 -23.635 0.165 ;
        RECT -23.965 -2.885 -23.635 -2.555 ;
        RECT -23.965 -8.325 -23.635 -7.995 ;
        RECT -23.965 -9.685 -23.635 -9.355 ;
        RECT -23.965 -14.95 -23.635 -14.62 ;
        RECT -23.965 -17.845 -23.635 -17.515 ;
        RECT -23.965 -19.79 -23.635 -19.46 ;
        RECT -23.965 -20.565 -23.635 -20.235 ;
        RECT -23.965 -32.805 -23.635 -32.475 ;
        RECT -23.965 -35.525 -23.635 -35.195 ;
        RECT -23.965 -36.885 -23.635 -36.555 ;
        RECT -23.965 -37.93 -23.635 -37.6 ;
        RECT -23.965 -40.965 -23.635 -40.635 ;
        RECT -23.965 -42.77 -23.635 -42.44 ;
        RECT -23.965 -43.685 -23.635 -43.355 ;
        RECT -23.965 -50.485 -23.635 -50.155 ;
        RECT -23.965 -51.845 -23.635 -51.515 ;
        RECT -23.965 -53.205 -23.635 -52.875 ;
        RECT -23.965 -54.565 -23.635 -54.235 ;
        RECT -23.965 -55.925 -23.635 -55.595 ;
        RECT -23.965 -57.285 -23.635 -56.955 ;
        RECT -23.965 -58.645 -23.635 -58.315 ;
        RECT -23.965 -60.005 -23.635 -59.675 ;
        RECT -23.965 -61.365 -23.635 -61.035 ;
        RECT -23.965 -62.725 -23.635 -62.395 ;
        RECT -23.965 -64.085 -23.635 -63.755 ;
        RECT -23.965 -65.445 -23.635 -65.115 ;
        RECT -23.965 -68.165 -23.635 -67.835 ;
        RECT -23.965 -69.525 -23.635 -69.195 ;
        RECT -23.965 -70.885 -23.635 -70.555 ;
        RECT -23.965 -72.245 -23.635 -71.915 ;
        RECT -23.965 -74.965 -23.635 -74.635 ;
        RECT -23.965 -76.71 -23.635 -76.38 ;
        RECT -23.965 -77.685 -23.635 -77.355 ;
        RECT -23.965 -79.045 -23.635 -78.715 ;
        RECT -23.965 -81.765 -23.635 -81.435 ;
        RECT -23.965 -83.125 -23.635 -82.795 ;
        RECT -23.965 -84.485 -23.635 -84.155 ;
        RECT -23.965 -85.25 -23.635 -84.92 ;
        RECT -23.965 -87.205 -23.635 -86.875 ;
        RECT -23.965 -89.925 -23.635 -89.595 ;
        RECT -23.965 -91.285 -23.635 -90.955 ;
        RECT -23.965 -92.645 -23.635 -92.315 ;
        RECT -23.965 -94.005 -23.635 -93.675 ;
        RECT -23.965 -96.725 -23.635 -96.395 ;
        RECT -23.965 -98.085 -23.635 -97.755 ;
        RECT -23.965 -98.89 -23.635 -98.56 ;
        RECT -23.965 -100.805 -23.635 -100.475 ;
        RECT -23.965 -102.165 -23.635 -101.835 ;
        RECT -23.965 -104.885 -23.635 -104.555 ;
        RECT -23.965 -106.245 -23.635 -105.915 ;
        RECT -23.965 -107.43 -23.635 -107.1 ;
        RECT -23.965 -115.765 -23.635 -115.435 ;
        RECT -23.965 -117.125 -23.635 -116.795 ;
        RECT -23.965 -118.485 -23.635 -118.155 ;
        RECT -23.965 -123.925 -23.635 -123.595 ;
        RECT -23.965 -125.285 -23.635 -124.955 ;
        RECT -23.965 -126.645 -23.635 -126.315 ;
        RECT -23.965 -128.005 -23.635 -127.675 ;
        RECT -23.965 -130.725 -23.635 -130.395 ;
        RECT -23.965 -136.165 -23.635 -135.835 ;
        RECT -23.965 -137.525 -23.635 -137.195 ;
        RECT -23.965 -141.605 -23.635 -141.275 ;
        RECT -23.965 -142.965 -23.635 -142.635 ;
        RECT -23.965 -147.045 -23.635 -146.715 ;
        RECT -23.965 -148.405 -23.635 -148.075 ;
        RECT -23.965 -149.765 -23.635 -149.435 ;
        RECT -23.965 -152.485 -23.635 -152.155 ;
        RECT -23.965 -153.845 -23.635 -153.515 ;
        RECT -23.965 -159.285 -23.635 -158.955 ;
        RECT -23.965 -160.645 -23.635 -160.315 ;
        RECT -23.965 -162.005 -23.635 -161.675 ;
        RECT -23.965 -163.365 -23.635 -163.035 ;
        RECT -23.965 -164.725 -23.635 -164.395 ;
        RECT -23.965 -166.085 -23.635 -165.755 ;
        RECT -23.965 -167.445 -23.635 -167.115 ;
        RECT -23.965 -168.805 -23.635 -168.475 ;
        RECT -23.965 -171.525 -23.635 -171.195 ;
        RECT -23.965 -172.885 -23.635 -172.555 ;
        RECT -23.965 -175.605 -23.635 -175.275 ;
        RECT -23.965 -176.685 -23.635 -176.355 ;
        RECT -23.965 -178.325 -23.635 -177.995 ;
        RECT -23.965 -179.685 -23.635 -179.355 ;
        RECT -23.965 -181.93 -23.635 -180.8 ;
        RECT -23.96 -182.045 -23.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -22.605 241.32 -22.275 242.45 ;
        RECT -22.605 239.195 -22.275 239.525 ;
        RECT -22.605 237.835 -22.275 238.165 ;
        RECT -22.605 236.475 -22.275 236.805 ;
        RECT -22.605 235.115 -22.275 235.445 ;
        RECT -22.605 233.755 -22.275 234.085 ;
        RECT -22.605 232.395 -22.275 232.725 ;
        RECT -22.605 231.035 -22.275 231.365 ;
        RECT -22.605 229.675 -22.275 230.005 ;
        RECT -22.605 228.315 -22.275 228.645 ;
        RECT -22.605 226.955 -22.275 227.285 ;
        RECT -22.605 225.595 -22.275 225.925 ;
        RECT -22.605 224.235 -22.275 224.565 ;
        RECT -22.605 222.875 -22.275 223.205 ;
        RECT -22.605 221.515 -22.275 221.845 ;
        RECT -22.605 220.155 -22.275 220.485 ;
        RECT -22.605 218.795 -22.275 219.125 ;
        RECT -22.605 217.435 -22.275 217.765 ;
        RECT -22.605 216.075 -22.275 216.405 ;
        RECT -22.605 214.715 -22.275 215.045 ;
        RECT -22.605 213.355 -22.275 213.685 ;
        RECT -22.605 211.995 -22.275 212.325 ;
        RECT -22.605 210.635 -22.275 210.965 ;
        RECT -22.605 209.275 -22.275 209.605 ;
        RECT -22.605 207.915 -22.275 208.245 ;
        RECT -22.605 206.555 -22.275 206.885 ;
        RECT -22.605 205.195 -22.275 205.525 ;
        RECT -22.605 203.835 -22.275 204.165 ;
        RECT -22.605 202.475 -22.275 202.805 ;
        RECT -22.605 201.115 -22.275 201.445 ;
        RECT -22.605 199.755 -22.275 200.085 ;
        RECT -22.605 198.395 -22.275 198.725 ;
        RECT -22.605 197.035 -22.275 197.365 ;
        RECT -22.605 195.675 -22.275 196.005 ;
        RECT -22.605 194.315 -22.275 194.645 ;
        RECT -22.605 192.955 -22.275 193.285 ;
        RECT -22.605 191.595 -22.275 191.925 ;
        RECT -22.605 190.235 -22.275 190.565 ;
        RECT -22.605 188.875 -22.275 189.205 ;
        RECT -22.605 187.515 -22.275 187.845 ;
        RECT -22.605 186.155 -22.275 186.485 ;
        RECT -22.605 184.795 -22.275 185.125 ;
        RECT -22.605 183.435 -22.275 183.765 ;
        RECT -22.605 182.075 -22.275 182.405 ;
        RECT -22.605 180.715 -22.275 181.045 ;
        RECT -22.605 179.355 -22.275 179.685 ;
        RECT -22.605 177.995 -22.275 178.325 ;
        RECT -22.605 176.635 -22.275 176.965 ;
        RECT -22.605 175.275 -22.275 175.605 ;
        RECT -22.605 173.915 -22.275 174.245 ;
        RECT -22.605 172.555 -22.275 172.885 ;
        RECT -22.605 171.195 -22.275 171.525 ;
        RECT -22.605 169.835 -22.275 170.165 ;
        RECT -22.605 168.475 -22.275 168.805 ;
        RECT -22.605 167.115 -22.275 167.445 ;
        RECT -22.605 165.755 -22.275 166.085 ;
        RECT -22.605 164.395 -22.275 164.725 ;
        RECT -22.605 163.035 -22.275 163.365 ;
        RECT -22.605 161.675 -22.275 162.005 ;
        RECT -22.605 160.315 -22.275 160.645 ;
        RECT -22.605 158.955 -22.275 159.285 ;
        RECT -22.605 157.595 -22.275 157.925 ;
        RECT -22.605 156.235 -22.275 156.565 ;
        RECT -22.605 154.875 -22.275 155.205 ;
        RECT -22.605 153.515 -22.275 153.845 ;
        RECT -22.605 152.155 -22.275 152.485 ;
        RECT -22.605 150.795 -22.275 151.125 ;
        RECT -22.605 149.435 -22.275 149.765 ;
        RECT -22.605 148.075 -22.275 148.405 ;
        RECT -22.605 146.715 -22.275 147.045 ;
        RECT -22.605 145.355 -22.275 145.685 ;
        RECT -22.605 143.995 -22.275 144.325 ;
        RECT -22.605 142.635 -22.275 142.965 ;
        RECT -22.605 141.275 -22.275 141.605 ;
        RECT -22.605 139.915 -22.275 140.245 ;
        RECT -22.605 138.555 -22.275 138.885 ;
        RECT -22.605 137.195 -22.275 137.525 ;
        RECT -22.605 135.835 -22.275 136.165 ;
        RECT -22.605 134.475 -22.275 134.805 ;
        RECT -22.605 133.115 -22.275 133.445 ;
        RECT -22.605 131.755 -22.275 132.085 ;
        RECT -22.605 130.395 -22.275 130.725 ;
        RECT -22.605 129.035 -22.275 129.365 ;
        RECT -22.605 127.675 -22.275 128.005 ;
        RECT -22.605 126.315 -22.275 126.645 ;
        RECT -22.605 124.955 -22.275 125.285 ;
        RECT -22.605 123.595 -22.275 123.925 ;
        RECT -22.605 122.235 -22.275 122.565 ;
        RECT -22.605 120.875 -22.275 121.205 ;
        RECT -22.605 119.515 -22.275 119.845 ;
        RECT -22.605 118.155 -22.275 118.485 ;
        RECT -22.605 116.795 -22.275 117.125 ;
        RECT -22.605 115.435 -22.275 115.765 ;
        RECT -22.605 114.075 -22.275 114.405 ;
        RECT -22.605 112.715 -22.275 113.045 ;
        RECT -22.605 111.355 -22.275 111.685 ;
        RECT -22.605 109.995 -22.275 110.325 ;
        RECT -22.605 108.635 -22.275 108.965 ;
        RECT -22.605 107.275 -22.275 107.605 ;
        RECT -22.605 105.915 -22.275 106.245 ;
        RECT -22.605 104.555 -22.275 104.885 ;
        RECT -22.605 103.195 -22.275 103.525 ;
        RECT -22.605 101.835 -22.275 102.165 ;
        RECT -22.605 100.475 -22.275 100.805 ;
        RECT -22.605 99.115 -22.275 99.445 ;
        RECT -22.605 97.755 -22.275 98.085 ;
        RECT -22.605 96.395 -22.275 96.725 ;
        RECT -22.605 95.035 -22.275 95.365 ;
        RECT -22.605 93.675 -22.275 94.005 ;
        RECT -22.605 92.315 -22.275 92.645 ;
        RECT -22.605 90.955 -22.275 91.285 ;
        RECT -22.605 89.595 -22.275 89.925 ;
        RECT -22.605 88.235 -22.275 88.565 ;
        RECT -22.605 86.875 -22.275 87.205 ;
        RECT -22.605 85.515 -22.275 85.845 ;
        RECT -22.605 84.155 -22.275 84.485 ;
        RECT -22.605 82.795 -22.275 83.125 ;
        RECT -22.605 81.435 -22.275 81.765 ;
        RECT -22.605 80.075 -22.275 80.405 ;
        RECT -22.605 78.715 -22.275 79.045 ;
        RECT -22.605 77.355 -22.275 77.685 ;
        RECT -22.605 75.995 -22.275 76.325 ;
        RECT -22.605 74.635 -22.275 74.965 ;
        RECT -22.605 73.275 -22.275 73.605 ;
        RECT -22.605 71.915 -22.275 72.245 ;
        RECT -22.605 70.555 -22.275 70.885 ;
        RECT -22.605 69.195 -22.275 69.525 ;
        RECT -22.605 67.835 -22.275 68.165 ;
        RECT -22.605 66.475 -22.275 66.805 ;
        RECT -22.605 65.115 -22.275 65.445 ;
        RECT -22.605 63.755 -22.275 64.085 ;
        RECT -22.605 62.395 -22.275 62.725 ;
        RECT -22.605 61.035 -22.275 61.365 ;
        RECT -22.605 59.675 -22.275 60.005 ;
        RECT -22.605 58.315 -22.275 58.645 ;
        RECT -22.605 56.955 -22.275 57.285 ;
        RECT -22.605 55.595 -22.275 55.925 ;
        RECT -22.605 54.235 -22.275 54.565 ;
        RECT -22.605 52.875 -22.275 53.205 ;
        RECT -22.605 51.515 -22.275 51.845 ;
        RECT -22.605 50.155 -22.275 50.485 ;
        RECT -22.605 48.795 -22.275 49.125 ;
        RECT -22.605 47.435 -22.275 47.765 ;
        RECT -22.605 46.075 -22.275 46.405 ;
        RECT -22.605 44.715 -22.275 45.045 ;
        RECT -22.605 43.355 -22.275 43.685 ;
        RECT -22.605 41.995 -22.275 42.325 ;
        RECT -22.605 40.635 -22.275 40.965 ;
        RECT -22.605 39.275 -22.275 39.605 ;
        RECT -22.605 37.915 -22.275 38.245 ;
        RECT -22.605 36.555 -22.275 36.885 ;
        RECT -22.605 35.195 -22.275 35.525 ;
        RECT -22.605 33.835 -22.275 34.165 ;
        RECT -22.605 32.475 -22.275 32.805 ;
        RECT -22.605 31.115 -22.275 31.445 ;
        RECT -22.605 29.755 -22.275 30.085 ;
        RECT -22.605 28.395 -22.275 28.725 ;
        RECT -22.605 27.035 -22.275 27.365 ;
        RECT -22.605 25.675 -22.275 26.005 ;
        RECT -22.605 24.315 -22.275 24.645 ;
        RECT -22.605 22.955 -22.275 23.285 ;
        RECT -22.605 21.595 -22.275 21.925 ;
        RECT -22.605 20.235 -22.275 20.565 ;
        RECT -22.605 18.875 -22.275 19.205 ;
        RECT -22.605 17.515 -22.275 17.845 ;
        RECT -22.605 16.155 -22.275 16.485 ;
        RECT -22.605 14.795 -22.275 15.125 ;
        RECT -22.605 13.435 -22.275 13.765 ;
        RECT -22.605 12.075 -22.275 12.405 ;
        RECT -22.605 10.715 -22.275 11.045 ;
        RECT -22.605 9.355 -22.275 9.685 ;
        RECT -22.605 7.995 -22.275 8.325 ;
        RECT -22.605 6.635 -22.275 6.965 ;
        RECT -22.605 5.275 -22.275 5.605 ;
        RECT -22.605 3.915 -22.275 4.245 ;
        RECT -22.605 2.555 -22.275 2.885 ;
        RECT -22.605 1.195 -22.275 1.525 ;
        RECT -22.605 -0.165 -22.275 0.165 ;
        RECT -22.605 -2.885 -22.275 -2.555 ;
        RECT -22.605 -8.325 -22.275 -7.995 ;
        RECT -22.605 -9.685 -22.275 -9.355 ;
        RECT -22.605 -14.95 -22.275 -14.62 ;
        RECT -22.605 -17.845 -22.275 -17.515 ;
        RECT -22.605 -19.79 -22.275 -19.46 ;
        RECT -22.605 -20.565 -22.275 -20.235 ;
        RECT -22.605 -32.805 -22.275 -32.475 ;
        RECT -22.605 -35.525 -22.275 -35.195 ;
        RECT -22.605 -36.885 -22.275 -36.555 ;
        RECT -22.605 -37.93 -22.275 -37.6 ;
        RECT -22.605 -40.965 -22.275 -40.635 ;
        RECT -22.605 -42.77 -22.275 -42.44 ;
        RECT -22.605 -43.685 -22.275 -43.355 ;
        RECT -22.605 -50.485 -22.275 -50.155 ;
        RECT -22.605 -51.845 -22.275 -51.515 ;
        RECT -22.605 -53.205 -22.275 -52.875 ;
        RECT -22.605 -54.565 -22.275 -54.235 ;
        RECT -22.605 -55.925 -22.275 -55.595 ;
        RECT -22.605 -57.285 -22.275 -56.955 ;
        RECT -22.605 -58.645 -22.275 -58.315 ;
        RECT -22.605 -60.005 -22.275 -59.675 ;
        RECT -22.605 -61.365 -22.275 -61.035 ;
        RECT -22.605 -62.725 -22.275 -62.395 ;
        RECT -22.605 -64.085 -22.275 -63.755 ;
        RECT -22.605 -65.445 -22.275 -65.115 ;
        RECT -22.605 -68.165 -22.275 -67.835 ;
        RECT -22.605 -69.525 -22.275 -69.195 ;
        RECT -22.605 -70.885 -22.275 -70.555 ;
        RECT -22.605 -72.245 -22.275 -71.915 ;
        RECT -22.605 -74.965 -22.275 -74.635 ;
        RECT -22.605 -76.71 -22.275 -76.38 ;
        RECT -22.605 -77.685 -22.275 -77.355 ;
        RECT -22.605 -79.045 -22.275 -78.715 ;
        RECT -22.605 -81.765 -22.275 -81.435 ;
        RECT -22.605 -83.125 -22.275 -82.795 ;
        RECT -22.605 -84.485 -22.275 -84.155 ;
        RECT -22.605 -85.25 -22.275 -84.92 ;
        RECT -22.605 -87.205 -22.275 -86.875 ;
        RECT -22.605 -89.925 -22.275 -89.595 ;
        RECT -22.605 -91.285 -22.275 -90.955 ;
        RECT -22.605 -92.645 -22.275 -92.315 ;
        RECT -22.605 -94.005 -22.275 -93.675 ;
        RECT -22.605 -96.725 -22.275 -96.395 ;
        RECT -22.605 -98.085 -22.275 -97.755 ;
        RECT -22.605 -98.89 -22.275 -98.56 ;
        RECT -22.605 -100.805 -22.275 -100.475 ;
        RECT -22.605 -102.165 -22.275 -101.835 ;
        RECT -22.605 -104.885 -22.275 -104.555 ;
        RECT -22.605 -107.43 -22.275 -107.1 ;
        RECT -22.605 -115.765 -22.275 -115.435 ;
        RECT -22.605 -117.125 -22.275 -116.795 ;
        RECT -22.605 -118.485 -22.275 -118.155 ;
        RECT -22.605 -123.925 -22.275 -123.595 ;
        RECT -22.605 -125.285 -22.275 -124.955 ;
        RECT -22.605 -126.645 -22.275 -126.315 ;
        RECT -22.605 -128.005 -22.275 -127.675 ;
        RECT -22.605 -130.725 -22.275 -130.395 ;
        RECT -22.605 -136.165 -22.275 -135.835 ;
        RECT -22.605 -137.525 -22.275 -137.195 ;
        RECT -22.605 -141.605 -22.275 -141.275 ;
        RECT -22.605 -142.965 -22.275 -142.635 ;
        RECT -22.605 -144.325 -22.275 -143.995 ;
        RECT -22.605 -147.045 -22.275 -146.715 ;
        RECT -22.605 -148.405 -22.275 -148.075 ;
        RECT -22.605 -149.765 -22.275 -149.435 ;
        RECT -22.605 -152.485 -22.275 -152.155 ;
        RECT -22.605 -153.845 -22.275 -153.515 ;
        RECT -22.605 -159.285 -22.275 -158.955 ;
        RECT -22.605 -160.645 -22.275 -160.315 ;
        RECT -22.605 -162.005 -22.275 -161.675 ;
        RECT -22.605 -163.365 -22.275 -163.035 ;
        RECT -22.605 -164.725 -22.275 -164.395 ;
        RECT -22.605 -166.085 -22.275 -165.755 ;
        RECT -22.605 -167.445 -22.275 -167.115 ;
        RECT -22.605 -168.805 -22.275 -168.475 ;
        RECT -22.605 -171.525 -22.275 -171.195 ;
        RECT -22.605 -175.605 -22.275 -175.275 ;
        RECT -22.605 -178.325 -22.275 -177.995 ;
        RECT -22.605 -179.685 -22.275 -179.355 ;
        RECT -22.605 -181.93 -22.275 -180.8 ;
        RECT -22.6 -182.045 -22.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 241.32 -20.915 242.45 ;
        RECT -21.245 239.195 -20.915 239.525 ;
        RECT -21.245 237.835 -20.915 238.165 ;
        RECT -21.245 236.475 -20.915 236.805 ;
        RECT -21.245 235.115 -20.915 235.445 ;
        RECT -21.245 233.755 -20.915 234.085 ;
        RECT -21.245 232.395 -20.915 232.725 ;
        RECT -21.245 231.035 -20.915 231.365 ;
        RECT -21.245 229.675 -20.915 230.005 ;
        RECT -21.245 228.315 -20.915 228.645 ;
        RECT -21.245 226.955 -20.915 227.285 ;
        RECT -21.245 225.595 -20.915 225.925 ;
        RECT -21.245 224.235 -20.915 224.565 ;
        RECT -21.245 222.875 -20.915 223.205 ;
        RECT -21.245 221.515 -20.915 221.845 ;
        RECT -21.245 220.155 -20.915 220.485 ;
        RECT -21.245 218.795 -20.915 219.125 ;
        RECT -21.245 217.435 -20.915 217.765 ;
        RECT -21.245 216.075 -20.915 216.405 ;
        RECT -21.245 214.715 -20.915 215.045 ;
        RECT -21.245 213.355 -20.915 213.685 ;
        RECT -21.245 211.995 -20.915 212.325 ;
        RECT -21.245 210.635 -20.915 210.965 ;
        RECT -21.245 209.275 -20.915 209.605 ;
        RECT -21.245 207.915 -20.915 208.245 ;
        RECT -21.245 206.555 -20.915 206.885 ;
        RECT -21.245 205.195 -20.915 205.525 ;
        RECT -21.245 203.835 -20.915 204.165 ;
        RECT -21.245 202.475 -20.915 202.805 ;
        RECT -21.245 201.115 -20.915 201.445 ;
        RECT -21.245 199.755 -20.915 200.085 ;
        RECT -21.245 198.395 -20.915 198.725 ;
        RECT -21.245 197.035 -20.915 197.365 ;
        RECT -21.245 195.675 -20.915 196.005 ;
        RECT -21.245 194.315 -20.915 194.645 ;
        RECT -21.245 192.955 -20.915 193.285 ;
        RECT -21.245 191.595 -20.915 191.925 ;
        RECT -21.245 190.235 -20.915 190.565 ;
        RECT -21.245 188.875 -20.915 189.205 ;
        RECT -21.245 187.515 -20.915 187.845 ;
        RECT -21.245 186.155 -20.915 186.485 ;
        RECT -21.245 184.795 -20.915 185.125 ;
        RECT -21.245 183.435 -20.915 183.765 ;
        RECT -21.245 182.075 -20.915 182.405 ;
        RECT -21.245 180.715 -20.915 181.045 ;
        RECT -21.245 179.355 -20.915 179.685 ;
        RECT -21.245 177.995 -20.915 178.325 ;
        RECT -21.245 176.635 -20.915 176.965 ;
        RECT -21.245 175.275 -20.915 175.605 ;
        RECT -21.245 173.915 -20.915 174.245 ;
        RECT -21.245 172.555 -20.915 172.885 ;
        RECT -21.245 171.195 -20.915 171.525 ;
        RECT -21.245 169.835 -20.915 170.165 ;
        RECT -21.245 168.475 -20.915 168.805 ;
        RECT -21.245 167.115 -20.915 167.445 ;
        RECT -21.245 165.755 -20.915 166.085 ;
        RECT -21.245 164.395 -20.915 164.725 ;
        RECT -21.245 163.035 -20.915 163.365 ;
        RECT -21.245 161.675 -20.915 162.005 ;
        RECT -21.245 160.315 -20.915 160.645 ;
        RECT -21.245 158.955 -20.915 159.285 ;
        RECT -21.245 157.595 -20.915 157.925 ;
        RECT -21.245 156.235 -20.915 156.565 ;
        RECT -21.245 154.875 -20.915 155.205 ;
        RECT -21.245 153.515 -20.915 153.845 ;
        RECT -21.245 152.155 -20.915 152.485 ;
        RECT -21.245 150.795 -20.915 151.125 ;
        RECT -21.245 149.435 -20.915 149.765 ;
        RECT -21.245 148.075 -20.915 148.405 ;
        RECT -21.245 146.715 -20.915 147.045 ;
        RECT -21.245 145.355 -20.915 145.685 ;
        RECT -21.245 143.995 -20.915 144.325 ;
        RECT -21.245 142.635 -20.915 142.965 ;
        RECT -21.245 141.275 -20.915 141.605 ;
        RECT -21.245 139.915 -20.915 140.245 ;
        RECT -21.245 138.555 -20.915 138.885 ;
        RECT -21.245 137.195 -20.915 137.525 ;
        RECT -21.245 135.835 -20.915 136.165 ;
        RECT -21.245 134.475 -20.915 134.805 ;
        RECT -21.245 133.115 -20.915 133.445 ;
        RECT -21.245 131.755 -20.915 132.085 ;
        RECT -21.245 130.395 -20.915 130.725 ;
        RECT -21.245 129.035 -20.915 129.365 ;
        RECT -21.245 127.675 -20.915 128.005 ;
        RECT -21.245 126.315 -20.915 126.645 ;
        RECT -21.245 124.955 -20.915 125.285 ;
        RECT -21.245 123.595 -20.915 123.925 ;
        RECT -21.245 122.235 -20.915 122.565 ;
        RECT -21.245 120.875 -20.915 121.205 ;
        RECT -21.245 119.515 -20.915 119.845 ;
        RECT -21.245 118.155 -20.915 118.485 ;
        RECT -21.245 116.795 -20.915 117.125 ;
        RECT -21.245 115.435 -20.915 115.765 ;
        RECT -21.245 114.075 -20.915 114.405 ;
        RECT -21.245 112.715 -20.915 113.045 ;
        RECT -21.245 111.355 -20.915 111.685 ;
        RECT -21.245 109.995 -20.915 110.325 ;
        RECT -21.245 108.635 -20.915 108.965 ;
        RECT -21.245 107.275 -20.915 107.605 ;
        RECT -21.245 105.915 -20.915 106.245 ;
        RECT -21.245 104.555 -20.915 104.885 ;
        RECT -21.245 103.195 -20.915 103.525 ;
        RECT -21.245 101.835 -20.915 102.165 ;
        RECT -21.245 100.475 -20.915 100.805 ;
        RECT -21.245 99.115 -20.915 99.445 ;
        RECT -21.245 97.755 -20.915 98.085 ;
        RECT -21.245 96.395 -20.915 96.725 ;
        RECT -21.245 95.035 -20.915 95.365 ;
        RECT -21.245 93.675 -20.915 94.005 ;
        RECT -21.245 92.315 -20.915 92.645 ;
        RECT -21.245 90.955 -20.915 91.285 ;
        RECT -21.245 89.595 -20.915 89.925 ;
        RECT -21.245 88.235 -20.915 88.565 ;
        RECT -21.245 86.875 -20.915 87.205 ;
        RECT -21.245 85.515 -20.915 85.845 ;
        RECT -21.245 84.155 -20.915 84.485 ;
        RECT -21.245 82.795 -20.915 83.125 ;
        RECT -21.245 81.435 -20.915 81.765 ;
        RECT -21.245 80.075 -20.915 80.405 ;
        RECT -21.245 78.715 -20.915 79.045 ;
        RECT -21.245 77.355 -20.915 77.685 ;
        RECT -21.245 75.995 -20.915 76.325 ;
        RECT -21.245 74.635 -20.915 74.965 ;
        RECT -21.245 73.275 -20.915 73.605 ;
        RECT -21.245 71.915 -20.915 72.245 ;
        RECT -21.245 70.555 -20.915 70.885 ;
        RECT -21.245 69.195 -20.915 69.525 ;
        RECT -21.245 67.835 -20.915 68.165 ;
        RECT -21.245 66.475 -20.915 66.805 ;
        RECT -21.245 65.115 -20.915 65.445 ;
        RECT -21.245 63.755 -20.915 64.085 ;
        RECT -21.245 62.395 -20.915 62.725 ;
        RECT -21.245 61.035 -20.915 61.365 ;
        RECT -21.245 59.675 -20.915 60.005 ;
        RECT -21.245 58.315 -20.915 58.645 ;
        RECT -21.245 56.955 -20.915 57.285 ;
        RECT -21.245 55.595 -20.915 55.925 ;
        RECT -21.245 54.235 -20.915 54.565 ;
        RECT -21.245 52.875 -20.915 53.205 ;
        RECT -21.245 51.515 -20.915 51.845 ;
        RECT -21.245 50.155 -20.915 50.485 ;
        RECT -21.245 48.795 -20.915 49.125 ;
        RECT -21.245 47.435 -20.915 47.765 ;
        RECT -21.245 46.075 -20.915 46.405 ;
        RECT -21.245 44.715 -20.915 45.045 ;
        RECT -21.245 43.355 -20.915 43.685 ;
        RECT -21.245 41.995 -20.915 42.325 ;
        RECT -21.245 40.635 -20.915 40.965 ;
        RECT -21.245 39.275 -20.915 39.605 ;
        RECT -21.245 37.915 -20.915 38.245 ;
        RECT -21.245 36.555 -20.915 36.885 ;
        RECT -21.245 35.195 -20.915 35.525 ;
        RECT -21.245 33.835 -20.915 34.165 ;
        RECT -21.245 32.475 -20.915 32.805 ;
        RECT -21.245 31.115 -20.915 31.445 ;
        RECT -21.245 29.755 -20.915 30.085 ;
        RECT -21.245 28.395 -20.915 28.725 ;
        RECT -21.245 27.035 -20.915 27.365 ;
        RECT -21.245 25.675 -20.915 26.005 ;
        RECT -21.245 24.315 -20.915 24.645 ;
        RECT -21.245 22.955 -20.915 23.285 ;
        RECT -21.245 21.595 -20.915 21.925 ;
        RECT -21.245 20.235 -20.915 20.565 ;
        RECT -21.245 18.875 -20.915 19.205 ;
        RECT -21.245 17.515 -20.915 17.845 ;
        RECT -21.245 16.155 -20.915 16.485 ;
        RECT -21.245 14.795 -20.915 15.125 ;
        RECT -21.245 13.435 -20.915 13.765 ;
        RECT -21.245 12.075 -20.915 12.405 ;
        RECT -21.245 10.715 -20.915 11.045 ;
        RECT -21.245 9.355 -20.915 9.685 ;
        RECT -21.245 7.995 -20.915 8.325 ;
        RECT -21.245 6.635 -20.915 6.965 ;
        RECT -21.245 5.275 -20.915 5.605 ;
        RECT -21.245 3.915 -20.915 4.245 ;
        RECT -21.245 2.555 -20.915 2.885 ;
        RECT -21.245 1.195 -20.915 1.525 ;
        RECT -21.245 -0.165 -20.915 0.165 ;
        RECT -21.245 -2.885 -20.915 -2.555 ;
        RECT -21.245 -4.245 -20.915 -3.915 ;
        RECT -21.245 -8.325 -20.915 -7.995 ;
        RECT -21.245 -9.685 -20.915 -9.355 ;
        RECT -21.245 -14.95 -20.915 -14.62 ;
        RECT -21.245 -17.845 -20.915 -17.515 ;
        RECT -21.245 -19.79 -20.915 -19.46 ;
        RECT -21.245 -20.565 -20.915 -20.235 ;
        RECT -21.24 -23.28 -20.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 -30.085 -20.915 -29.755 ;
        RECT -21.245 -31.445 -20.915 -31.115 ;
        RECT -21.245 -32.805 -20.915 -32.475 ;
        RECT -21.245 -35.525 -20.915 -35.195 ;
        RECT -21.245 -36.885 -20.915 -36.555 ;
        RECT -21.245 -37.93 -20.915 -37.6 ;
        RECT -21.245 -40.965 -20.915 -40.635 ;
        RECT -21.245 -42.77 -20.915 -42.44 ;
        RECT -21.245 -43.685 -20.915 -43.355 ;
        RECT -21.245 -50.485 -20.915 -50.155 ;
        RECT -21.245 -51.845 -20.915 -51.515 ;
        RECT -21.245 -53.205 -20.915 -52.875 ;
        RECT -21.245 -54.565 -20.915 -54.235 ;
        RECT -21.245 -55.925 -20.915 -55.595 ;
        RECT -21.245 -57.285 -20.915 -56.955 ;
        RECT -21.245 -58.645 -20.915 -58.315 ;
        RECT -21.245 -60.005 -20.915 -59.675 ;
        RECT -21.245 -61.365 -20.915 -61.035 ;
        RECT -21.245 -62.725 -20.915 -62.395 ;
        RECT -21.245 -64.085 -20.915 -63.755 ;
        RECT -21.245 -65.445 -20.915 -65.115 ;
        RECT -21.245 -68.165 -20.915 -67.835 ;
        RECT -21.245 -69.525 -20.915 -69.195 ;
        RECT -21.245 -70.885 -20.915 -70.555 ;
        RECT -21.245 -72.245 -20.915 -71.915 ;
        RECT -21.245 -74.965 -20.915 -74.635 ;
        RECT -21.245 -76.71 -20.915 -76.38 ;
        RECT -21.245 -77.685 -20.915 -77.355 ;
        RECT -21.245 -79.045 -20.915 -78.715 ;
        RECT -21.245 -81.765 -20.915 -81.435 ;
        RECT -21.245 -83.125 -20.915 -82.795 ;
        RECT -21.245 -84.485 -20.915 -84.155 ;
        RECT -21.245 -85.25 -20.915 -84.92 ;
        RECT -21.245 -87.205 -20.915 -86.875 ;
        RECT -21.245 -89.925 -20.915 -89.595 ;
        RECT -21.245 -91.285 -20.915 -90.955 ;
        RECT -21.245 -92.645 -20.915 -92.315 ;
        RECT -21.245 -94.005 -20.915 -93.675 ;
        RECT -21.245 -96.725 -20.915 -96.395 ;
        RECT -21.245 -98.085 -20.915 -97.755 ;
        RECT -21.245 -98.89 -20.915 -98.56 ;
        RECT -21.245 -100.805 -20.915 -100.475 ;
        RECT -21.245 -102.165 -20.915 -101.835 ;
        RECT -21.245 -104.885 -20.915 -104.555 ;
        RECT -21.245 -107.43 -20.915 -107.1 ;
        RECT -21.24 -111 -20.92 -29.08 ;
    END
    PORT
      LAYER met3 ;
        RECT -21.245 -117.125 -20.915 -116.795 ;
        RECT -21.245 -118.485 -20.915 -118.155 ;
        RECT -21.245 -125.285 -20.915 -124.955 ;
        RECT -21.245 -126.645 -20.915 -126.315 ;
        RECT -21.245 -128.005 -20.915 -127.675 ;
        RECT -21.245 -130.725 -20.915 -130.395 ;
        RECT -21.245 -136.165 -20.915 -135.835 ;
        RECT -21.245 -141.605 -20.915 -141.275 ;
        RECT -21.245 -144.325 -20.915 -143.995 ;
        RECT -21.245 -147.045 -20.915 -146.715 ;
        RECT -21.245 -148.405 -20.915 -148.075 ;
        RECT -21.245 -149.765 -20.915 -149.435 ;
        RECT -21.245 -152.485 -20.915 -152.155 ;
        RECT -21.245 -153.845 -20.915 -153.515 ;
        RECT -21.245 -159.285 -20.915 -158.955 ;
        RECT -21.245 -160.645 -20.915 -160.315 ;
        RECT -21.245 -162.005 -20.915 -161.675 ;
        RECT -21.245 -163.365 -20.915 -163.035 ;
        RECT -21.245 -164.725 -20.915 -164.395 ;
        RECT -21.245 -166.085 -20.915 -165.755 ;
        RECT -21.245 -167.445 -20.915 -167.115 ;
        RECT -21.245 -168.805 -20.915 -168.475 ;
        RECT -21.245 -171.525 -20.915 -171.195 ;
        RECT -21.245 -172.885 -20.915 -172.555 ;
        RECT -21.24 -172.885 -20.92 -116.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -19.885 101.835 -19.555 102.165 ;
        RECT -19.885 100.475 -19.555 100.805 ;
        RECT -19.885 99.115 -19.555 99.445 ;
        RECT -19.885 97.755 -19.555 98.085 ;
        RECT -19.885 96.395 -19.555 96.725 ;
        RECT -19.885 95.035 -19.555 95.365 ;
        RECT -19.885 93.675 -19.555 94.005 ;
        RECT -19.885 92.315 -19.555 92.645 ;
        RECT -19.885 90.955 -19.555 91.285 ;
        RECT -19.885 89.595 -19.555 89.925 ;
        RECT -19.885 88.235 -19.555 88.565 ;
        RECT -19.885 86.875 -19.555 87.205 ;
        RECT -19.885 85.515 -19.555 85.845 ;
        RECT -19.885 84.155 -19.555 84.485 ;
        RECT -19.885 82.795 -19.555 83.125 ;
        RECT -19.885 81.435 -19.555 81.765 ;
        RECT -19.885 80.075 -19.555 80.405 ;
        RECT -19.885 78.715 -19.555 79.045 ;
        RECT -19.885 77.355 -19.555 77.685 ;
        RECT -19.885 75.995 -19.555 76.325 ;
        RECT -19.885 74.635 -19.555 74.965 ;
        RECT -19.885 73.275 -19.555 73.605 ;
        RECT -19.885 71.915 -19.555 72.245 ;
        RECT -19.885 70.555 -19.555 70.885 ;
        RECT -19.885 69.195 -19.555 69.525 ;
        RECT -19.885 67.835 -19.555 68.165 ;
        RECT -19.885 66.475 -19.555 66.805 ;
        RECT -19.885 65.115 -19.555 65.445 ;
        RECT -19.885 63.755 -19.555 64.085 ;
        RECT -19.885 62.395 -19.555 62.725 ;
        RECT -19.885 61.035 -19.555 61.365 ;
        RECT -19.885 59.675 -19.555 60.005 ;
        RECT -19.885 58.315 -19.555 58.645 ;
        RECT -19.885 56.955 -19.555 57.285 ;
        RECT -19.885 55.595 -19.555 55.925 ;
        RECT -19.885 54.235 -19.555 54.565 ;
        RECT -19.885 52.875 -19.555 53.205 ;
        RECT -19.885 51.515 -19.555 51.845 ;
        RECT -19.885 50.155 -19.555 50.485 ;
        RECT -19.885 48.795 -19.555 49.125 ;
        RECT -19.885 47.435 -19.555 47.765 ;
        RECT -19.885 46.075 -19.555 46.405 ;
        RECT -19.885 44.715 -19.555 45.045 ;
        RECT -19.885 43.355 -19.555 43.685 ;
        RECT -19.885 41.995 -19.555 42.325 ;
        RECT -19.885 40.635 -19.555 40.965 ;
        RECT -19.885 39.275 -19.555 39.605 ;
        RECT -19.885 37.915 -19.555 38.245 ;
        RECT -19.885 36.555 -19.555 36.885 ;
        RECT -19.885 35.195 -19.555 35.525 ;
        RECT -19.885 33.835 -19.555 34.165 ;
        RECT -19.885 32.475 -19.555 32.805 ;
        RECT -19.885 31.115 -19.555 31.445 ;
        RECT -19.885 29.755 -19.555 30.085 ;
        RECT -19.885 28.395 -19.555 28.725 ;
        RECT -19.885 27.035 -19.555 27.365 ;
        RECT -19.885 25.675 -19.555 26.005 ;
        RECT -19.885 24.315 -19.555 24.645 ;
        RECT -19.885 22.955 -19.555 23.285 ;
        RECT -19.885 21.595 -19.555 21.925 ;
        RECT -19.885 20.235 -19.555 20.565 ;
        RECT -19.885 18.875 -19.555 19.205 ;
        RECT -19.885 17.515 -19.555 17.845 ;
        RECT -19.885 16.155 -19.555 16.485 ;
        RECT -19.885 14.795 -19.555 15.125 ;
        RECT -19.885 13.435 -19.555 13.765 ;
        RECT -19.885 12.075 -19.555 12.405 ;
        RECT -19.885 10.715 -19.555 11.045 ;
        RECT -19.885 9.355 -19.555 9.685 ;
        RECT -19.885 7.995 -19.555 8.325 ;
        RECT -19.885 6.635 -19.555 6.965 ;
        RECT -19.885 5.275 -19.555 5.605 ;
        RECT -19.885 3.915 -19.555 4.245 ;
        RECT -19.885 2.555 -19.555 2.885 ;
        RECT -19.885 1.195 -19.555 1.525 ;
        RECT -19.885 -0.165 -19.555 0.165 ;
        RECT -19.885 -2.885 -19.555 -2.555 ;
        RECT -19.885 -4.245 -19.555 -3.915 ;
        RECT -19.885 -8.325 -19.555 -7.995 ;
        RECT -19.885 -9.685 -19.555 -9.355 ;
        RECT -19.885 -14.95 -19.555 -14.62 ;
        RECT -19.885 -17.845 -19.555 -17.515 ;
        RECT -19.885 -19.79 -19.555 -19.46 ;
        RECT -19.885 -20.565 -19.555 -20.235 ;
        RECT -19.88 -22.6 -19.56 242.565 ;
        RECT -19.885 241.32 -19.555 242.45 ;
        RECT -19.885 239.195 -19.555 239.525 ;
        RECT -19.885 237.835 -19.555 238.165 ;
        RECT -19.885 236.475 -19.555 236.805 ;
        RECT -19.885 235.115 -19.555 235.445 ;
        RECT -19.885 233.755 -19.555 234.085 ;
        RECT -19.885 232.395 -19.555 232.725 ;
        RECT -19.885 231.035 -19.555 231.365 ;
        RECT -19.885 229.675 -19.555 230.005 ;
        RECT -19.885 228.315 -19.555 228.645 ;
        RECT -19.885 226.955 -19.555 227.285 ;
        RECT -19.885 225.595 -19.555 225.925 ;
        RECT -19.885 224.235 -19.555 224.565 ;
        RECT -19.885 222.875 -19.555 223.205 ;
        RECT -19.885 221.515 -19.555 221.845 ;
        RECT -19.885 220.155 -19.555 220.485 ;
        RECT -19.885 218.795 -19.555 219.125 ;
        RECT -19.885 217.435 -19.555 217.765 ;
        RECT -19.885 216.075 -19.555 216.405 ;
        RECT -19.885 214.715 -19.555 215.045 ;
        RECT -19.885 213.355 -19.555 213.685 ;
        RECT -19.885 211.995 -19.555 212.325 ;
        RECT -19.885 210.635 -19.555 210.965 ;
        RECT -19.885 209.275 -19.555 209.605 ;
        RECT -19.885 207.915 -19.555 208.245 ;
        RECT -19.885 206.555 -19.555 206.885 ;
        RECT -19.885 205.195 -19.555 205.525 ;
        RECT -19.885 203.835 -19.555 204.165 ;
        RECT -19.885 202.475 -19.555 202.805 ;
        RECT -19.885 201.115 -19.555 201.445 ;
        RECT -19.885 199.755 -19.555 200.085 ;
        RECT -19.885 198.395 -19.555 198.725 ;
        RECT -19.885 197.035 -19.555 197.365 ;
        RECT -19.885 195.675 -19.555 196.005 ;
        RECT -19.885 194.315 -19.555 194.645 ;
        RECT -19.885 192.955 -19.555 193.285 ;
        RECT -19.885 191.595 -19.555 191.925 ;
        RECT -19.885 190.235 -19.555 190.565 ;
        RECT -19.885 188.875 -19.555 189.205 ;
        RECT -19.885 187.515 -19.555 187.845 ;
        RECT -19.885 186.155 -19.555 186.485 ;
        RECT -19.885 184.795 -19.555 185.125 ;
        RECT -19.885 183.435 -19.555 183.765 ;
        RECT -19.885 182.075 -19.555 182.405 ;
        RECT -19.885 180.715 -19.555 181.045 ;
        RECT -19.885 179.355 -19.555 179.685 ;
        RECT -19.885 177.995 -19.555 178.325 ;
        RECT -19.885 176.635 -19.555 176.965 ;
        RECT -19.885 175.275 -19.555 175.605 ;
        RECT -19.885 173.915 -19.555 174.245 ;
        RECT -19.885 172.555 -19.555 172.885 ;
        RECT -19.885 171.195 -19.555 171.525 ;
        RECT -19.885 169.835 -19.555 170.165 ;
        RECT -19.885 168.475 -19.555 168.805 ;
        RECT -19.885 167.115 -19.555 167.445 ;
        RECT -19.885 165.755 -19.555 166.085 ;
        RECT -19.885 164.395 -19.555 164.725 ;
        RECT -19.885 163.035 -19.555 163.365 ;
        RECT -19.885 161.675 -19.555 162.005 ;
        RECT -19.885 160.315 -19.555 160.645 ;
        RECT -19.885 158.955 -19.555 159.285 ;
        RECT -19.885 157.595 -19.555 157.925 ;
        RECT -19.885 156.235 -19.555 156.565 ;
        RECT -19.885 154.875 -19.555 155.205 ;
        RECT -19.885 153.515 -19.555 153.845 ;
        RECT -19.885 152.155 -19.555 152.485 ;
        RECT -19.885 150.795 -19.555 151.125 ;
        RECT -19.885 149.435 -19.555 149.765 ;
        RECT -19.885 148.075 -19.555 148.405 ;
        RECT -19.885 146.715 -19.555 147.045 ;
        RECT -19.885 145.355 -19.555 145.685 ;
        RECT -19.885 143.995 -19.555 144.325 ;
        RECT -19.885 142.635 -19.555 142.965 ;
        RECT -19.885 141.275 -19.555 141.605 ;
        RECT -19.885 139.915 -19.555 140.245 ;
        RECT -19.885 138.555 -19.555 138.885 ;
        RECT -19.885 137.195 -19.555 137.525 ;
        RECT -19.885 135.835 -19.555 136.165 ;
        RECT -19.885 134.475 -19.555 134.805 ;
        RECT -19.885 133.115 -19.555 133.445 ;
        RECT -19.885 131.755 -19.555 132.085 ;
        RECT -19.885 130.395 -19.555 130.725 ;
        RECT -19.885 129.035 -19.555 129.365 ;
        RECT -19.885 127.675 -19.555 128.005 ;
        RECT -19.885 126.315 -19.555 126.645 ;
        RECT -19.885 124.955 -19.555 125.285 ;
        RECT -19.885 123.595 -19.555 123.925 ;
        RECT -19.885 122.235 -19.555 122.565 ;
        RECT -19.885 120.875 -19.555 121.205 ;
        RECT -19.885 119.515 -19.555 119.845 ;
        RECT -19.885 118.155 -19.555 118.485 ;
        RECT -19.885 116.795 -19.555 117.125 ;
        RECT -19.885 115.435 -19.555 115.765 ;
        RECT -19.885 114.075 -19.555 114.405 ;
        RECT -19.885 112.715 -19.555 113.045 ;
        RECT -19.885 111.355 -19.555 111.685 ;
        RECT -19.885 109.995 -19.555 110.325 ;
        RECT -19.885 108.635 -19.555 108.965 ;
        RECT -19.885 107.275 -19.555 107.605 ;
        RECT -19.885 105.915 -19.555 106.245 ;
        RECT -19.885 104.555 -19.555 104.885 ;
        RECT -19.885 103.195 -19.555 103.525 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.765 -69.525 -30.435 -69.195 ;
        RECT -30.765 -70.885 -30.435 -70.555 ;
        RECT -30.765 -72.245 -30.435 -71.915 ;
        RECT -30.765 -73.605 -30.435 -73.275 ;
        RECT -30.765 -74.965 -30.435 -74.635 ;
        RECT -30.765 -76.325 -30.435 -75.995 ;
        RECT -30.765 -77.685 -30.435 -77.355 ;
        RECT -30.765 -79.045 -30.435 -78.715 ;
        RECT -30.765 -80.405 -30.435 -80.075 ;
        RECT -30.765 -81.765 -30.435 -81.435 ;
        RECT -30.765 -83.125 -30.435 -82.795 ;
        RECT -30.765 -84.485 -30.435 -84.155 ;
        RECT -30.765 -85.845 -30.435 -85.515 ;
        RECT -30.765 -87.205 -30.435 -86.875 ;
        RECT -30.76 -87.88 -30.44 -67.84 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.765 -123.925 -30.435 -123.595 ;
        RECT -30.765 -125.285 -30.435 -124.955 ;
        RECT -30.765 -126.645 -30.435 -126.315 ;
        RECT -30.765 -128.005 -30.435 -127.675 ;
        RECT -30.765 -129.365 -30.435 -129.035 ;
        RECT -30.765 -130.725 -30.435 -130.395 ;
        RECT -30.765 -133.445 -30.435 -133.115 ;
        RECT -30.765 -134.805 -30.435 -134.475 ;
        RECT -30.765 -136.165 -30.435 -135.835 ;
        RECT -30.765 -137.525 -30.435 -137.195 ;
        RECT -30.765 -141.605 -30.435 -141.275 ;
        RECT -30.765 -142.965 -30.435 -142.635 ;
        RECT -30.765 -144.325 -30.435 -143.995 ;
        RECT -30.765 -145.685 -30.435 -145.355 ;
        RECT -30.765 -147.045 -30.435 -146.715 ;
        RECT -30.765 -148.405 -30.435 -148.075 ;
        RECT -30.765 -149.765 -30.435 -149.435 ;
        RECT -30.765 -152.485 -30.435 -152.155 ;
        RECT -30.765 -153.845 -30.435 -153.515 ;
        RECT -30.765 -157.925 -30.435 -157.595 ;
        RECT -30.765 -159.285 -30.435 -158.955 ;
        RECT -30.765 -160.645 -30.435 -160.315 ;
        RECT -30.765 -162.005 -30.435 -161.675 ;
        RECT -30.765 -163.365 -30.435 -163.035 ;
        RECT -30.765 -164.725 -30.435 -164.395 ;
        RECT -30.765 -166.085 -30.435 -165.755 ;
        RECT -30.765 -167.445 -30.435 -167.115 ;
        RECT -30.765 -168.805 -30.435 -168.475 ;
        RECT -30.765 -171.525 -30.435 -171.195 ;
        RECT -30.765 -172.885 -30.435 -172.555 ;
        RECT -30.765 -174.245 -30.435 -173.915 ;
        RECT -30.765 -175.605 -30.435 -175.275 ;
        RECT -30.765 -176.685 -30.435 -176.355 ;
        RECT -30.765 -178.325 -30.435 -177.995 ;
        RECT -30.765 -179.685 -30.435 -179.355 ;
        RECT -30.765 -181.93 -30.435 -180.8 ;
        RECT -30.76 -182.045 -30.44 -121.56 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 241.32 -29.075 242.45 ;
        RECT -29.405 239.195 -29.075 239.525 ;
        RECT -29.405 237.835 -29.075 238.165 ;
        RECT -29.405 236.475 -29.075 236.805 ;
        RECT -29.405 235.115 -29.075 235.445 ;
        RECT -29.405 233.755 -29.075 234.085 ;
        RECT -29.405 232.395 -29.075 232.725 ;
        RECT -29.405 231.035 -29.075 231.365 ;
        RECT -29.405 229.675 -29.075 230.005 ;
        RECT -29.405 228.315 -29.075 228.645 ;
        RECT -29.405 226.955 -29.075 227.285 ;
        RECT -29.405 225.595 -29.075 225.925 ;
        RECT -29.405 224.235 -29.075 224.565 ;
        RECT -29.405 222.875 -29.075 223.205 ;
        RECT -29.405 221.515 -29.075 221.845 ;
        RECT -29.405 220.155 -29.075 220.485 ;
        RECT -29.405 218.795 -29.075 219.125 ;
        RECT -29.405 217.435 -29.075 217.765 ;
        RECT -29.405 216.075 -29.075 216.405 ;
        RECT -29.405 214.715 -29.075 215.045 ;
        RECT -29.405 213.355 -29.075 213.685 ;
        RECT -29.405 211.995 -29.075 212.325 ;
        RECT -29.405 210.635 -29.075 210.965 ;
        RECT -29.405 209.275 -29.075 209.605 ;
        RECT -29.405 207.915 -29.075 208.245 ;
        RECT -29.405 206.555 -29.075 206.885 ;
        RECT -29.405 205.195 -29.075 205.525 ;
        RECT -29.405 203.835 -29.075 204.165 ;
        RECT -29.405 202.475 -29.075 202.805 ;
        RECT -29.405 201.115 -29.075 201.445 ;
        RECT -29.405 199.755 -29.075 200.085 ;
        RECT -29.405 198.395 -29.075 198.725 ;
        RECT -29.405 197.035 -29.075 197.365 ;
        RECT -29.405 195.675 -29.075 196.005 ;
        RECT -29.405 194.315 -29.075 194.645 ;
        RECT -29.405 192.955 -29.075 193.285 ;
        RECT -29.405 191.595 -29.075 191.925 ;
        RECT -29.405 190.235 -29.075 190.565 ;
        RECT -29.405 188.875 -29.075 189.205 ;
        RECT -29.405 187.515 -29.075 187.845 ;
        RECT -29.405 186.155 -29.075 186.485 ;
        RECT -29.405 184.795 -29.075 185.125 ;
        RECT -29.405 183.435 -29.075 183.765 ;
        RECT -29.405 182.075 -29.075 182.405 ;
        RECT -29.405 180.715 -29.075 181.045 ;
        RECT -29.405 179.355 -29.075 179.685 ;
        RECT -29.405 177.995 -29.075 178.325 ;
        RECT -29.405 176.635 -29.075 176.965 ;
        RECT -29.405 175.275 -29.075 175.605 ;
        RECT -29.405 173.915 -29.075 174.245 ;
        RECT -29.405 172.555 -29.075 172.885 ;
        RECT -29.405 171.195 -29.075 171.525 ;
        RECT -29.405 169.835 -29.075 170.165 ;
        RECT -29.405 168.475 -29.075 168.805 ;
        RECT -29.405 167.115 -29.075 167.445 ;
        RECT -29.405 165.755 -29.075 166.085 ;
        RECT -29.405 164.395 -29.075 164.725 ;
        RECT -29.405 163.035 -29.075 163.365 ;
        RECT -29.405 161.675 -29.075 162.005 ;
        RECT -29.405 160.315 -29.075 160.645 ;
        RECT -29.405 158.955 -29.075 159.285 ;
        RECT -29.405 157.595 -29.075 157.925 ;
        RECT -29.405 156.235 -29.075 156.565 ;
        RECT -29.405 154.875 -29.075 155.205 ;
        RECT -29.405 153.515 -29.075 153.845 ;
        RECT -29.405 152.155 -29.075 152.485 ;
        RECT -29.405 150.795 -29.075 151.125 ;
        RECT -29.405 149.435 -29.075 149.765 ;
        RECT -29.405 148.075 -29.075 148.405 ;
        RECT -29.405 146.715 -29.075 147.045 ;
        RECT -29.405 145.355 -29.075 145.685 ;
        RECT -29.405 143.995 -29.075 144.325 ;
        RECT -29.405 142.635 -29.075 142.965 ;
        RECT -29.405 141.275 -29.075 141.605 ;
        RECT -29.405 139.915 -29.075 140.245 ;
        RECT -29.405 138.555 -29.075 138.885 ;
        RECT -29.405 137.195 -29.075 137.525 ;
        RECT -29.405 135.835 -29.075 136.165 ;
        RECT -29.405 134.475 -29.075 134.805 ;
        RECT -29.405 133.115 -29.075 133.445 ;
        RECT -29.405 131.755 -29.075 132.085 ;
        RECT -29.405 130.395 -29.075 130.725 ;
        RECT -29.405 129.035 -29.075 129.365 ;
        RECT -29.405 127.675 -29.075 128.005 ;
        RECT -29.405 126.315 -29.075 126.645 ;
        RECT -29.405 124.955 -29.075 125.285 ;
        RECT -29.405 123.595 -29.075 123.925 ;
        RECT -29.405 122.235 -29.075 122.565 ;
        RECT -29.405 120.875 -29.075 121.205 ;
        RECT -29.405 119.515 -29.075 119.845 ;
        RECT -29.405 118.155 -29.075 118.485 ;
        RECT -29.405 116.795 -29.075 117.125 ;
        RECT -29.405 115.435 -29.075 115.765 ;
        RECT -29.405 114.075 -29.075 114.405 ;
        RECT -29.405 112.715 -29.075 113.045 ;
        RECT -29.405 111.355 -29.075 111.685 ;
        RECT -29.405 109.995 -29.075 110.325 ;
        RECT -29.405 108.635 -29.075 108.965 ;
        RECT -29.405 107.275 -29.075 107.605 ;
        RECT -29.405 105.915 -29.075 106.245 ;
        RECT -29.405 104.555 -29.075 104.885 ;
        RECT -29.405 103.195 -29.075 103.525 ;
        RECT -29.405 101.835 -29.075 102.165 ;
        RECT -29.405 100.475 -29.075 100.805 ;
        RECT -29.405 99.115 -29.075 99.445 ;
        RECT -29.405 97.755 -29.075 98.085 ;
        RECT -29.405 96.395 -29.075 96.725 ;
        RECT -29.405 95.035 -29.075 95.365 ;
        RECT -29.405 93.675 -29.075 94.005 ;
        RECT -29.405 92.315 -29.075 92.645 ;
        RECT -29.405 90.955 -29.075 91.285 ;
        RECT -29.405 89.595 -29.075 89.925 ;
        RECT -29.405 88.235 -29.075 88.565 ;
        RECT -29.405 86.875 -29.075 87.205 ;
        RECT -29.405 85.515 -29.075 85.845 ;
        RECT -29.405 84.155 -29.075 84.485 ;
        RECT -29.405 82.795 -29.075 83.125 ;
        RECT -29.405 81.435 -29.075 81.765 ;
        RECT -29.405 80.075 -29.075 80.405 ;
        RECT -29.405 78.715 -29.075 79.045 ;
        RECT -29.405 77.355 -29.075 77.685 ;
        RECT -29.405 75.995 -29.075 76.325 ;
        RECT -29.405 74.635 -29.075 74.965 ;
        RECT -29.405 73.275 -29.075 73.605 ;
        RECT -29.405 71.915 -29.075 72.245 ;
        RECT -29.405 70.555 -29.075 70.885 ;
        RECT -29.405 69.195 -29.075 69.525 ;
        RECT -29.405 67.835 -29.075 68.165 ;
        RECT -29.405 66.475 -29.075 66.805 ;
        RECT -29.405 65.115 -29.075 65.445 ;
        RECT -29.405 63.755 -29.075 64.085 ;
        RECT -29.405 62.395 -29.075 62.725 ;
        RECT -29.405 61.035 -29.075 61.365 ;
        RECT -29.405 59.675 -29.075 60.005 ;
        RECT -29.405 58.315 -29.075 58.645 ;
        RECT -29.405 56.955 -29.075 57.285 ;
        RECT -29.405 55.595 -29.075 55.925 ;
        RECT -29.405 54.235 -29.075 54.565 ;
        RECT -29.405 52.875 -29.075 53.205 ;
        RECT -29.405 51.515 -29.075 51.845 ;
        RECT -29.405 50.155 -29.075 50.485 ;
        RECT -29.405 48.795 -29.075 49.125 ;
        RECT -29.405 47.435 -29.075 47.765 ;
        RECT -29.405 46.075 -29.075 46.405 ;
        RECT -29.405 44.715 -29.075 45.045 ;
        RECT -29.405 43.355 -29.075 43.685 ;
        RECT -29.405 41.995 -29.075 42.325 ;
        RECT -29.405 40.635 -29.075 40.965 ;
        RECT -29.405 39.275 -29.075 39.605 ;
        RECT -29.405 37.915 -29.075 38.245 ;
        RECT -29.405 36.555 -29.075 36.885 ;
        RECT -29.405 35.195 -29.075 35.525 ;
        RECT -29.405 33.835 -29.075 34.165 ;
        RECT -29.405 32.475 -29.075 32.805 ;
        RECT -29.405 31.115 -29.075 31.445 ;
        RECT -29.405 29.755 -29.075 30.085 ;
        RECT -29.405 28.395 -29.075 28.725 ;
        RECT -29.405 27.035 -29.075 27.365 ;
        RECT -29.405 25.675 -29.075 26.005 ;
        RECT -29.405 24.315 -29.075 24.645 ;
        RECT -29.405 22.955 -29.075 23.285 ;
        RECT -29.405 21.595 -29.075 21.925 ;
        RECT -29.405 20.235 -29.075 20.565 ;
        RECT -29.405 18.875 -29.075 19.205 ;
        RECT -29.405 17.515 -29.075 17.845 ;
        RECT -29.405 16.155 -29.075 16.485 ;
        RECT -29.405 14.795 -29.075 15.125 ;
        RECT -29.405 13.435 -29.075 13.765 ;
        RECT -29.405 12.075 -29.075 12.405 ;
        RECT -29.405 10.715 -29.075 11.045 ;
        RECT -29.405 9.355 -29.075 9.685 ;
        RECT -29.405 7.995 -29.075 8.325 ;
        RECT -29.405 6.635 -29.075 6.965 ;
        RECT -29.405 5.275 -29.075 5.605 ;
        RECT -29.405 3.915 -29.075 4.245 ;
        RECT -29.405 2.555 -29.075 2.885 ;
        RECT -29.405 1.195 -29.075 1.525 ;
        RECT -29.405 -0.165 -29.075 0.165 ;
        RECT -29.405 -8.325 -29.075 -7.995 ;
        RECT -29.405 -9.685 -29.075 -9.355 ;
        RECT -29.405 -14.95 -29.075 -14.62 ;
        RECT -29.405 -17.845 -29.075 -17.515 ;
        RECT -29.405 -19.79 -29.075 -19.46 ;
        RECT -29.405 -20.565 -29.075 -20.235 ;
        RECT -29.405 -32.805 -29.075 -32.475 ;
        RECT -29.405 -35.525 -29.075 -35.195 ;
        RECT -29.405 -36.885 -29.075 -36.555 ;
        RECT -29.405 -37.93 -29.075 -37.6 ;
        RECT -29.405 -40.965 -29.075 -40.635 ;
        RECT -29.405 -42.77 -29.075 -42.44 ;
        RECT -29.405 -43.685 -29.075 -43.355 ;
        RECT -29.405 -50.485 -29.075 -50.155 ;
        RECT -29.405 -51.845 -29.075 -51.515 ;
        RECT -29.405 -54.565 -29.075 -54.235 ;
        RECT -29.405 -55.925 -29.075 -55.595 ;
        RECT -29.405 -60.005 -29.075 -59.675 ;
        RECT -29.405 -62.725 -29.075 -62.395 ;
        RECT -29.4 -64.08 -29.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 -69.525 -29.075 -69.195 ;
        RECT -29.405 -70.885 -29.075 -70.555 ;
        RECT -29.405 -72.245 -29.075 -71.915 ;
        RECT -29.405 -74.965 -29.075 -74.635 ;
        RECT -29.405 -76.71 -29.075 -76.38 ;
        RECT -29.405 -77.685 -29.075 -77.355 ;
        RECT -29.405 -79.045 -29.075 -78.715 ;
        RECT -29.405 -81.765 -29.075 -81.435 ;
        RECT -29.405 -83.125 -29.075 -82.795 ;
        RECT -29.405 -84.485 -29.075 -84.155 ;
        RECT -29.405 -85.25 -29.075 -84.92 ;
        RECT -29.405 -87.205 -29.075 -86.875 ;
        RECT -29.405 -89.925 -29.075 -89.595 ;
        RECT -29.405 -91.285 -29.075 -90.955 ;
        RECT -29.405 -92.645 -29.075 -92.315 ;
        RECT -29.405 -94.005 -29.075 -93.675 ;
        RECT -29.405 -96.725 -29.075 -96.395 ;
        RECT -29.405 -98.085 -29.075 -97.755 ;
        RECT -29.405 -98.89 -29.075 -98.56 ;
        RECT -29.405 -100.805 -29.075 -100.475 ;
        RECT -29.405 -102.165 -29.075 -101.835 ;
        RECT -29.405 -104.885 -29.075 -104.555 ;
        RECT -29.405 -106.245 -29.075 -105.915 ;
        RECT -29.405 -107.43 -29.075 -107.1 ;
        RECT -29.405 -108.965 -29.075 -108.635 ;
        RECT -29.4 -113.04 -29.08 -68.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -29.405 -175.605 -29.075 -175.275 ;
        RECT -29.405 -176.685 -29.075 -176.355 ;
        RECT -29.405 -178.325 -29.075 -177.995 ;
        RECT -29.405 -179.685 -29.075 -179.355 ;
        RECT -29.405 -181.93 -29.075 -180.8 ;
        RECT -29.4 -182.045 -29.08 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -28.045 241.32 -27.715 242.45 ;
        RECT -28.045 239.195 -27.715 239.525 ;
        RECT -28.045 237.835 -27.715 238.165 ;
        RECT -28.045 236.475 -27.715 236.805 ;
        RECT -28.045 235.115 -27.715 235.445 ;
        RECT -28.045 233.755 -27.715 234.085 ;
        RECT -28.045 232.395 -27.715 232.725 ;
        RECT -28.045 231.035 -27.715 231.365 ;
        RECT -28.045 229.675 -27.715 230.005 ;
        RECT -28.045 228.315 -27.715 228.645 ;
        RECT -28.045 226.955 -27.715 227.285 ;
        RECT -28.045 225.595 -27.715 225.925 ;
        RECT -28.045 224.235 -27.715 224.565 ;
        RECT -28.045 222.875 -27.715 223.205 ;
        RECT -28.045 221.515 -27.715 221.845 ;
        RECT -28.045 220.155 -27.715 220.485 ;
        RECT -28.045 218.795 -27.715 219.125 ;
        RECT -28.045 217.435 -27.715 217.765 ;
        RECT -28.045 216.075 -27.715 216.405 ;
        RECT -28.045 214.715 -27.715 215.045 ;
        RECT -28.045 213.355 -27.715 213.685 ;
        RECT -28.045 211.995 -27.715 212.325 ;
        RECT -28.045 210.635 -27.715 210.965 ;
        RECT -28.045 209.275 -27.715 209.605 ;
        RECT -28.045 207.915 -27.715 208.245 ;
        RECT -28.045 206.555 -27.715 206.885 ;
        RECT -28.045 205.195 -27.715 205.525 ;
        RECT -28.045 203.835 -27.715 204.165 ;
        RECT -28.045 202.475 -27.715 202.805 ;
        RECT -28.045 201.115 -27.715 201.445 ;
        RECT -28.045 199.755 -27.715 200.085 ;
        RECT -28.045 198.395 -27.715 198.725 ;
        RECT -28.045 197.035 -27.715 197.365 ;
        RECT -28.045 195.675 -27.715 196.005 ;
        RECT -28.045 194.315 -27.715 194.645 ;
        RECT -28.045 192.955 -27.715 193.285 ;
        RECT -28.045 191.595 -27.715 191.925 ;
        RECT -28.045 190.235 -27.715 190.565 ;
        RECT -28.045 188.875 -27.715 189.205 ;
        RECT -28.045 187.515 -27.715 187.845 ;
        RECT -28.045 186.155 -27.715 186.485 ;
        RECT -28.045 184.795 -27.715 185.125 ;
        RECT -28.045 183.435 -27.715 183.765 ;
        RECT -28.045 182.075 -27.715 182.405 ;
        RECT -28.045 180.715 -27.715 181.045 ;
        RECT -28.045 179.355 -27.715 179.685 ;
        RECT -28.045 177.995 -27.715 178.325 ;
        RECT -28.045 176.635 -27.715 176.965 ;
        RECT -28.045 175.275 -27.715 175.605 ;
        RECT -28.045 173.915 -27.715 174.245 ;
        RECT -28.045 172.555 -27.715 172.885 ;
        RECT -28.045 171.195 -27.715 171.525 ;
        RECT -28.045 169.835 -27.715 170.165 ;
        RECT -28.045 168.475 -27.715 168.805 ;
        RECT -28.045 167.115 -27.715 167.445 ;
        RECT -28.045 165.755 -27.715 166.085 ;
        RECT -28.045 164.395 -27.715 164.725 ;
        RECT -28.045 163.035 -27.715 163.365 ;
        RECT -28.045 161.675 -27.715 162.005 ;
        RECT -28.045 160.315 -27.715 160.645 ;
        RECT -28.045 158.955 -27.715 159.285 ;
        RECT -28.045 157.595 -27.715 157.925 ;
        RECT -28.045 156.235 -27.715 156.565 ;
        RECT -28.045 154.875 -27.715 155.205 ;
        RECT -28.045 153.515 -27.715 153.845 ;
        RECT -28.045 152.155 -27.715 152.485 ;
        RECT -28.045 150.795 -27.715 151.125 ;
        RECT -28.045 149.435 -27.715 149.765 ;
        RECT -28.045 148.075 -27.715 148.405 ;
        RECT -28.045 146.715 -27.715 147.045 ;
        RECT -28.045 145.355 -27.715 145.685 ;
        RECT -28.045 143.995 -27.715 144.325 ;
        RECT -28.045 142.635 -27.715 142.965 ;
        RECT -28.045 141.275 -27.715 141.605 ;
        RECT -28.045 139.915 -27.715 140.245 ;
        RECT -28.045 138.555 -27.715 138.885 ;
        RECT -28.045 137.195 -27.715 137.525 ;
        RECT -28.045 135.835 -27.715 136.165 ;
        RECT -28.045 134.475 -27.715 134.805 ;
        RECT -28.045 133.115 -27.715 133.445 ;
        RECT -28.045 131.755 -27.715 132.085 ;
        RECT -28.045 130.395 -27.715 130.725 ;
        RECT -28.045 129.035 -27.715 129.365 ;
        RECT -28.045 127.675 -27.715 128.005 ;
        RECT -28.045 126.315 -27.715 126.645 ;
        RECT -28.045 124.955 -27.715 125.285 ;
        RECT -28.045 123.595 -27.715 123.925 ;
        RECT -28.045 122.235 -27.715 122.565 ;
        RECT -28.045 120.875 -27.715 121.205 ;
        RECT -28.045 119.515 -27.715 119.845 ;
        RECT -28.045 118.155 -27.715 118.485 ;
        RECT -28.045 116.795 -27.715 117.125 ;
        RECT -28.045 115.435 -27.715 115.765 ;
        RECT -28.045 114.075 -27.715 114.405 ;
        RECT -28.045 112.715 -27.715 113.045 ;
        RECT -28.045 111.355 -27.715 111.685 ;
        RECT -28.045 109.995 -27.715 110.325 ;
        RECT -28.045 108.635 -27.715 108.965 ;
        RECT -28.045 107.275 -27.715 107.605 ;
        RECT -28.045 105.915 -27.715 106.245 ;
        RECT -28.045 104.555 -27.715 104.885 ;
        RECT -28.045 103.195 -27.715 103.525 ;
        RECT -28.045 101.835 -27.715 102.165 ;
        RECT -28.045 100.475 -27.715 100.805 ;
        RECT -28.045 99.115 -27.715 99.445 ;
        RECT -28.045 97.755 -27.715 98.085 ;
        RECT -28.045 96.395 -27.715 96.725 ;
        RECT -28.045 95.035 -27.715 95.365 ;
        RECT -28.045 93.675 -27.715 94.005 ;
        RECT -28.045 92.315 -27.715 92.645 ;
        RECT -28.045 90.955 -27.715 91.285 ;
        RECT -28.045 89.595 -27.715 89.925 ;
        RECT -28.045 88.235 -27.715 88.565 ;
        RECT -28.045 86.875 -27.715 87.205 ;
        RECT -28.045 85.515 -27.715 85.845 ;
        RECT -28.045 84.155 -27.715 84.485 ;
        RECT -28.045 82.795 -27.715 83.125 ;
        RECT -28.045 81.435 -27.715 81.765 ;
        RECT -28.045 80.075 -27.715 80.405 ;
        RECT -28.045 78.715 -27.715 79.045 ;
        RECT -28.045 77.355 -27.715 77.685 ;
        RECT -28.045 75.995 -27.715 76.325 ;
        RECT -28.045 74.635 -27.715 74.965 ;
        RECT -28.045 73.275 -27.715 73.605 ;
        RECT -28.045 71.915 -27.715 72.245 ;
        RECT -28.045 70.555 -27.715 70.885 ;
        RECT -28.045 69.195 -27.715 69.525 ;
        RECT -28.045 67.835 -27.715 68.165 ;
        RECT -28.045 66.475 -27.715 66.805 ;
        RECT -28.045 65.115 -27.715 65.445 ;
        RECT -28.045 63.755 -27.715 64.085 ;
        RECT -28.045 62.395 -27.715 62.725 ;
        RECT -28.045 61.035 -27.715 61.365 ;
        RECT -28.045 59.675 -27.715 60.005 ;
        RECT -28.045 58.315 -27.715 58.645 ;
        RECT -28.045 56.955 -27.715 57.285 ;
        RECT -28.045 55.595 -27.715 55.925 ;
        RECT -28.045 54.235 -27.715 54.565 ;
        RECT -28.045 52.875 -27.715 53.205 ;
        RECT -28.045 51.515 -27.715 51.845 ;
        RECT -28.045 50.155 -27.715 50.485 ;
        RECT -28.045 48.795 -27.715 49.125 ;
        RECT -28.045 47.435 -27.715 47.765 ;
        RECT -28.045 46.075 -27.715 46.405 ;
        RECT -28.045 44.715 -27.715 45.045 ;
        RECT -28.045 43.355 -27.715 43.685 ;
        RECT -28.045 41.995 -27.715 42.325 ;
        RECT -28.045 40.635 -27.715 40.965 ;
        RECT -28.045 39.275 -27.715 39.605 ;
        RECT -28.045 37.915 -27.715 38.245 ;
        RECT -28.045 36.555 -27.715 36.885 ;
        RECT -28.045 35.195 -27.715 35.525 ;
        RECT -28.045 33.835 -27.715 34.165 ;
        RECT -28.045 32.475 -27.715 32.805 ;
        RECT -28.045 31.115 -27.715 31.445 ;
        RECT -28.045 29.755 -27.715 30.085 ;
        RECT -28.045 28.395 -27.715 28.725 ;
        RECT -28.045 27.035 -27.715 27.365 ;
        RECT -28.045 25.675 -27.715 26.005 ;
        RECT -28.045 24.315 -27.715 24.645 ;
        RECT -28.045 22.955 -27.715 23.285 ;
        RECT -28.045 21.595 -27.715 21.925 ;
        RECT -28.045 20.235 -27.715 20.565 ;
        RECT -28.045 18.875 -27.715 19.205 ;
        RECT -28.045 17.515 -27.715 17.845 ;
        RECT -28.045 16.155 -27.715 16.485 ;
        RECT -28.045 14.795 -27.715 15.125 ;
        RECT -28.045 13.435 -27.715 13.765 ;
        RECT -28.045 12.075 -27.715 12.405 ;
        RECT -28.045 10.715 -27.715 11.045 ;
        RECT -28.045 9.355 -27.715 9.685 ;
        RECT -28.045 7.995 -27.715 8.325 ;
        RECT -28.045 6.635 -27.715 6.965 ;
        RECT -28.045 5.275 -27.715 5.605 ;
        RECT -28.045 3.915 -27.715 4.245 ;
        RECT -28.045 2.555 -27.715 2.885 ;
        RECT -28.045 1.195 -27.715 1.525 ;
        RECT -28.045 -0.165 -27.715 0.165 ;
        RECT -28.045 -8.325 -27.715 -7.995 ;
        RECT -28.045 -9.685 -27.715 -9.355 ;
        RECT -28.045 -14.95 -27.715 -14.62 ;
        RECT -28.045 -17.845 -27.715 -17.515 ;
        RECT -28.045 -19.79 -27.715 -19.46 ;
        RECT -28.045 -20.565 -27.715 -20.235 ;
        RECT -28.045 -32.805 -27.715 -32.475 ;
        RECT -28.045 -35.525 -27.715 -35.195 ;
        RECT -28.045 -36.885 -27.715 -36.555 ;
        RECT -28.045 -37.93 -27.715 -37.6 ;
        RECT -28.045 -40.965 -27.715 -40.635 ;
        RECT -28.045 -42.77 -27.715 -42.44 ;
        RECT -28.045 -43.685 -27.715 -43.355 ;
        RECT -28.045 -50.485 -27.715 -50.155 ;
        RECT -28.045 -51.845 -27.715 -51.515 ;
        RECT -28.045 -54.565 -27.715 -54.235 ;
        RECT -28.045 -55.925 -27.715 -55.595 ;
        RECT -28.045 -60.005 -27.715 -59.675 ;
        RECT -28.045 -62.725 -27.715 -62.395 ;
        RECT -28.045 -68.165 -27.715 -67.835 ;
        RECT -28.045 -69.525 -27.715 -69.195 ;
        RECT -28.045 -70.885 -27.715 -70.555 ;
        RECT -28.045 -72.245 -27.715 -71.915 ;
        RECT -28.045 -74.965 -27.715 -74.635 ;
        RECT -28.045 -76.71 -27.715 -76.38 ;
        RECT -28.045 -77.685 -27.715 -77.355 ;
        RECT -28.045 -79.045 -27.715 -78.715 ;
        RECT -28.045 -81.765 -27.715 -81.435 ;
        RECT -28.045 -83.125 -27.715 -82.795 ;
        RECT -28.045 -84.485 -27.715 -84.155 ;
        RECT -28.045 -85.25 -27.715 -84.92 ;
        RECT -28.045 -87.205 -27.715 -86.875 ;
        RECT -28.045 -89.925 -27.715 -89.595 ;
        RECT -28.045 -91.285 -27.715 -90.955 ;
        RECT -28.045 -92.645 -27.715 -92.315 ;
        RECT -28.045 -94.005 -27.715 -93.675 ;
        RECT -28.045 -96.725 -27.715 -96.395 ;
        RECT -28.045 -98.085 -27.715 -97.755 ;
        RECT -28.045 -98.89 -27.715 -98.56 ;
        RECT -28.045 -100.805 -27.715 -100.475 ;
        RECT -28.045 -102.165 -27.715 -101.835 ;
        RECT -28.045 -104.885 -27.715 -104.555 ;
        RECT -28.045 -106.245 -27.715 -105.915 ;
        RECT -28.045 -107.43 -27.715 -107.1 ;
        RECT -28.045 -114.405 -27.715 -114.075 ;
        RECT -28.045 -115.765 -27.715 -115.435 ;
        RECT -28.045 -117.125 -27.715 -116.795 ;
        RECT -28.045 -118.485 -27.715 -118.155 ;
        RECT -28.045 -123.925 -27.715 -123.595 ;
        RECT -28.045 -126.645 -27.715 -126.315 ;
        RECT -28.045 -128.005 -27.715 -127.675 ;
        RECT -28.045 -129.365 -27.715 -129.035 ;
        RECT -28.045 -130.725 -27.715 -130.395 ;
        RECT -28.045 -133.445 -27.715 -133.115 ;
        RECT -28.045 -134.805 -27.715 -134.475 ;
        RECT -28.045 -136.165 -27.715 -135.835 ;
        RECT -28.045 -137.525 -27.715 -137.195 ;
        RECT -28.045 -141.605 -27.715 -141.275 ;
        RECT -28.045 -142.965 -27.715 -142.635 ;
        RECT -28.045 -144.325 -27.715 -143.995 ;
        RECT -28.045 -145.685 -27.715 -145.355 ;
        RECT -28.045 -147.045 -27.715 -146.715 ;
        RECT -28.045 -148.405 -27.715 -148.075 ;
        RECT -28.045 -149.765 -27.715 -149.435 ;
        RECT -28.045 -152.485 -27.715 -152.155 ;
        RECT -28.045 -153.845 -27.715 -153.515 ;
        RECT -28.045 -157.925 -27.715 -157.595 ;
        RECT -28.045 -159.285 -27.715 -158.955 ;
        RECT -28.045 -160.645 -27.715 -160.315 ;
        RECT -28.045 -162.005 -27.715 -161.675 ;
        RECT -28.045 -163.365 -27.715 -163.035 ;
        RECT -28.045 -164.725 -27.715 -164.395 ;
        RECT -28.045 -166.085 -27.715 -165.755 ;
        RECT -28.045 -167.445 -27.715 -167.115 ;
        RECT -28.045 -168.805 -27.715 -168.475 ;
        RECT -28.045 -171.525 -27.715 -171.195 ;
        RECT -28.045 -172.885 -27.715 -172.555 ;
        RECT -28.04 -172.885 -27.72 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.685 241.32 -26.355 242.45 ;
        RECT -26.685 239.195 -26.355 239.525 ;
        RECT -26.685 237.835 -26.355 238.165 ;
        RECT -26.685 236.475 -26.355 236.805 ;
        RECT -26.685 235.115 -26.355 235.445 ;
        RECT -26.685 233.755 -26.355 234.085 ;
        RECT -26.685 232.395 -26.355 232.725 ;
        RECT -26.685 231.035 -26.355 231.365 ;
        RECT -26.685 229.675 -26.355 230.005 ;
        RECT -26.685 228.315 -26.355 228.645 ;
        RECT -26.685 226.955 -26.355 227.285 ;
        RECT -26.685 225.595 -26.355 225.925 ;
        RECT -26.685 224.235 -26.355 224.565 ;
        RECT -26.685 222.875 -26.355 223.205 ;
        RECT -26.685 221.515 -26.355 221.845 ;
        RECT -26.685 220.155 -26.355 220.485 ;
        RECT -26.685 218.795 -26.355 219.125 ;
        RECT -26.685 217.435 -26.355 217.765 ;
        RECT -26.685 216.075 -26.355 216.405 ;
        RECT -26.685 214.715 -26.355 215.045 ;
        RECT -26.685 213.355 -26.355 213.685 ;
        RECT -26.685 211.995 -26.355 212.325 ;
        RECT -26.685 210.635 -26.355 210.965 ;
        RECT -26.685 209.275 -26.355 209.605 ;
        RECT -26.685 207.915 -26.355 208.245 ;
        RECT -26.685 206.555 -26.355 206.885 ;
        RECT -26.685 205.195 -26.355 205.525 ;
        RECT -26.685 203.835 -26.355 204.165 ;
        RECT -26.685 202.475 -26.355 202.805 ;
        RECT -26.685 201.115 -26.355 201.445 ;
        RECT -26.685 199.755 -26.355 200.085 ;
        RECT -26.685 198.395 -26.355 198.725 ;
        RECT -26.685 197.035 -26.355 197.365 ;
        RECT -26.685 195.675 -26.355 196.005 ;
        RECT -26.685 194.315 -26.355 194.645 ;
        RECT -26.685 192.955 -26.355 193.285 ;
        RECT -26.685 191.595 -26.355 191.925 ;
        RECT -26.685 190.235 -26.355 190.565 ;
        RECT -26.685 188.875 -26.355 189.205 ;
        RECT -26.685 187.515 -26.355 187.845 ;
        RECT -26.685 186.155 -26.355 186.485 ;
        RECT -26.685 184.795 -26.355 185.125 ;
        RECT -26.685 183.435 -26.355 183.765 ;
        RECT -26.685 182.075 -26.355 182.405 ;
        RECT -26.685 180.715 -26.355 181.045 ;
        RECT -26.685 179.355 -26.355 179.685 ;
        RECT -26.685 177.995 -26.355 178.325 ;
        RECT -26.685 176.635 -26.355 176.965 ;
        RECT -26.685 175.275 -26.355 175.605 ;
        RECT -26.685 173.915 -26.355 174.245 ;
        RECT -26.685 172.555 -26.355 172.885 ;
        RECT -26.685 171.195 -26.355 171.525 ;
        RECT -26.685 169.835 -26.355 170.165 ;
        RECT -26.685 168.475 -26.355 168.805 ;
        RECT -26.685 167.115 -26.355 167.445 ;
        RECT -26.685 165.755 -26.355 166.085 ;
        RECT -26.685 164.395 -26.355 164.725 ;
        RECT -26.685 163.035 -26.355 163.365 ;
        RECT -26.685 161.675 -26.355 162.005 ;
        RECT -26.685 160.315 -26.355 160.645 ;
        RECT -26.685 158.955 -26.355 159.285 ;
        RECT -26.685 157.595 -26.355 157.925 ;
        RECT -26.685 156.235 -26.355 156.565 ;
        RECT -26.685 154.875 -26.355 155.205 ;
        RECT -26.685 153.515 -26.355 153.845 ;
        RECT -26.685 152.155 -26.355 152.485 ;
        RECT -26.685 150.795 -26.355 151.125 ;
        RECT -26.685 149.435 -26.355 149.765 ;
        RECT -26.685 148.075 -26.355 148.405 ;
        RECT -26.685 146.715 -26.355 147.045 ;
        RECT -26.685 145.355 -26.355 145.685 ;
        RECT -26.685 143.995 -26.355 144.325 ;
        RECT -26.685 142.635 -26.355 142.965 ;
        RECT -26.685 141.275 -26.355 141.605 ;
        RECT -26.685 139.915 -26.355 140.245 ;
        RECT -26.685 138.555 -26.355 138.885 ;
        RECT -26.685 137.195 -26.355 137.525 ;
        RECT -26.685 135.835 -26.355 136.165 ;
        RECT -26.685 134.475 -26.355 134.805 ;
        RECT -26.685 133.115 -26.355 133.445 ;
        RECT -26.685 131.755 -26.355 132.085 ;
        RECT -26.685 130.395 -26.355 130.725 ;
        RECT -26.685 129.035 -26.355 129.365 ;
        RECT -26.685 127.675 -26.355 128.005 ;
        RECT -26.685 126.315 -26.355 126.645 ;
        RECT -26.685 124.955 -26.355 125.285 ;
        RECT -26.685 123.595 -26.355 123.925 ;
        RECT -26.685 122.235 -26.355 122.565 ;
        RECT -26.685 120.875 -26.355 121.205 ;
        RECT -26.685 119.515 -26.355 119.845 ;
        RECT -26.685 118.155 -26.355 118.485 ;
        RECT -26.685 116.795 -26.355 117.125 ;
        RECT -26.685 115.435 -26.355 115.765 ;
        RECT -26.685 114.075 -26.355 114.405 ;
        RECT -26.685 112.715 -26.355 113.045 ;
        RECT -26.685 111.355 -26.355 111.685 ;
        RECT -26.685 109.995 -26.355 110.325 ;
        RECT -26.685 108.635 -26.355 108.965 ;
        RECT -26.685 107.275 -26.355 107.605 ;
        RECT -26.685 105.915 -26.355 106.245 ;
        RECT -26.685 104.555 -26.355 104.885 ;
        RECT -26.685 103.195 -26.355 103.525 ;
        RECT -26.685 101.835 -26.355 102.165 ;
        RECT -26.685 100.475 -26.355 100.805 ;
        RECT -26.685 99.115 -26.355 99.445 ;
        RECT -26.685 97.755 -26.355 98.085 ;
        RECT -26.685 96.395 -26.355 96.725 ;
        RECT -26.685 95.035 -26.355 95.365 ;
        RECT -26.685 93.675 -26.355 94.005 ;
        RECT -26.685 92.315 -26.355 92.645 ;
        RECT -26.685 90.955 -26.355 91.285 ;
        RECT -26.685 89.595 -26.355 89.925 ;
        RECT -26.685 88.235 -26.355 88.565 ;
        RECT -26.685 86.875 -26.355 87.205 ;
        RECT -26.685 85.515 -26.355 85.845 ;
        RECT -26.685 84.155 -26.355 84.485 ;
        RECT -26.685 82.795 -26.355 83.125 ;
        RECT -26.685 81.435 -26.355 81.765 ;
        RECT -26.685 80.075 -26.355 80.405 ;
        RECT -26.685 78.715 -26.355 79.045 ;
        RECT -26.685 77.355 -26.355 77.685 ;
        RECT -26.685 75.995 -26.355 76.325 ;
        RECT -26.685 74.635 -26.355 74.965 ;
        RECT -26.685 73.275 -26.355 73.605 ;
        RECT -26.685 71.915 -26.355 72.245 ;
        RECT -26.685 70.555 -26.355 70.885 ;
        RECT -26.685 69.195 -26.355 69.525 ;
        RECT -26.685 67.835 -26.355 68.165 ;
        RECT -26.685 66.475 -26.355 66.805 ;
        RECT -26.685 65.115 -26.355 65.445 ;
        RECT -26.685 63.755 -26.355 64.085 ;
        RECT -26.685 62.395 -26.355 62.725 ;
        RECT -26.685 61.035 -26.355 61.365 ;
        RECT -26.685 59.675 -26.355 60.005 ;
        RECT -26.685 58.315 -26.355 58.645 ;
        RECT -26.685 56.955 -26.355 57.285 ;
        RECT -26.685 55.595 -26.355 55.925 ;
        RECT -26.685 54.235 -26.355 54.565 ;
        RECT -26.685 52.875 -26.355 53.205 ;
        RECT -26.685 51.515 -26.355 51.845 ;
        RECT -26.685 50.155 -26.355 50.485 ;
        RECT -26.685 48.795 -26.355 49.125 ;
        RECT -26.685 47.435 -26.355 47.765 ;
        RECT -26.685 46.075 -26.355 46.405 ;
        RECT -26.685 44.715 -26.355 45.045 ;
        RECT -26.685 43.355 -26.355 43.685 ;
        RECT -26.685 41.995 -26.355 42.325 ;
        RECT -26.685 40.635 -26.355 40.965 ;
        RECT -26.685 39.275 -26.355 39.605 ;
        RECT -26.685 37.915 -26.355 38.245 ;
        RECT -26.685 36.555 -26.355 36.885 ;
        RECT -26.685 35.195 -26.355 35.525 ;
        RECT -26.685 33.835 -26.355 34.165 ;
        RECT -26.685 32.475 -26.355 32.805 ;
        RECT -26.685 31.115 -26.355 31.445 ;
        RECT -26.685 29.755 -26.355 30.085 ;
        RECT -26.685 28.395 -26.355 28.725 ;
        RECT -26.685 27.035 -26.355 27.365 ;
        RECT -26.685 25.675 -26.355 26.005 ;
        RECT -26.685 24.315 -26.355 24.645 ;
        RECT -26.685 22.955 -26.355 23.285 ;
        RECT -26.685 21.595 -26.355 21.925 ;
        RECT -26.685 20.235 -26.355 20.565 ;
        RECT -26.685 18.875 -26.355 19.205 ;
        RECT -26.685 17.515 -26.355 17.845 ;
        RECT -26.685 16.155 -26.355 16.485 ;
        RECT -26.685 14.795 -26.355 15.125 ;
        RECT -26.685 13.435 -26.355 13.765 ;
        RECT -26.685 12.075 -26.355 12.405 ;
        RECT -26.685 10.715 -26.355 11.045 ;
        RECT -26.685 9.355 -26.355 9.685 ;
        RECT -26.685 7.995 -26.355 8.325 ;
        RECT -26.685 6.635 -26.355 6.965 ;
        RECT -26.685 5.275 -26.355 5.605 ;
        RECT -26.685 3.915 -26.355 4.245 ;
        RECT -26.685 2.555 -26.355 2.885 ;
        RECT -26.685 1.195 -26.355 1.525 ;
        RECT -26.685 -0.165 -26.355 0.165 ;
        RECT -26.685 -8.325 -26.355 -7.995 ;
        RECT -26.685 -9.685 -26.355 -9.355 ;
        RECT -26.685 -14.95 -26.355 -14.62 ;
        RECT -26.685 -17.845 -26.355 -17.515 ;
        RECT -26.685 -19.79 -26.355 -19.46 ;
        RECT -26.685 -20.565 -26.355 -20.235 ;
        RECT -26.685 -32.805 -26.355 -32.475 ;
        RECT -26.685 -35.525 -26.355 -35.195 ;
        RECT -26.685 -36.885 -26.355 -36.555 ;
        RECT -26.685 -37.93 -26.355 -37.6 ;
        RECT -26.685 -40.965 -26.355 -40.635 ;
        RECT -26.685 -42.77 -26.355 -42.44 ;
        RECT -26.685 -43.685 -26.355 -43.355 ;
        RECT -26.685 -50.485 -26.355 -50.155 ;
        RECT -26.685 -51.845 -26.355 -51.515 ;
        RECT -26.685 -54.565 -26.355 -54.235 ;
        RECT -26.685 -55.925 -26.355 -55.595 ;
        RECT -26.685 -60.005 -26.355 -59.675 ;
        RECT -26.685 -62.725 -26.355 -62.395 ;
        RECT -26.685 -68.165 -26.355 -67.835 ;
        RECT -26.685 -69.525 -26.355 -69.195 ;
        RECT -26.685 -70.885 -26.355 -70.555 ;
        RECT -26.685 -72.245 -26.355 -71.915 ;
        RECT -26.685 -74.965 -26.355 -74.635 ;
        RECT -26.685 -76.71 -26.355 -76.38 ;
        RECT -26.685 -77.685 -26.355 -77.355 ;
        RECT -26.685 -79.045 -26.355 -78.715 ;
        RECT -26.685 -81.765 -26.355 -81.435 ;
        RECT -26.685 -83.125 -26.355 -82.795 ;
        RECT -26.685 -84.485 -26.355 -84.155 ;
        RECT -26.685 -85.25 -26.355 -84.92 ;
        RECT -26.685 -87.205 -26.355 -86.875 ;
        RECT -26.685 -89.925 -26.355 -89.595 ;
        RECT -26.685 -91.285 -26.355 -90.955 ;
        RECT -26.685 -92.645 -26.355 -92.315 ;
        RECT -26.685 -94.005 -26.355 -93.675 ;
        RECT -26.685 -96.725 -26.355 -96.395 ;
        RECT -26.685 -98.085 -26.355 -97.755 ;
        RECT -26.685 -98.89 -26.355 -98.56 ;
        RECT -26.685 -100.805 -26.355 -100.475 ;
        RECT -26.685 -102.165 -26.355 -101.835 ;
        RECT -26.685 -104.885 -26.355 -104.555 ;
        RECT -26.685 -106.245 -26.355 -105.915 ;
        RECT -26.685 -107.43 -26.355 -107.1 ;
        RECT -26.685 -114.405 -26.355 -114.075 ;
        RECT -26.685 -115.765 -26.355 -115.435 ;
        RECT -26.685 -117.125 -26.355 -116.795 ;
        RECT -26.685 -118.485 -26.355 -118.155 ;
        RECT -26.685 -123.925 -26.355 -123.595 ;
        RECT -26.685 -126.645 -26.355 -126.315 ;
        RECT -26.685 -128.005 -26.355 -127.675 ;
        RECT -26.685 -129.365 -26.355 -129.035 ;
        RECT -26.685 -130.725 -26.355 -130.395 ;
        RECT -26.685 -136.165 -26.355 -135.835 ;
        RECT -26.685 -137.525 -26.355 -137.195 ;
        RECT -26.685 -141.605 -26.355 -141.275 ;
        RECT -26.685 -142.965 -26.355 -142.635 ;
        RECT -26.685 -144.325 -26.355 -143.995 ;
        RECT -26.685 -147.045 -26.355 -146.715 ;
        RECT -26.685 -148.405 -26.355 -148.075 ;
        RECT -26.685 -149.765 -26.355 -149.435 ;
        RECT -26.685 -152.485 -26.355 -152.155 ;
        RECT -26.685 -153.845 -26.355 -153.515 ;
        RECT -26.685 -157.925 -26.355 -157.595 ;
        RECT -26.685 -159.285 -26.355 -158.955 ;
        RECT -26.685 -160.645 -26.355 -160.315 ;
        RECT -26.685 -162.005 -26.355 -161.675 ;
        RECT -26.685 -163.365 -26.355 -163.035 ;
        RECT -26.685 -164.725 -26.355 -164.395 ;
        RECT -26.685 -166.085 -26.355 -165.755 ;
        RECT -26.685 -167.445 -26.355 -167.115 ;
        RECT -26.68 -167.445 -26.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -26.685 -174.245 -26.355 -173.915 ;
        RECT -26.685 -175.605 -26.355 -175.275 ;
        RECT -26.685 -176.685 -26.355 -176.355 ;
        RECT -26.685 -178.325 -26.355 -177.995 ;
        RECT -26.685 -179.685 -26.355 -179.355 ;
        RECT -26.685 -181.93 -26.355 -180.8 ;
        RECT -26.68 -182.045 -26.36 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -25.325 56.955 -24.995 57.285 ;
        RECT -25.325 55.595 -24.995 55.925 ;
        RECT -25.325 54.235 -24.995 54.565 ;
        RECT -25.325 52.875 -24.995 53.205 ;
        RECT -25.325 51.515 -24.995 51.845 ;
        RECT -25.325 50.155 -24.995 50.485 ;
        RECT -25.325 48.795 -24.995 49.125 ;
        RECT -25.325 47.435 -24.995 47.765 ;
        RECT -25.325 46.075 -24.995 46.405 ;
        RECT -25.325 44.715 -24.995 45.045 ;
        RECT -25.325 43.355 -24.995 43.685 ;
        RECT -25.325 41.995 -24.995 42.325 ;
        RECT -25.325 40.635 -24.995 40.965 ;
        RECT -25.325 39.275 -24.995 39.605 ;
        RECT -25.325 37.915 -24.995 38.245 ;
        RECT -25.325 36.555 -24.995 36.885 ;
        RECT -25.325 35.195 -24.995 35.525 ;
        RECT -25.325 33.835 -24.995 34.165 ;
        RECT -25.325 32.475 -24.995 32.805 ;
        RECT -25.325 31.115 -24.995 31.445 ;
        RECT -25.325 29.755 -24.995 30.085 ;
        RECT -25.325 28.395 -24.995 28.725 ;
        RECT -25.325 27.035 -24.995 27.365 ;
        RECT -25.325 25.675 -24.995 26.005 ;
        RECT -25.325 24.315 -24.995 24.645 ;
        RECT -25.325 22.955 -24.995 23.285 ;
        RECT -25.325 21.595 -24.995 21.925 ;
        RECT -25.325 20.235 -24.995 20.565 ;
        RECT -25.325 18.875 -24.995 19.205 ;
        RECT -25.325 17.515 -24.995 17.845 ;
        RECT -25.325 16.155 -24.995 16.485 ;
        RECT -25.325 14.795 -24.995 15.125 ;
        RECT -25.325 13.435 -24.995 13.765 ;
        RECT -25.325 12.075 -24.995 12.405 ;
        RECT -25.325 10.715 -24.995 11.045 ;
        RECT -25.325 9.355 -24.995 9.685 ;
        RECT -25.325 7.995 -24.995 8.325 ;
        RECT -25.325 6.635 -24.995 6.965 ;
        RECT -25.325 5.275 -24.995 5.605 ;
        RECT -25.325 3.915 -24.995 4.245 ;
        RECT -25.325 2.555 -24.995 2.885 ;
        RECT -25.325 1.195 -24.995 1.525 ;
        RECT -25.325 -0.165 -24.995 0.165 ;
        RECT -25.325 -2.885 -24.995 -2.555 ;
        RECT -25.325 -8.325 -24.995 -7.995 ;
        RECT -25.325 -9.685 -24.995 -9.355 ;
        RECT -25.325 -14.95 -24.995 -14.62 ;
        RECT -25.325 -17.845 -24.995 -17.515 ;
        RECT -25.325 -19.79 -24.995 -19.46 ;
        RECT -25.325 -20.565 -24.995 -20.235 ;
        RECT -25.325 -32.805 -24.995 -32.475 ;
        RECT -25.325 -35.525 -24.995 -35.195 ;
        RECT -25.325 -36.885 -24.995 -36.555 ;
        RECT -25.325 -37.93 -24.995 -37.6 ;
        RECT -25.325 -40.965 -24.995 -40.635 ;
        RECT -25.325 -42.77 -24.995 -42.44 ;
        RECT -25.325 -43.685 -24.995 -43.355 ;
        RECT -25.325 -50.485 -24.995 -50.155 ;
        RECT -25.325 -51.845 -24.995 -51.515 ;
        RECT -25.325 -54.565 -24.995 -54.235 ;
        RECT -25.325 -55.925 -24.995 -55.595 ;
        RECT -25.325 -60.005 -24.995 -59.675 ;
        RECT -25.325 -62.725 -24.995 -62.395 ;
        RECT -25.325 -68.165 -24.995 -67.835 ;
        RECT -25.325 -69.525 -24.995 -69.195 ;
        RECT -25.325 -70.885 -24.995 -70.555 ;
        RECT -25.325 -72.245 -24.995 -71.915 ;
        RECT -25.325 -74.965 -24.995 -74.635 ;
        RECT -25.325 -76.71 -24.995 -76.38 ;
        RECT -25.325 -77.685 -24.995 -77.355 ;
        RECT -25.325 -79.045 -24.995 -78.715 ;
        RECT -25.325 -81.765 -24.995 -81.435 ;
        RECT -25.325 -83.125 -24.995 -82.795 ;
        RECT -25.325 -84.485 -24.995 -84.155 ;
        RECT -25.325 -85.25 -24.995 -84.92 ;
        RECT -25.325 -87.205 -24.995 -86.875 ;
        RECT -25.325 -89.925 -24.995 -89.595 ;
        RECT -25.325 -91.285 -24.995 -90.955 ;
        RECT -25.325 -92.645 -24.995 -92.315 ;
        RECT -25.325 -94.005 -24.995 -93.675 ;
        RECT -25.325 -96.725 -24.995 -96.395 ;
        RECT -25.325 -98.085 -24.995 -97.755 ;
        RECT -25.325 -98.89 -24.995 -98.56 ;
        RECT -25.325 -100.805 -24.995 -100.475 ;
        RECT -25.325 -102.165 -24.995 -101.835 ;
        RECT -25.325 -104.885 -24.995 -104.555 ;
        RECT -25.325 -106.245 -24.995 -105.915 ;
        RECT -25.325 -107.43 -24.995 -107.1 ;
        RECT -25.325 -114.405 -24.995 -114.075 ;
        RECT -25.325 -115.765 -24.995 -115.435 ;
        RECT -25.325 -117.125 -24.995 -116.795 ;
        RECT -25.325 -118.485 -24.995 -118.155 ;
        RECT -25.325 -123.925 -24.995 -123.595 ;
        RECT -25.325 -125.285 -24.995 -124.955 ;
        RECT -25.325 -126.645 -24.995 -126.315 ;
        RECT -25.325 -128.005 -24.995 -127.675 ;
        RECT -25.325 -129.365 -24.995 -129.035 ;
        RECT -25.325 -130.725 -24.995 -130.395 ;
        RECT -25.325 -136.165 -24.995 -135.835 ;
        RECT -25.325 -137.525 -24.995 -137.195 ;
        RECT -25.325 -141.605 -24.995 -141.275 ;
        RECT -25.325 -142.965 -24.995 -142.635 ;
        RECT -25.325 -144.325 -24.995 -143.995 ;
        RECT -25.325 -147.045 -24.995 -146.715 ;
        RECT -25.325 -148.405 -24.995 -148.075 ;
        RECT -25.325 -149.765 -24.995 -149.435 ;
        RECT -25.325 -152.485 -24.995 -152.155 ;
        RECT -25.325 -153.845 -24.995 -153.515 ;
        RECT -25.325 -157.925 -24.995 -157.595 ;
        RECT -25.325 -159.285 -24.995 -158.955 ;
        RECT -25.325 -160.645 -24.995 -160.315 ;
        RECT -25.325 -162.005 -24.995 -161.675 ;
        RECT -25.325 -163.365 -24.995 -163.035 ;
        RECT -25.325 -164.725 -24.995 -164.395 ;
        RECT -25.325 -166.085 -24.995 -165.755 ;
        RECT -25.325 -167.445 -24.995 -167.115 ;
        RECT -25.325 -168.805 -24.995 -168.475 ;
        RECT -25.325 -171.525 -24.995 -171.195 ;
        RECT -25.325 -172.885 -24.995 -172.555 ;
        RECT -25.325 -174.245 -24.995 -173.915 ;
        RECT -25.325 -175.605 -24.995 -175.275 ;
        RECT -25.325 -176.685 -24.995 -176.355 ;
        RECT -25.325 -178.325 -24.995 -177.995 ;
        RECT -25.325 -179.685 -24.995 -179.355 ;
        RECT -25.325 -181.93 -24.995 -180.8 ;
        RECT -25.32 -182.045 -25 242.565 ;
        RECT -25.325 241.32 -24.995 242.45 ;
        RECT -25.325 239.195 -24.995 239.525 ;
        RECT -25.325 237.835 -24.995 238.165 ;
        RECT -25.325 236.475 -24.995 236.805 ;
        RECT -25.325 235.115 -24.995 235.445 ;
        RECT -25.325 233.755 -24.995 234.085 ;
        RECT -25.325 232.395 -24.995 232.725 ;
        RECT -25.325 231.035 -24.995 231.365 ;
        RECT -25.325 229.675 -24.995 230.005 ;
        RECT -25.325 228.315 -24.995 228.645 ;
        RECT -25.325 226.955 -24.995 227.285 ;
        RECT -25.325 225.595 -24.995 225.925 ;
        RECT -25.325 224.235 -24.995 224.565 ;
        RECT -25.325 222.875 -24.995 223.205 ;
        RECT -25.325 221.515 -24.995 221.845 ;
        RECT -25.325 220.155 -24.995 220.485 ;
        RECT -25.325 218.795 -24.995 219.125 ;
        RECT -25.325 217.435 -24.995 217.765 ;
        RECT -25.325 216.075 -24.995 216.405 ;
        RECT -25.325 214.715 -24.995 215.045 ;
        RECT -25.325 213.355 -24.995 213.685 ;
        RECT -25.325 211.995 -24.995 212.325 ;
        RECT -25.325 210.635 -24.995 210.965 ;
        RECT -25.325 209.275 -24.995 209.605 ;
        RECT -25.325 207.915 -24.995 208.245 ;
        RECT -25.325 206.555 -24.995 206.885 ;
        RECT -25.325 205.195 -24.995 205.525 ;
        RECT -25.325 203.835 -24.995 204.165 ;
        RECT -25.325 202.475 -24.995 202.805 ;
        RECT -25.325 201.115 -24.995 201.445 ;
        RECT -25.325 199.755 -24.995 200.085 ;
        RECT -25.325 198.395 -24.995 198.725 ;
        RECT -25.325 197.035 -24.995 197.365 ;
        RECT -25.325 195.675 -24.995 196.005 ;
        RECT -25.325 194.315 -24.995 194.645 ;
        RECT -25.325 192.955 -24.995 193.285 ;
        RECT -25.325 191.595 -24.995 191.925 ;
        RECT -25.325 190.235 -24.995 190.565 ;
        RECT -25.325 188.875 -24.995 189.205 ;
        RECT -25.325 187.515 -24.995 187.845 ;
        RECT -25.325 186.155 -24.995 186.485 ;
        RECT -25.325 184.795 -24.995 185.125 ;
        RECT -25.325 183.435 -24.995 183.765 ;
        RECT -25.325 182.075 -24.995 182.405 ;
        RECT -25.325 180.715 -24.995 181.045 ;
        RECT -25.325 179.355 -24.995 179.685 ;
        RECT -25.325 177.995 -24.995 178.325 ;
        RECT -25.325 176.635 -24.995 176.965 ;
        RECT -25.325 175.275 -24.995 175.605 ;
        RECT -25.325 173.915 -24.995 174.245 ;
        RECT -25.325 172.555 -24.995 172.885 ;
        RECT -25.325 171.195 -24.995 171.525 ;
        RECT -25.325 169.835 -24.995 170.165 ;
        RECT -25.325 168.475 -24.995 168.805 ;
        RECT -25.325 167.115 -24.995 167.445 ;
        RECT -25.325 165.755 -24.995 166.085 ;
        RECT -25.325 164.395 -24.995 164.725 ;
        RECT -25.325 163.035 -24.995 163.365 ;
        RECT -25.325 161.675 -24.995 162.005 ;
        RECT -25.325 160.315 -24.995 160.645 ;
        RECT -25.325 158.955 -24.995 159.285 ;
        RECT -25.325 157.595 -24.995 157.925 ;
        RECT -25.325 156.235 -24.995 156.565 ;
        RECT -25.325 154.875 -24.995 155.205 ;
        RECT -25.325 153.515 -24.995 153.845 ;
        RECT -25.325 152.155 -24.995 152.485 ;
        RECT -25.325 150.795 -24.995 151.125 ;
        RECT -25.325 149.435 -24.995 149.765 ;
        RECT -25.325 148.075 -24.995 148.405 ;
        RECT -25.325 146.715 -24.995 147.045 ;
        RECT -25.325 145.355 -24.995 145.685 ;
        RECT -25.325 143.995 -24.995 144.325 ;
        RECT -25.325 142.635 -24.995 142.965 ;
        RECT -25.325 141.275 -24.995 141.605 ;
        RECT -25.325 139.915 -24.995 140.245 ;
        RECT -25.325 138.555 -24.995 138.885 ;
        RECT -25.325 137.195 -24.995 137.525 ;
        RECT -25.325 135.835 -24.995 136.165 ;
        RECT -25.325 134.475 -24.995 134.805 ;
        RECT -25.325 133.115 -24.995 133.445 ;
        RECT -25.325 131.755 -24.995 132.085 ;
        RECT -25.325 130.395 -24.995 130.725 ;
        RECT -25.325 129.035 -24.995 129.365 ;
        RECT -25.325 127.675 -24.995 128.005 ;
        RECT -25.325 126.315 -24.995 126.645 ;
        RECT -25.325 124.955 -24.995 125.285 ;
        RECT -25.325 123.595 -24.995 123.925 ;
        RECT -25.325 122.235 -24.995 122.565 ;
        RECT -25.325 120.875 -24.995 121.205 ;
        RECT -25.325 119.515 -24.995 119.845 ;
        RECT -25.325 118.155 -24.995 118.485 ;
        RECT -25.325 116.795 -24.995 117.125 ;
        RECT -25.325 115.435 -24.995 115.765 ;
        RECT -25.325 114.075 -24.995 114.405 ;
        RECT -25.325 112.715 -24.995 113.045 ;
        RECT -25.325 111.355 -24.995 111.685 ;
        RECT -25.325 109.995 -24.995 110.325 ;
        RECT -25.325 108.635 -24.995 108.965 ;
        RECT -25.325 107.275 -24.995 107.605 ;
        RECT -25.325 105.915 -24.995 106.245 ;
        RECT -25.325 104.555 -24.995 104.885 ;
        RECT -25.325 103.195 -24.995 103.525 ;
        RECT -25.325 101.835 -24.995 102.165 ;
        RECT -25.325 100.475 -24.995 100.805 ;
        RECT -25.325 99.115 -24.995 99.445 ;
        RECT -25.325 97.755 -24.995 98.085 ;
        RECT -25.325 96.395 -24.995 96.725 ;
        RECT -25.325 95.035 -24.995 95.365 ;
        RECT -25.325 93.675 -24.995 94.005 ;
        RECT -25.325 92.315 -24.995 92.645 ;
        RECT -25.325 90.955 -24.995 91.285 ;
        RECT -25.325 89.595 -24.995 89.925 ;
        RECT -25.325 88.235 -24.995 88.565 ;
        RECT -25.325 86.875 -24.995 87.205 ;
        RECT -25.325 85.515 -24.995 85.845 ;
        RECT -25.325 84.155 -24.995 84.485 ;
        RECT -25.325 82.795 -24.995 83.125 ;
        RECT -25.325 81.435 -24.995 81.765 ;
        RECT -25.325 80.075 -24.995 80.405 ;
        RECT -25.325 78.715 -24.995 79.045 ;
        RECT -25.325 77.355 -24.995 77.685 ;
        RECT -25.325 75.995 -24.995 76.325 ;
        RECT -25.325 74.635 -24.995 74.965 ;
        RECT -25.325 73.275 -24.995 73.605 ;
        RECT -25.325 71.915 -24.995 72.245 ;
        RECT -25.325 70.555 -24.995 70.885 ;
        RECT -25.325 69.195 -24.995 69.525 ;
        RECT -25.325 67.835 -24.995 68.165 ;
        RECT -25.325 66.475 -24.995 66.805 ;
        RECT -25.325 65.115 -24.995 65.445 ;
        RECT -25.325 63.755 -24.995 64.085 ;
        RECT -25.325 62.395 -24.995 62.725 ;
        RECT -25.325 61.035 -24.995 61.365 ;
        RECT -25.325 59.675 -24.995 60.005 ;
        RECT -25.325 58.315 -24.995 58.645 ;
    END
    PORT
      LAYER met3 ;
        RECT -34.845 241.32 -34.515 242.45 ;
        RECT -34.845 239.195 -34.515 239.525 ;
        RECT -34.845 237.835 -34.515 238.165 ;
        RECT -34.845 236.475 -34.515 236.805 ;
        RECT -34.845 235.115 -34.515 235.445 ;
        RECT -34.845 233.755 -34.515 234.085 ;
        RECT -34.845 232.395 -34.515 232.725 ;
        RECT -34.845 231.035 -34.515 231.365 ;
        RECT -34.845 229.675 -34.515 230.005 ;
        RECT -34.845 228.315 -34.515 228.645 ;
        RECT -34.845 226.955 -34.515 227.285 ;
        RECT -34.845 225.595 -34.515 225.925 ;
        RECT -34.845 224.235 -34.515 224.565 ;
        RECT -34.845 222.875 -34.515 223.205 ;
        RECT -34.845 221.515 -34.515 221.845 ;
        RECT -34.845 220.155 -34.515 220.485 ;
        RECT -34.845 218.795 -34.515 219.125 ;
        RECT -34.845 217.435 -34.515 217.765 ;
        RECT -34.845 216.075 -34.515 216.405 ;
        RECT -34.845 214.715 -34.515 215.045 ;
        RECT -34.845 213.355 -34.515 213.685 ;
        RECT -34.845 211.995 -34.515 212.325 ;
        RECT -34.845 210.635 -34.515 210.965 ;
        RECT -34.845 209.275 -34.515 209.605 ;
        RECT -34.845 207.915 -34.515 208.245 ;
        RECT -34.845 206.555 -34.515 206.885 ;
        RECT -34.845 205.195 -34.515 205.525 ;
        RECT -34.845 203.835 -34.515 204.165 ;
        RECT -34.845 202.475 -34.515 202.805 ;
        RECT -34.845 201.115 -34.515 201.445 ;
        RECT -34.845 199.755 -34.515 200.085 ;
        RECT -34.845 198.395 -34.515 198.725 ;
        RECT -34.845 197.035 -34.515 197.365 ;
        RECT -34.845 195.675 -34.515 196.005 ;
        RECT -34.845 194.315 -34.515 194.645 ;
        RECT -34.845 192.955 -34.515 193.285 ;
        RECT -34.845 191.595 -34.515 191.925 ;
        RECT -34.845 190.235 -34.515 190.565 ;
        RECT -34.845 188.875 -34.515 189.205 ;
        RECT -34.845 187.515 -34.515 187.845 ;
        RECT -34.845 186.155 -34.515 186.485 ;
        RECT -34.845 184.795 -34.515 185.125 ;
        RECT -34.845 183.435 -34.515 183.765 ;
        RECT -34.845 182.075 -34.515 182.405 ;
        RECT -34.845 180.715 -34.515 181.045 ;
        RECT -34.845 179.355 -34.515 179.685 ;
        RECT -34.845 177.995 -34.515 178.325 ;
        RECT -34.845 176.635 -34.515 176.965 ;
        RECT -34.845 175.275 -34.515 175.605 ;
        RECT -34.845 173.915 -34.515 174.245 ;
        RECT -34.845 172.555 -34.515 172.885 ;
        RECT -34.845 171.195 -34.515 171.525 ;
        RECT -34.845 169.835 -34.515 170.165 ;
        RECT -34.845 168.475 -34.515 168.805 ;
        RECT -34.845 167.115 -34.515 167.445 ;
        RECT -34.845 165.755 -34.515 166.085 ;
        RECT -34.845 164.395 -34.515 164.725 ;
        RECT -34.845 163.035 -34.515 163.365 ;
        RECT -34.845 161.675 -34.515 162.005 ;
        RECT -34.845 160.315 -34.515 160.645 ;
        RECT -34.845 158.955 -34.515 159.285 ;
        RECT -34.845 157.595 -34.515 157.925 ;
        RECT -34.845 156.235 -34.515 156.565 ;
        RECT -34.845 154.875 -34.515 155.205 ;
        RECT -34.845 153.515 -34.515 153.845 ;
        RECT -34.845 152.155 -34.515 152.485 ;
        RECT -34.845 150.795 -34.515 151.125 ;
        RECT -34.845 149.435 -34.515 149.765 ;
        RECT -34.845 148.075 -34.515 148.405 ;
        RECT -34.845 146.715 -34.515 147.045 ;
        RECT -34.845 145.355 -34.515 145.685 ;
        RECT -34.845 143.995 -34.515 144.325 ;
        RECT -34.845 142.635 -34.515 142.965 ;
        RECT -34.845 141.275 -34.515 141.605 ;
        RECT -34.845 139.915 -34.515 140.245 ;
        RECT -34.845 138.555 -34.515 138.885 ;
        RECT -34.845 137.195 -34.515 137.525 ;
        RECT -34.845 135.835 -34.515 136.165 ;
        RECT -34.845 134.475 -34.515 134.805 ;
        RECT -34.845 133.115 -34.515 133.445 ;
        RECT -34.845 131.755 -34.515 132.085 ;
        RECT -34.845 130.395 -34.515 130.725 ;
        RECT -34.845 129.035 -34.515 129.365 ;
        RECT -34.845 127.675 -34.515 128.005 ;
        RECT -34.845 126.315 -34.515 126.645 ;
        RECT -34.845 124.955 -34.515 125.285 ;
        RECT -34.845 123.595 -34.515 123.925 ;
        RECT -34.845 122.235 -34.515 122.565 ;
        RECT -34.845 120.875 -34.515 121.205 ;
        RECT -34.845 119.515 -34.515 119.845 ;
        RECT -34.845 118.155 -34.515 118.485 ;
        RECT -34.845 116.795 -34.515 117.125 ;
        RECT -34.845 115.435 -34.515 115.765 ;
        RECT -34.845 114.075 -34.515 114.405 ;
        RECT -34.845 112.715 -34.515 113.045 ;
        RECT -34.845 111.355 -34.515 111.685 ;
        RECT -34.845 109.995 -34.515 110.325 ;
        RECT -34.845 108.635 -34.515 108.965 ;
        RECT -34.845 107.275 -34.515 107.605 ;
        RECT -34.845 105.915 -34.515 106.245 ;
        RECT -34.845 104.555 -34.515 104.885 ;
        RECT -34.845 103.195 -34.515 103.525 ;
        RECT -34.845 101.835 -34.515 102.165 ;
        RECT -34.845 100.475 -34.515 100.805 ;
        RECT -34.845 99.115 -34.515 99.445 ;
        RECT -34.845 97.755 -34.515 98.085 ;
        RECT -34.845 96.395 -34.515 96.725 ;
        RECT -34.845 95.035 -34.515 95.365 ;
        RECT -34.845 93.675 -34.515 94.005 ;
        RECT -34.845 92.315 -34.515 92.645 ;
        RECT -34.845 90.955 -34.515 91.285 ;
        RECT -34.845 89.595 -34.515 89.925 ;
        RECT -34.845 88.235 -34.515 88.565 ;
        RECT -34.845 86.875 -34.515 87.205 ;
        RECT -34.845 85.515 -34.515 85.845 ;
        RECT -34.845 84.155 -34.515 84.485 ;
        RECT -34.845 82.795 -34.515 83.125 ;
        RECT -34.845 81.435 -34.515 81.765 ;
        RECT -34.845 80.075 -34.515 80.405 ;
        RECT -34.845 78.715 -34.515 79.045 ;
        RECT -34.845 77.355 -34.515 77.685 ;
        RECT -34.845 75.995 -34.515 76.325 ;
        RECT -34.845 74.635 -34.515 74.965 ;
        RECT -34.845 73.275 -34.515 73.605 ;
        RECT -34.845 71.915 -34.515 72.245 ;
        RECT -34.845 70.555 -34.515 70.885 ;
        RECT -34.845 69.195 -34.515 69.525 ;
        RECT -34.845 67.835 -34.515 68.165 ;
        RECT -34.845 66.475 -34.515 66.805 ;
        RECT -34.845 65.115 -34.515 65.445 ;
        RECT -34.845 63.755 -34.515 64.085 ;
        RECT -34.845 62.395 -34.515 62.725 ;
        RECT -34.845 61.035 -34.515 61.365 ;
        RECT -34.845 59.675 -34.515 60.005 ;
        RECT -34.845 58.315 -34.515 58.645 ;
        RECT -34.845 56.955 -34.515 57.285 ;
        RECT -34.845 55.595 -34.515 55.925 ;
        RECT -34.845 54.235 -34.515 54.565 ;
        RECT -34.845 52.875 -34.515 53.205 ;
        RECT -34.845 51.515 -34.515 51.845 ;
        RECT -34.845 50.155 -34.515 50.485 ;
        RECT -34.845 48.795 -34.515 49.125 ;
        RECT -34.845 47.435 -34.515 47.765 ;
        RECT -34.845 46.075 -34.515 46.405 ;
        RECT -34.845 44.715 -34.515 45.045 ;
        RECT -34.845 43.355 -34.515 43.685 ;
        RECT -34.845 41.995 -34.515 42.325 ;
        RECT -34.845 40.635 -34.515 40.965 ;
        RECT -34.845 39.275 -34.515 39.605 ;
        RECT -34.845 37.915 -34.515 38.245 ;
        RECT -34.845 36.555 -34.515 36.885 ;
        RECT -34.845 35.195 -34.515 35.525 ;
        RECT -34.845 33.835 -34.515 34.165 ;
        RECT -34.845 32.475 -34.515 32.805 ;
        RECT -34.845 31.115 -34.515 31.445 ;
        RECT -34.845 29.755 -34.515 30.085 ;
        RECT -34.845 28.395 -34.515 28.725 ;
        RECT -34.845 27.035 -34.515 27.365 ;
        RECT -34.845 25.675 -34.515 26.005 ;
        RECT -34.845 24.315 -34.515 24.645 ;
        RECT -34.845 22.955 -34.515 23.285 ;
        RECT -34.845 21.595 -34.515 21.925 ;
        RECT -34.845 20.235 -34.515 20.565 ;
        RECT -34.845 18.875 -34.515 19.205 ;
        RECT -34.845 17.515 -34.515 17.845 ;
        RECT -34.845 16.155 -34.515 16.485 ;
        RECT -34.845 14.795 -34.515 15.125 ;
        RECT -34.845 13.435 -34.515 13.765 ;
        RECT -34.845 12.075 -34.515 12.405 ;
        RECT -34.845 10.715 -34.515 11.045 ;
        RECT -34.845 9.355 -34.515 9.685 ;
        RECT -34.845 7.995 -34.515 8.325 ;
        RECT -34.845 6.635 -34.515 6.965 ;
        RECT -34.845 5.275 -34.515 5.605 ;
        RECT -34.845 3.915 -34.515 4.245 ;
        RECT -34.845 2.555 -34.515 2.885 ;
        RECT -34.845 1.195 -34.515 1.525 ;
        RECT -34.845 -0.165 -34.515 0.165 ;
        RECT -34.845 -8.325 -34.515 -7.995 ;
        RECT -34.845 -11.045 -34.515 -10.715 ;
        RECT -34.845 -15.125 -34.515 -14.795 ;
        RECT -34.845 -16.485 -34.515 -16.155 ;
        RECT -34.845 -17.845 -34.515 -17.515 ;
        RECT -34.845 -19.205 -34.515 -18.875 ;
        RECT -34.845 -20.565 -34.515 -20.235 ;
        RECT -34.845 -21.925 -34.515 -21.595 ;
        RECT -34.845 -23.285 -34.515 -22.955 ;
        RECT -34.845 -24.645 -34.515 -24.315 ;
        RECT -34.845 -32.805 -34.515 -32.475 ;
        RECT -34.845 -35.525 -34.515 -35.195 ;
        RECT -34.845 -36.885 -34.515 -36.555 ;
        RECT -34.845 -37.93 -34.515 -37.6 ;
        RECT -34.845 -40.965 -34.515 -40.635 ;
        RECT -34.845 -42.77 -34.515 -42.44 ;
        RECT -34.845 -43.685 -34.515 -43.355 ;
        RECT -34.845 -50.485 -34.515 -50.155 ;
        RECT -34.845 -51.845 -34.515 -51.515 ;
        RECT -34.845 -54.565 -34.515 -54.235 ;
        RECT -34.845 -55.925 -34.515 -55.595 ;
        RECT -34.845 -60.005 -34.515 -59.675 ;
        RECT -34.845 -62.725 -34.515 -62.395 ;
        RECT -34.845 -69.525 -34.515 -69.195 ;
        RECT -34.845 -70.885 -34.515 -70.555 ;
        RECT -34.845 -72.245 -34.515 -71.915 ;
        RECT -34.845 -73.605 -34.515 -73.275 ;
        RECT -34.845 -74.965 -34.515 -74.635 ;
        RECT -34.845 -76.325 -34.515 -75.995 ;
        RECT -34.845 -77.685 -34.515 -77.355 ;
        RECT -34.845 -79.045 -34.515 -78.715 ;
        RECT -34.845 -80.405 -34.515 -80.075 ;
        RECT -34.845 -81.765 -34.515 -81.435 ;
        RECT -34.845 -83.125 -34.515 -82.795 ;
        RECT -34.845 -84.485 -34.515 -84.155 ;
        RECT -34.845 -85.845 -34.515 -85.515 ;
        RECT -34.845 -87.205 -34.515 -86.875 ;
        RECT -34.845 -88.565 -34.515 -88.235 ;
        RECT -34.845 -89.925 -34.515 -89.595 ;
        RECT -34.845 -91.285 -34.515 -90.955 ;
        RECT -34.845 -92.645 -34.515 -92.315 ;
        RECT -34.845 -94.005 -34.515 -93.675 ;
        RECT -34.845 -95.365 -34.515 -95.035 ;
        RECT -34.845 -96.725 -34.515 -96.395 ;
        RECT -34.845 -98.085 -34.515 -97.755 ;
        RECT -34.845 -99.445 -34.515 -99.115 ;
        RECT -34.845 -100.805 -34.515 -100.475 ;
        RECT -34.845 -102.165 -34.515 -101.835 ;
        RECT -34.845 -103.525 -34.515 -103.195 ;
        RECT -34.845 -104.885 -34.515 -104.555 ;
        RECT -34.845 -106.245 -34.515 -105.915 ;
        RECT -34.845 -107.605 -34.515 -107.275 ;
        RECT -34.845 -108.965 -34.515 -108.635 ;
        RECT -34.845 -110.325 -34.515 -109.995 ;
        RECT -34.845 -111.685 -34.515 -111.355 ;
        RECT -34.845 -113.045 -34.515 -112.715 ;
        RECT -34.845 -114.405 -34.515 -114.075 ;
        RECT -34.845 -115.765 -34.515 -115.435 ;
        RECT -34.845 -117.125 -34.515 -116.795 ;
        RECT -34.845 -118.485 -34.515 -118.155 ;
        RECT -34.845 -121.205 -34.515 -120.875 ;
        RECT -34.845 -123.925 -34.515 -123.595 ;
        RECT -34.845 -126.645 -34.515 -126.315 ;
        RECT -34.845 -128.005 -34.515 -127.675 ;
        RECT -34.845 -129.365 -34.515 -129.035 ;
        RECT -34.845 -130.725 -34.515 -130.395 ;
        RECT -34.845 -133.445 -34.515 -133.115 ;
        RECT -34.845 -134.805 -34.515 -134.475 ;
        RECT -34.845 -136.165 -34.515 -135.835 ;
        RECT -34.845 -137.525 -34.515 -137.195 ;
        RECT -34.845 -138.885 -34.515 -138.555 ;
        RECT -34.845 -141.605 -34.515 -141.275 ;
        RECT -34.845 -142.965 -34.515 -142.635 ;
        RECT -34.845 -144.325 -34.515 -143.995 ;
        RECT -34.845 -145.685 -34.515 -145.355 ;
        RECT -34.845 -147.045 -34.515 -146.715 ;
        RECT -34.845 -148.405 -34.515 -148.075 ;
        RECT -34.845 -149.765 -34.515 -149.435 ;
        RECT -34.845 -152.485 -34.515 -152.155 ;
        RECT -34.845 -153.845 -34.515 -153.515 ;
        RECT -34.845 -157.925 -34.515 -157.595 ;
        RECT -34.845 -159.285 -34.515 -158.955 ;
        RECT -34.845 -160.645 -34.515 -160.315 ;
        RECT -34.845 -162.005 -34.515 -161.675 ;
        RECT -34.845 -163.365 -34.515 -163.035 ;
        RECT -34.845 -164.725 -34.515 -164.395 ;
        RECT -34.845 -166.085 -34.515 -165.755 ;
        RECT -34.845 -167.445 -34.515 -167.115 ;
        RECT -34.845 -168.805 -34.515 -168.475 ;
        RECT -34.845 -171.525 -34.515 -171.195 ;
        RECT -34.845 -175.605 -34.515 -175.275 ;
        RECT -34.845 -178.325 -34.515 -177.995 ;
        RECT -34.845 -179.685 -34.515 -179.355 ;
        RECT -34.845 -181.93 -34.515 -180.8 ;
        RECT -34.84 -182.045 -34.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -33.485 241.32 -33.155 242.45 ;
        RECT -33.485 239.195 -33.155 239.525 ;
        RECT -33.485 237.835 -33.155 238.165 ;
        RECT -33.485 236.475 -33.155 236.805 ;
        RECT -33.485 235.115 -33.155 235.445 ;
        RECT -33.485 233.755 -33.155 234.085 ;
        RECT -33.485 232.395 -33.155 232.725 ;
        RECT -33.485 231.035 -33.155 231.365 ;
        RECT -33.485 229.675 -33.155 230.005 ;
        RECT -33.485 228.315 -33.155 228.645 ;
        RECT -33.485 226.955 -33.155 227.285 ;
        RECT -33.485 225.595 -33.155 225.925 ;
        RECT -33.485 224.235 -33.155 224.565 ;
        RECT -33.485 222.875 -33.155 223.205 ;
        RECT -33.485 221.515 -33.155 221.845 ;
        RECT -33.485 220.155 -33.155 220.485 ;
        RECT -33.485 218.795 -33.155 219.125 ;
        RECT -33.485 217.435 -33.155 217.765 ;
        RECT -33.485 216.075 -33.155 216.405 ;
        RECT -33.485 214.715 -33.155 215.045 ;
        RECT -33.485 213.355 -33.155 213.685 ;
        RECT -33.485 211.995 -33.155 212.325 ;
        RECT -33.485 210.635 -33.155 210.965 ;
        RECT -33.485 209.275 -33.155 209.605 ;
        RECT -33.485 207.915 -33.155 208.245 ;
        RECT -33.485 206.555 -33.155 206.885 ;
        RECT -33.485 205.195 -33.155 205.525 ;
        RECT -33.485 203.835 -33.155 204.165 ;
        RECT -33.485 202.475 -33.155 202.805 ;
        RECT -33.485 201.115 -33.155 201.445 ;
        RECT -33.485 199.755 -33.155 200.085 ;
        RECT -33.485 198.395 -33.155 198.725 ;
        RECT -33.485 197.035 -33.155 197.365 ;
        RECT -33.485 195.675 -33.155 196.005 ;
        RECT -33.485 194.315 -33.155 194.645 ;
        RECT -33.485 192.955 -33.155 193.285 ;
        RECT -33.485 191.595 -33.155 191.925 ;
        RECT -33.485 190.235 -33.155 190.565 ;
        RECT -33.485 188.875 -33.155 189.205 ;
        RECT -33.485 187.515 -33.155 187.845 ;
        RECT -33.485 186.155 -33.155 186.485 ;
        RECT -33.485 184.795 -33.155 185.125 ;
        RECT -33.485 183.435 -33.155 183.765 ;
        RECT -33.485 182.075 -33.155 182.405 ;
        RECT -33.485 180.715 -33.155 181.045 ;
        RECT -33.485 179.355 -33.155 179.685 ;
        RECT -33.485 177.995 -33.155 178.325 ;
        RECT -33.485 176.635 -33.155 176.965 ;
        RECT -33.485 175.275 -33.155 175.605 ;
        RECT -33.485 173.915 -33.155 174.245 ;
        RECT -33.485 172.555 -33.155 172.885 ;
        RECT -33.485 171.195 -33.155 171.525 ;
        RECT -33.485 169.835 -33.155 170.165 ;
        RECT -33.485 168.475 -33.155 168.805 ;
        RECT -33.485 167.115 -33.155 167.445 ;
        RECT -33.485 165.755 -33.155 166.085 ;
        RECT -33.485 164.395 -33.155 164.725 ;
        RECT -33.485 163.035 -33.155 163.365 ;
        RECT -33.485 161.675 -33.155 162.005 ;
        RECT -33.485 160.315 -33.155 160.645 ;
        RECT -33.485 158.955 -33.155 159.285 ;
        RECT -33.485 157.595 -33.155 157.925 ;
        RECT -33.485 156.235 -33.155 156.565 ;
        RECT -33.485 154.875 -33.155 155.205 ;
        RECT -33.485 153.515 -33.155 153.845 ;
        RECT -33.485 152.155 -33.155 152.485 ;
        RECT -33.485 150.795 -33.155 151.125 ;
        RECT -33.485 149.435 -33.155 149.765 ;
        RECT -33.485 148.075 -33.155 148.405 ;
        RECT -33.485 146.715 -33.155 147.045 ;
        RECT -33.485 145.355 -33.155 145.685 ;
        RECT -33.485 143.995 -33.155 144.325 ;
        RECT -33.485 142.635 -33.155 142.965 ;
        RECT -33.485 141.275 -33.155 141.605 ;
        RECT -33.485 139.915 -33.155 140.245 ;
        RECT -33.485 138.555 -33.155 138.885 ;
        RECT -33.485 137.195 -33.155 137.525 ;
        RECT -33.485 135.835 -33.155 136.165 ;
        RECT -33.485 134.475 -33.155 134.805 ;
        RECT -33.485 133.115 -33.155 133.445 ;
        RECT -33.485 131.755 -33.155 132.085 ;
        RECT -33.485 130.395 -33.155 130.725 ;
        RECT -33.485 129.035 -33.155 129.365 ;
        RECT -33.485 127.675 -33.155 128.005 ;
        RECT -33.485 126.315 -33.155 126.645 ;
        RECT -33.485 124.955 -33.155 125.285 ;
        RECT -33.485 123.595 -33.155 123.925 ;
        RECT -33.485 122.235 -33.155 122.565 ;
        RECT -33.485 120.875 -33.155 121.205 ;
        RECT -33.485 119.515 -33.155 119.845 ;
        RECT -33.485 118.155 -33.155 118.485 ;
        RECT -33.485 116.795 -33.155 117.125 ;
        RECT -33.485 115.435 -33.155 115.765 ;
        RECT -33.485 114.075 -33.155 114.405 ;
        RECT -33.485 112.715 -33.155 113.045 ;
        RECT -33.485 111.355 -33.155 111.685 ;
        RECT -33.485 109.995 -33.155 110.325 ;
        RECT -33.485 108.635 -33.155 108.965 ;
        RECT -33.485 107.275 -33.155 107.605 ;
        RECT -33.485 105.915 -33.155 106.245 ;
        RECT -33.485 104.555 -33.155 104.885 ;
        RECT -33.485 103.195 -33.155 103.525 ;
        RECT -33.485 101.835 -33.155 102.165 ;
        RECT -33.485 100.475 -33.155 100.805 ;
        RECT -33.485 99.115 -33.155 99.445 ;
        RECT -33.485 97.755 -33.155 98.085 ;
        RECT -33.485 96.395 -33.155 96.725 ;
        RECT -33.485 95.035 -33.155 95.365 ;
        RECT -33.485 93.675 -33.155 94.005 ;
        RECT -33.485 92.315 -33.155 92.645 ;
        RECT -33.485 90.955 -33.155 91.285 ;
        RECT -33.485 89.595 -33.155 89.925 ;
        RECT -33.485 88.235 -33.155 88.565 ;
        RECT -33.485 86.875 -33.155 87.205 ;
        RECT -33.485 85.515 -33.155 85.845 ;
        RECT -33.485 84.155 -33.155 84.485 ;
        RECT -33.485 82.795 -33.155 83.125 ;
        RECT -33.485 81.435 -33.155 81.765 ;
        RECT -33.485 80.075 -33.155 80.405 ;
        RECT -33.485 78.715 -33.155 79.045 ;
        RECT -33.485 77.355 -33.155 77.685 ;
        RECT -33.485 75.995 -33.155 76.325 ;
        RECT -33.485 74.635 -33.155 74.965 ;
        RECT -33.485 73.275 -33.155 73.605 ;
        RECT -33.485 71.915 -33.155 72.245 ;
        RECT -33.485 70.555 -33.155 70.885 ;
        RECT -33.485 69.195 -33.155 69.525 ;
        RECT -33.485 67.835 -33.155 68.165 ;
        RECT -33.485 66.475 -33.155 66.805 ;
        RECT -33.485 65.115 -33.155 65.445 ;
        RECT -33.485 63.755 -33.155 64.085 ;
        RECT -33.485 62.395 -33.155 62.725 ;
        RECT -33.485 61.035 -33.155 61.365 ;
        RECT -33.485 59.675 -33.155 60.005 ;
        RECT -33.485 58.315 -33.155 58.645 ;
        RECT -33.485 56.955 -33.155 57.285 ;
        RECT -33.485 55.595 -33.155 55.925 ;
        RECT -33.485 54.235 -33.155 54.565 ;
        RECT -33.485 52.875 -33.155 53.205 ;
        RECT -33.485 51.515 -33.155 51.845 ;
        RECT -33.485 50.155 -33.155 50.485 ;
        RECT -33.485 48.795 -33.155 49.125 ;
        RECT -33.485 47.435 -33.155 47.765 ;
        RECT -33.485 46.075 -33.155 46.405 ;
        RECT -33.485 44.715 -33.155 45.045 ;
        RECT -33.485 43.355 -33.155 43.685 ;
        RECT -33.485 41.995 -33.155 42.325 ;
        RECT -33.485 40.635 -33.155 40.965 ;
        RECT -33.485 39.275 -33.155 39.605 ;
        RECT -33.485 37.915 -33.155 38.245 ;
        RECT -33.485 36.555 -33.155 36.885 ;
        RECT -33.485 35.195 -33.155 35.525 ;
        RECT -33.485 33.835 -33.155 34.165 ;
        RECT -33.485 32.475 -33.155 32.805 ;
        RECT -33.485 31.115 -33.155 31.445 ;
        RECT -33.485 29.755 -33.155 30.085 ;
        RECT -33.485 28.395 -33.155 28.725 ;
        RECT -33.485 27.035 -33.155 27.365 ;
        RECT -33.485 25.675 -33.155 26.005 ;
        RECT -33.485 24.315 -33.155 24.645 ;
        RECT -33.485 22.955 -33.155 23.285 ;
        RECT -33.485 21.595 -33.155 21.925 ;
        RECT -33.485 20.235 -33.155 20.565 ;
        RECT -33.485 18.875 -33.155 19.205 ;
        RECT -33.485 17.515 -33.155 17.845 ;
        RECT -33.485 16.155 -33.155 16.485 ;
        RECT -33.485 14.795 -33.155 15.125 ;
        RECT -33.485 13.435 -33.155 13.765 ;
        RECT -33.485 12.075 -33.155 12.405 ;
        RECT -33.485 10.715 -33.155 11.045 ;
        RECT -33.485 9.355 -33.155 9.685 ;
        RECT -33.485 7.995 -33.155 8.325 ;
        RECT -33.485 6.635 -33.155 6.965 ;
        RECT -33.485 5.275 -33.155 5.605 ;
        RECT -33.485 3.915 -33.155 4.245 ;
        RECT -33.485 2.555 -33.155 2.885 ;
        RECT -33.485 1.195 -33.155 1.525 ;
        RECT -33.485 -0.165 -33.155 0.165 ;
        RECT -33.485 -8.325 -33.155 -7.995 ;
        RECT -33.485 -11.045 -33.155 -10.715 ;
        RECT -33.485 -15.125 -33.155 -14.795 ;
        RECT -33.485 -16.485 -33.155 -16.155 ;
        RECT -33.485 -17.845 -33.155 -17.515 ;
        RECT -33.485 -19.205 -33.155 -18.875 ;
        RECT -33.485 -20.565 -33.155 -20.235 ;
        RECT -33.485 -21.925 -33.155 -21.595 ;
        RECT -33.485 -23.285 -33.155 -22.955 ;
        RECT -33.485 -24.645 -33.155 -24.315 ;
        RECT -33.485 -32.805 -33.155 -32.475 ;
        RECT -33.485 -35.525 -33.155 -35.195 ;
        RECT -33.485 -36.885 -33.155 -36.555 ;
        RECT -33.485 -37.93 -33.155 -37.6 ;
        RECT -33.485 -40.965 -33.155 -40.635 ;
        RECT -33.485 -42.77 -33.155 -42.44 ;
        RECT -33.485 -43.685 -33.155 -43.355 ;
        RECT -33.485 -50.485 -33.155 -50.155 ;
        RECT -33.485 -51.845 -33.155 -51.515 ;
        RECT -33.485 -54.565 -33.155 -54.235 ;
        RECT -33.485 -55.925 -33.155 -55.595 ;
        RECT -33.485 -60.005 -33.155 -59.675 ;
        RECT -33.485 -62.725 -33.155 -62.395 ;
        RECT -33.485 -69.525 -33.155 -69.195 ;
        RECT -33.485 -70.885 -33.155 -70.555 ;
        RECT -33.485 -72.245 -33.155 -71.915 ;
        RECT -33.485 -73.605 -33.155 -73.275 ;
        RECT -33.485 -74.965 -33.155 -74.635 ;
        RECT -33.485 -76.325 -33.155 -75.995 ;
        RECT -33.485 -77.685 -33.155 -77.355 ;
        RECT -33.485 -79.045 -33.155 -78.715 ;
        RECT -33.485 -80.405 -33.155 -80.075 ;
        RECT -33.485 -81.765 -33.155 -81.435 ;
        RECT -33.485 -83.125 -33.155 -82.795 ;
        RECT -33.485 -84.485 -33.155 -84.155 ;
        RECT -33.485 -85.845 -33.155 -85.515 ;
        RECT -33.485 -87.205 -33.155 -86.875 ;
        RECT -33.485 -88.565 -33.155 -88.235 ;
        RECT -33.485 -89.925 -33.155 -89.595 ;
        RECT -33.485 -91.285 -33.155 -90.955 ;
        RECT -33.485 -92.645 -33.155 -92.315 ;
        RECT -33.485 -94.005 -33.155 -93.675 ;
        RECT -33.485 -95.365 -33.155 -95.035 ;
        RECT -33.485 -96.725 -33.155 -96.395 ;
        RECT -33.485 -98.085 -33.155 -97.755 ;
        RECT -33.485 -99.445 -33.155 -99.115 ;
        RECT -33.485 -100.805 -33.155 -100.475 ;
        RECT -33.485 -102.165 -33.155 -101.835 ;
        RECT -33.485 -103.525 -33.155 -103.195 ;
        RECT -33.485 -104.885 -33.155 -104.555 ;
        RECT -33.485 -106.245 -33.155 -105.915 ;
        RECT -33.485 -107.605 -33.155 -107.275 ;
        RECT -33.485 -108.965 -33.155 -108.635 ;
        RECT -33.485 -110.325 -33.155 -109.995 ;
        RECT -33.485 -111.685 -33.155 -111.355 ;
        RECT -33.485 -113.045 -33.155 -112.715 ;
        RECT -33.485 -114.405 -33.155 -114.075 ;
        RECT -33.485 -115.765 -33.155 -115.435 ;
        RECT -33.485 -117.125 -33.155 -116.795 ;
        RECT -33.485 -118.485 -33.155 -118.155 ;
        RECT -33.485 -121.205 -33.155 -120.875 ;
        RECT -33.485 -123.925 -33.155 -123.595 ;
        RECT -33.485 -126.645 -33.155 -126.315 ;
        RECT -33.485 -128.005 -33.155 -127.675 ;
        RECT -33.485 -129.365 -33.155 -129.035 ;
        RECT -33.485 -130.725 -33.155 -130.395 ;
        RECT -33.485 -133.445 -33.155 -133.115 ;
        RECT -33.485 -134.805 -33.155 -134.475 ;
        RECT -33.485 -136.165 -33.155 -135.835 ;
        RECT -33.485 -137.525 -33.155 -137.195 ;
        RECT -33.485 -138.885 -33.155 -138.555 ;
        RECT -33.485 -141.605 -33.155 -141.275 ;
        RECT -33.485 -142.965 -33.155 -142.635 ;
        RECT -33.485 -144.325 -33.155 -143.995 ;
        RECT -33.485 -145.685 -33.155 -145.355 ;
        RECT -33.485 -147.045 -33.155 -146.715 ;
        RECT -33.485 -148.405 -33.155 -148.075 ;
        RECT -33.485 -149.765 -33.155 -149.435 ;
        RECT -33.485 -152.485 -33.155 -152.155 ;
        RECT -33.485 -153.845 -33.155 -153.515 ;
        RECT -33.485 -157.925 -33.155 -157.595 ;
        RECT -33.485 -159.285 -33.155 -158.955 ;
        RECT -33.485 -160.645 -33.155 -160.315 ;
        RECT -33.485 -162.005 -33.155 -161.675 ;
        RECT -33.485 -163.365 -33.155 -163.035 ;
        RECT -33.485 -164.725 -33.155 -164.395 ;
        RECT -33.485 -166.085 -33.155 -165.755 ;
        RECT -33.485 -167.445 -33.155 -167.115 ;
        RECT -33.485 -168.805 -33.155 -168.475 ;
        RECT -33.485 -171.525 -33.155 -171.195 ;
        RECT -33.485 -172.885 -33.155 -172.555 ;
        RECT -33.485 -175.605 -33.155 -175.275 ;
        RECT -33.485 -176.685 -33.155 -176.355 ;
        RECT -33.485 -178.325 -33.155 -177.995 ;
        RECT -33.485 -179.685 -33.155 -179.355 ;
        RECT -33.485 -181.93 -33.155 -180.8 ;
        RECT -33.48 -182.045 -33.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -32.125 241.32 -31.795 242.45 ;
        RECT -32.125 239.195 -31.795 239.525 ;
        RECT -32.125 237.835 -31.795 238.165 ;
        RECT -32.125 236.475 -31.795 236.805 ;
        RECT -32.125 235.115 -31.795 235.445 ;
        RECT -32.125 233.755 -31.795 234.085 ;
        RECT -32.125 232.395 -31.795 232.725 ;
        RECT -32.125 231.035 -31.795 231.365 ;
        RECT -32.125 229.675 -31.795 230.005 ;
        RECT -32.125 228.315 -31.795 228.645 ;
        RECT -32.125 226.955 -31.795 227.285 ;
        RECT -32.125 225.595 -31.795 225.925 ;
        RECT -32.125 224.235 -31.795 224.565 ;
        RECT -32.125 222.875 -31.795 223.205 ;
        RECT -32.125 221.515 -31.795 221.845 ;
        RECT -32.125 220.155 -31.795 220.485 ;
        RECT -32.125 218.795 -31.795 219.125 ;
        RECT -32.125 217.435 -31.795 217.765 ;
        RECT -32.125 216.075 -31.795 216.405 ;
        RECT -32.125 214.715 -31.795 215.045 ;
        RECT -32.125 213.355 -31.795 213.685 ;
        RECT -32.125 211.995 -31.795 212.325 ;
        RECT -32.125 210.635 -31.795 210.965 ;
        RECT -32.125 209.275 -31.795 209.605 ;
        RECT -32.125 207.915 -31.795 208.245 ;
        RECT -32.125 206.555 -31.795 206.885 ;
        RECT -32.125 205.195 -31.795 205.525 ;
        RECT -32.125 203.835 -31.795 204.165 ;
        RECT -32.125 202.475 -31.795 202.805 ;
        RECT -32.125 201.115 -31.795 201.445 ;
        RECT -32.125 199.755 -31.795 200.085 ;
        RECT -32.125 198.395 -31.795 198.725 ;
        RECT -32.125 197.035 -31.795 197.365 ;
        RECT -32.125 195.675 -31.795 196.005 ;
        RECT -32.125 194.315 -31.795 194.645 ;
        RECT -32.125 192.955 -31.795 193.285 ;
        RECT -32.125 191.595 -31.795 191.925 ;
        RECT -32.125 190.235 -31.795 190.565 ;
        RECT -32.125 188.875 -31.795 189.205 ;
        RECT -32.125 187.515 -31.795 187.845 ;
        RECT -32.125 186.155 -31.795 186.485 ;
        RECT -32.125 184.795 -31.795 185.125 ;
        RECT -32.125 183.435 -31.795 183.765 ;
        RECT -32.125 182.075 -31.795 182.405 ;
        RECT -32.125 180.715 -31.795 181.045 ;
        RECT -32.125 179.355 -31.795 179.685 ;
        RECT -32.125 177.995 -31.795 178.325 ;
        RECT -32.125 176.635 -31.795 176.965 ;
        RECT -32.125 175.275 -31.795 175.605 ;
        RECT -32.125 173.915 -31.795 174.245 ;
        RECT -32.125 172.555 -31.795 172.885 ;
        RECT -32.125 171.195 -31.795 171.525 ;
        RECT -32.125 169.835 -31.795 170.165 ;
        RECT -32.125 168.475 -31.795 168.805 ;
        RECT -32.125 167.115 -31.795 167.445 ;
        RECT -32.125 165.755 -31.795 166.085 ;
        RECT -32.125 164.395 -31.795 164.725 ;
        RECT -32.125 163.035 -31.795 163.365 ;
        RECT -32.125 161.675 -31.795 162.005 ;
        RECT -32.125 160.315 -31.795 160.645 ;
        RECT -32.125 158.955 -31.795 159.285 ;
        RECT -32.125 157.595 -31.795 157.925 ;
        RECT -32.125 156.235 -31.795 156.565 ;
        RECT -32.125 154.875 -31.795 155.205 ;
        RECT -32.125 153.515 -31.795 153.845 ;
        RECT -32.125 152.155 -31.795 152.485 ;
        RECT -32.125 150.795 -31.795 151.125 ;
        RECT -32.125 149.435 -31.795 149.765 ;
        RECT -32.125 148.075 -31.795 148.405 ;
        RECT -32.125 146.715 -31.795 147.045 ;
        RECT -32.125 145.355 -31.795 145.685 ;
        RECT -32.125 143.995 -31.795 144.325 ;
        RECT -32.125 142.635 -31.795 142.965 ;
        RECT -32.125 141.275 -31.795 141.605 ;
        RECT -32.125 139.915 -31.795 140.245 ;
        RECT -32.125 138.555 -31.795 138.885 ;
        RECT -32.125 137.195 -31.795 137.525 ;
        RECT -32.125 135.835 -31.795 136.165 ;
        RECT -32.125 134.475 -31.795 134.805 ;
        RECT -32.125 133.115 -31.795 133.445 ;
        RECT -32.125 131.755 -31.795 132.085 ;
        RECT -32.125 130.395 -31.795 130.725 ;
        RECT -32.125 129.035 -31.795 129.365 ;
        RECT -32.125 127.675 -31.795 128.005 ;
        RECT -32.125 126.315 -31.795 126.645 ;
        RECT -32.125 124.955 -31.795 125.285 ;
        RECT -32.125 123.595 -31.795 123.925 ;
        RECT -32.125 122.235 -31.795 122.565 ;
        RECT -32.125 120.875 -31.795 121.205 ;
        RECT -32.125 119.515 -31.795 119.845 ;
        RECT -32.125 118.155 -31.795 118.485 ;
        RECT -32.125 116.795 -31.795 117.125 ;
        RECT -32.125 115.435 -31.795 115.765 ;
        RECT -32.125 114.075 -31.795 114.405 ;
        RECT -32.125 112.715 -31.795 113.045 ;
        RECT -32.125 111.355 -31.795 111.685 ;
        RECT -32.125 109.995 -31.795 110.325 ;
        RECT -32.125 108.635 -31.795 108.965 ;
        RECT -32.125 107.275 -31.795 107.605 ;
        RECT -32.125 105.915 -31.795 106.245 ;
        RECT -32.125 104.555 -31.795 104.885 ;
        RECT -32.125 103.195 -31.795 103.525 ;
        RECT -32.125 101.835 -31.795 102.165 ;
        RECT -32.125 100.475 -31.795 100.805 ;
        RECT -32.125 99.115 -31.795 99.445 ;
        RECT -32.125 97.755 -31.795 98.085 ;
        RECT -32.125 96.395 -31.795 96.725 ;
        RECT -32.125 95.035 -31.795 95.365 ;
        RECT -32.125 93.675 -31.795 94.005 ;
        RECT -32.125 92.315 -31.795 92.645 ;
        RECT -32.125 90.955 -31.795 91.285 ;
        RECT -32.125 89.595 -31.795 89.925 ;
        RECT -32.125 88.235 -31.795 88.565 ;
        RECT -32.125 86.875 -31.795 87.205 ;
        RECT -32.125 85.515 -31.795 85.845 ;
        RECT -32.125 84.155 -31.795 84.485 ;
        RECT -32.125 82.795 -31.795 83.125 ;
        RECT -32.125 81.435 -31.795 81.765 ;
        RECT -32.125 80.075 -31.795 80.405 ;
        RECT -32.125 78.715 -31.795 79.045 ;
        RECT -32.125 77.355 -31.795 77.685 ;
        RECT -32.125 75.995 -31.795 76.325 ;
        RECT -32.125 74.635 -31.795 74.965 ;
        RECT -32.125 73.275 -31.795 73.605 ;
        RECT -32.125 71.915 -31.795 72.245 ;
        RECT -32.125 70.555 -31.795 70.885 ;
        RECT -32.125 69.195 -31.795 69.525 ;
        RECT -32.125 67.835 -31.795 68.165 ;
        RECT -32.125 66.475 -31.795 66.805 ;
        RECT -32.125 65.115 -31.795 65.445 ;
        RECT -32.125 63.755 -31.795 64.085 ;
        RECT -32.125 62.395 -31.795 62.725 ;
        RECT -32.125 61.035 -31.795 61.365 ;
        RECT -32.125 59.675 -31.795 60.005 ;
        RECT -32.125 58.315 -31.795 58.645 ;
        RECT -32.125 56.955 -31.795 57.285 ;
        RECT -32.125 55.595 -31.795 55.925 ;
        RECT -32.125 54.235 -31.795 54.565 ;
        RECT -32.125 52.875 -31.795 53.205 ;
        RECT -32.125 51.515 -31.795 51.845 ;
        RECT -32.125 50.155 -31.795 50.485 ;
        RECT -32.125 48.795 -31.795 49.125 ;
        RECT -32.125 47.435 -31.795 47.765 ;
        RECT -32.125 46.075 -31.795 46.405 ;
        RECT -32.125 44.715 -31.795 45.045 ;
        RECT -32.125 43.355 -31.795 43.685 ;
        RECT -32.125 41.995 -31.795 42.325 ;
        RECT -32.125 40.635 -31.795 40.965 ;
        RECT -32.125 39.275 -31.795 39.605 ;
        RECT -32.125 37.915 -31.795 38.245 ;
        RECT -32.125 36.555 -31.795 36.885 ;
        RECT -32.125 35.195 -31.795 35.525 ;
        RECT -32.125 33.835 -31.795 34.165 ;
        RECT -32.125 32.475 -31.795 32.805 ;
        RECT -32.125 31.115 -31.795 31.445 ;
        RECT -32.125 29.755 -31.795 30.085 ;
        RECT -32.125 28.395 -31.795 28.725 ;
        RECT -32.125 27.035 -31.795 27.365 ;
        RECT -32.125 25.675 -31.795 26.005 ;
        RECT -32.125 24.315 -31.795 24.645 ;
        RECT -32.125 22.955 -31.795 23.285 ;
        RECT -32.125 21.595 -31.795 21.925 ;
        RECT -32.125 20.235 -31.795 20.565 ;
        RECT -32.125 18.875 -31.795 19.205 ;
        RECT -32.125 17.515 -31.795 17.845 ;
        RECT -32.125 16.155 -31.795 16.485 ;
        RECT -32.125 14.795 -31.795 15.125 ;
        RECT -32.125 13.435 -31.795 13.765 ;
        RECT -32.125 12.075 -31.795 12.405 ;
        RECT -32.125 10.715 -31.795 11.045 ;
        RECT -32.125 9.355 -31.795 9.685 ;
        RECT -32.125 7.995 -31.795 8.325 ;
        RECT -32.125 6.635 -31.795 6.965 ;
        RECT -32.125 5.275 -31.795 5.605 ;
        RECT -32.125 3.915 -31.795 4.245 ;
        RECT -32.125 2.555 -31.795 2.885 ;
        RECT -32.125 1.195 -31.795 1.525 ;
        RECT -32.125 -0.165 -31.795 0.165 ;
        RECT -32.125 -8.325 -31.795 -7.995 ;
        RECT -32.125 -11.045 -31.795 -10.715 ;
        RECT -32.125 -15.125 -31.795 -14.795 ;
        RECT -32.125 -16.485 -31.795 -16.155 ;
        RECT -32.125 -17.845 -31.795 -17.515 ;
        RECT -32.125 -19.205 -31.795 -18.875 ;
        RECT -32.125 -20.565 -31.795 -20.235 ;
        RECT -32.125 -21.925 -31.795 -21.595 ;
        RECT -32.125 -23.285 -31.795 -22.955 ;
        RECT -32.125 -24.645 -31.795 -24.315 ;
        RECT -32.125 -32.805 -31.795 -32.475 ;
        RECT -32.125 -35.525 -31.795 -35.195 ;
        RECT -32.125 -36.885 -31.795 -36.555 ;
        RECT -32.125 -37.93 -31.795 -37.6 ;
        RECT -32.125 -40.965 -31.795 -40.635 ;
        RECT -32.125 -42.77 -31.795 -42.44 ;
        RECT -32.125 -43.685 -31.795 -43.355 ;
        RECT -32.125 -50.485 -31.795 -50.155 ;
        RECT -32.125 -51.845 -31.795 -51.515 ;
        RECT -32.125 -54.565 -31.795 -54.235 ;
        RECT -32.125 -55.925 -31.795 -55.595 ;
        RECT -32.125 -60.005 -31.795 -59.675 ;
        RECT -32.125 -62.725 -31.795 -62.395 ;
        RECT -32.125 -69.525 -31.795 -69.195 ;
        RECT -32.125 -70.885 -31.795 -70.555 ;
        RECT -32.125 -72.245 -31.795 -71.915 ;
        RECT -32.125 -73.605 -31.795 -73.275 ;
        RECT -32.125 -74.965 -31.795 -74.635 ;
        RECT -32.125 -76.325 -31.795 -75.995 ;
        RECT -32.125 -77.685 -31.795 -77.355 ;
        RECT -32.125 -79.045 -31.795 -78.715 ;
        RECT -32.125 -80.405 -31.795 -80.075 ;
        RECT -32.125 -81.765 -31.795 -81.435 ;
        RECT -32.125 -83.125 -31.795 -82.795 ;
        RECT -32.125 -84.485 -31.795 -84.155 ;
        RECT -32.125 -85.845 -31.795 -85.515 ;
        RECT -32.125 -87.205 -31.795 -86.875 ;
        RECT -32.125 -88.565 -31.795 -88.235 ;
        RECT -32.125 -89.925 -31.795 -89.595 ;
        RECT -32.125 -91.285 -31.795 -90.955 ;
        RECT -32.125 -92.645 -31.795 -92.315 ;
        RECT -32.125 -94.005 -31.795 -93.675 ;
        RECT -32.125 -95.365 -31.795 -95.035 ;
        RECT -32.125 -96.725 -31.795 -96.395 ;
        RECT -32.125 -98.085 -31.795 -97.755 ;
        RECT -32.125 -99.445 -31.795 -99.115 ;
        RECT -32.125 -100.805 -31.795 -100.475 ;
        RECT -32.125 -102.165 -31.795 -101.835 ;
        RECT -32.125 -103.525 -31.795 -103.195 ;
        RECT -32.125 -104.885 -31.795 -104.555 ;
        RECT -32.125 -106.245 -31.795 -105.915 ;
        RECT -32.125 -107.605 -31.795 -107.275 ;
        RECT -32.125 -108.965 -31.795 -108.635 ;
        RECT -32.125 -110.325 -31.795 -109.995 ;
        RECT -32.125 -111.685 -31.795 -111.355 ;
        RECT -32.125 -113.045 -31.795 -112.715 ;
        RECT -32.125 -114.405 -31.795 -114.075 ;
        RECT -32.125 -115.765 -31.795 -115.435 ;
        RECT -32.125 -117.125 -31.795 -116.795 ;
        RECT -32.125 -118.485 -31.795 -118.155 ;
        RECT -32.125 -121.205 -31.795 -120.875 ;
        RECT -32.125 -123.925 -31.795 -123.595 ;
        RECT -32.125 -126.645 -31.795 -126.315 ;
        RECT -32.125 -128.005 -31.795 -127.675 ;
        RECT -32.125 -129.365 -31.795 -129.035 ;
        RECT -32.125 -130.725 -31.795 -130.395 ;
        RECT -32.125 -133.445 -31.795 -133.115 ;
        RECT -32.125 -134.805 -31.795 -134.475 ;
        RECT -32.125 -136.165 -31.795 -135.835 ;
        RECT -32.125 -137.525 -31.795 -137.195 ;
        RECT -32.125 -141.605 -31.795 -141.275 ;
        RECT -32.125 -142.965 -31.795 -142.635 ;
        RECT -32.125 -144.325 -31.795 -143.995 ;
        RECT -32.125 -145.685 -31.795 -145.355 ;
        RECT -32.125 -147.045 -31.795 -146.715 ;
        RECT -32.125 -148.405 -31.795 -148.075 ;
        RECT -32.125 -149.765 -31.795 -149.435 ;
        RECT -32.125 -152.485 -31.795 -152.155 ;
        RECT -32.125 -153.845 -31.795 -153.515 ;
        RECT -32.125 -157.925 -31.795 -157.595 ;
        RECT -32.125 -159.285 -31.795 -158.955 ;
        RECT -32.125 -160.645 -31.795 -160.315 ;
        RECT -32.125 -162.005 -31.795 -161.675 ;
        RECT -32.125 -163.365 -31.795 -163.035 ;
        RECT -32.125 -164.725 -31.795 -164.395 ;
        RECT -32.125 -166.085 -31.795 -165.755 ;
        RECT -32.125 -167.445 -31.795 -167.115 ;
        RECT -32.125 -168.805 -31.795 -168.475 ;
        RECT -32.125 -171.525 -31.795 -171.195 ;
        RECT -32.125 -172.885 -31.795 -172.555 ;
        RECT -32.125 -174.245 -31.795 -173.915 ;
        RECT -32.125 -175.605 -31.795 -175.275 ;
        RECT -32.125 -176.685 -31.795 -176.355 ;
        RECT -32.125 -178.325 -31.795 -177.995 ;
        RECT -32.125 -179.685 -31.795 -179.355 ;
        RECT -32.125 -181.93 -31.795 -180.8 ;
        RECT -32.12 -182.045 -31.8 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -30.765 133.115 -30.435 133.445 ;
        RECT -30.765 131.755 -30.435 132.085 ;
        RECT -30.765 130.395 -30.435 130.725 ;
        RECT -30.765 129.035 -30.435 129.365 ;
        RECT -30.765 127.675 -30.435 128.005 ;
        RECT -30.765 126.315 -30.435 126.645 ;
        RECT -30.765 124.955 -30.435 125.285 ;
        RECT -30.765 123.595 -30.435 123.925 ;
        RECT -30.765 122.235 -30.435 122.565 ;
        RECT -30.765 120.875 -30.435 121.205 ;
        RECT -30.765 119.515 -30.435 119.845 ;
        RECT -30.765 118.155 -30.435 118.485 ;
        RECT -30.765 116.795 -30.435 117.125 ;
        RECT -30.765 115.435 -30.435 115.765 ;
        RECT -30.765 114.075 -30.435 114.405 ;
        RECT -30.765 112.715 -30.435 113.045 ;
        RECT -30.765 111.355 -30.435 111.685 ;
        RECT -30.765 109.995 -30.435 110.325 ;
        RECT -30.765 108.635 -30.435 108.965 ;
        RECT -30.765 107.275 -30.435 107.605 ;
        RECT -30.765 105.915 -30.435 106.245 ;
        RECT -30.765 104.555 -30.435 104.885 ;
        RECT -30.765 103.195 -30.435 103.525 ;
        RECT -30.765 101.835 -30.435 102.165 ;
        RECT -30.765 100.475 -30.435 100.805 ;
        RECT -30.765 99.115 -30.435 99.445 ;
        RECT -30.765 97.755 -30.435 98.085 ;
        RECT -30.765 96.395 -30.435 96.725 ;
        RECT -30.765 95.035 -30.435 95.365 ;
        RECT -30.765 93.675 -30.435 94.005 ;
        RECT -30.765 92.315 -30.435 92.645 ;
        RECT -30.765 90.955 -30.435 91.285 ;
        RECT -30.765 89.595 -30.435 89.925 ;
        RECT -30.765 88.235 -30.435 88.565 ;
        RECT -30.765 86.875 -30.435 87.205 ;
        RECT -30.765 85.515 -30.435 85.845 ;
        RECT -30.765 84.155 -30.435 84.485 ;
        RECT -30.765 82.795 -30.435 83.125 ;
        RECT -30.765 81.435 -30.435 81.765 ;
        RECT -30.765 80.075 -30.435 80.405 ;
        RECT -30.765 78.715 -30.435 79.045 ;
        RECT -30.765 77.355 -30.435 77.685 ;
        RECT -30.765 75.995 -30.435 76.325 ;
        RECT -30.765 74.635 -30.435 74.965 ;
        RECT -30.765 73.275 -30.435 73.605 ;
        RECT -30.765 71.915 -30.435 72.245 ;
        RECT -30.765 70.555 -30.435 70.885 ;
        RECT -30.765 69.195 -30.435 69.525 ;
        RECT -30.765 67.835 -30.435 68.165 ;
        RECT -30.765 66.475 -30.435 66.805 ;
        RECT -30.765 65.115 -30.435 65.445 ;
        RECT -30.765 63.755 -30.435 64.085 ;
        RECT -30.765 62.395 -30.435 62.725 ;
        RECT -30.765 61.035 -30.435 61.365 ;
        RECT -30.765 59.675 -30.435 60.005 ;
        RECT -30.765 58.315 -30.435 58.645 ;
        RECT -30.765 56.955 -30.435 57.285 ;
        RECT -30.765 55.595 -30.435 55.925 ;
        RECT -30.765 54.235 -30.435 54.565 ;
        RECT -30.765 52.875 -30.435 53.205 ;
        RECT -30.765 51.515 -30.435 51.845 ;
        RECT -30.765 50.155 -30.435 50.485 ;
        RECT -30.765 48.795 -30.435 49.125 ;
        RECT -30.765 47.435 -30.435 47.765 ;
        RECT -30.765 46.075 -30.435 46.405 ;
        RECT -30.765 44.715 -30.435 45.045 ;
        RECT -30.765 43.355 -30.435 43.685 ;
        RECT -30.765 41.995 -30.435 42.325 ;
        RECT -30.765 40.635 -30.435 40.965 ;
        RECT -30.765 39.275 -30.435 39.605 ;
        RECT -30.765 37.915 -30.435 38.245 ;
        RECT -30.765 36.555 -30.435 36.885 ;
        RECT -30.765 35.195 -30.435 35.525 ;
        RECT -30.765 33.835 -30.435 34.165 ;
        RECT -30.765 32.475 -30.435 32.805 ;
        RECT -30.765 31.115 -30.435 31.445 ;
        RECT -30.765 29.755 -30.435 30.085 ;
        RECT -30.765 28.395 -30.435 28.725 ;
        RECT -30.765 27.035 -30.435 27.365 ;
        RECT -30.765 25.675 -30.435 26.005 ;
        RECT -30.765 24.315 -30.435 24.645 ;
        RECT -30.765 22.955 -30.435 23.285 ;
        RECT -30.765 21.595 -30.435 21.925 ;
        RECT -30.765 20.235 -30.435 20.565 ;
        RECT -30.765 18.875 -30.435 19.205 ;
        RECT -30.765 17.515 -30.435 17.845 ;
        RECT -30.765 16.155 -30.435 16.485 ;
        RECT -30.765 14.795 -30.435 15.125 ;
        RECT -30.765 13.435 -30.435 13.765 ;
        RECT -30.765 12.075 -30.435 12.405 ;
        RECT -30.765 10.715 -30.435 11.045 ;
        RECT -30.765 9.355 -30.435 9.685 ;
        RECT -30.765 7.995 -30.435 8.325 ;
        RECT -30.765 6.635 -30.435 6.965 ;
        RECT -30.765 5.275 -30.435 5.605 ;
        RECT -30.765 3.915 -30.435 4.245 ;
        RECT -30.765 2.555 -30.435 2.885 ;
        RECT -30.765 1.195 -30.435 1.525 ;
        RECT -30.765 -0.165 -30.435 0.165 ;
        RECT -30.765 -8.325 -30.435 -7.995 ;
        RECT -30.765 -9.685 -30.435 -9.355 ;
        RECT -30.765 -11.045 -30.435 -10.715 ;
        RECT -30.765 -15.125 -30.435 -14.795 ;
        RECT -30.765 -16.485 -30.435 -16.155 ;
        RECT -30.765 -17.845 -30.435 -17.515 ;
        RECT -30.765 -19.205 -30.435 -18.875 ;
        RECT -30.765 -20.565 -30.435 -20.235 ;
        RECT -30.765 -21.925 -30.435 -21.595 ;
        RECT -30.765 -23.285 -30.435 -22.955 ;
        RECT -30.765 -24.645 -30.435 -24.315 ;
        RECT -30.765 -32.805 -30.435 -32.475 ;
        RECT -30.765 -35.525 -30.435 -35.195 ;
        RECT -30.765 -36.885 -30.435 -36.555 ;
        RECT -30.765 -37.93 -30.435 -37.6 ;
        RECT -30.765 -40.965 -30.435 -40.635 ;
        RECT -30.765 -42.77 -30.435 -42.44 ;
        RECT -30.765 -43.685 -30.435 -43.355 ;
        RECT -30.765 -50.485 -30.435 -50.155 ;
        RECT -30.765 -51.845 -30.435 -51.515 ;
        RECT -30.765 -54.565 -30.435 -54.235 ;
        RECT -30.765 -55.925 -30.435 -55.595 ;
        RECT -30.765 -60.005 -30.435 -59.675 ;
        RECT -30.765 -62.725 -30.435 -62.395 ;
        RECT -30.76 -64.76 -30.44 242.565 ;
        RECT -30.765 241.32 -30.435 242.45 ;
        RECT -30.765 239.195 -30.435 239.525 ;
        RECT -30.765 237.835 -30.435 238.165 ;
        RECT -30.765 236.475 -30.435 236.805 ;
        RECT -30.765 235.115 -30.435 235.445 ;
        RECT -30.765 233.755 -30.435 234.085 ;
        RECT -30.765 232.395 -30.435 232.725 ;
        RECT -30.765 231.035 -30.435 231.365 ;
        RECT -30.765 229.675 -30.435 230.005 ;
        RECT -30.765 228.315 -30.435 228.645 ;
        RECT -30.765 226.955 -30.435 227.285 ;
        RECT -30.765 225.595 -30.435 225.925 ;
        RECT -30.765 224.235 -30.435 224.565 ;
        RECT -30.765 222.875 -30.435 223.205 ;
        RECT -30.765 221.515 -30.435 221.845 ;
        RECT -30.765 220.155 -30.435 220.485 ;
        RECT -30.765 218.795 -30.435 219.125 ;
        RECT -30.765 217.435 -30.435 217.765 ;
        RECT -30.765 216.075 -30.435 216.405 ;
        RECT -30.765 214.715 -30.435 215.045 ;
        RECT -30.765 213.355 -30.435 213.685 ;
        RECT -30.765 211.995 -30.435 212.325 ;
        RECT -30.765 210.635 -30.435 210.965 ;
        RECT -30.765 209.275 -30.435 209.605 ;
        RECT -30.765 207.915 -30.435 208.245 ;
        RECT -30.765 206.555 -30.435 206.885 ;
        RECT -30.765 205.195 -30.435 205.525 ;
        RECT -30.765 203.835 -30.435 204.165 ;
        RECT -30.765 202.475 -30.435 202.805 ;
        RECT -30.765 201.115 -30.435 201.445 ;
        RECT -30.765 199.755 -30.435 200.085 ;
        RECT -30.765 198.395 -30.435 198.725 ;
        RECT -30.765 197.035 -30.435 197.365 ;
        RECT -30.765 195.675 -30.435 196.005 ;
        RECT -30.765 194.315 -30.435 194.645 ;
        RECT -30.765 192.955 -30.435 193.285 ;
        RECT -30.765 191.595 -30.435 191.925 ;
        RECT -30.765 190.235 -30.435 190.565 ;
        RECT -30.765 188.875 -30.435 189.205 ;
        RECT -30.765 187.515 -30.435 187.845 ;
        RECT -30.765 186.155 -30.435 186.485 ;
        RECT -30.765 184.795 -30.435 185.125 ;
        RECT -30.765 183.435 -30.435 183.765 ;
        RECT -30.765 182.075 -30.435 182.405 ;
        RECT -30.765 180.715 -30.435 181.045 ;
        RECT -30.765 179.355 -30.435 179.685 ;
        RECT -30.765 177.995 -30.435 178.325 ;
        RECT -30.765 176.635 -30.435 176.965 ;
        RECT -30.765 175.275 -30.435 175.605 ;
        RECT -30.765 173.915 -30.435 174.245 ;
        RECT -30.765 172.555 -30.435 172.885 ;
        RECT -30.765 171.195 -30.435 171.525 ;
        RECT -30.765 169.835 -30.435 170.165 ;
        RECT -30.765 168.475 -30.435 168.805 ;
        RECT -30.765 167.115 -30.435 167.445 ;
        RECT -30.765 165.755 -30.435 166.085 ;
        RECT -30.765 164.395 -30.435 164.725 ;
        RECT -30.765 163.035 -30.435 163.365 ;
        RECT -30.765 161.675 -30.435 162.005 ;
        RECT -30.765 160.315 -30.435 160.645 ;
        RECT -30.765 158.955 -30.435 159.285 ;
        RECT -30.765 157.595 -30.435 157.925 ;
        RECT -30.765 156.235 -30.435 156.565 ;
        RECT -30.765 154.875 -30.435 155.205 ;
        RECT -30.765 153.515 -30.435 153.845 ;
        RECT -30.765 152.155 -30.435 152.485 ;
        RECT -30.765 150.795 -30.435 151.125 ;
        RECT -30.765 149.435 -30.435 149.765 ;
        RECT -30.765 148.075 -30.435 148.405 ;
        RECT -30.765 146.715 -30.435 147.045 ;
        RECT -30.765 145.355 -30.435 145.685 ;
        RECT -30.765 143.995 -30.435 144.325 ;
        RECT -30.765 142.635 -30.435 142.965 ;
        RECT -30.765 141.275 -30.435 141.605 ;
        RECT -30.765 139.915 -30.435 140.245 ;
        RECT -30.765 138.555 -30.435 138.885 ;
        RECT -30.765 137.195 -30.435 137.525 ;
        RECT -30.765 135.835 -30.435 136.165 ;
        RECT -30.765 134.475 -30.435 134.805 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.925 241.32 -38.595 242.45 ;
        RECT -38.925 239.195 -38.595 239.525 ;
        RECT -38.925 237.835 -38.595 238.165 ;
        RECT -38.925 236.475 -38.595 236.805 ;
        RECT -38.925 235.115 -38.595 235.445 ;
        RECT -38.925 233.755 -38.595 234.085 ;
        RECT -38.925 232.395 -38.595 232.725 ;
        RECT -38.925 231.035 -38.595 231.365 ;
        RECT -38.925 229.675 -38.595 230.005 ;
        RECT -38.925 228.315 -38.595 228.645 ;
        RECT -38.925 226.955 -38.595 227.285 ;
        RECT -38.925 225.595 -38.595 225.925 ;
        RECT -38.925 224.235 -38.595 224.565 ;
        RECT -38.925 222.875 -38.595 223.205 ;
        RECT -38.925 221.515 -38.595 221.845 ;
        RECT -38.925 220.155 -38.595 220.485 ;
        RECT -38.925 218.795 -38.595 219.125 ;
        RECT -38.925 217.435 -38.595 217.765 ;
        RECT -38.925 216.075 -38.595 216.405 ;
        RECT -38.925 214.715 -38.595 215.045 ;
        RECT -38.925 213.355 -38.595 213.685 ;
        RECT -38.925 211.995 -38.595 212.325 ;
        RECT -38.925 210.635 -38.595 210.965 ;
        RECT -38.925 209.275 -38.595 209.605 ;
        RECT -38.925 207.915 -38.595 208.245 ;
        RECT -38.925 206.555 -38.595 206.885 ;
        RECT -38.925 205.195 -38.595 205.525 ;
        RECT -38.925 203.835 -38.595 204.165 ;
        RECT -38.925 202.475 -38.595 202.805 ;
        RECT -38.925 201.115 -38.595 201.445 ;
        RECT -38.925 199.755 -38.595 200.085 ;
        RECT -38.925 198.395 -38.595 198.725 ;
        RECT -38.925 197.035 -38.595 197.365 ;
        RECT -38.925 195.675 -38.595 196.005 ;
        RECT -38.925 194.315 -38.595 194.645 ;
        RECT -38.925 192.955 -38.595 193.285 ;
        RECT -38.925 191.595 -38.595 191.925 ;
        RECT -38.925 190.235 -38.595 190.565 ;
        RECT -38.925 188.875 -38.595 189.205 ;
        RECT -38.925 187.515 -38.595 187.845 ;
        RECT -38.925 186.155 -38.595 186.485 ;
        RECT -38.925 184.795 -38.595 185.125 ;
        RECT -38.925 183.435 -38.595 183.765 ;
        RECT -38.925 182.075 -38.595 182.405 ;
        RECT -38.925 180.715 -38.595 181.045 ;
        RECT -38.925 179.355 -38.595 179.685 ;
        RECT -38.925 177.995 -38.595 178.325 ;
        RECT -38.925 176.635 -38.595 176.965 ;
        RECT -38.925 175.275 -38.595 175.605 ;
        RECT -38.925 173.915 -38.595 174.245 ;
        RECT -38.925 172.555 -38.595 172.885 ;
        RECT -38.925 171.195 -38.595 171.525 ;
        RECT -38.925 169.835 -38.595 170.165 ;
        RECT -38.925 168.475 -38.595 168.805 ;
        RECT -38.925 167.115 -38.595 167.445 ;
        RECT -38.925 165.755 -38.595 166.085 ;
        RECT -38.925 164.395 -38.595 164.725 ;
        RECT -38.925 163.035 -38.595 163.365 ;
        RECT -38.925 161.675 -38.595 162.005 ;
        RECT -38.925 160.315 -38.595 160.645 ;
        RECT -38.925 158.955 -38.595 159.285 ;
        RECT -38.925 157.595 -38.595 157.925 ;
        RECT -38.925 156.235 -38.595 156.565 ;
        RECT -38.925 154.875 -38.595 155.205 ;
        RECT -38.925 153.515 -38.595 153.845 ;
        RECT -38.925 152.155 -38.595 152.485 ;
        RECT -38.925 150.795 -38.595 151.125 ;
        RECT -38.925 149.435 -38.595 149.765 ;
        RECT -38.925 148.075 -38.595 148.405 ;
        RECT -38.925 146.715 -38.595 147.045 ;
        RECT -38.925 145.355 -38.595 145.685 ;
        RECT -38.925 143.995 -38.595 144.325 ;
        RECT -38.925 142.635 -38.595 142.965 ;
        RECT -38.925 141.275 -38.595 141.605 ;
        RECT -38.925 139.915 -38.595 140.245 ;
        RECT -38.925 138.555 -38.595 138.885 ;
        RECT -38.925 137.195 -38.595 137.525 ;
        RECT -38.925 135.835 -38.595 136.165 ;
        RECT -38.925 134.475 -38.595 134.805 ;
        RECT -38.925 133.115 -38.595 133.445 ;
        RECT -38.925 131.755 -38.595 132.085 ;
        RECT -38.925 130.395 -38.595 130.725 ;
        RECT -38.925 129.035 -38.595 129.365 ;
        RECT -38.925 127.675 -38.595 128.005 ;
        RECT -38.925 126.315 -38.595 126.645 ;
        RECT -38.925 124.955 -38.595 125.285 ;
        RECT -38.925 123.595 -38.595 123.925 ;
        RECT -38.925 122.235 -38.595 122.565 ;
        RECT -38.925 120.875 -38.595 121.205 ;
        RECT -38.925 119.515 -38.595 119.845 ;
        RECT -38.925 118.155 -38.595 118.485 ;
        RECT -38.925 116.795 -38.595 117.125 ;
        RECT -38.925 115.435 -38.595 115.765 ;
        RECT -38.925 114.075 -38.595 114.405 ;
        RECT -38.925 112.715 -38.595 113.045 ;
        RECT -38.925 111.355 -38.595 111.685 ;
        RECT -38.925 109.995 -38.595 110.325 ;
        RECT -38.925 108.635 -38.595 108.965 ;
        RECT -38.925 107.275 -38.595 107.605 ;
        RECT -38.925 105.915 -38.595 106.245 ;
        RECT -38.925 104.555 -38.595 104.885 ;
        RECT -38.925 103.195 -38.595 103.525 ;
        RECT -38.925 101.835 -38.595 102.165 ;
        RECT -38.925 100.475 -38.595 100.805 ;
        RECT -38.925 99.115 -38.595 99.445 ;
        RECT -38.925 97.755 -38.595 98.085 ;
        RECT -38.925 96.395 -38.595 96.725 ;
        RECT -38.925 95.035 -38.595 95.365 ;
        RECT -38.925 93.675 -38.595 94.005 ;
        RECT -38.925 92.315 -38.595 92.645 ;
        RECT -38.925 90.955 -38.595 91.285 ;
        RECT -38.925 89.595 -38.595 89.925 ;
        RECT -38.925 88.235 -38.595 88.565 ;
        RECT -38.925 86.875 -38.595 87.205 ;
        RECT -38.925 85.515 -38.595 85.845 ;
        RECT -38.925 84.155 -38.595 84.485 ;
        RECT -38.925 82.795 -38.595 83.125 ;
        RECT -38.925 81.435 -38.595 81.765 ;
        RECT -38.925 80.075 -38.595 80.405 ;
        RECT -38.925 78.715 -38.595 79.045 ;
        RECT -38.925 77.355 -38.595 77.685 ;
        RECT -38.925 75.995 -38.595 76.325 ;
        RECT -38.925 74.635 -38.595 74.965 ;
        RECT -38.925 73.275 -38.595 73.605 ;
        RECT -38.925 71.915 -38.595 72.245 ;
        RECT -38.925 70.555 -38.595 70.885 ;
        RECT -38.925 69.195 -38.595 69.525 ;
        RECT -38.925 67.835 -38.595 68.165 ;
        RECT -38.925 66.475 -38.595 66.805 ;
        RECT -38.925 65.115 -38.595 65.445 ;
        RECT -38.925 63.755 -38.595 64.085 ;
        RECT -38.925 62.395 -38.595 62.725 ;
        RECT -38.925 61.035 -38.595 61.365 ;
        RECT -38.925 59.675 -38.595 60.005 ;
        RECT -38.925 58.315 -38.595 58.645 ;
        RECT -38.925 56.955 -38.595 57.285 ;
        RECT -38.925 55.595 -38.595 55.925 ;
        RECT -38.925 54.235 -38.595 54.565 ;
        RECT -38.925 52.875 -38.595 53.205 ;
        RECT -38.925 51.515 -38.595 51.845 ;
        RECT -38.925 50.155 -38.595 50.485 ;
        RECT -38.925 48.795 -38.595 49.125 ;
        RECT -38.925 47.435 -38.595 47.765 ;
        RECT -38.925 46.075 -38.595 46.405 ;
        RECT -38.925 44.715 -38.595 45.045 ;
        RECT -38.925 43.355 -38.595 43.685 ;
        RECT -38.925 41.995 -38.595 42.325 ;
        RECT -38.925 40.635 -38.595 40.965 ;
        RECT -38.925 39.275 -38.595 39.605 ;
        RECT -38.925 37.915 -38.595 38.245 ;
        RECT -38.925 36.555 -38.595 36.885 ;
        RECT -38.925 35.195 -38.595 35.525 ;
        RECT -38.925 33.835 -38.595 34.165 ;
        RECT -38.925 32.475 -38.595 32.805 ;
        RECT -38.925 31.115 -38.595 31.445 ;
        RECT -38.925 29.755 -38.595 30.085 ;
        RECT -38.925 28.395 -38.595 28.725 ;
        RECT -38.925 27.035 -38.595 27.365 ;
        RECT -38.925 25.675 -38.595 26.005 ;
        RECT -38.925 24.315 -38.595 24.645 ;
        RECT -38.925 22.955 -38.595 23.285 ;
        RECT -38.925 21.595 -38.595 21.925 ;
        RECT -38.925 20.235 -38.595 20.565 ;
        RECT -38.925 18.875 -38.595 19.205 ;
        RECT -38.925 17.515 -38.595 17.845 ;
        RECT -38.925 16.155 -38.595 16.485 ;
        RECT -38.925 14.795 -38.595 15.125 ;
        RECT -38.925 13.435 -38.595 13.765 ;
        RECT -38.925 12.075 -38.595 12.405 ;
        RECT -38.925 10.715 -38.595 11.045 ;
        RECT -38.925 9.355 -38.595 9.685 ;
        RECT -38.925 7.995 -38.595 8.325 ;
        RECT -38.925 6.635 -38.595 6.965 ;
        RECT -38.925 5.275 -38.595 5.605 ;
        RECT -38.925 3.915 -38.595 4.245 ;
        RECT -38.925 2.555 -38.595 2.885 ;
        RECT -38.925 1.195 -38.595 1.525 ;
        RECT -38.925 -0.165 -38.595 0.165 ;
        RECT -38.925 -2.885 -38.595 -2.555 ;
        RECT -38.925 -4.245 -38.595 -3.915 ;
        RECT -38.925 -11.045 -38.595 -10.715 ;
        RECT -38.925 -15.125 -38.595 -14.795 ;
        RECT -38.925 -16.485 -38.595 -16.155 ;
        RECT -38.925 -17.845 -38.595 -17.515 ;
        RECT -38.925 -19.205 -38.595 -18.875 ;
        RECT -38.925 -20.565 -38.595 -20.235 ;
        RECT -38.925 -21.925 -38.595 -21.595 ;
        RECT -38.925 -23.285 -38.595 -22.955 ;
        RECT -38.925 -24.645 -38.595 -24.315 ;
        RECT -38.925 -32.805 -38.595 -32.475 ;
        RECT -38.925 -35.525 -38.595 -35.195 ;
        RECT -38.925 -36.885 -38.595 -36.555 ;
        RECT -38.925 -37.93 -38.595 -37.6 ;
        RECT -38.925 -40.965 -38.595 -40.635 ;
        RECT -38.925 -42.77 -38.595 -42.44 ;
        RECT -38.925 -43.685 -38.595 -43.355 ;
        RECT -38.925 -50.485 -38.595 -50.155 ;
        RECT -38.925 -51.845 -38.595 -51.515 ;
        RECT -38.925 -54.565 -38.595 -54.235 ;
        RECT -38.925 -55.925 -38.595 -55.595 ;
        RECT -38.925 -60.005 -38.595 -59.675 ;
        RECT -38.925 -62.725 -38.595 -62.395 ;
        RECT -38.925 -69.525 -38.595 -69.195 ;
        RECT -38.925 -70.885 -38.595 -70.555 ;
        RECT -38.925 -72.245 -38.595 -71.915 ;
        RECT -38.925 -73.605 -38.595 -73.275 ;
        RECT -38.925 -74.965 -38.595 -74.635 ;
        RECT -38.925 -76.325 -38.595 -75.995 ;
        RECT -38.925 -77.685 -38.595 -77.355 ;
        RECT -38.925 -79.045 -38.595 -78.715 ;
        RECT -38.925 -80.405 -38.595 -80.075 ;
        RECT -38.925 -81.765 -38.595 -81.435 ;
        RECT -38.925 -83.125 -38.595 -82.795 ;
        RECT -38.925 -84.485 -38.595 -84.155 ;
        RECT -38.925 -85.845 -38.595 -85.515 ;
        RECT -38.925 -87.205 -38.595 -86.875 ;
        RECT -38.925 -88.565 -38.595 -88.235 ;
        RECT -38.925 -89.925 -38.595 -89.595 ;
        RECT -38.925 -92.645 -38.595 -92.315 ;
        RECT -38.925 -94.005 -38.595 -93.675 ;
        RECT -38.925 -95.365 -38.595 -95.035 ;
        RECT -38.925 -96.725 -38.595 -96.395 ;
        RECT -38.925 -98.085 -38.595 -97.755 ;
        RECT -38.925 -99.69 -38.595 -99.36 ;
        RECT -38.925 -100.805 -38.595 -100.475 ;
        RECT -38.925 -103.525 -38.595 -103.195 ;
        RECT -38.925 -104.885 -38.595 -104.555 ;
        RECT -38.925 -106.245 -38.595 -105.915 ;
        RECT -38.925 -107.83 -38.595 -107.5 ;
        RECT -38.925 -108.965 -38.595 -108.635 ;
        RECT -38.925 -110.325 -38.595 -109.995 ;
        RECT -38.925 -111.685 -38.595 -111.355 ;
        RECT -38.925 -115.765 -38.595 -115.435 ;
        RECT -38.925 -117.125 -38.595 -116.795 ;
        RECT -38.925 -118.485 -38.595 -118.155 ;
        RECT -38.925 -121.205 -38.595 -120.875 ;
        RECT -38.925 -123.925 -38.595 -123.595 ;
        RECT -38.925 -125.285 -38.595 -124.955 ;
        RECT -38.925 -126.645 -38.595 -126.315 ;
        RECT -38.925 -128.005 -38.595 -127.675 ;
        RECT -38.925 -129.365 -38.595 -129.035 ;
        RECT -38.925 -130.725 -38.595 -130.395 ;
        RECT -38.925 -133.445 -38.595 -133.115 ;
        RECT -38.925 -134.805 -38.595 -134.475 ;
        RECT -38.925 -136.165 -38.595 -135.835 ;
        RECT -38.925 -137.525 -38.595 -137.195 ;
        RECT -38.925 -138.885 -38.595 -138.555 ;
        RECT -38.925 -140.245 -38.595 -139.915 ;
        RECT -38.925 -141.605 -38.595 -141.275 ;
        RECT -38.925 -142.965 -38.595 -142.635 ;
        RECT -38.925 -144.325 -38.595 -143.995 ;
        RECT -38.925 -145.685 -38.595 -145.355 ;
        RECT -38.925 -147.045 -38.595 -146.715 ;
        RECT -38.925 -148.405 -38.595 -148.075 ;
        RECT -38.925 -149.765 -38.595 -149.435 ;
        RECT -38.925 -152.485 -38.595 -152.155 ;
        RECT -38.925 -153.845 -38.595 -153.515 ;
        RECT -38.925 -156.565 -38.595 -156.235 ;
        RECT -38.925 -157.925 -38.595 -157.595 ;
        RECT -38.925 -159.285 -38.595 -158.955 ;
        RECT -38.925 -160.645 -38.595 -160.315 ;
        RECT -38.925 -162.005 -38.595 -161.675 ;
        RECT -38.925 -163.365 -38.595 -163.035 ;
        RECT -38.925 -164.725 -38.595 -164.395 ;
        RECT -38.925 -166.085 -38.595 -165.755 ;
        RECT -38.925 -167.445 -38.595 -167.115 ;
        RECT -38.92 -167.445 -38.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -38.925 -174.245 -38.595 -173.915 ;
        RECT -38.925 -175.605 -38.595 -175.275 ;
        RECT -38.925 -176.685 -38.595 -176.355 ;
        RECT -38.925 -178.325 -38.595 -177.995 ;
        RECT -38.925 -179.685 -38.595 -179.355 ;
        RECT -38.925 -181.93 -38.595 -180.8 ;
        RECT -38.92 -182.045 -38.6 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -37.565 241.32 -37.235 242.45 ;
        RECT -37.565 239.195 -37.235 239.525 ;
        RECT -37.565 237.835 -37.235 238.165 ;
        RECT -37.565 236.475 -37.235 236.805 ;
        RECT -37.565 235.115 -37.235 235.445 ;
        RECT -37.565 233.755 -37.235 234.085 ;
        RECT -37.565 232.395 -37.235 232.725 ;
        RECT -37.565 231.035 -37.235 231.365 ;
        RECT -37.565 229.675 -37.235 230.005 ;
        RECT -37.565 228.315 -37.235 228.645 ;
        RECT -37.565 226.955 -37.235 227.285 ;
        RECT -37.565 225.595 -37.235 225.925 ;
        RECT -37.565 224.235 -37.235 224.565 ;
        RECT -37.565 222.875 -37.235 223.205 ;
        RECT -37.565 221.515 -37.235 221.845 ;
        RECT -37.565 220.155 -37.235 220.485 ;
        RECT -37.565 218.795 -37.235 219.125 ;
        RECT -37.565 217.435 -37.235 217.765 ;
        RECT -37.565 216.075 -37.235 216.405 ;
        RECT -37.565 214.715 -37.235 215.045 ;
        RECT -37.565 213.355 -37.235 213.685 ;
        RECT -37.565 211.995 -37.235 212.325 ;
        RECT -37.565 210.635 -37.235 210.965 ;
        RECT -37.565 209.275 -37.235 209.605 ;
        RECT -37.565 207.915 -37.235 208.245 ;
        RECT -37.565 206.555 -37.235 206.885 ;
        RECT -37.565 205.195 -37.235 205.525 ;
        RECT -37.565 203.835 -37.235 204.165 ;
        RECT -37.565 202.475 -37.235 202.805 ;
        RECT -37.565 201.115 -37.235 201.445 ;
        RECT -37.565 199.755 -37.235 200.085 ;
        RECT -37.565 198.395 -37.235 198.725 ;
        RECT -37.565 197.035 -37.235 197.365 ;
        RECT -37.565 195.675 -37.235 196.005 ;
        RECT -37.565 194.315 -37.235 194.645 ;
        RECT -37.565 192.955 -37.235 193.285 ;
        RECT -37.565 191.595 -37.235 191.925 ;
        RECT -37.565 190.235 -37.235 190.565 ;
        RECT -37.565 188.875 -37.235 189.205 ;
        RECT -37.565 187.515 -37.235 187.845 ;
        RECT -37.565 186.155 -37.235 186.485 ;
        RECT -37.565 184.795 -37.235 185.125 ;
        RECT -37.565 183.435 -37.235 183.765 ;
        RECT -37.565 182.075 -37.235 182.405 ;
        RECT -37.565 180.715 -37.235 181.045 ;
        RECT -37.565 179.355 -37.235 179.685 ;
        RECT -37.565 177.995 -37.235 178.325 ;
        RECT -37.565 176.635 -37.235 176.965 ;
        RECT -37.565 175.275 -37.235 175.605 ;
        RECT -37.565 173.915 -37.235 174.245 ;
        RECT -37.565 172.555 -37.235 172.885 ;
        RECT -37.565 171.195 -37.235 171.525 ;
        RECT -37.565 169.835 -37.235 170.165 ;
        RECT -37.565 168.475 -37.235 168.805 ;
        RECT -37.565 167.115 -37.235 167.445 ;
        RECT -37.565 165.755 -37.235 166.085 ;
        RECT -37.565 164.395 -37.235 164.725 ;
        RECT -37.565 163.035 -37.235 163.365 ;
        RECT -37.565 161.675 -37.235 162.005 ;
        RECT -37.565 160.315 -37.235 160.645 ;
        RECT -37.565 158.955 -37.235 159.285 ;
        RECT -37.565 157.595 -37.235 157.925 ;
        RECT -37.565 156.235 -37.235 156.565 ;
        RECT -37.565 154.875 -37.235 155.205 ;
        RECT -37.565 153.515 -37.235 153.845 ;
        RECT -37.565 152.155 -37.235 152.485 ;
        RECT -37.565 150.795 -37.235 151.125 ;
        RECT -37.565 149.435 -37.235 149.765 ;
        RECT -37.565 148.075 -37.235 148.405 ;
        RECT -37.565 146.715 -37.235 147.045 ;
        RECT -37.565 145.355 -37.235 145.685 ;
        RECT -37.565 143.995 -37.235 144.325 ;
        RECT -37.565 142.635 -37.235 142.965 ;
        RECT -37.565 141.275 -37.235 141.605 ;
        RECT -37.565 139.915 -37.235 140.245 ;
        RECT -37.565 138.555 -37.235 138.885 ;
        RECT -37.565 137.195 -37.235 137.525 ;
        RECT -37.565 135.835 -37.235 136.165 ;
        RECT -37.565 134.475 -37.235 134.805 ;
        RECT -37.565 133.115 -37.235 133.445 ;
        RECT -37.565 131.755 -37.235 132.085 ;
        RECT -37.565 130.395 -37.235 130.725 ;
        RECT -37.565 129.035 -37.235 129.365 ;
        RECT -37.565 127.675 -37.235 128.005 ;
        RECT -37.565 126.315 -37.235 126.645 ;
        RECT -37.565 124.955 -37.235 125.285 ;
        RECT -37.565 123.595 -37.235 123.925 ;
        RECT -37.565 122.235 -37.235 122.565 ;
        RECT -37.565 120.875 -37.235 121.205 ;
        RECT -37.565 119.515 -37.235 119.845 ;
        RECT -37.565 118.155 -37.235 118.485 ;
        RECT -37.565 116.795 -37.235 117.125 ;
        RECT -37.565 115.435 -37.235 115.765 ;
        RECT -37.565 114.075 -37.235 114.405 ;
        RECT -37.565 112.715 -37.235 113.045 ;
        RECT -37.565 111.355 -37.235 111.685 ;
        RECT -37.565 109.995 -37.235 110.325 ;
        RECT -37.565 108.635 -37.235 108.965 ;
        RECT -37.565 107.275 -37.235 107.605 ;
        RECT -37.565 105.915 -37.235 106.245 ;
        RECT -37.565 104.555 -37.235 104.885 ;
        RECT -37.565 103.195 -37.235 103.525 ;
        RECT -37.565 101.835 -37.235 102.165 ;
        RECT -37.565 100.475 -37.235 100.805 ;
        RECT -37.565 99.115 -37.235 99.445 ;
        RECT -37.565 97.755 -37.235 98.085 ;
        RECT -37.565 96.395 -37.235 96.725 ;
        RECT -37.565 95.035 -37.235 95.365 ;
        RECT -37.565 93.675 -37.235 94.005 ;
        RECT -37.565 92.315 -37.235 92.645 ;
        RECT -37.565 90.955 -37.235 91.285 ;
        RECT -37.565 89.595 -37.235 89.925 ;
        RECT -37.565 88.235 -37.235 88.565 ;
        RECT -37.565 86.875 -37.235 87.205 ;
        RECT -37.565 85.515 -37.235 85.845 ;
        RECT -37.565 84.155 -37.235 84.485 ;
        RECT -37.565 82.795 -37.235 83.125 ;
        RECT -37.565 81.435 -37.235 81.765 ;
        RECT -37.565 80.075 -37.235 80.405 ;
        RECT -37.565 78.715 -37.235 79.045 ;
        RECT -37.565 77.355 -37.235 77.685 ;
        RECT -37.565 75.995 -37.235 76.325 ;
        RECT -37.565 74.635 -37.235 74.965 ;
        RECT -37.565 73.275 -37.235 73.605 ;
        RECT -37.565 71.915 -37.235 72.245 ;
        RECT -37.565 70.555 -37.235 70.885 ;
        RECT -37.565 69.195 -37.235 69.525 ;
        RECT -37.565 67.835 -37.235 68.165 ;
        RECT -37.565 66.475 -37.235 66.805 ;
        RECT -37.565 65.115 -37.235 65.445 ;
        RECT -37.565 63.755 -37.235 64.085 ;
        RECT -37.565 62.395 -37.235 62.725 ;
        RECT -37.565 61.035 -37.235 61.365 ;
        RECT -37.565 59.675 -37.235 60.005 ;
        RECT -37.565 58.315 -37.235 58.645 ;
        RECT -37.565 56.955 -37.235 57.285 ;
        RECT -37.565 55.595 -37.235 55.925 ;
        RECT -37.565 54.235 -37.235 54.565 ;
        RECT -37.565 52.875 -37.235 53.205 ;
        RECT -37.565 51.515 -37.235 51.845 ;
        RECT -37.565 50.155 -37.235 50.485 ;
        RECT -37.565 48.795 -37.235 49.125 ;
        RECT -37.565 47.435 -37.235 47.765 ;
        RECT -37.565 46.075 -37.235 46.405 ;
        RECT -37.565 44.715 -37.235 45.045 ;
        RECT -37.565 43.355 -37.235 43.685 ;
        RECT -37.565 41.995 -37.235 42.325 ;
        RECT -37.565 40.635 -37.235 40.965 ;
        RECT -37.565 39.275 -37.235 39.605 ;
        RECT -37.565 37.915 -37.235 38.245 ;
        RECT -37.565 36.555 -37.235 36.885 ;
        RECT -37.565 35.195 -37.235 35.525 ;
        RECT -37.565 33.835 -37.235 34.165 ;
        RECT -37.565 32.475 -37.235 32.805 ;
        RECT -37.565 31.115 -37.235 31.445 ;
        RECT -37.565 29.755 -37.235 30.085 ;
        RECT -37.565 28.395 -37.235 28.725 ;
        RECT -37.565 27.035 -37.235 27.365 ;
        RECT -37.565 25.675 -37.235 26.005 ;
        RECT -37.565 24.315 -37.235 24.645 ;
        RECT -37.565 22.955 -37.235 23.285 ;
        RECT -37.565 21.595 -37.235 21.925 ;
        RECT -37.565 20.235 -37.235 20.565 ;
        RECT -37.565 18.875 -37.235 19.205 ;
        RECT -37.565 17.515 -37.235 17.845 ;
        RECT -37.565 16.155 -37.235 16.485 ;
        RECT -37.565 14.795 -37.235 15.125 ;
        RECT -37.565 13.435 -37.235 13.765 ;
        RECT -37.565 12.075 -37.235 12.405 ;
        RECT -37.565 10.715 -37.235 11.045 ;
        RECT -37.565 9.355 -37.235 9.685 ;
        RECT -37.565 7.995 -37.235 8.325 ;
        RECT -37.565 6.635 -37.235 6.965 ;
        RECT -37.565 5.275 -37.235 5.605 ;
        RECT -37.565 3.915 -37.235 4.245 ;
        RECT -37.565 2.555 -37.235 2.885 ;
        RECT -37.565 1.195 -37.235 1.525 ;
        RECT -37.565 -0.165 -37.235 0.165 ;
        RECT -37.565 -2.885 -37.235 -2.555 ;
        RECT -37.565 -11.045 -37.235 -10.715 ;
        RECT -37.565 -15.125 -37.235 -14.795 ;
        RECT -37.565 -16.485 -37.235 -16.155 ;
        RECT -37.565 -17.845 -37.235 -17.515 ;
        RECT -37.565 -19.205 -37.235 -18.875 ;
        RECT -37.565 -20.565 -37.235 -20.235 ;
        RECT -37.565 -21.925 -37.235 -21.595 ;
        RECT -37.565 -23.285 -37.235 -22.955 ;
        RECT -37.565 -24.645 -37.235 -24.315 ;
        RECT -37.565 -32.805 -37.235 -32.475 ;
        RECT -37.565 -35.525 -37.235 -35.195 ;
        RECT -37.565 -36.885 -37.235 -36.555 ;
        RECT -37.565 -37.93 -37.235 -37.6 ;
        RECT -37.565 -40.965 -37.235 -40.635 ;
        RECT -37.565 -42.77 -37.235 -42.44 ;
        RECT -37.565 -43.685 -37.235 -43.355 ;
        RECT -37.565 -50.485 -37.235 -50.155 ;
        RECT -37.565 -51.845 -37.235 -51.515 ;
        RECT -37.565 -53.205 -37.235 -52.875 ;
        RECT -37.565 -54.565 -37.235 -54.235 ;
        RECT -37.565 -55.925 -37.235 -55.595 ;
        RECT -37.565 -57.285 -37.235 -56.955 ;
        RECT -37.565 -58.645 -37.235 -58.315 ;
        RECT -37.565 -60.005 -37.235 -59.675 ;
        RECT -37.565 -61.365 -37.235 -61.035 ;
        RECT -37.565 -62.725 -37.235 -62.395 ;
        RECT -37.565 -64.085 -37.235 -63.755 ;
        RECT -37.565 -65.445 -37.235 -65.115 ;
        RECT -37.565 -69.525 -37.235 -69.195 ;
        RECT -37.565 -70.885 -37.235 -70.555 ;
        RECT -37.565 -72.245 -37.235 -71.915 ;
        RECT -37.565 -73.605 -37.235 -73.275 ;
        RECT -37.565 -74.965 -37.235 -74.635 ;
        RECT -37.565 -76.325 -37.235 -75.995 ;
        RECT -37.565 -77.685 -37.235 -77.355 ;
        RECT -37.565 -79.045 -37.235 -78.715 ;
        RECT -37.565 -80.405 -37.235 -80.075 ;
        RECT -37.565 -81.765 -37.235 -81.435 ;
        RECT -37.565 -83.125 -37.235 -82.795 ;
        RECT -37.565 -84.485 -37.235 -84.155 ;
        RECT -37.565 -85.845 -37.235 -85.515 ;
        RECT -37.565 -87.205 -37.235 -86.875 ;
        RECT -37.565 -88.565 -37.235 -88.235 ;
        RECT -37.565 -89.925 -37.235 -89.595 ;
        RECT -37.565 -92.645 -37.235 -92.315 ;
        RECT -37.565 -94.005 -37.235 -93.675 ;
        RECT -37.565 -95.365 -37.235 -95.035 ;
        RECT -37.565 -96.725 -37.235 -96.395 ;
        RECT -37.565 -98.085 -37.235 -97.755 ;
        RECT -37.565 -99.69 -37.235 -99.36 ;
        RECT -37.565 -100.805 -37.235 -100.475 ;
        RECT -37.565 -103.525 -37.235 -103.195 ;
        RECT -37.565 -104.885 -37.235 -104.555 ;
        RECT -37.565 -106.245 -37.235 -105.915 ;
        RECT -37.565 -107.83 -37.235 -107.5 ;
        RECT -37.565 -108.965 -37.235 -108.635 ;
        RECT -37.565 -110.325 -37.235 -109.995 ;
        RECT -37.565 -111.685 -37.235 -111.355 ;
        RECT -37.565 -115.765 -37.235 -115.435 ;
        RECT -37.565 -117.125 -37.235 -116.795 ;
        RECT -37.565 -118.485 -37.235 -118.155 ;
        RECT -37.565 -121.205 -37.235 -120.875 ;
        RECT -37.565 -123.925 -37.235 -123.595 ;
        RECT -37.565 -125.285 -37.235 -124.955 ;
        RECT -37.565 -126.645 -37.235 -126.315 ;
        RECT -37.565 -128.005 -37.235 -127.675 ;
        RECT -37.565 -129.365 -37.235 -129.035 ;
        RECT -37.565 -130.725 -37.235 -130.395 ;
        RECT -37.565 -133.445 -37.235 -133.115 ;
        RECT -37.565 -134.805 -37.235 -134.475 ;
        RECT -37.565 -136.165 -37.235 -135.835 ;
        RECT -37.565 -137.525 -37.235 -137.195 ;
        RECT -37.565 -138.885 -37.235 -138.555 ;
        RECT -37.565 -140.245 -37.235 -139.915 ;
        RECT -37.565 -141.605 -37.235 -141.275 ;
        RECT -37.565 -142.965 -37.235 -142.635 ;
        RECT -37.565 -144.325 -37.235 -143.995 ;
        RECT -37.565 -145.685 -37.235 -145.355 ;
        RECT -37.565 -147.045 -37.235 -146.715 ;
        RECT -37.565 -148.405 -37.235 -148.075 ;
        RECT -37.565 -149.765 -37.235 -149.435 ;
        RECT -37.565 -152.485 -37.235 -152.155 ;
        RECT -37.565 -153.845 -37.235 -153.515 ;
        RECT -37.565 -157.925 -37.235 -157.595 ;
        RECT -37.565 -159.285 -37.235 -158.955 ;
        RECT -37.565 -160.645 -37.235 -160.315 ;
        RECT -37.565 -162.005 -37.235 -161.675 ;
        RECT -37.565 -163.365 -37.235 -163.035 ;
        RECT -37.565 -164.725 -37.235 -164.395 ;
        RECT -37.565 -166.085 -37.235 -165.755 ;
        RECT -37.565 -167.445 -37.235 -167.115 ;
        RECT -37.565 -168.805 -37.235 -168.475 ;
        RECT -37.565 -171.525 -37.235 -171.195 ;
        RECT -37.565 -174.245 -37.235 -173.915 ;
        RECT -37.565 -175.605 -37.235 -175.275 ;
        RECT -37.565 -176.685 -37.235 -176.355 ;
        RECT -37.565 -178.325 -37.235 -177.995 ;
        RECT -37.565 -179.685 -37.235 -179.355 ;
        RECT -37.565 -181.93 -37.235 -180.8 ;
        RECT -37.56 -182.045 -37.24 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -36.205 168.475 -35.875 168.805 ;
        RECT -36.205 167.115 -35.875 167.445 ;
        RECT -36.205 165.755 -35.875 166.085 ;
        RECT -36.205 164.395 -35.875 164.725 ;
        RECT -36.205 163.035 -35.875 163.365 ;
        RECT -36.205 161.675 -35.875 162.005 ;
        RECT -36.205 160.315 -35.875 160.645 ;
        RECT -36.205 158.955 -35.875 159.285 ;
        RECT -36.205 157.595 -35.875 157.925 ;
        RECT -36.205 156.235 -35.875 156.565 ;
        RECT -36.205 154.875 -35.875 155.205 ;
        RECT -36.205 153.515 -35.875 153.845 ;
        RECT -36.205 152.155 -35.875 152.485 ;
        RECT -36.205 150.795 -35.875 151.125 ;
        RECT -36.205 149.435 -35.875 149.765 ;
        RECT -36.205 148.075 -35.875 148.405 ;
        RECT -36.205 146.715 -35.875 147.045 ;
        RECT -36.205 145.355 -35.875 145.685 ;
        RECT -36.205 143.995 -35.875 144.325 ;
        RECT -36.205 142.635 -35.875 142.965 ;
        RECT -36.205 141.275 -35.875 141.605 ;
        RECT -36.205 139.915 -35.875 140.245 ;
        RECT -36.205 138.555 -35.875 138.885 ;
        RECT -36.205 137.195 -35.875 137.525 ;
        RECT -36.205 135.835 -35.875 136.165 ;
        RECT -36.205 134.475 -35.875 134.805 ;
        RECT -36.205 133.115 -35.875 133.445 ;
        RECT -36.205 131.755 -35.875 132.085 ;
        RECT -36.205 130.395 -35.875 130.725 ;
        RECT -36.205 129.035 -35.875 129.365 ;
        RECT -36.205 127.675 -35.875 128.005 ;
        RECT -36.205 126.315 -35.875 126.645 ;
        RECT -36.205 124.955 -35.875 125.285 ;
        RECT -36.205 123.595 -35.875 123.925 ;
        RECT -36.205 122.235 -35.875 122.565 ;
        RECT -36.205 120.875 -35.875 121.205 ;
        RECT -36.205 119.515 -35.875 119.845 ;
        RECT -36.205 118.155 -35.875 118.485 ;
        RECT -36.205 116.795 -35.875 117.125 ;
        RECT -36.205 115.435 -35.875 115.765 ;
        RECT -36.205 114.075 -35.875 114.405 ;
        RECT -36.205 112.715 -35.875 113.045 ;
        RECT -36.205 111.355 -35.875 111.685 ;
        RECT -36.205 109.995 -35.875 110.325 ;
        RECT -36.205 108.635 -35.875 108.965 ;
        RECT -36.205 107.275 -35.875 107.605 ;
        RECT -36.205 105.915 -35.875 106.245 ;
        RECT -36.205 104.555 -35.875 104.885 ;
        RECT -36.205 103.195 -35.875 103.525 ;
        RECT -36.205 101.835 -35.875 102.165 ;
        RECT -36.205 100.475 -35.875 100.805 ;
        RECT -36.205 99.115 -35.875 99.445 ;
        RECT -36.205 97.755 -35.875 98.085 ;
        RECT -36.205 96.395 -35.875 96.725 ;
        RECT -36.205 95.035 -35.875 95.365 ;
        RECT -36.205 93.675 -35.875 94.005 ;
        RECT -36.205 92.315 -35.875 92.645 ;
        RECT -36.205 90.955 -35.875 91.285 ;
        RECT -36.205 89.595 -35.875 89.925 ;
        RECT -36.205 88.235 -35.875 88.565 ;
        RECT -36.205 86.875 -35.875 87.205 ;
        RECT -36.205 85.515 -35.875 85.845 ;
        RECT -36.205 84.155 -35.875 84.485 ;
        RECT -36.205 82.795 -35.875 83.125 ;
        RECT -36.205 81.435 -35.875 81.765 ;
        RECT -36.205 80.075 -35.875 80.405 ;
        RECT -36.205 78.715 -35.875 79.045 ;
        RECT -36.205 77.355 -35.875 77.685 ;
        RECT -36.205 75.995 -35.875 76.325 ;
        RECT -36.205 74.635 -35.875 74.965 ;
        RECT -36.205 73.275 -35.875 73.605 ;
        RECT -36.205 71.915 -35.875 72.245 ;
        RECT -36.205 70.555 -35.875 70.885 ;
        RECT -36.205 69.195 -35.875 69.525 ;
        RECT -36.205 67.835 -35.875 68.165 ;
        RECT -36.205 66.475 -35.875 66.805 ;
        RECT -36.205 65.115 -35.875 65.445 ;
        RECT -36.205 63.755 -35.875 64.085 ;
        RECT -36.205 62.395 -35.875 62.725 ;
        RECT -36.205 61.035 -35.875 61.365 ;
        RECT -36.205 59.675 -35.875 60.005 ;
        RECT -36.205 58.315 -35.875 58.645 ;
        RECT -36.205 56.955 -35.875 57.285 ;
        RECT -36.205 55.595 -35.875 55.925 ;
        RECT -36.205 54.235 -35.875 54.565 ;
        RECT -36.205 52.875 -35.875 53.205 ;
        RECT -36.205 51.515 -35.875 51.845 ;
        RECT -36.205 50.155 -35.875 50.485 ;
        RECT -36.205 48.795 -35.875 49.125 ;
        RECT -36.205 47.435 -35.875 47.765 ;
        RECT -36.205 46.075 -35.875 46.405 ;
        RECT -36.205 44.715 -35.875 45.045 ;
        RECT -36.205 43.355 -35.875 43.685 ;
        RECT -36.205 41.995 -35.875 42.325 ;
        RECT -36.205 40.635 -35.875 40.965 ;
        RECT -36.205 39.275 -35.875 39.605 ;
        RECT -36.205 37.915 -35.875 38.245 ;
        RECT -36.205 36.555 -35.875 36.885 ;
        RECT -36.205 35.195 -35.875 35.525 ;
        RECT -36.205 33.835 -35.875 34.165 ;
        RECT -36.205 32.475 -35.875 32.805 ;
        RECT -36.205 31.115 -35.875 31.445 ;
        RECT -36.205 29.755 -35.875 30.085 ;
        RECT -36.205 28.395 -35.875 28.725 ;
        RECT -36.205 27.035 -35.875 27.365 ;
        RECT -36.205 25.675 -35.875 26.005 ;
        RECT -36.205 24.315 -35.875 24.645 ;
        RECT -36.205 22.955 -35.875 23.285 ;
        RECT -36.205 21.595 -35.875 21.925 ;
        RECT -36.205 20.235 -35.875 20.565 ;
        RECT -36.205 18.875 -35.875 19.205 ;
        RECT -36.205 17.515 -35.875 17.845 ;
        RECT -36.205 16.155 -35.875 16.485 ;
        RECT -36.205 14.795 -35.875 15.125 ;
        RECT -36.205 13.435 -35.875 13.765 ;
        RECT -36.205 12.075 -35.875 12.405 ;
        RECT -36.205 10.715 -35.875 11.045 ;
        RECT -36.205 9.355 -35.875 9.685 ;
        RECT -36.205 7.995 -35.875 8.325 ;
        RECT -36.205 6.635 -35.875 6.965 ;
        RECT -36.205 5.275 -35.875 5.605 ;
        RECT -36.205 3.915 -35.875 4.245 ;
        RECT -36.205 2.555 -35.875 2.885 ;
        RECT -36.205 1.195 -35.875 1.525 ;
        RECT -36.205 -0.165 -35.875 0.165 ;
        RECT -36.205 -8.325 -35.875 -7.995 ;
        RECT -36.205 -11.045 -35.875 -10.715 ;
        RECT -36.205 -15.125 -35.875 -14.795 ;
        RECT -36.205 -16.485 -35.875 -16.155 ;
        RECT -36.205 -17.845 -35.875 -17.515 ;
        RECT -36.205 -19.205 -35.875 -18.875 ;
        RECT -36.205 -20.565 -35.875 -20.235 ;
        RECT -36.205 -21.925 -35.875 -21.595 ;
        RECT -36.205 -23.285 -35.875 -22.955 ;
        RECT -36.205 -24.645 -35.875 -24.315 ;
        RECT -36.205 -32.805 -35.875 -32.475 ;
        RECT -36.205 -35.525 -35.875 -35.195 ;
        RECT -36.205 -36.885 -35.875 -36.555 ;
        RECT -36.205 -37.93 -35.875 -37.6 ;
        RECT -36.205 -40.965 -35.875 -40.635 ;
        RECT -36.205 -42.77 -35.875 -42.44 ;
        RECT -36.205 -43.685 -35.875 -43.355 ;
        RECT -36.205 -50.485 -35.875 -50.155 ;
        RECT -36.205 -51.845 -35.875 -51.515 ;
        RECT -36.205 -53.205 -35.875 -52.875 ;
        RECT -36.205 -54.565 -35.875 -54.235 ;
        RECT -36.205 -55.925 -35.875 -55.595 ;
        RECT -36.205 -57.285 -35.875 -56.955 ;
        RECT -36.205 -58.645 -35.875 -58.315 ;
        RECT -36.205 -60.005 -35.875 -59.675 ;
        RECT -36.205 -61.365 -35.875 -61.035 ;
        RECT -36.205 -62.725 -35.875 -62.395 ;
        RECT -36.205 -64.085 -35.875 -63.755 ;
        RECT -36.205 -65.445 -35.875 -65.115 ;
        RECT -36.205 -69.525 -35.875 -69.195 ;
        RECT -36.205 -70.885 -35.875 -70.555 ;
        RECT -36.205 -72.245 -35.875 -71.915 ;
        RECT -36.205 -73.605 -35.875 -73.275 ;
        RECT -36.205 -74.965 -35.875 -74.635 ;
        RECT -36.205 -76.325 -35.875 -75.995 ;
        RECT -36.205 -77.685 -35.875 -77.355 ;
        RECT -36.205 -79.045 -35.875 -78.715 ;
        RECT -36.205 -80.405 -35.875 -80.075 ;
        RECT -36.205 -81.765 -35.875 -81.435 ;
        RECT -36.205 -83.125 -35.875 -82.795 ;
        RECT -36.205 -84.485 -35.875 -84.155 ;
        RECT -36.205 -85.845 -35.875 -85.515 ;
        RECT -36.205 -87.205 -35.875 -86.875 ;
        RECT -36.205 -88.565 -35.875 -88.235 ;
        RECT -36.205 -89.925 -35.875 -89.595 ;
        RECT -36.205 -92.645 -35.875 -92.315 ;
        RECT -36.205 -94.005 -35.875 -93.675 ;
        RECT -36.205 -95.365 -35.875 -95.035 ;
        RECT -36.205 -96.725 -35.875 -96.395 ;
        RECT -36.205 -98.085 -35.875 -97.755 ;
        RECT -36.205 -100.805 -35.875 -100.475 ;
        RECT -36.205 -103.525 -35.875 -103.195 ;
        RECT -36.205 -104.885 -35.875 -104.555 ;
        RECT -36.205 -106.245 -35.875 -105.915 ;
        RECT -36.205 -108.965 -35.875 -108.635 ;
        RECT -36.205 -110.325 -35.875 -109.995 ;
        RECT -36.205 -111.685 -35.875 -111.355 ;
        RECT -36.205 -115.765 -35.875 -115.435 ;
        RECT -36.205 -117.125 -35.875 -116.795 ;
        RECT -36.205 -118.485 -35.875 -118.155 ;
        RECT -36.205 -121.205 -35.875 -120.875 ;
        RECT -36.205 -123.925 -35.875 -123.595 ;
        RECT -36.205 -125.285 -35.875 -124.955 ;
        RECT -36.205 -126.645 -35.875 -126.315 ;
        RECT -36.205 -128.005 -35.875 -127.675 ;
        RECT -36.205 -129.365 -35.875 -129.035 ;
        RECT -36.205 -130.725 -35.875 -130.395 ;
        RECT -36.205 -133.445 -35.875 -133.115 ;
        RECT -36.205 -134.805 -35.875 -134.475 ;
        RECT -36.205 -136.165 -35.875 -135.835 ;
        RECT -36.205 -137.525 -35.875 -137.195 ;
        RECT -36.205 -138.885 -35.875 -138.555 ;
        RECT -36.205 -140.245 -35.875 -139.915 ;
        RECT -36.205 -141.605 -35.875 -141.275 ;
        RECT -36.205 -142.965 -35.875 -142.635 ;
        RECT -36.205 -144.325 -35.875 -143.995 ;
        RECT -36.205 -145.685 -35.875 -145.355 ;
        RECT -36.205 -147.045 -35.875 -146.715 ;
        RECT -36.205 -148.405 -35.875 -148.075 ;
        RECT -36.205 -149.765 -35.875 -149.435 ;
        RECT -36.205 -152.485 -35.875 -152.155 ;
        RECT -36.205 -153.845 -35.875 -153.515 ;
        RECT -36.205 -157.925 -35.875 -157.595 ;
        RECT -36.205 -159.285 -35.875 -158.955 ;
        RECT -36.205 -160.645 -35.875 -160.315 ;
        RECT -36.205 -162.005 -35.875 -161.675 ;
        RECT -36.205 -163.365 -35.875 -163.035 ;
        RECT -36.205 -164.725 -35.875 -164.395 ;
        RECT -36.205 -166.085 -35.875 -165.755 ;
        RECT -36.205 -167.445 -35.875 -167.115 ;
        RECT -36.205 -168.805 -35.875 -168.475 ;
        RECT -36.205 -171.525 -35.875 -171.195 ;
        RECT -36.205 -175.605 -35.875 -175.275 ;
        RECT -36.205 -176.685 -35.875 -176.355 ;
        RECT -36.205 -178.325 -35.875 -177.995 ;
        RECT -36.205 -179.685 -35.875 -179.355 ;
        RECT -36.205 -181.93 -35.875 -180.8 ;
        RECT -36.2 -182.045 -35.88 242.565 ;
        RECT -36.205 241.32 -35.875 242.45 ;
        RECT -36.205 239.195 -35.875 239.525 ;
        RECT -36.205 237.835 -35.875 238.165 ;
        RECT -36.205 236.475 -35.875 236.805 ;
        RECT -36.205 235.115 -35.875 235.445 ;
        RECT -36.205 233.755 -35.875 234.085 ;
        RECT -36.205 232.395 -35.875 232.725 ;
        RECT -36.205 231.035 -35.875 231.365 ;
        RECT -36.205 229.675 -35.875 230.005 ;
        RECT -36.205 228.315 -35.875 228.645 ;
        RECT -36.205 226.955 -35.875 227.285 ;
        RECT -36.205 225.595 -35.875 225.925 ;
        RECT -36.205 224.235 -35.875 224.565 ;
        RECT -36.205 222.875 -35.875 223.205 ;
        RECT -36.205 221.515 -35.875 221.845 ;
        RECT -36.205 220.155 -35.875 220.485 ;
        RECT -36.205 218.795 -35.875 219.125 ;
        RECT -36.205 217.435 -35.875 217.765 ;
        RECT -36.205 216.075 -35.875 216.405 ;
        RECT -36.205 214.715 -35.875 215.045 ;
        RECT -36.205 213.355 -35.875 213.685 ;
        RECT -36.205 211.995 -35.875 212.325 ;
        RECT -36.205 210.635 -35.875 210.965 ;
        RECT -36.205 209.275 -35.875 209.605 ;
        RECT -36.205 207.915 -35.875 208.245 ;
        RECT -36.205 206.555 -35.875 206.885 ;
        RECT -36.205 205.195 -35.875 205.525 ;
        RECT -36.205 203.835 -35.875 204.165 ;
        RECT -36.205 202.475 -35.875 202.805 ;
        RECT -36.205 201.115 -35.875 201.445 ;
        RECT -36.205 199.755 -35.875 200.085 ;
        RECT -36.205 198.395 -35.875 198.725 ;
        RECT -36.205 197.035 -35.875 197.365 ;
        RECT -36.205 195.675 -35.875 196.005 ;
        RECT -36.205 194.315 -35.875 194.645 ;
        RECT -36.205 192.955 -35.875 193.285 ;
        RECT -36.205 191.595 -35.875 191.925 ;
        RECT -36.205 190.235 -35.875 190.565 ;
        RECT -36.205 188.875 -35.875 189.205 ;
        RECT -36.205 187.515 -35.875 187.845 ;
        RECT -36.205 186.155 -35.875 186.485 ;
        RECT -36.205 184.795 -35.875 185.125 ;
        RECT -36.205 183.435 -35.875 183.765 ;
        RECT -36.205 182.075 -35.875 182.405 ;
        RECT -36.205 180.715 -35.875 181.045 ;
        RECT -36.205 179.355 -35.875 179.685 ;
        RECT -36.205 177.995 -35.875 178.325 ;
        RECT -36.205 176.635 -35.875 176.965 ;
        RECT -36.205 175.275 -35.875 175.605 ;
        RECT -36.205 173.915 -35.875 174.245 ;
        RECT -36.205 172.555 -35.875 172.885 ;
        RECT -36.205 171.195 -35.875 171.525 ;
        RECT -36.205 169.835 -35.875 170.165 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.365 241.32 -44.035 242.45 ;
        RECT -44.365 239.195 -44.035 239.525 ;
        RECT -44.365 237.835 -44.035 238.165 ;
        RECT -44.365 236.475 -44.035 236.805 ;
        RECT -44.365 235.115 -44.035 235.445 ;
        RECT -44.365 233.755 -44.035 234.085 ;
        RECT -44.365 232.395 -44.035 232.725 ;
        RECT -44.365 231.035 -44.035 231.365 ;
        RECT -44.365 229.675 -44.035 230.005 ;
        RECT -44.365 228.315 -44.035 228.645 ;
        RECT -44.365 226.955 -44.035 227.285 ;
        RECT -44.365 225.595 -44.035 225.925 ;
        RECT -44.365 224.235 -44.035 224.565 ;
        RECT -44.365 222.875 -44.035 223.205 ;
        RECT -44.365 221.515 -44.035 221.845 ;
        RECT -44.365 220.155 -44.035 220.485 ;
        RECT -44.365 218.795 -44.035 219.125 ;
        RECT -44.365 217.435 -44.035 217.765 ;
        RECT -44.365 216.075 -44.035 216.405 ;
        RECT -44.365 214.715 -44.035 215.045 ;
        RECT -44.365 213.355 -44.035 213.685 ;
        RECT -44.365 211.995 -44.035 212.325 ;
        RECT -44.365 210.635 -44.035 210.965 ;
        RECT -44.365 209.275 -44.035 209.605 ;
        RECT -44.365 207.915 -44.035 208.245 ;
        RECT -44.365 206.555 -44.035 206.885 ;
        RECT -44.365 205.195 -44.035 205.525 ;
        RECT -44.365 203.835 -44.035 204.165 ;
        RECT -44.365 202.475 -44.035 202.805 ;
        RECT -44.365 201.115 -44.035 201.445 ;
        RECT -44.365 199.755 -44.035 200.085 ;
        RECT -44.365 198.395 -44.035 198.725 ;
        RECT -44.365 197.035 -44.035 197.365 ;
        RECT -44.365 195.675 -44.035 196.005 ;
        RECT -44.365 194.315 -44.035 194.645 ;
        RECT -44.365 192.955 -44.035 193.285 ;
        RECT -44.365 191.595 -44.035 191.925 ;
        RECT -44.365 190.235 -44.035 190.565 ;
        RECT -44.365 188.875 -44.035 189.205 ;
        RECT -44.365 187.515 -44.035 187.845 ;
        RECT -44.365 186.155 -44.035 186.485 ;
        RECT -44.365 184.795 -44.035 185.125 ;
        RECT -44.365 183.435 -44.035 183.765 ;
        RECT -44.365 182.075 -44.035 182.405 ;
        RECT -44.365 180.715 -44.035 181.045 ;
        RECT -44.365 179.355 -44.035 179.685 ;
        RECT -44.365 177.995 -44.035 178.325 ;
        RECT -44.365 176.635 -44.035 176.965 ;
        RECT -44.365 175.275 -44.035 175.605 ;
        RECT -44.365 173.915 -44.035 174.245 ;
        RECT -44.365 172.555 -44.035 172.885 ;
        RECT -44.365 171.195 -44.035 171.525 ;
        RECT -44.365 169.835 -44.035 170.165 ;
        RECT -44.365 168.475 -44.035 168.805 ;
        RECT -44.365 167.115 -44.035 167.445 ;
        RECT -44.365 165.755 -44.035 166.085 ;
        RECT -44.365 164.395 -44.035 164.725 ;
        RECT -44.365 163.035 -44.035 163.365 ;
        RECT -44.365 161.675 -44.035 162.005 ;
        RECT -44.365 160.315 -44.035 160.645 ;
        RECT -44.365 158.955 -44.035 159.285 ;
        RECT -44.365 157.595 -44.035 157.925 ;
        RECT -44.365 156.235 -44.035 156.565 ;
        RECT -44.365 154.875 -44.035 155.205 ;
        RECT -44.365 153.515 -44.035 153.845 ;
        RECT -44.365 152.155 -44.035 152.485 ;
        RECT -44.365 150.795 -44.035 151.125 ;
        RECT -44.365 149.435 -44.035 149.765 ;
        RECT -44.365 148.075 -44.035 148.405 ;
        RECT -44.365 146.715 -44.035 147.045 ;
        RECT -44.365 145.355 -44.035 145.685 ;
        RECT -44.365 143.995 -44.035 144.325 ;
        RECT -44.365 142.635 -44.035 142.965 ;
        RECT -44.365 141.275 -44.035 141.605 ;
        RECT -44.365 139.915 -44.035 140.245 ;
        RECT -44.365 138.555 -44.035 138.885 ;
        RECT -44.365 137.195 -44.035 137.525 ;
        RECT -44.365 135.835 -44.035 136.165 ;
        RECT -44.365 134.475 -44.035 134.805 ;
        RECT -44.365 133.115 -44.035 133.445 ;
        RECT -44.365 131.755 -44.035 132.085 ;
        RECT -44.365 130.395 -44.035 130.725 ;
        RECT -44.365 129.035 -44.035 129.365 ;
        RECT -44.365 127.675 -44.035 128.005 ;
        RECT -44.365 126.315 -44.035 126.645 ;
        RECT -44.365 124.955 -44.035 125.285 ;
        RECT -44.365 123.595 -44.035 123.925 ;
        RECT -44.365 122.235 -44.035 122.565 ;
        RECT -44.365 120.875 -44.035 121.205 ;
        RECT -44.365 119.515 -44.035 119.845 ;
        RECT -44.365 118.155 -44.035 118.485 ;
        RECT -44.365 116.795 -44.035 117.125 ;
        RECT -44.365 115.435 -44.035 115.765 ;
        RECT -44.365 114.075 -44.035 114.405 ;
        RECT -44.365 112.715 -44.035 113.045 ;
        RECT -44.365 111.355 -44.035 111.685 ;
        RECT -44.365 109.995 -44.035 110.325 ;
        RECT -44.365 108.635 -44.035 108.965 ;
        RECT -44.365 107.275 -44.035 107.605 ;
        RECT -44.365 105.915 -44.035 106.245 ;
        RECT -44.365 104.555 -44.035 104.885 ;
        RECT -44.365 103.195 -44.035 103.525 ;
        RECT -44.365 101.835 -44.035 102.165 ;
        RECT -44.365 100.475 -44.035 100.805 ;
        RECT -44.365 99.115 -44.035 99.445 ;
        RECT -44.365 97.755 -44.035 98.085 ;
        RECT -44.365 96.395 -44.035 96.725 ;
        RECT -44.365 95.035 -44.035 95.365 ;
        RECT -44.365 93.675 -44.035 94.005 ;
        RECT -44.365 92.315 -44.035 92.645 ;
        RECT -44.365 90.955 -44.035 91.285 ;
        RECT -44.365 89.595 -44.035 89.925 ;
        RECT -44.365 88.235 -44.035 88.565 ;
        RECT -44.365 86.875 -44.035 87.205 ;
        RECT -44.365 85.515 -44.035 85.845 ;
        RECT -44.365 84.155 -44.035 84.485 ;
        RECT -44.365 82.795 -44.035 83.125 ;
        RECT -44.365 81.435 -44.035 81.765 ;
        RECT -44.365 80.075 -44.035 80.405 ;
        RECT -44.365 78.715 -44.035 79.045 ;
        RECT -44.365 77.355 -44.035 77.685 ;
        RECT -44.365 75.995 -44.035 76.325 ;
        RECT -44.365 74.635 -44.035 74.965 ;
        RECT -44.365 73.275 -44.035 73.605 ;
        RECT -44.365 71.915 -44.035 72.245 ;
        RECT -44.365 70.555 -44.035 70.885 ;
        RECT -44.365 69.195 -44.035 69.525 ;
        RECT -44.365 67.835 -44.035 68.165 ;
        RECT -44.365 66.475 -44.035 66.805 ;
        RECT -44.365 65.115 -44.035 65.445 ;
        RECT -44.365 63.755 -44.035 64.085 ;
        RECT -44.365 62.395 -44.035 62.725 ;
        RECT -44.365 61.035 -44.035 61.365 ;
        RECT -44.365 59.675 -44.035 60.005 ;
        RECT -44.365 58.315 -44.035 58.645 ;
        RECT -44.365 56.955 -44.035 57.285 ;
        RECT -44.365 55.595 -44.035 55.925 ;
        RECT -44.365 54.235 -44.035 54.565 ;
        RECT -44.365 52.875 -44.035 53.205 ;
        RECT -44.365 51.515 -44.035 51.845 ;
        RECT -44.365 50.155 -44.035 50.485 ;
        RECT -44.365 48.795 -44.035 49.125 ;
        RECT -44.365 47.435 -44.035 47.765 ;
        RECT -44.365 46.075 -44.035 46.405 ;
        RECT -44.365 44.715 -44.035 45.045 ;
        RECT -44.365 43.355 -44.035 43.685 ;
        RECT -44.365 41.995 -44.035 42.325 ;
        RECT -44.365 40.635 -44.035 40.965 ;
        RECT -44.365 39.275 -44.035 39.605 ;
        RECT -44.365 37.915 -44.035 38.245 ;
        RECT -44.365 36.555 -44.035 36.885 ;
        RECT -44.365 35.195 -44.035 35.525 ;
        RECT -44.365 33.835 -44.035 34.165 ;
        RECT -44.365 32.475 -44.035 32.805 ;
        RECT -44.365 31.115 -44.035 31.445 ;
        RECT -44.365 29.755 -44.035 30.085 ;
        RECT -44.365 28.395 -44.035 28.725 ;
        RECT -44.365 27.035 -44.035 27.365 ;
        RECT -44.365 25.675 -44.035 26.005 ;
        RECT -44.365 24.315 -44.035 24.645 ;
        RECT -44.365 22.955 -44.035 23.285 ;
        RECT -44.365 21.595 -44.035 21.925 ;
        RECT -44.365 20.235 -44.035 20.565 ;
        RECT -44.365 18.875 -44.035 19.205 ;
        RECT -44.365 17.515 -44.035 17.845 ;
        RECT -44.365 16.155 -44.035 16.485 ;
        RECT -44.365 14.795 -44.035 15.125 ;
        RECT -44.365 13.435 -44.035 13.765 ;
        RECT -44.365 12.075 -44.035 12.405 ;
        RECT -44.365 10.715 -44.035 11.045 ;
        RECT -44.365 9.355 -44.035 9.685 ;
        RECT -44.365 7.995 -44.035 8.325 ;
        RECT -44.365 6.635 -44.035 6.965 ;
        RECT -44.365 5.275 -44.035 5.605 ;
        RECT -44.365 3.915 -44.035 4.245 ;
        RECT -44.365 2.555 -44.035 2.885 ;
        RECT -44.365 1.195 -44.035 1.525 ;
        RECT -44.365 -0.165 -44.035 0.165 ;
        RECT -44.365 -4.245 -44.035 -3.915 ;
        RECT -44.365 -5.605 -44.035 -5.275 ;
        RECT -44.365 -6.965 -44.035 -6.635 ;
        RECT -44.365 -11.045 -44.035 -10.715 ;
        RECT -44.365 -15.125 -44.035 -14.795 ;
        RECT -44.365 -16.485 -44.035 -16.155 ;
        RECT -44.365 -17.845 -44.035 -17.515 ;
        RECT -44.365 -19.205 -44.035 -18.875 ;
        RECT -44.365 -20.565 -44.035 -20.235 ;
        RECT -44.365 -21.925 -44.035 -21.595 ;
        RECT -44.365 -23.285 -44.035 -22.955 ;
        RECT -44.365 -24.645 -44.035 -24.315 ;
        RECT -44.365 -32.805 -44.035 -32.475 ;
        RECT -44.365 -35.525 -44.035 -35.195 ;
        RECT -44.365 -36.885 -44.035 -36.555 ;
        RECT -44.365 -37.93 -44.035 -37.6 ;
        RECT -44.365 -40.965 -44.035 -40.635 ;
        RECT -44.365 -42.77 -44.035 -42.44 ;
        RECT -44.365 -43.685 -44.035 -43.355 ;
        RECT -44.365 -50.485 -44.035 -50.155 ;
        RECT -44.365 -51.845 -44.035 -51.515 ;
        RECT -44.365 -54.565 -44.035 -54.235 ;
        RECT -44.365 -55.925 -44.035 -55.595 ;
        RECT -44.365 -60.005 -44.035 -59.675 ;
        RECT -44.365 -62.725 -44.035 -62.395 ;
        RECT -44.36 -64.08 -44.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.365 -69.525 -44.035 -69.195 ;
        RECT -44.365 -70.885 -44.035 -70.555 ;
        RECT -44.365 -72.245 -44.035 -71.915 ;
        RECT -44.365 -73.605 -44.035 -73.275 ;
        RECT -44.365 -74.965 -44.035 -74.635 ;
        RECT -44.365 -76.325 -44.035 -75.995 ;
        RECT -44.365 -77.685 -44.035 -77.355 ;
        RECT -44.365 -79.045 -44.035 -78.715 ;
        RECT -44.365 -80.405 -44.035 -80.075 ;
        RECT -44.365 -81.765 -44.035 -81.435 ;
        RECT -44.365 -83.125 -44.035 -82.795 ;
        RECT -44.365 -84.485 -44.035 -84.155 ;
        RECT -44.365 -85.845 -44.035 -85.515 ;
        RECT -44.365 -87.205 -44.035 -86.875 ;
        RECT -44.365 -88.565 -44.035 -88.235 ;
        RECT -44.365 -89.925 -44.035 -89.595 ;
        RECT -44.365 -92.645 -44.035 -92.315 ;
        RECT -44.365 -94.005 -44.035 -93.675 ;
        RECT -44.365 -95.365 -44.035 -95.035 ;
        RECT -44.365 -96.725 -44.035 -96.395 ;
        RECT -44.365 -98.085 -44.035 -97.755 ;
        RECT -44.365 -99.69 -44.035 -99.36 ;
        RECT -44.365 -100.805 -44.035 -100.475 ;
        RECT -44.365 -103.525 -44.035 -103.195 ;
        RECT -44.365 -104.885 -44.035 -104.555 ;
        RECT -44.365 -106.245 -44.035 -105.915 ;
        RECT -44.365 -107.83 -44.035 -107.5 ;
        RECT -44.365 -108.965 -44.035 -108.635 ;
        RECT -44.365 -110.325 -44.035 -109.995 ;
        RECT -44.365 -111.685 -44.035 -111.355 ;
        RECT -44.36 -113.04 -44.04 -68.52 ;
    END
    PORT
      LAYER met3 ;
        RECT -44.365 -174.245 -44.035 -173.915 ;
        RECT -44.365 -175.605 -44.035 -175.275 ;
        RECT -44.365 -176.685 -44.035 -176.355 ;
        RECT -44.365 -178.325 -44.035 -177.995 ;
        RECT -44.365 -179.685 -44.035 -179.355 ;
        RECT -44.365 -181.93 -44.035 -180.8 ;
        RECT -44.36 -182.045 -44.04 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.005 241.32 -42.675 242.45 ;
        RECT -43.005 239.195 -42.675 239.525 ;
        RECT -43.005 237.835 -42.675 238.165 ;
        RECT -43.005 236.475 -42.675 236.805 ;
        RECT -43.005 235.115 -42.675 235.445 ;
        RECT -43.005 233.755 -42.675 234.085 ;
        RECT -43.005 232.395 -42.675 232.725 ;
        RECT -43.005 231.035 -42.675 231.365 ;
        RECT -43.005 229.675 -42.675 230.005 ;
        RECT -43.005 228.315 -42.675 228.645 ;
        RECT -43.005 226.955 -42.675 227.285 ;
        RECT -43.005 225.595 -42.675 225.925 ;
        RECT -43.005 224.235 -42.675 224.565 ;
        RECT -43.005 222.875 -42.675 223.205 ;
        RECT -43.005 221.515 -42.675 221.845 ;
        RECT -43.005 220.155 -42.675 220.485 ;
        RECT -43.005 218.795 -42.675 219.125 ;
        RECT -43.005 217.435 -42.675 217.765 ;
        RECT -43.005 216.075 -42.675 216.405 ;
        RECT -43.005 214.715 -42.675 215.045 ;
        RECT -43.005 213.355 -42.675 213.685 ;
        RECT -43.005 211.995 -42.675 212.325 ;
        RECT -43.005 210.635 -42.675 210.965 ;
        RECT -43.005 209.275 -42.675 209.605 ;
        RECT -43.005 207.915 -42.675 208.245 ;
        RECT -43.005 206.555 -42.675 206.885 ;
        RECT -43.005 205.195 -42.675 205.525 ;
        RECT -43.005 203.835 -42.675 204.165 ;
        RECT -43.005 202.475 -42.675 202.805 ;
        RECT -43.005 201.115 -42.675 201.445 ;
        RECT -43.005 199.755 -42.675 200.085 ;
        RECT -43.005 198.395 -42.675 198.725 ;
        RECT -43.005 197.035 -42.675 197.365 ;
        RECT -43.005 195.675 -42.675 196.005 ;
        RECT -43.005 194.315 -42.675 194.645 ;
        RECT -43.005 192.955 -42.675 193.285 ;
        RECT -43.005 191.595 -42.675 191.925 ;
        RECT -43.005 190.235 -42.675 190.565 ;
        RECT -43.005 188.875 -42.675 189.205 ;
        RECT -43.005 187.515 -42.675 187.845 ;
        RECT -43.005 186.155 -42.675 186.485 ;
        RECT -43.005 184.795 -42.675 185.125 ;
        RECT -43.005 183.435 -42.675 183.765 ;
        RECT -43.005 182.075 -42.675 182.405 ;
        RECT -43.005 180.715 -42.675 181.045 ;
        RECT -43.005 179.355 -42.675 179.685 ;
        RECT -43.005 177.995 -42.675 178.325 ;
        RECT -43.005 176.635 -42.675 176.965 ;
        RECT -43.005 175.275 -42.675 175.605 ;
        RECT -43.005 173.915 -42.675 174.245 ;
        RECT -43.005 172.555 -42.675 172.885 ;
        RECT -43.005 171.195 -42.675 171.525 ;
        RECT -43.005 169.835 -42.675 170.165 ;
        RECT -43.005 168.475 -42.675 168.805 ;
        RECT -43.005 167.115 -42.675 167.445 ;
        RECT -43.005 165.755 -42.675 166.085 ;
        RECT -43.005 164.395 -42.675 164.725 ;
        RECT -43.005 163.035 -42.675 163.365 ;
        RECT -43.005 161.675 -42.675 162.005 ;
        RECT -43.005 160.315 -42.675 160.645 ;
        RECT -43.005 158.955 -42.675 159.285 ;
        RECT -43.005 157.595 -42.675 157.925 ;
        RECT -43.005 156.235 -42.675 156.565 ;
        RECT -43.005 154.875 -42.675 155.205 ;
        RECT -43.005 153.515 -42.675 153.845 ;
        RECT -43.005 152.155 -42.675 152.485 ;
        RECT -43.005 150.795 -42.675 151.125 ;
        RECT -43.005 149.435 -42.675 149.765 ;
        RECT -43.005 148.075 -42.675 148.405 ;
        RECT -43.005 146.715 -42.675 147.045 ;
        RECT -43.005 145.355 -42.675 145.685 ;
        RECT -43.005 143.995 -42.675 144.325 ;
        RECT -43.005 142.635 -42.675 142.965 ;
        RECT -43.005 141.275 -42.675 141.605 ;
        RECT -43.005 139.915 -42.675 140.245 ;
        RECT -43.005 138.555 -42.675 138.885 ;
        RECT -43.005 137.195 -42.675 137.525 ;
        RECT -43.005 135.835 -42.675 136.165 ;
        RECT -43.005 134.475 -42.675 134.805 ;
        RECT -43.005 133.115 -42.675 133.445 ;
        RECT -43.005 131.755 -42.675 132.085 ;
        RECT -43.005 130.395 -42.675 130.725 ;
        RECT -43.005 129.035 -42.675 129.365 ;
        RECT -43.005 127.675 -42.675 128.005 ;
        RECT -43.005 126.315 -42.675 126.645 ;
        RECT -43.005 124.955 -42.675 125.285 ;
        RECT -43.005 123.595 -42.675 123.925 ;
        RECT -43.005 122.235 -42.675 122.565 ;
        RECT -43.005 120.875 -42.675 121.205 ;
        RECT -43.005 119.515 -42.675 119.845 ;
        RECT -43.005 118.155 -42.675 118.485 ;
        RECT -43.005 116.795 -42.675 117.125 ;
        RECT -43.005 115.435 -42.675 115.765 ;
        RECT -43.005 114.075 -42.675 114.405 ;
        RECT -43.005 112.715 -42.675 113.045 ;
        RECT -43.005 111.355 -42.675 111.685 ;
        RECT -43.005 109.995 -42.675 110.325 ;
        RECT -43.005 108.635 -42.675 108.965 ;
        RECT -43.005 107.275 -42.675 107.605 ;
        RECT -43.005 105.915 -42.675 106.245 ;
        RECT -43.005 104.555 -42.675 104.885 ;
        RECT -43.005 103.195 -42.675 103.525 ;
        RECT -43.005 101.835 -42.675 102.165 ;
        RECT -43.005 100.475 -42.675 100.805 ;
        RECT -43.005 99.115 -42.675 99.445 ;
        RECT -43.005 97.755 -42.675 98.085 ;
        RECT -43.005 96.395 -42.675 96.725 ;
        RECT -43.005 95.035 -42.675 95.365 ;
        RECT -43.005 93.675 -42.675 94.005 ;
        RECT -43.005 92.315 -42.675 92.645 ;
        RECT -43.005 90.955 -42.675 91.285 ;
        RECT -43.005 89.595 -42.675 89.925 ;
        RECT -43.005 88.235 -42.675 88.565 ;
        RECT -43.005 86.875 -42.675 87.205 ;
        RECT -43.005 85.515 -42.675 85.845 ;
        RECT -43.005 84.155 -42.675 84.485 ;
        RECT -43.005 82.795 -42.675 83.125 ;
        RECT -43.005 81.435 -42.675 81.765 ;
        RECT -43.005 80.075 -42.675 80.405 ;
        RECT -43.005 78.715 -42.675 79.045 ;
        RECT -43.005 77.355 -42.675 77.685 ;
        RECT -43.005 75.995 -42.675 76.325 ;
        RECT -43.005 74.635 -42.675 74.965 ;
        RECT -43.005 73.275 -42.675 73.605 ;
        RECT -43.005 71.915 -42.675 72.245 ;
        RECT -43.005 70.555 -42.675 70.885 ;
        RECT -43.005 69.195 -42.675 69.525 ;
        RECT -43.005 67.835 -42.675 68.165 ;
        RECT -43.005 66.475 -42.675 66.805 ;
        RECT -43.005 65.115 -42.675 65.445 ;
        RECT -43.005 63.755 -42.675 64.085 ;
        RECT -43.005 62.395 -42.675 62.725 ;
        RECT -43.005 61.035 -42.675 61.365 ;
        RECT -43.005 59.675 -42.675 60.005 ;
        RECT -43.005 58.315 -42.675 58.645 ;
        RECT -43.005 56.955 -42.675 57.285 ;
        RECT -43.005 55.595 -42.675 55.925 ;
        RECT -43.005 54.235 -42.675 54.565 ;
        RECT -43.005 52.875 -42.675 53.205 ;
        RECT -43.005 51.515 -42.675 51.845 ;
        RECT -43.005 50.155 -42.675 50.485 ;
        RECT -43.005 48.795 -42.675 49.125 ;
        RECT -43.005 47.435 -42.675 47.765 ;
        RECT -43.005 46.075 -42.675 46.405 ;
        RECT -43.005 44.715 -42.675 45.045 ;
        RECT -43.005 43.355 -42.675 43.685 ;
        RECT -43.005 41.995 -42.675 42.325 ;
        RECT -43.005 40.635 -42.675 40.965 ;
        RECT -43.005 39.275 -42.675 39.605 ;
        RECT -43.005 37.915 -42.675 38.245 ;
        RECT -43.005 36.555 -42.675 36.885 ;
        RECT -43.005 35.195 -42.675 35.525 ;
        RECT -43.005 33.835 -42.675 34.165 ;
        RECT -43.005 32.475 -42.675 32.805 ;
        RECT -43.005 31.115 -42.675 31.445 ;
        RECT -43.005 29.755 -42.675 30.085 ;
        RECT -43.005 28.395 -42.675 28.725 ;
        RECT -43.005 27.035 -42.675 27.365 ;
        RECT -43.005 25.675 -42.675 26.005 ;
        RECT -43.005 24.315 -42.675 24.645 ;
        RECT -43.005 22.955 -42.675 23.285 ;
        RECT -43.005 21.595 -42.675 21.925 ;
        RECT -43.005 20.235 -42.675 20.565 ;
        RECT -43.005 18.875 -42.675 19.205 ;
        RECT -43.005 17.515 -42.675 17.845 ;
        RECT -43.005 16.155 -42.675 16.485 ;
        RECT -43.005 14.795 -42.675 15.125 ;
        RECT -43.005 13.435 -42.675 13.765 ;
        RECT -43.005 12.075 -42.675 12.405 ;
        RECT -43.005 10.715 -42.675 11.045 ;
        RECT -43.005 9.355 -42.675 9.685 ;
        RECT -43.005 7.995 -42.675 8.325 ;
        RECT -43.005 6.635 -42.675 6.965 ;
        RECT -43.005 5.275 -42.675 5.605 ;
        RECT -43.005 3.915 -42.675 4.245 ;
        RECT -43.005 2.555 -42.675 2.885 ;
        RECT -43.005 1.195 -42.675 1.525 ;
        RECT -43.005 -0.165 -42.675 0.165 ;
        RECT -43.005 -5.605 -42.675 -5.275 ;
        RECT -43.005 -6.965 -42.675 -6.635 ;
        RECT -43.005 -11.045 -42.675 -10.715 ;
        RECT -43.005 -15.125 -42.675 -14.795 ;
        RECT -43.005 -16.485 -42.675 -16.155 ;
        RECT -43.005 -17.845 -42.675 -17.515 ;
        RECT -43.005 -19.205 -42.675 -18.875 ;
        RECT -43.005 -20.565 -42.675 -20.235 ;
        RECT -43.005 -21.925 -42.675 -21.595 ;
        RECT -43.005 -23.285 -42.675 -22.955 ;
        RECT -43.005 -24.645 -42.675 -24.315 ;
        RECT -43.005 -32.805 -42.675 -32.475 ;
        RECT -43.005 -35.525 -42.675 -35.195 ;
        RECT -43.005 -36.885 -42.675 -36.555 ;
        RECT -43.005 -37.93 -42.675 -37.6 ;
        RECT -43.005 -40.965 -42.675 -40.635 ;
        RECT -43.005 -42.77 -42.675 -42.44 ;
        RECT -43.005 -43.685 -42.675 -43.355 ;
        RECT -43.005 -50.485 -42.675 -50.155 ;
        RECT -43.005 -51.845 -42.675 -51.515 ;
        RECT -43.005 -54.565 -42.675 -54.235 ;
        RECT -43.005 -55.925 -42.675 -55.595 ;
        RECT -43.005 -60.005 -42.675 -59.675 ;
        RECT -43.005 -62.725 -42.675 -62.395 ;
        RECT -43 -63.4 -42.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -43.005 -69.525 -42.675 -69.195 ;
        RECT -43.005 -70.885 -42.675 -70.555 ;
        RECT -43.005 -72.245 -42.675 -71.915 ;
        RECT -43.005 -73.605 -42.675 -73.275 ;
        RECT -43.005 -74.965 -42.675 -74.635 ;
        RECT -43.005 -76.325 -42.675 -75.995 ;
        RECT -43.005 -77.685 -42.675 -77.355 ;
        RECT -43.005 -79.045 -42.675 -78.715 ;
        RECT -43.005 -80.405 -42.675 -80.075 ;
        RECT -43.005 -81.765 -42.675 -81.435 ;
        RECT -43.005 -83.125 -42.675 -82.795 ;
        RECT -43.005 -84.485 -42.675 -84.155 ;
        RECT -43.005 -85.845 -42.675 -85.515 ;
        RECT -43.005 -87.205 -42.675 -86.875 ;
        RECT -43.005 -88.565 -42.675 -88.235 ;
        RECT -43.005 -89.925 -42.675 -89.595 ;
        RECT -43.005 -92.645 -42.675 -92.315 ;
        RECT -43.005 -94.005 -42.675 -93.675 ;
        RECT -43.005 -95.365 -42.675 -95.035 ;
        RECT -43.005 -96.725 -42.675 -96.395 ;
        RECT -43.005 -98.085 -42.675 -97.755 ;
        RECT -43.005 -99.69 -42.675 -99.36 ;
        RECT -43.005 -100.805 -42.675 -100.475 ;
        RECT -43.005 -103.525 -42.675 -103.195 ;
        RECT -43.005 -104.885 -42.675 -104.555 ;
        RECT -43.005 -106.245 -42.675 -105.915 ;
        RECT -43.005 -107.83 -42.675 -107.5 ;
        RECT -43.005 -108.965 -42.675 -108.635 ;
        RECT -43.005 -110.325 -42.675 -109.995 ;
        RECT -43.005 -111.685 -42.675 -111.355 ;
        RECT -43.005 -114.405 -42.675 -114.075 ;
        RECT -43.005 -115.765 -42.675 -115.435 ;
        RECT -43.005 -117.125 -42.675 -116.795 ;
        RECT -43.005 -118.485 -42.675 -118.155 ;
        RECT -43.005 -121.205 -42.675 -120.875 ;
        RECT -43.005 -123.925 -42.675 -123.595 ;
        RECT -43.005 -125.285 -42.675 -124.955 ;
        RECT -43.005 -126.645 -42.675 -126.315 ;
        RECT -43.005 -128.005 -42.675 -127.675 ;
        RECT -43.005 -129.365 -42.675 -129.035 ;
        RECT -43.005 -130.725 -42.675 -130.395 ;
        RECT -43.005 -132.085 -42.675 -131.755 ;
        RECT -43.005 -133.445 -42.675 -133.115 ;
        RECT -43.005 -134.805 -42.675 -134.475 ;
        RECT -43.005 -136.165 -42.675 -135.835 ;
        RECT -43.005 -137.525 -42.675 -137.195 ;
        RECT -43.005 -138.885 -42.675 -138.555 ;
        RECT -43.005 -140.245 -42.675 -139.915 ;
        RECT -43.005 -141.605 -42.675 -141.275 ;
        RECT -43.005 -142.965 -42.675 -142.635 ;
        RECT -43.005 -144.325 -42.675 -143.995 ;
        RECT -43.005 -145.685 -42.675 -145.355 ;
        RECT -43.005 -147.045 -42.675 -146.715 ;
        RECT -43.005 -148.405 -42.675 -148.075 ;
        RECT -43.005 -149.765 -42.675 -149.435 ;
        RECT -43.005 -151.125 -42.675 -150.795 ;
        RECT -43.005 -152.485 -42.675 -152.155 ;
        RECT -43.005 -153.845 -42.675 -153.515 ;
        RECT -43.005 -155.205 -42.675 -154.875 ;
        RECT -43.005 -156.565 -42.675 -156.235 ;
        RECT -43.005 -157.925 -42.675 -157.595 ;
        RECT -43.005 -159.285 -42.675 -158.955 ;
        RECT -43.005 -160.645 -42.675 -160.315 ;
        RECT -43.005 -162.005 -42.675 -161.675 ;
        RECT -43.005 -163.365 -42.675 -163.035 ;
        RECT -43.005 -164.725 -42.675 -164.395 ;
        RECT -43.005 -166.085 -42.675 -165.755 ;
        RECT -43.005 -167.445 -42.675 -167.115 ;
        RECT -43.005 -168.805 -42.675 -168.475 ;
        RECT -43.005 -171.525 -42.675 -171.195 ;
        RECT -43.005 -174.245 -42.675 -173.915 ;
        RECT -43.005 -175.605 -42.675 -175.275 ;
        RECT -43.005 -176.685 -42.675 -176.355 ;
        RECT -43.005 -178.325 -42.675 -177.995 ;
        RECT -43.005 -179.685 -42.675 -179.355 ;
        RECT -43.005 -181.93 -42.675 -180.8 ;
        RECT -43 -182.045 -42.68 -67.16 ;
    END
    PORT
      LAYER met3 ;
        RECT -41.645 241.32 -41.315 242.45 ;
        RECT -41.645 239.195 -41.315 239.525 ;
        RECT -41.645 237.835 -41.315 238.165 ;
        RECT -41.645 236.475 -41.315 236.805 ;
        RECT -41.645 235.115 -41.315 235.445 ;
        RECT -41.645 233.755 -41.315 234.085 ;
        RECT -41.645 232.395 -41.315 232.725 ;
        RECT -41.645 231.035 -41.315 231.365 ;
        RECT -41.645 229.675 -41.315 230.005 ;
        RECT -41.645 228.315 -41.315 228.645 ;
        RECT -41.645 226.955 -41.315 227.285 ;
        RECT -41.645 225.595 -41.315 225.925 ;
        RECT -41.645 224.235 -41.315 224.565 ;
        RECT -41.645 222.875 -41.315 223.205 ;
        RECT -41.645 221.515 -41.315 221.845 ;
        RECT -41.645 220.155 -41.315 220.485 ;
        RECT -41.645 218.795 -41.315 219.125 ;
        RECT -41.645 217.435 -41.315 217.765 ;
        RECT -41.645 216.075 -41.315 216.405 ;
        RECT -41.645 214.715 -41.315 215.045 ;
        RECT -41.645 213.355 -41.315 213.685 ;
        RECT -41.645 211.995 -41.315 212.325 ;
        RECT -41.645 210.635 -41.315 210.965 ;
        RECT -41.645 209.275 -41.315 209.605 ;
        RECT -41.645 207.915 -41.315 208.245 ;
        RECT -41.645 206.555 -41.315 206.885 ;
        RECT -41.645 205.195 -41.315 205.525 ;
        RECT -41.645 203.835 -41.315 204.165 ;
        RECT -41.645 202.475 -41.315 202.805 ;
        RECT -41.645 201.115 -41.315 201.445 ;
        RECT -41.645 199.755 -41.315 200.085 ;
        RECT -41.645 198.395 -41.315 198.725 ;
        RECT -41.645 197.035 -41.315 197.365 ;
        RECT -41.645 195.675 -41.315 196.005 ;
        RECT -41.645 194.315 -41.315 194.645 ;
        RECT -41.645 192.955 -41.315 193.285 ;
        RECT -41.645 191.595 -41.315 191.925 ;
        RECT -41.645 190.235 -41.315 190.565 ;
        RECT -41.645 188.875 -41.315 189.205 ;
        RECT -41.645 187.515 -41.315 187.845 ;
        RECT -41.645 186.155 -41.315 186.485 ;
        RECT -41.645 184.795 -41.315 185.125 ;
        RECT -41.645 183.435 -41.315 183.765 ;
        RECT -41.645 182.075 -41.315 182.405 ;
        RECT -41.645 180.715 -41.315 181.045 ;
        RECT -41.645 179.355 -41.315 179.685 ;
        RECT -41.645 177.995 -41.315 178.325 ;
        RECT -41.645 176.635 -41.315 176.965 ;
        RECT -41.645 175.275 -41.315 175.605 ;
        RECT -41.645 173.915 -41.315 174.245 ;
        RECT -41.645 172.555 -41.315 172.885 ;
        RECT -41.645 171.195 -41.315 171.525 ;
        RECT -41.645 169.835 -41.315 170.165 ;
        RECT -41.645 168.475 -41.315 168.805 ;
        RECT -41.645 167.115 -41.315 167.445 ;
        RECT -41.645 165.755 -41.315 166.085 ;
        RECT -41.645 164.395 -41.315 164.725 ;
        RECT -41.645 163.035 -41.315 163.365 ;
        RECT -41.645 161.675 -41.315 162.005 ;
        RECT -41.645 160.315 -41.315 160.645 ;
        RECT -41.645 158.955 -41.315 159.285 ;
        RECT -41.645 157.595 -41.315 157.925 ;
        RECT -41.645 156.235 -41.315 156.565 ;
        RECT -41.645 154.875 -41.315 155.205 ;
        RECT -41.645 153.515 -41.315 153.845 ;
        RECT -41.645 152.155 -41.315 152.485 ;
        RECT -41.645 150.795 -41.315 151.125 ;
        RECT -41.645 149.435 -41.315 149.765 ;
        RECT -41.645 148.075 -41.315 148.405 ;
        RECT -41.645 146.715 -41.315 147.045 ;
        RECT -41.645 145.355 -41.315 145.685 ;
        RECT -41.645 143.995 -41.315 144.325 ;
        RECT -41.645 142.635 -41.315 142.965 ;
        RECT -41.645 141.275 -41.315 141.605 ;
        RECT -41.645 139.915 -41.315 140.245 ;
        RECT -41.645 138.555 -41.315 138.885 ;
        RECT -41.645 137.195 -41.315 137.525 ;
        RECT -41.645 135.835 -41.315 136.165 ;
        RECT -41.645 134.475 -41.315 134.805 ;
        RECT -41.645 133.115 -41.315 133.445 ;
        RECT -41.645 131.755 -41.315 132.085 ;
        RECT -41.645 130.395 -41.315 130.725 ;
        RECT -41.645 129.035 -41.315 129.365 ;
        RECT -41.645 127.675 -41.315 128.005 ;
        RECT -41.645 126.315 -41.315 126.645 ;
        RECT -41.645 124.955 -41.315 125.285 ;
        RECT -41.645 123.595 -41.315 123.925 ;
        RECT -41.645 122.235 -41.315 122.565 ;
        RECT -41.645 120.875 -41.315 121.205 ;
        RECT -41.645 119.515 -41.315 119.845 ;
        RECT -41.645 118.155 -41.315 118.485 ;
        RECT -41.645 116.795 -41.315 117.125 ;
        RECT -41.645 115.435 -41.315 115.765 ;
        RECT -41.645 114.075 -41.315 114.405 ;
        RECT -41.645 112.715 -41.315 113.045 ;
        RECT -41.645 111.355 -41.315 111.685 ;
        RECT -41.645 109.995 -41.315 110.325 ;
        RECT -41.645 108.635 -41.315 108.965 ;
        RECT -41.645 107.275 -41.315 107.605 ;
        RECT -41.645 105.915 -41.315 106.245 ;
        RECT -41.645 104.555 -41.315 104.885 ;
        RECT -41.645 103.195 -41.315 103.525 ;
        RECT -41.645 101.835 -41.315 102.165 ;
        RECT -41.645 100.475 -41.315 100.805 ;
        RECT -41.645 99.115 -41.315 99.445 ;
        RECT -41.645 97.755 -41.315 98.085 ;
        RECT -41.645 96.395 -41.315 96.725 ;
        RECT -41.645 95.035 -41.315 95.365 ;
        RECT -41.645 93.675 -41.315 94.005 ;
        RECT -41.645 92.315 -41.315 92.645 ;
        RECT -41.645 90.955 -41.315 91.285 ;
        RECT -41.645 89.595 -41.315 89.925 ;
        RECT -41.645 88.235 -41.315 88.565 ;
        RECT -41.645 86.875 -41.315 87.205 ;
        RECT -41.645 85.515 -41.315 85.845 ;
        RECT -41.645 84.155 -41.315 84.485 ;
        RECT -41.645 82.795 -41.315 83.125 ;
        RECT -41.645 81.435 -41.315 81.765 ;
        RECT -41.645 80.075 -41.315 80.405 ;
        RECT -41.645 78.715 -41.315 79.045 ;
        RECT -41.645 77.355 -41.315 77.685 ;
        RECT -41.645 75.995 -41.315 76.325 ;
        RECT -41.645 74.635 -41.315 74.965 ;
        RECT -41.645 73.275 -41.315 73.605 ;
        RECT -41.645 71.915 -41.315 72.245 ;
        RECT -41.645 70.555 -41.315 70.885 ;
        RECT -41.645 69.195 -41.315 69.525 ;
        RECT -41.645 67.835 -41.315 68.165 ;
        RECT -41.645 66.475 -41.315 66.805 ;
        RECT -41.645 65.115 -41.315 65.445 ;
        RECT -41.645 63.755 -41.315 64.085 ;
        RECT -41.645 62.395 -41.315 62.725 ;
        RECT -41.645 61.035 -41.315 61.365 ;
        RECT -41.645 59.675 -41.315 60.005 ;
        RECT -41.645 58.315 -41.315 58.645 ;
        RECT -41.645 56.955 -41.315 57.285 ;
        RECT -41.645 55.595 -41.315 55.925 ;
        RECT -41.645 54.235 -41.315 54.565 ;
        RECT -41.645 52.875 -41.315 53.205 ;
        RECT -41.645 51.515 -41.315 51.845 ;
        RECT -41.645 50.155 -41.315 50.485 ;
        RECT -41.645 48.795 -41.315 49.125 ;
        RECT -41.645 47.435 -41.315 47.765 ;
        RECT -41.645 46.075 -41.315 46.405 ;
        RECT -41.645 44.715 -41.315 45.045 ;
        RECT -41.645 43.355 -41.315 43.685 ;
        RECT -41.645 41.995 -41.315 42.325 ;
        RECT -41.645 40.635 -41.315 40.965 ;
        RECT -41.645 39.275 -41.315 39.605 ;
        RECT -41.645 37.915 -41.315 38.245 ;
        RECT -41.645 36.555 -41.315 36.885 ;
        RECT -41.645 35.195 -41.315 35.525 ;
        RECT -41.645 33.835 -41.315 34.165 ;
        RECT -41.645 32.475 -41.315 32.805 ;
        RECT -41.645 31.115 -41.315 31.445 ;
        RECT -41.645 29.755 -41.315 30.085 ;
        RECT -41.645 28.395 -41.315 28.725 ;
        RECT -41.645 27.035 -41.315 27.365 ;
        RECT -41.645 25.675 -41.315 26.005 ;
        RECT -41.645 24.315 -41.315 24.645 ;
        RECT -41.645 22.955 -41.315 23.285 ;
        RECT -41.645 21.595 -41.315 21.925 ;
        RECT -41.645 20.235 -41.315 20.565 ;
        RECT -41.645 18.875 -41.315 19.205 ;
        RECT -41.645 17.515 -41.315 17.845 ;
        RECT -41.645 16.155 -41.315 16.485 ;
        RECT -41.645 14.795 -41.315 15.125 ;
        RECT -41.645 13.435 -41.315 13.765 ;
        RECT -41.645 12.075 -41.315 12.405 ;
        RECT -41.645 10.715 -41.315 11.045 ;
        RECT -41.645 9.355 -41.315 9.685 ;
        RECT -41.645 7.995 -41.315 8.325 ;
        RECT -41.645 6.635 -41.315 6.965 ;
        RECT -41.645 5.275 -41.315 5.605 ;
        RECT -41.645 3.915 -41.315 4.245 ;
        RECT -41.645 2.555 -41.315 2.885 ;
        RECT -41.645 1.195 -41.315 1.525 ;
        RECT -41.645 -0.165 -41.315 0.165 ;
        RECT -41.645 -5.605 -41.315 -5.275 ;
        RECT -41.645 -6.965 -41.315 -6.635 ;
        RECT -41.645 -11.045 -41.315 -10.715 ;
        RECT -41.645 -15.125 -41.315 -14.795 ;
        RECT -41.645 -16.485 -41.315 -16.155 ;
        RECT -41.645 -17.845 -41.315 -17.515 ;
        RECT -41.645 -19.205 -41.315 -18.875 ;
        RECT -41.645 -20.565 -41.315 -20.235 ;
        RECT -41.645 -21.925 -41.315 -21.595 ;
        RECT -41.645 -23.285 -41.315 -22.955 ;
        RECT -41.645 -24.645 -41.315 -24.315 ;
        RECT -41.645 -32.805 -41.315 -32.475 ;
        RECT -41.645 -35.525 -41.315 -35.195 ;
        RECT -41.645 -36.885 -41.315 -36.555 ;
        RECT -41.645 -37.93 -41.315 -37.6 ;
        RECT -41.645 -40.965 -41.315 -40.635 ;
        RECT -41.645 -42.77 -41.315 -42.44 ;
        RECT -41.645 -43.685 -41.315 -43.355 ;
        RECT -41.645 -50.485 -41.315 -50.155 ;
        RECT -41.645 -51.845 -41.315 -51.515 ;
        RECT -41.645 -54.565 -41.315 -54.235 ;
        RECT -41.645 -55.925 -41.315 -55.595 ;
        RECT -41.645 -60.005 -41.315 -59.675 ;
        RECT -41.645 -62.725 -41.315 -62.395 ;
        RECT -41.645 -66.805 -41.315 -66.475 ;
        RECT -41.645 -69.525 -41.315 -69.195 ;
        RECT -41.645 -70.885 -41.315 -70.555 ;
        RECT -41.645 -72.245 -41.315 -71.915 ;
        RECT -41.645 -73.605 -41.315 -73.275 ;
        RECT -41.645 -74.965 -41.315 -74.635 ;
        RECT -41.645 -76.325 -41.315 -75.995 ;
        RECT -41.645 -77.685 -41.315 -77.355 ;
        RECT -41.645 -79.045 -41.315 -78.715 ;
        RECT -41.645 -80.405 -41.315 -80.075 ;
        RECT -41.645 -81.765 -41.315 -81.435 ;
        RECT -41.645 -83.125 -41.315 -82.795 ;
        RECT -41.645 -84.485 -41.315 -84.155 ;
        RECT -41.645 -85.845 -41.315 -85.515 ;
        RECT -41.645 -87.205 -41.315 -86.875 ;
        RECT -41.645 -88.565 -41.315 -88.235 ;
        RECT -41.645 -89.925 -41.315 -89.595 ;
        RECT -41.645 -92.645 -41.315 -92.315 ;
        RECT -41.645 -94.005 -41.315 -93.675 ;
        RECT -41.645 -95.365 -41.315 -95.035 ;
        RECT -41.645 -96.725 -41.315 -96.395 ;
        RECT -41.645 -98.085 -41.315 -97.755 ;
        RECT -41.645 -99.69 -41.315 -99.36 ;
        RECT -41.645 -100.805 -41.315 -100.475 ;
        RECT -41.645 -103.525 -41.315 -103.195 ;
        RECT -41.645 -104.885 -41.315 -104.555 ;
        RECT -41.645 -106.245 -41.315 -105.915 ;
        RECT -41.645 -107.83 -41.315 -107.5 ;
        RECT -41.645 -108.965 -41.315 -108.635 ;
        RECT -41.645 -110.325 -41.315 -109.995 ;
        RECT -41.645 -111.685 -41.315 -111.355 ;
        RECT -41.645 -114.405 -41.315 -114.075 ;
        RECT -41.645 -115.765 -41.315 -115.435 ;
        RECT -41.645 -117.125 -41.315 -116.795 ;
        RECT -41.645 -118.485 -41.315 -118.155 ;
        RECT -41.645 -121.205 -41.315 -120.875 ;
        RECT -41.645 -123.925 -41.315 -123.595 ;
        RECT -41.645 -125.285 -41.315 -124.955 ;
        RECT -41.645 -126.645 -41.315 -126.315 ;
        RECT -41.645 -128.005 -41.315 -127.675 ;
        RECT -41.645 -129.365 -41.315 -129.035 ;
        RECT -41.645 -130.725 -41.315 -130.395 ;
        RECT -41.645 -132.085 -41.315 -131.755 ;
        RECT -41.645 -133.445 -41.315 -133.115 ;
        RECT -41.645 -134.805 -41.315 -134.475 ;
        RECT -41.645 -136.165 -41.315 -135.835 ;
        RECT -41.645 -137.525 -41.315 -137.195 ;
        RECT -41.645 -138.885 -41.315 -138.555 ;
        RECT -41.645 -140.245 -41.315 -139.915 ;
        RECT -41.645 -141.605 -41.315 -141.275 ;
        RECT -41.645 -142.965 -41.315 -142.635 ;
        RECT -41.645 -144.325 -41.315 -143.995 ;
        RECT -41.645 -145.685 -41.315 -145.355 ;
        RECT -41.645 -147.045 -41.315 -146.715 ;
        RECT -41.645 -148.405 -41.315 -148.075 ;
        RECT -41.645 -149.765 -41.315 -149.435 ;
        RECT -41.645 -151.125 -41.315 -150.795 ;
        RECT -41.645 -152.485 -41.315 -152.155 ;
        RECT -41.645 -153.845 -41.315 -153.515 ;
        RECT -41.645 -155.205 -41.315 -154.875 ;
        RECT -41.645 -156.565 -41.315 -156.235 ;
        RECT -41.645 -157.925 -41.315 -157.595 ;
        RECT -41.645 -159.285 -41.315 -158.955 ;
        RECT -41.645 -160.645 -41.315 -160.315 ;
        RECT -41.645 -162.005 -41.315 -161.675 ;
        RECT -41.645 -163.365 -41.315 -163.035 ;
        RECT -41.645 -164.725 -41.315 -164.395 ;
        RECT -41.645 -166.085 -41.315 -165.755 ;
        RECT -41.645 -167.445 -41.315 -167.115 ;
        RECT -41.645 -168.805 -41.315 -168.475 ;
        RECT -41.645 -171.525 -41.315 -171.195 ;
        RECT -41.645 -175.605 -41.315 -175.275 ;
        RECT -41.645 -176.685 -41.315 -176.355 ;
        RECT -41.645 -178.325 -41.315 -177.995 ;
        RECT -41.645 -179.685 -41.315 -179.355 ;
        RECT -41.645 -181.93 -41.315 -180.8 ;
        RECT -41.64 -182.045 -41.32 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -40.285 -98.085 -39.955 -97.755 ;
        RECT -40.285 -99.69 -39.955 -99.36 ;
        RECT -40.285 -100.805 -39.955 -100.475 ;
        RECT -40.285 -103.525 -39.955 -103.195 ;
        RECT -40.285 -104.885 -39.955 -104.555 ;
        RECT -40.285 -106.245 -39.955 -105.915 ;
        RECT -40.285 -107.83 -39.955 -107.5 ;
        RECT -40.285 -108.965 -39.955 -108.635 ;
        RECT -40.285 -110.325 -39.955 -109.995 ;
        RECT -40.285 -111.685 -39.955 -111.355 ;
        RECT -40.285 -114.405 -39.955 -114.075 ;
        RECT -40.285 -115.765 -39.955 -115.435 ;
        RECT -40.285 -117.125 -39.955 -116.795 ;
        RECT -40.285 -118.485 -39.955 -118.155 ;
        RECT -40.285 -121.205 -39.955 -120.875 ;
        RECT -40.285 -123.925 -39.955 -123.595 ;
        RECT -40.285 -125.285 -39.955 -124.955 ;
        RECT -40.285 -126.645 -39.955 -126.315 ;
        RECT -40.285 -128.005 -39.955 -127.675 ;
        RECT -40.285 -129.365 -39.955 -129.035 ;
        RECT -40.285 -130.725 -39.955 -130.395 ;
        RECT -40.285 -133.445 -39.955 -133.115 ;
        RECT -40.285 -134.805 -39.955 -134.475 ;
        RECT -40.285 -136.165 -39.955 -135.835 ;
        RECT -40.285 -137.525 -39.955 -137.195 ;
        RECT -40.285 -138.885 -39.955 -138.555 ;
        RECT -40.285 -140.245 -39.955 -139.915 ;
        RECT -40.285 -141.605 -39.955 -141.275 ;
        RECT -40.285 -142.965 -39.955 -142.635 ;
        RECT -40.285 -144.325 -39.955 -143.995 ;
        RECT -40.285 -145.685 -39.955 -145.355 ;
        RECT -40.285 -147.045 -39.955 -146.715 ;
        RECT -40.285 -148.405 -39.955 -148.075 ;
        RECT -40.285 -149.765 -39.955 -149.435 ;
        RECT -40.285 -152.485 -39.955 -152.155 ;
        RECT -40.285 -153.845 -39.955 -153.515 ;
        RECT -40.285 -156.565 -39.955 -156.235 ;
        RECT -40.285 -159.285 -39.955 -158.955 ;
        RECT -40.285 -160.645 -39.955 -160.315 ;
        RECT -40.285 -162.005 -39.955 -161.675 ;
        RECT -40.285 -163.365 -39.955 -163.035 ;
        RECT -40.285 -164.725 -39.955 -164.395 ;
        RECT -40.285 -166.085 -39.955 -165.755 ;
        RECT -40.285 -167.445 -39.955 -167.115 ;
        RECT -40.285 -168.805 -39.955 -168.475 ;
        RECT -40.285 -171.525 -39.955 -171.195 ;
        RECT -40.28 -172.88 -39.96 242.565 ;
        RECT -40.285 241.32 -39.955 242.45 ;
        RECT -40.285 239.195 -39.955 239.525 ;
        RECT -40.285 237.835 -39.955 238.165 ;
        RECT -40.285 236.475 -39.955 236.805 ;
        RECT -40.285 235.115 -39.955 235.445 ;
        RECT -40.285 233.755 -39.955 234.085 ;
        RECT -40.285 232.395 -39.955 232.725 ;
        RECT -40.285 231.035 -39.955 231.365 ;
        RECT -40.285 229.675 -39.955 230.005 ;
        RECT -40.285 228.315 -39.955 228.645 ;
        RECT -40.285 226.955 -39.955 227.285 ;
        RECT -40.285 225.595 -39.955 225.925 ;
        RECT -40.285 224.235 -39.955 224.565 ;
        RECT -40.285 222.875 -39.955 223.205 ;
        RECT -40.285 221.515 -39.955 221.845 ;
        RECT -40.285 220.155 -39.955 220.485 ;
        RECT -40.285 218.795 -39.955 219.125 ;
        RECT -40.285 217.435 -39.955 217.765 ;
        RECT -40.285 216.075 -39.955 216.405 ;
        RECT -40.285 214.715 -39.955 215.045 ;
        RECT -40.285 213.355 -39.955 213.685 ;
        RECT -40.285 211.995 -39.955 212.325 ;
        RECT -40.285 210.635 -39.955 210.965 ;
        RECT -40.285 209.275 -39.955 209.605 ;
        RECT -40.285 207.915 -39.955 208.245 ;
        RECT -40.285 206.555 -39.955 206.885 ;
        RECT -40.285 205.195 -39.955 205.525 ;
        RECT -40.285 203.835 -39.955 204.165 ;
        RECT -40.285 202.475 -39.955 202.805 ;
        RECT -40.285 201.115 -39.955 201.445 ;
        RECT -40.285 199.755 -39.955 200.085 ;
        RECT -40.285 198.395 -39.955 198.725 ;
        RECT -40.285 197.035 -39.955 197.365 ;
        RECT -40.285 195.675 -39.955 196.005 ;
        RECT -40.285 194.315 -39.955 194.645 ;
        RECT -40.285 192.955 -39.955 193.285 ;
        RECT -40.285 191.595 -39.955 191.925 ;
        RECT -40.285 190.235 -39.955 190.565 ;
        RECT -40.285 188.875 -39.955 189.205 ;
        RECT -40.285 187.515 -39.955 187.845 ;
        RECT -40.285 186.155 -39.955 186.485 ;
        RECT -40.285 184.795 -39.955 185.125 ;
        RECT -40.285 183.435 -39.955 183.765 ;
        RECT -40.285 182.075 -39.955 182.405 ;
        RECT -40.285 180.715 -39.955 181.045 ;
        RECT -40.285 179.355 -39.955 179.685 ;
        RECT -40.285 177.995 -39.955 178.325 ;
        RECT -40.285 176.635 -39.955 176.965 ;
        RECT -40.285 175.275 -39.955 175.605 ;
        RECT -40.285 173.915 -39.955 174.245 ;
        RECT -40.285 172.555 -39.955 172.885 ;
        RECT -40.285 171.195 -39.955 171.525 ;
        RECT -40.285 169.835 -39.955 170.165 ;
        RECT -40.285 168.475 -39.955 168.805 ;
        RECT -40.285 167.115 -39.955 167.445 ;
        RECT -40.285 165.755 -39.955 166.085 ;
        RECT -40.285 164.395 -39.955 164.725 ;
        RECT -40.285 163.035 -39.955 163.365 ;
        RECT -40.285 161.675 -39.955 162.005 ;
        RECT -40.285 160.315 -39.955 160.645 ;
        RECT -40.285 158.955 -39.955 159.285 ;
        RECT -40.285 157.595 -39.955 157.925 ;
        RECT -40.285 156.235 -39.955 156.565 ;
        RECT -40.285 154.875 -39.955 155.205 ;
        RECT -40.285 153.515 -39.955 153.845 ;
        RECT -40.285 152.155 -39.955 152.485 ;
        RECT -40.285 150.795 -39.955 151.125 ;
        RECT -40.285 149.435 -39.955 149.765 ;
        RECT -40.285 148.075 -39.955 148.405 ;
        RECT -40.285 146.715 -39.955 147.045 ;
        RECT -40.285 145.355 -39.955 145.685 ;
        RECT -40.285 143.995 -39.955 144.325 ;
        RECT -40.285 142.635 -39.955 142.965 ;
        RECT -40.285 141.275 -39.955 141.605 ;
        RECT -40.285 139.915 -39.955 140.245 ;
        RECT -40.285 138.555 -39.955 138.885 ;
        RECT -40.285 137.195 -39.955 137.525 ;
        RECT -40.285 135.835 -39.955 136.165 ;
        RECT -40.285 134.475 -39.955 134.805 ;
        RECT -40.285 133.115 -39.955 133.445 ;
        RECT -40.285 131.755 -39.955 132.085 ;
        RECT -40.285 130.395 -39.955 130.725 ;
        RECT -40.285 129.035 -39.955 129.365 ;
        RECT -40.285 127.675 -39.955 128.005 ;
        RECT -40.285 126.315 -39.955 126.645 ;
        RECT -40.285 124.955 -39.955 125.285 ;
        RECT -40.285 123.595 -39.955 123.925 ;
        RECT -40.285 122.235 -39.955 122.565 ;
        RECT -40.285 120.875 -39.955 121.205 ;
        RECT -40.285 119.515 -39.955 119.845 ;
        RECT -40.285 118.155 -39.955 118.485 ;
        RECT -40.285 116.795 -39.955 117.125 ;
        RECT -40.285 115.435 -39.955 115.765 ;
        RECT -40.285 114.075 -39.955 114.405 ;
        RECT -40.285 112.715 -39.955 113.045 ;
        RECT -40.285 111.355 -39.955 111.685 ;
        RECT -40.285 109.995 -39.955 110.325 ;
        RECT -40.285 108.635 -39.955 108.965 ;
        RECT -40.285 107.275 -39.955 107.605 ;
        RECT -40.285 105.915 -39.955 106.245 ;
        RECT -40.285 104.555 -39.955 104.885 ;
        RECT -40.285 103.195 -39.955 103.525 ;
        RECT -40.285 101.835 -39.955 102.165 ;
        RECT -40.285 100.475 -39.955 100.805 ;
        RECT -40.285 99.115 -39.955 99.445 ;
        RECT -40.285 97.755 -39.955 98.085 ;
        RECT -40.285 96.395 -39.955 96.725 ;
        RECT -40.285 95.035 -39.955 95.365 ;
        RECT -40.285 93.675 -39.955 94.005 ;
        RECT -40.285 92.315 -39.955 92.645 ;
        RECT -40.285 90.955 -39.955 91.285 ;
        RECT -40.285 89.595 -39.955 89.925 ;
        RECT -40.285 88.235 -39.955 88.565 ;
        RECT -40.285 86.875 -39.955 87.205 ;
        RECT -40.285 85.515 -39.955 85.845 ;
        RECT -40.285 84.155 -39.955 84.485 ;
        RECT -40.285 82.795 -39.955 83.125 ;
        RECT -40.285 81.435 -39.955 81.765 ;
        RECT -40.285 80.075 -39.955 80.405 ;
        RECT -40.285 78.715 -39.955 79.045 ;
        RECT -40.285 77.355 -39.955 77.685 ;
        RECT -40.285 75.995 -39.955 76.325 ;
        RECT -40.285 74.635 -39.955 74.965 ;
        RECT -40.285 73.275 -39.955 73.605 ;
        RECT -40.285 71.915 -39.955 72.245 ;
        RECT -40.285 70.555 -39.955 70.885 ;
        RECT -40.285 69.195 -39.955 69.525 ;
        RECT -40.285 67.835 -39.955 68.165 ;
        RECT -40.285 66.475 -39.955 66.805 ;
        RECT -40.285 65.115 -39.955 65.445 ;
        RECT -40.285 63.755 -39.955 64.085 ;
        RECT -40.285 62.395 -39.955 62.725 ;
        RECT -40.285 61.035 -39.955 61.365 ;
        RECT -40.285 59.675 -39.955 60.005 ;
        RECT -40.285 58.315 -39.955 58.645 ;
        RECT -40.285 56.955 -39.955 57.285 ;
        RECT -40.285 55.595 -39.955 55.925 ;
        RECT -40.285 54.235 -39.955 54.565 ;
        RECT -40.285 52.875 -39.955 53.205 ;
        RECT -40.285 51.515 -39.955 51.845 ;
        RECT -40.285 50.155 -39.955 50.485 ;
        RECT -40.285 48.795 -39.955 49.125 ;
        RECT -40.285 47.435 -39.955 47.765 ;
        RECT -40.285 46.075 -39.955 46.405 ;
        RECT -40.285 44.715 -39.955 45.045 ;
        RECT -40.285 43.355 -39.955 43.685 ;
        RECT -40.285 41.995 -39.955 42.325 ;
        RECT -40.285 40.635 -39.955 40.965 ;
        RECT -40.285 39.275 -39.955 39.605 ;
        RECT -40.285 37.915 -39.955 38.245 ;
        RECT -40.285 36.555 -39.955 36.885 ;
        RECT -40.285 35.195 -39.955 35.525 ;
        RECT -40.285 33.835 -39.955 34.165 ;
        RECT -40.285 32.475 -39.955 32.805 ;
        RECT -40.285 31.115 -39.955 31.445 ;
        RECT -40.285 29.755 -39.955 30.085 ;
        RECT -40.285 28.395 -39.955 28.725 ;
        RECT -40.285 27.035 -39.955 27.365 ;
        RECT -40.285 25.675 -39.955 26.005 ;
        RECT -40.285 24.315 -39.955 24.645 ;
        RECT -40.285 22.955 -39.955 23.285 ;
        RECT -40.285 21.595 -39.955 21.925 ;
        RECT -40.285 20.235 -39.955 20.565 ;
        RECT -40.285 18.875 -39.955 19.205 ;
        RECT -40.285 17.515 -39.955 17.845 ;
        RECT -40.285 16.155 -39.955 16.485 ;
        RECT -40.285 14.795 -39.955 15.125 ;
        RECT -40.285 13.435 -39.955 13.765 ;
        RECT -40.285 12.075 -39.955 12.405 ;
        RECT -40.285 10.715 -39.955 11.045 ;
        RECT -40.285 9.355 -39.955 9.685 ;
        RECT -40.285 7.995 -39.955 8.325 ;
        RECT -40.285 6.635 -39.955 6.965 ;
        RECT -40.285 5.275 -39.955 5.605 ;
        RECT -40.285 3.915 -39.955 4.245 ;
        RECT -40.285 2.555 -39.955 2.885 ;
        RECT -40.285 1.195 -39.955 1.525 ;
        RECT -40.285 -0.165 -39.955 0.165 ;
        RECT -40.285 -2.885 -39.955 -2.555 ;
        RECT -40.285 -4.245 -39.955 -3.915 ;
        RECT -40.285 -5.605 -39.955 -5.275 ;
        RECT -40.285 -11.045 -39.955 -10.715 ;
        RECT -40.285 -15.125 -39.955 -14.795 ;
        RECT -40.285 -16.485 -39.955 -16.155 ;
        RECT -40.285 -17.845 -39.955 -17.515 ;
        RECT -40.285 -19.205 -39.955 -18.875 ;
        RECT -40.285 -20.565 -39.955 -20.235 ;
        RECT -40.285 -21.925 -39.955 -21.595 ;
        RECT -40.285 -23.285 -39.955 -22.955 ;
        RECT -40.285 -24.645 -39.955 -24.315 ;
        RECT -40.285 -32.805 -39.955 -32.475 ;
        RECT -40.285 -35.525 -39.955 -35.195 ;
        RECT -40.285 -36.885 -39.955 -36.555 ;
        RECT -40.285 -37.93 -39.955 -37.6 ;
        RECT -40.285 -40.965 -39.955 -40.635 ;
        RECT -40.285 -42.77 -39.955 -42.44 ;
        RECT -40.285 -43.685 -39.955 -43.355 ;
        RECT -40.285 -50.485 -39.955 -50.155 ;
        RECT -40.285 -51.845 -39.955 -51.515 ;
        RECT -40.285 -54.565 -39.955 -54.235 ;
        RECT -40.285 -55.925 -39.955 -55.595 ;
        RECT -40.285 -60.005 -39.955 -59.675 ;
        RECT -40.285 -62.725 -39.955 -62.395 ;
        RECT -40.285 -66.805 -39.955 -66.475 ;
        RECT -40.285 -69.525 -39.955 -69.195 ;
        RECT -40.285 -70.885 -39.955 -70.555 ;
        RECT -40.285 -72.245 -39.955 -71.915 ;
        RECT -40.285 -73.605 -39.955 -73.275 ;
        RECT -40.285 -74.965 -39.955 -74.635 ;
        RECT -40.285 -76.325 -39.955 -75.995 ;
        RECT -40.285 -77.685 -39.955 -77.355 ;
        RECT -40.285 -79.045 -39.955 -78.715 ;
        RECT -40.285 -80.405 -39.955 -80.075 ;
        RECT -40.285 -81.765 -39.955 -81.435 ;
        RECT -40.285 -83.125 -39.955 -82.795 ;
        RECT -40.285 -84.485 -39.955 -84.155 ;
        RECT -40.285 -85.845 -39.955 -85.515 ;
        RECT -40.285 -87.205 -39.955 -86.875 ;
        RECT -40.285 -88.565 -39.955 -88.235 ;
        RECT -40.285 -89.925 -39.955 -89.595 ;
        RECT -40.285 -92.645 -39.955 -92.315 ;
        RECT -40.285 -94.005 -39.955 -93.675 ;
        RECT -40.285 -95.365 -39.955 -95.035 ;
        RECT -40.285 -96.725 -39.955 -96.395 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.165 -174.245 -50.835 -173.915 ;
        RECT -51.165 -175.605 -50.835 -175.275 ;
        RECT -51.165 -176.685 -50.835 -176.355 ;
        RECT -51.165 -178.325 -50.835 -177.995 ;
        RECT -51.165 -179.685 -50.835 -179.355 ;
        RECT -51.165 -181.93 -50.835 -180.8 ;
        RECT -51.16 -182.045 -50.84 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -49.805 241.32 -49.475 242.45 ;
        RECT -49.805 239.195 -49.475 239.525 ;
        RECT -49.805 237.835 -49.475 238.165 ;
        RECT -49.805 236.475 -49.475 236.805 ;
        RECT -49.805 235.115 -49.475 235.445 ;
        RECT -49.805 233.755 -49.475 234.085 ;
        RECT -49.805 232.395 -49.475 232.725 ;
        RECT -49.805 231.035 -49.475 231.365 ;
        RECT -49.805 229.675 -49.475 230.005 ;
        RECT -49.805 228.315 -49.475 228.645 ;
        RECT -49.805 226.955 -49.475 227.285 ;
        RECT -49.805 225.595 -49.475 225.925 ;
        RECT -49.805 224.235 -49.475 224.565 ;
        RECT -49.805 222.875 -49.475 223.205 ;
        RECT -49.805 221.515 -49.475 221.845 ;
        RECT -49.805 220.155 -49.475 220.485 ;
        RECT -49.805 218.795 -49.475 219.125 ;
        RECT -49.805 217.435 -49.475 217.765 ;
        RECT -49.805 216.075 -49.475 216.405 ;
        RECT -49.805 214.715 -49.475 215.045 ;
        RECT -49.805 213.355 -49.475 213.685 ;
        RECT -49.805 211.995 -49.475 212.325 ;
        RECT -49.805 210.635 -49.475 210.965 ;
        RECT -49.805 209.275 -49.475 209.605 ;
        RECT -49.805 207.915 -49.475 208.245 ;
        RECT -49.805 206.555 -49.475 206.885 ;
        RECT -49.805 205.195 -49.475 205.525 ;
        RECT -49.805 203.835 -49.475 204.165 ;
        RECT -49.805 202.475 -49.475 202.805 ;
        RECT -49.805 201.115 -49.475 201.445 ;
        RECT -49.805 199.755 -49.475 200.085 ;
        RECT -49.805 198.395 -49.475 198.725 ;
        RECT -49.805 197.035 -49.475 197.365 ;
        RECT -49.805 195.675 -49.475 196.005 ;
        RECT -49.805 194.315 -49.475 194.645 ;
        RECT -49.805 192.955 -49.475 193.285 ;
        RECT -49.805 191.595 -49.475 191.925 ;
        RECT -49.805 190.235 -49.475 190.565 ;
        RECT -49.805 188.875 -49.475 189.205 ;
        RECT -49.805 187.515 -49.475 187.845 ;
        RECT -49.805 186.155 -49.475 186.485 ;
        RECT -49.805 184.795 -49.475 185.125 ;
        RECT -49.805 183.435 -49.475 183.765 ;
        RECT -49.805 182.075 -49.475 182.405 ;
        RECT -49.805 180.715 -49.475 181.045 ;
        RECT -49.805 179.355 -49.475 179.685 ;
        RECT -49.805 177.995 -49.475 178.325 ;
        RECT -49.805 176.635 -49.475 176.965 ;
        RECT -49.805 175.275 -49.475 175.605 ;
        RECT -49.805 173.915 -49.475 174.245 ;
        RECT -49.805 172.555 -49.475 172.885 ;
        RECT -49.805 171.195 -49.475 171.525 ;
        RECT -49.805 169.835 -49.475 170.165 ;
        RECT -49.805 168.475 -49.475 168.805 ;
        RECT -49.805 167.115 -49.475 167.445 ;
        RECT -49.805 165.755 -49.475 166.085 ;
        RECT -49.805 164.395 -49.475 164.725 ;
        RECT -49.805 163.035 -49.475 163.365 ;
        RECT -49.805 161.675 -49.475 162.005 ;
        RECT -49.805 160.315 -49.475 160.645 ;
        RECT -49.805 158.955 -49.475 159.285 ;
        RECT -49.805 157.595 -49.475 157.925 ;
        RECT -49.805 156.235 -49.475 156.565 ;
        RECT -49.805 154.875 -49.475 155.205 ;
        RECT -49.805 153.515 -49.475 153.845 ;
        RECT -49.805 152.155 -49.475 152.485 ;
        RECT -49.805 150.795 -49.475 151.125 ;
        RECT -49.805 149.435 -49.475 149.765 ;
        RECT -49.805 148.075 -49.475 148.405 ;
        RECT -49.805 146.715 -49.475 147.045 ;
        RECT -49.805 145.355 -49.475 145.685 ;
        RECT -49.805 143.995 -49.475 144.325 ;
        RECT -49.805 142.635 -49.475 142.965 ;
        RECT -49.805 141.275 -49.475 141.605 ;
        RECT -49.805 139.915 -49.475 140.245 ;
        RECT -49.805 138.555 -49.475 138.885 ;
        RECT -49.805 137.225 -49.475 137.555 ;
        RECT -49.805 135.175 -49.475 135.505 ;
        RECT -49.805 132.815 -49.475 133.145 ;
        RECT -49.805 131.665 -49.475 131.995 ;
        RECT -49.805 129.655 -49.475 129.985 ;
        RECT -49.805 128.505 -49.475 128.835 ;
        RECT -49.805 126.495 -49.475 126.825 ;
        RECT -49.805 125.345 -49.475 125.675 ;
        RECT -49.805 123.335 -49.475 123.665 ;
        RECT -49.805 122.185 -49.475 122.515 ;
        RECT -49.805 120.175 -49.475 120.505 ;
        RECT -49.805 119.025 -49.475 119.355 ;
        RECT -49.805 117.185 -49.475 117.515 ;
        RECT -49.805 115.865 -49.475 116.195 ;
        RECT -49.805 113.855 -49.475 114.185 ;
        RECT -49.805 112.705 -49.475 113.035 ;
        RECT -49.805 110.695 -49.475 111.025 ;
        RECT -49.805 109.545 -49.475 109.875 ;
        RECT -49.805 107.535 -49.475 107.865 ;
        RECT -49.805 106.385 -49.475 106.715 ;
        RECT -49.805 104.375 -49.475 104.705 ;
        RECT -49.805 103.225 -49.475 103.555 ;
        RECT -49.805 100.865 -49.475 101.195 ;
        RECT -49.805 98.81 -49.475 99.14 ;
        RECT -49.805 97.755 -49.475 98.085 ;
        RECT -49.805 96.395 -49.475 96.725 ;
        RECT -49.805 95.035 -49.475 95.365 ;
        RECT -49.805 93.675 -49.475 94.005 ;
        RECT -49.805 92.315 -49.475 92.645 ;
        RECT -49.805 90.955 -49.475 91.285 ;
        RECT -49.805 89.595 -49.475 89.925 ;
        RECT -49.805 88.235 -49.475 88.565 ;
        RECT -49.805 86.875 -49.475 87.205 ;
        RECT -49.805 85.515 -49.475 85.845 ;
        RECT -49.805 84.155 -49.475 84.485 ;
        RECT -49.805 82.795 -49.475 83.125 ;
        RECT -49.805 81.435 -49.475 81.765 ;
        RECT -49.805 80.075 -49.475 80.405 ;
        RECT -49.805 78.715 -49.475 79.045 ;
        RECT -49.805 77.355 -49.475 77.685 ;
        RECT -49.805 75.995 -49.475 76.325 ;
        RECT -49.805 74.635 -49.475 74.965 ;
        RECT -49.805 73.275 -49.475 73.605 ;
        RECT -49.805 71.915 -49.475 72.245 ;
        RECT -49.805 70.555 -49.475 70.885 ;
        RECT -49.805 69.195 -49.475 69.525 ;
        RECT -49.805 67.835 -49.475 68.165 ;
        RECT -49.805 66.475 -49.475 66.805 ;
        RECT -49.805 65.115 -49.475 65.445 ;
        RECT -49.805 63.755 -49.475 64.085 ;
        RECT -49.805 62.395 -49.475 62.725 ;
        RECT -49.805 61.035 -49.475 61.365 ;
        RECT -49.805 59.675 -49.475 60.005 ;
        RECT -49.805 58.315 -49.475 58.645 ;
        RECT -49.805 56.955 -49.475 57.285 ;
        RECT -49.805 55.595 -49.475 55.925 ;
        RECT -49.805 54.235 -49.475 54.565 ;
        RECT -49.805 52.875 -49.475 53.205 ;
        RECT -49.805 51.515 -49.475 51.845 ;
        RECT -49.805 50.155 -49.475 50.485 ;
        RECT -49.805 48.795 -49.475 49.125 ;
        RECT -49.805 47.435 -49.475 47.765 ;
        RECT -49.805 46.075 -49.475 46.405 ;
        RECT -49.805 44.715 -49.475 45.045 ;
        RECT -49.805 43.355 -49.475 43.685 ;
        RECT -49.805 41.995 -49.475 42.325 ;
        RECT -49.805 40.635 -49.475 40.965 ;
        RECT -49.805 39.275 -49.475 39.605 ;
        RECT -49.805 37.915 -49.475 38.245 ;
        RECT -49.805 36.555 -49.475 36.885 ;
        RECT -49.805 35.195 -49.475 35.525 ;
        RECT -49.805 33.835 -49.475 34.165 ;
        RECT -49.805 32.475 -49.475 32.805 ;
        RECT -49.805 31.115 -49.475 31.445 ;
        RECT -49.805 29.755 -49.475 30.085 ;
        RECT -49.805 28.395 -49.475 28.725 ;
        RECT -49.805 27.035 -49.475 27.365 ;
        RECT -49.805 25.675 -49.475 26.005 ;
        RECT -49.805 24.315 -49.475 24.645 ;
        RECT -49.805 22.955 -49.475 23.285 ;
        RECT -49.805 21.595 -49.475 21.925 ;
        RECT -49.805 20.235 -49.475 20.565 ;
        RECT -49.805 18.875 -49.475 19.205 ;
        RECT -49.805 17.515 -49.475 17.845 ;
        RECT -49.805 16.155 -49.475 16.485 ;
        RECT -49.805 14.795 -49.475 15.125 ;
        RECT -49.805 13.435 -49.475 13.765 ;
        RECT -49.805 12.075 -49.475 12.405 ;
        RECT -49.805 10.715 -49.475 11.045 ;
        RECT -49.805 9.355 -49.475 9.685 ;
        RECT -49.805 7.995 -49.475 8.325 ;
        RECT -49.805 6.635 -49.475 6.965 ;
        RECT -49.805 5.275 -49.475 5.605 ;
        RECT -49.805 3.915 -49.475 4.245 ;
        RECT -49.805 2.555 -49.475 2.885 ;
        RECT -49.805 1.195 -49.475 1.525 ;
        RECT -49.805 -0.165 -49.475 0.165 ;
        RECT -49.805 -2.885 -49.475 -2.555 ;
        RECT -49.805 -4.245 -49.475 -3.915 ;
        RECT -49.805 -5.605 -49.475 -5.275 ;
        RECT -49.805 -6.965 -49.475 -6.635 ;
        RECT -49.805 -8.325 -49.475 -7.995 ;
        RECT -49.805 -9.685 -49.475 -9.355 ;
        RECT -49.805 -11.045 -49.475 -10.715 ;
        RECT -49.805 -12.405 -49.475 -12.075 ;
        RECT -49.805 -15.125 -49.475 -14.795 ;
        RECT -49.805 -16.485 -49.475 -16.155 ;
        RECT -49.805 -17.845 -49.475 -17.515 ;
        RECT -49.805 -19.205 -49.475 -18.875 ;
        RECT -49.805 -20.565 -49.475 -20.235 ;
        RECT -49.805 -21.925 -49.475 -21.595 ;
        RECT -49.805 -23.285 -49.475 -22.955 ;
        RECT -49.805 -24.645 -49.475 -24.315 ;
        RECT -49.805 -30.085 -49.475 -29.755 ;
        RECT -49.805 -31.445 -49.475 -31.115 ;
        RECT -49.805 -32.805 -49.475 -32.475 ;
        RECT -49.805 -35.525 -49.475 -35.195 ;
        RECT -49.805 -36.885 -49.475 -36.555 ;
        RECT -49.805 -40.965 -49.475 -40.635 ;
        RECT -49.805 -43.685 -49.475 -43.355 ;
        RECT -49.805 -50.485 -49.475 -50.155 ;
        RECT -49.805 -51.845 -49.475 -51.515 ;
        RECT -49.805 -54.565 -49.475 -54.235 ;
        RECT -49.805 -55.925 -49.475 -55.595 ;
        RECT -49.805 -60.005 -49.475 -59.675 ;
        RECT -49.805 -62.725 -49.475 -62.395 ;
        RECT -49.805 -68.165 -49.475 -67.835 ;
        RECT -49.805 -69.525 -49.475 -69.195 ;
        RECT -49.805 -70.885 -49.475 -70.555 ;
        RECT -49.805 -72.245 -49.475 -71.915 ;
        RECT -49.805 -73.605 -49.475 -73.275 ;
        RECT -49.805 -74.965 -49.475 -74.635 ;
        RECT -49.805 -76.325 -49.475 -75.995 ;
        RECT -49.805 -77.685 -49.475 -77.355 ;
        RECT -49.805 -79.045 -49.475 -78.715 ;
        RECT -49.805 -80.405 -49.475 -80.075 ;
        RECT -49.805 -81.765 -49.475 -81.435 ;
        RECT -49.805 -83.125 -49.475 -82.795 ;
        RECT -49.805 -84.485 -49.475 -84.155 ;
        RECT -49.805 -85.845 -49.475 -85.515 ;
        RECT -49.805 -87.205 -49.475 -86.875 ;
        RECT -49.805 -88.565 -49.475 -88.235 ;
        RECT -49.805 -89.925 -49.475 -89.595 ;
        RECT -49.805 -92.645 -49.475 -92.315 ;
        RECT -49.805 -94.005 -49.475 -93.675 ;
        RECT -49.805 -95.365 -49.475 -95.035 ;
        RECT -49.805 -96.725 -49.475 -96.395 ;
        RECT -49.805 -98.085 -49.475 -97.755 ;
        RECT -49.805 -99.69 -49.475 -99.36 ;
        RECT -49.805 -100.805 -49.475 -100.475 ;
        RECT -49.805 -103.525 -49.475 -103.195 ;
        RECT -49.805 -104.885 -49.475 -104.555 ;
        RECT -49.805 -106.245 -49.475 -105.915 ;
        RECT -49.805 -107.83 -49.475 -107.5 ;
        RECT -49.805 -108.965 -49.475 -108.635 ;
        RECT -49.805 -110.325 -49.475 -109.995 ;
        RECT -49.805 -111.685 -49.475 -111.355 ;
        RECT -49.805 -114.405 -49.475 -114.075 ;
        RECT -49.805 -115.765 -49.475 -115.435 ;
        RECT -49.805 -117.125 -49.475 -116.795 ;
        RECT -49.805 -118.485 -49.475 -118.155 ;
        RECT -49.805 -121.205 -49.475 -120.875 ;
        RECT -49.805 -123.925 -49.475 -123.595 ;
        RECT -49.805 -125.285 -49.475 -124.955 ;
        RECT -49.805 -126.645 -49.475 -126.315 ;
        RECT -49.805 -128.005 -49.475 -127.675 ;
        RECT -49.805 -129.365 -49.475 -129.035 ;
        RECT -49.805 -130.725 -49.475 -130.395 ;
        RECT -49.805 -132.085 -49.475 -131.755 ;
        RECT -49.805 -133.445 -49.475 -133.115 ;
        RECT -49.805 -134.805 -49.475 -134.475 ;
        RECT -49.805 -136.165 -49.475 -135.835 ;
        RECT -49.805 -137.525 -49.475 -137.195 ;
        RECT -49.805 -138.885 -49.475 -138.555 ;
        RECT -49.805 -140.245 -49.475 -139.915 ;
        RECT -49.805 -141.605 -49.475 -141.275 ;
        RECT -49.805 -142.965 -49.475 -142.635 ;
        RECT -49.805 -144.325 -49.475 -143.995 ;
        RECT -49.805 -145.685 -49.475 -145.355 ;
        RECT -49.805 -147.045 -49.475 -146.715 ;
        RECT -49.805 -148.405 -49.475 -148.075 ;
        RECT -49.805 -149.765 -49.475 -149.435 ;
        RECT -49.805 -151.125 -49.475 -150.795 ;
        RECT -49.805 -152.485 -49.475 -152.155 ;
        RECT -49.805 -153.845 -49.475 -153.515 ;
        RECT -49.805 -155.205 -49.475 -154.875 ;
        RECT -49.805 -156.565 -49.475 -156.235 ;
        RECT -49.805 -157.925 -49.475 -157.595 ;
        RECT -49.805 -159.285 -49.475 -158.955 ;
        RECT -49.805 -160.645 -49.475 -160.315 ;
        RECT -49.805 -162.005 -49.475 -161.675 ;
        RECT -49.805 -163.365 -49.475 -163.035 ;
        RECT -49.805 -164.725 -49.475 -164.395 ;
        RECT -49.805 -166.085 -49.475 -165.755 ;
        RECT -49.805 -167.445 -49.475 -167.115 ;
        RECT -49.805 -168.805 -49.475 -168.475 ;
        RECT -49.805 -171.525 -49.475 -171.195 ;
        RECT -49.805 -172.885 -49.475 -172.555 ;
        RECT -49.805 -174.245 -49.475 -173.915 ;
        RECT -49.805 -175.605 -49.475 -175.275 ;
        RECT -49.805 -176.685 -49.475 -176.355 ;
        RECT -49.805 -178.325 -49.475 -177.995 ;
        RECT -49.805 -179.685 -49.475 -179.355 ;
        RECT -49.805 -181.93 -49.475 -180.8 ;
        RECT -49.8 -182.045 -49.48 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 241.32 -48.115 242.45 ;
        RECT -48.445 239.195 -48.115 239.525 ;
        RECT -48.445 237.835 -48.115 238.165 ;
        RECT -48.445 236.475 -48.115 236.805 ;
        RECT -48.445 235.115 -48.115 235.445 ;
        RECT -48.445 233.755 -48.115 234.085 ;
        RECT -48.445 232.395 -48.115 232.725 ;
        RECT -48.445 231.035 -48.115 231.365 ;
        RECT -48.445 229.675 -48.115 230.005 ;
        RECT -48.445 228.315 -48.115 228.645 ;
        RECT -48.445 226.955 -48.115 227.285 ;
        RECT -48.445 225.595 -48.115 225.925 ;
        RECT -48.445 224.235 -48.115 224.565 ;
        RECT -48.445 222.875 -48.115 223.205 ;
        RECT -48.445 221.515 -48.115 221.845 ;
        RECT -48.445 220.155 -48.115 220.485 ;
        RECT -48.445 218.795 -48.115 219.125 ;
        RECT -48.445 217.435 -48.115 217.765 ;
        RECT -48.445 216.075 -48.115 216.405 ;
        RECT -48.445 214.715 -48.115 215.045 ;
        RECT -48.445 213.355 -48.115 213.685 ;
        RECT -48.445 211.995 -48.115 212.325 ;
        RECT -48.445 210.635 -48.115 210.965 ;
        RECT -48.445 209.275 -48.115 209.605 ;
        RECT -48.445 207.915 -48.115 208.245 ;
        RECT -48.445 206.555 -48.115 206.885 ;
        RECT -48.445 205.195 -48.115 205.525 ;
        RECT -48.445 203.835 -48.115 204.165 ;
        RECT -48.445 202.475 -48.115 202.805 ;
        RECT -48.445 201.115 -48.115 201.445 ;
        RECT -48.445 199.755 -48.115 200.085 ;
        RECT -48.445 198.395 -48.115 198.725 ;
        RECT -48.445 197.035 -48.115 197.365 ;
        RECT -48.445 195.675 -48.115 196.005 ;
        RECT -48.445 194.315 -48.115 194.645 ;
        RECT -48.445 192.955 -48.115 193.285 ;
        RECT -48.445 191.595 -48.115 191.925 ;
        RECT -48.445 190.235 -48.115 190.565 ;
        RECT -48.445 188.875 -48.115 189.205 ;
        RECT -48.445 187.515 -48.115 187.845 ;
        RECT -48.445 186.155 -48.115 186.485 ;
        RECT -48.445 184.795 -48.115 185.125 ;
        RECT -48.445 183.435 -48.115 183.765 ;
        RECT -48.445 182.075 -48.115 182.405 ;
        RECT -48.445 180.715 -48.115 181.045 ;
        RECT -48.445 179.355 -48.115 179.685 ;
        RECT -48.445 177.995 -48.115 178.325 ;
        RECT -48.445 176.635 -48.115 176.965 ;
        RECT -48.445 175.275 -48.115 175.605 ;
        RECT -48.445 173.915 -48.115 174.245 ;
        RECT -48.445 172.555 -48.115 172.885 ;
        RECT -48.445 171.195 -48.115 171.525 ;
        RECT -48.445 169.835 -48.115 170.165 ;
        RECT -48.445 168.475 -48.115 168.805 ;
        RECT -48.445 167.115 -48.115 167.445 ;
        RECT -48.445 165.755 -48.115 166.085 ;
        RECT -48.445 164.395 -48.115 164.725 ;
        RECT -48.445 163.035 -48.115 163.365 ;
        RECT -48.445 161.675 -48.115 162.005 ;
        RECT -48.445 160.315 -48.115 160.645 ;
        RECT -48.445 158.955 -48.115 159.285 ;
        RECT -48.445 157.595 -48.115 157.925 ;
        RECT -48.445 156.235 -48.115 156.565 ;
        RECT -48.445 154.875 -48.115 155.205 ;
        RECT -48.445 153.515 -48.115 153.845 ;
        RECT -48.445 152.155 -48.115 152.485 ;
        RECT -48.445 150.795 -48.115 151.125 ;
        RECT -48.445 149.435 -48.115 149.765 ;
        RECT -48.445 148.075 -48.115 148.405 ;
        RECT -48.445 146.715 -48.115 147.045 ;
        RECT -48.445 145.355 -48.115 145.685 ;
        RECT -48.445 143.995 -48.115 144.325 ;
        RECT -48.445 142.635 -48.115 142.965 ;
        RECT -48.445 141.275 -48.115 141.605 ;
        RECT -48.445 139.915 -48.115 140.245 ;
        RECT -48.445 138.555 -48.115 138.885 ;
        RECT -48.445 137.225 -48.115 137.555 ;
        RECT -48.445 135.175 -48.115 135.505 ;
        RECT -48.445 132.815 -48.115 133.145 ;
        RECT -48.445 131.665 -48.115 131.995 ;
        RECT -48.445 129.655 -48.115 129.985 ;
        RECT -48.445 128.505 -48.115 128.835 ;
        RECT -48.445 126.495 -48.115 126.825 ;
        RECT -48.445 125.345 -48.115 125.675 ;
        RECT -48.445 123.335 -48.115 123.665 ;
        RECT -48.445 122.185 -48.115 122.515 ;
        RECT -48.445 120.175 -48.115 120.505 ;
        RECT -48.445 119.025 -48.115 119.355 ;
        RECT -48.445 117.185 -48.115 117.515 ;
        RECT -48.445 115.865 -48.115 116.195 ;
        RECT -48.445 113.855 -48.115 114.185 ;
        RECT -48.445 112.705 -48.115 113.035 ;
        RECT -48.445 110.695 -48.115 111.025 ;
        RECT -48.445 109.545 -48.115 109.875 ;
        RECT -48.445 107.535 -48.115 107.865 ;
        RECT -48.445 106.385 -48.115 106.715 ;
        RECT -48.445 104.375 -48.115 104.705 ;
        RECT -48.445 103.225 -48.115 103.555 ;
        RECT -48.445 100.865 -48.115 101.195 ;
        RECT -48.445 98.81 -48.115 99.14 ;
        RECT -48.445 97.755 -48.115 98.085 ;
        RECT -48.445 96.395 -48.115 96.725 ;
        RECT -48.445 95.035 -48.115 95.365 ;
        RECT -48.445 93.675 -48.115 94.005 ;
        RECT -48.445 92.315 -48.115 92.645 ;
        RECT -48.445 90.955 -48.115 91.285 ;
        RECT -48.445 89.595 -48.115 89.925 ;
        RECT -48.445 88.235 -48.115 88.565 ;
        RECT -48.445 86.875 -48.115 87.205 ;
        RECT -48.445 85.515 -48.115 85.845 ;
        RECT -48.445 84.155 -48.115 84.485 ;
        RECT -48.445 82.795 -48.115 83.125 ;
        RECT -48.445 81.435 -48.115 81.765 ;
        RECT -48.445 80.075 -48.115 80.405 ;
        RECT -48.445 78.715 -48.115 79.045 ;
        RECT -48.445 77.355 -48.115 77.685 ;
        RECT -48.445 75.995 -48.115 76.325 ;
        RECT -48.445 74.635 -48.115 74.965 ;
        RECT -48.445 73.275 -48.115 73.605 ;
        RECT -48.445 71.915 -48.115 72.245 ;
        RECT -48.445 70.555 -48.115 70.885 ;
        RECT -48.445 69.195 -48.115 69.525 ;
        RECT -48.445 67.835 -48.115 68.165 ;
        RECT -48.445 66.475 -48.115 66.805 ;
        RECT -48.445 65.115 -48.115 65.445 ;
        RECT -48.445 63.755 -48.115 64.085 ;
        RECT -48.445 62.395 -48.115 62.725 ;
        RECT -48.445 61.035 -48.115 61.365 ;
        RECT -48.445 59.675 -48.115 60.005 ;
        RECT -48.445 58.315 -48.115 58.645 ;
        RECT -48.445 56.955 -48.115 57.285 ;
        RECT -48.445 55.595 -48.115 55.925 ;
        RECT -48.445 54.235 -48.115 54.565 ;
        RECT -48.445 52.875 -48.115 53.205 ;
        RECT -48.445 51.515 -48.115 51.845 ;
        RECT -48.445 50.155 -48.115 50.485 ;
        RECT -48.445 48.795 -48.115 49.125 ;
        RECT -48.445 47.435 -48.115 47.765 ;
        RECT -48.445 46.075 -48.115 46.405 ;
        RECT -48.445 44.715 -48.115 45.045 ;
        RECT -48.445 43.355 -48.115 43.685 ;
        RECT -48.445 41.995 -48.115 42.325 ;
        RECT -48.445 40.635 -48.115 40.965 ;
        RECT -48.445 39.275 -48.115 39.605 ;
        RECT -48.445 37.915 -48.115 38.245 ;
        RECT -48.445 36.555 -48.115 36.885 ;
        RECT -48.445 35.195 -48.115 35.525 ;
        RECT -48.445 33.835 -48.115 34.165 ;
        RECT -48.445 32.475 -48.115 32.805 ;
        RECT -48.445 31.115 -48.115 31.445 ;
        RECT -48.445 29.755 -48.115 30.085 ;
        RECT -48.445 28.395 -48.115 28.725 ;
        RECT -48.445 27.035 -48.115 27.365 ;
        RECT -48.445 25.675 -48.115 26.005 ;
        RECT -48.445 24.315 -48.115 24.645 ;
        RECT -48.445 22.955 -48.115 23.285 ;
        RECT -48.445 21.595 -48.115 21.925 ;
        RECT -48.445 20.235 -48.115 20.565 ;
        RECT -48.445 18.875 -48.115 19.205 ;
        RECT -48.445 17.515 -48.115 17.845 ;
        RECT -48.445 16.155 -48.115 16.485 ;
        RECT -48.445 14.795 -48.115 15.125 ;
        RECT -48.445 13.435 -48.115 13.765 ;
        RECT -48.445 12.075 -48.115 12.405 ;
        RECT -48.445 10.715 -48.115 11.045 ;
        RECT -48.445 9.355 -48.115 9.685 ;
        RECT -48.445 7.995 -48.115 8.325 ;
        RECT -48.445 6.635 -48.115 6.965 ;
        RECT -48.445 5.275 -48.115 5.605 ;
        RECT -48.445 3.915 -48.115 4.245 ;
        RECT -48.445 2.555 -48.115 2.885 ;
        RECT -48.445 1.195 -48.115 1.525 ;
        RECT -48.445 -0.165 -48.115 0.165 ;
        RECT -48.445 -2.885 -48.115 -2.555 ;
        RECT -48.445 -4.245 -48.115 -3.915 ;
        RECT -48.445 -5.605 -48.115 -5.275 ;
        RECT -48.445 -6.965 -48.115 -6.635 ;
        RECT -48.445 -8.325 -48.115 -7.995 ;
        RECT -48.445 -9.685 -48.115 -9.355 ;
        RECT -48.445 -11.045 -48.115 -10.715 ;
        RECT -48.445 -15.125 -48.115 -14.795 ;
        RECT -48.445 -16.485 -48.115 -16.155 ;
        RECT -48.445 -17.845 -48.115 -17.515 ;
        RECT -48.445 -19.205 -48.115 -18.875 ;
        RECT -48.445 -20.565 -48.115 -20.235 ;
        RECT -48.445 -21.925 -48.115 -21.595 ;
        RECT -48.445 -23.285 -48.115 -22.955 ;
        RECT -48.445 -24.645 -48.115 -24.315 ;
        RECT -48.445 -30.085 -48.115 -29.755 ;
        RECT -48.445 -32.805 -48.115 -32.475 ;
        RECT -48.445 -35.525 -48.115 -35.195 ;
        RECT -48.445 -36.885 -48.115 -36.555 ;
        RECT -48.445 -37.93 -48.115 -37.6 ;
        RECT -48.445 -40.965 -48.115 -40.635 ;
        RECT -48.445 -42.77 -48.115 -42.44 ;
        RECT -48.445 -43.685 -48.115 -43.355 ;
        RECT -48.445 -50.485 -48.115 -50.155 ;
        RECT -48.445 -51.845 -48.115 -51.515 ;
        RECT -48.445 -54.565 -48.115 -54.235 ;
        RECT -48.445 -55.925 -48.115 -55.595 ;
        RECT -48.445 -60.005 -48.115 -59.675 ;
        RECT -48.445 -62.725 -48.115 -62.395 ;
        RECT -48.445 -69.525 -48.115 -69.195 ;
        RECT -48.445 -70.885 -48.115 -70.555 ;
        RECT -48.445 -72.245 -48.115 -71.915 ;
        RECT -48.445 -73.605 -48.115 -73.275 ;
        RECT -48.445 -74.965 -48.115 -74.635 ;
        RECT -48.445 -76.325 -48.115 -75.995 ;
        RECT -48.445 -77.685 -48.115 -77.355 ;
        RECT -48.445 -79.045 -48.115 -78.715 ;
        RECT -48.445 -80.405 -48.115 -80.075 ;
        RECT -48.445 -81.765 -48.115 -81.435 ;
        RECT -48.445 -83.125 -48.115 -82.795 ;
        RECT -48.445 -84.485 -48.115 -84.155 ;
        RECT -48.445 -85.845 -48.115 -85.515 ;
        RECT -48.445 -87.205 -48.115 -86.875 ;
        RECT -48.445 -88.565 -48.115 -88.235 ;
        RECT -48.445 -89.925 -48.115 -89.595 ;
        RECT -48.445 -92.645 -48.115 -92.315 ;
        RECT -48.445 -94.005 -48.115 -93.675 ;
        RECT -48.445 -95.365 -48.115 -95.035 ;
        RECT -48.445 -96.725 -48.115 -96.395 ;
        RECT -48.445 -98.085 -48.115 -97.755 ;
        RECT -48.445 -99.69 -48.115 -99.36 ;
        RECT -48.445 -100.805 -48.115 -100.475 ;
        RECT -48.445 -103.525 -48.115 -103.195 ;
        RECT -48.445 -104.885 -48.115 -104.555 ;
        RECT -48.445 -106.245 -48.115 -105.915 ;
        RECT -48.445 -107.83 -48.115 -107.5 ;
        RECT -48.445 -108.965 -48.115 -108.635 ;
        RECT -48.445 -110.325 -48.115 -109.995 ;
        RECT -48.445 -111.685 -48.115 -111.355 ;
        RECT -48.44 -113.72 -48.12 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -48.445 -175.605 -48.115 -175.275 ;
        RECT -48.445 -176.685 -48.115 -176.355 ;
        RECT -48.445 -178.325 -48.115 -177.995 ;
        RECT -48.445 -179.685 -48.115 -179.355 ;
        RECT -48.445 -181.93 -48.115 -180.8 ;
        RECT -48.44 -182.045 -48.12 -175.275 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.085 241.32 -46.755 242.45 ;
        RECT -47.085 239.195 -46.755 239.525 ;
        RECT -47.085 237.835 -46.755 238.165 ;
        RECT -47.085 236.475 -46.755 236.805 ;
        RECT -47.085 235.115 -46.755 235.445 ;
        RECT -47.085 233.755 -46.755 234.085 ;
        RECT -47.085 232.395 -46.755 232.725 ;
        RECT -47.085 231.035 -46.755 231.365 ;
        RECT -47.085 229.675 -46.755 230.005 ;
        RECT -47.085 228.315 -46.755 228.645 ;
        RECT -47.085 226.955 -46.755 227.285 ;
        RECT -47.085 225.595 -46.755 225.925 ;
        RECT -47.085 224.235 -46.755 224.565 ;
        RECT -47.085 222.875 -46.755 223.205 ;
        RECT -47.085 221.515 -46.755 221.845 ;
        RECT -47.085 220.155 -46.755 220.485 ;
        RECT -47.085 218.795 -46.755 219.125 ;
        RECT -47.085 217.435 -46.755 217.765 ;
        RECT -47.085 216.075 -46.755 216.405 ;
        RECT -47.085 214.715 -46.755 215.045 ;
        RECT -47.085 213.355 -46.755 213.685 ;
        RECT -47.085 211.995 -46.755 212.325 ;
        RECT -47.085 210.635 -46.755 210.965 ;
        RECT -47.085 209.275 -46.755 209.605 ;
        RECT -47.085 207.915 -46.755 208.245 ;
        RECT -47.085 206.555 -46.755 206.885 ;
        RECT -47.085 205.195 -46.755 205.525 ;
        RECT -47.085 203.835 -46.755 204.165 ;
        RECT -47.085 202.475 -46.755 202.805 ;
        RECT -47.085 201.115 -46.755 201.445 ;
        RECT -47.085 199.755 -46.755 200.085 ;
        RECT -47.085 198.395 -46.755 198.725 ;
        RECT -47.085 197.035 -46.755 197.365 ;
        RECT -47.085 195.675 -46.755 196.005 ;
        RECT -47.085 194.315 -46.755 194.645 ;
        RECT -47.085 192.955 -46.755 193.285 ;
        RECT -47.085 191.595 -46.755 191.925 ;
        RECT -47.085 190.235 -46.755 190.565 ;
        RECT -47.085 188.875 -46.755 189.205 ;
        RECT -47.085 187.515 -46.755 187.845 ;
        RECT -47.085 186.155 -46.755 186.485 ;
        RECT -47.085 184.795 -46.755 185.125 ;
        RECT -47.085 183.435 -46.755 183.765 ;
        RECT -47.085 182.075 -46.755 182.405 ;
        RECT -47.085 180.715 -46.755 181.045 ;
        RECT -47.085 179.355 -46.755 179.685 ;
        RECT -47.085 177.995 -46.755 178.325 ;
        RECT -47.085 176.635 -46.755 176.965 ;
        RECT -47.085 175.275 -46.755 175.605 ;
        RECT -47.085 173.915 -46.755 174.245 ;
        RECT -47.085 172.555 -46.755 172.885 ;
        RECT -47.085 171.195 -46.755 171.525 ;
        RECT -47.085 169.835 -46.755 170.165 ;
        RECT -47.085 168.475 -46.755 168.805 ;
        RECT -47.085 167.115 -46.755 167.445 ;
        RECT -47.085 165.755 -46.755 166.085 ;
        RECT -47.085 164.395 -46.755 164.725 ;
        RECT -47.085 163.035 -46.755 163.365 ;
        RECT -47.085 161.675 -46.755 162.005 ;
        RECT -47.085 160.315 -46.755 160.645 ;
        RECT -47.085 158.955 -46.755 159.285 ;
        RECT -47.085 157.595 -46.755 157.925 ;
        RECT -47.085 156.235 -46.755 156.565 ;
        RECT -47.085 154.875 -46.755 155.205 ;
        RECT -47.085 153.515 -46.755 153.845 ;
        RECT -47.085 152.155 -46.755 152.485 ;
        RECT -47.085 150.795 -46.755 151.125 ;
        RECT -47.085 149.435 -46.755 149.765 ;
        RECT -47.085 148.075 -46.755 148.405 ;
        RECT -47.085 146.715 -46.755 147.045 ;
        RECT -47.085 145.355 -46.755 145.685 ;
        RECT -47.085 143.995 -46.755 144.325 ;
        RECT -47.085 142.635 -46.755 142.965 ;
        RECT -47.085 141.275 -46.755 141.605 ;
        RECT -47.085 139.915 -46.755 140.245 ;
        RECT -47.085 138.555 -46.755 138.885 ;
        RECT -47.085 137.195 -46.755 137.525 ;
        RECT -47.085 135.835 -46.755 136.165 ;
        RECT -47.085 134.475 -46.755 134.805 ;
        RECT -47.085 133.115 -46.755 133.445 ;
        RECT -47.085 131.755 -46.755 132.085 ;
        RECT -47.085 130.395 -46.755 130.725 ;
        RECT -47.085 129.035 -46.755 129.365 ;
        RECT -47.085 127.675 -46.755 128.005 ;
        RECT -47.085 126.315 -46.755 126.645 ;
        RECT -47.085 124.955 -46.755 125.285 ;
        RECT -47.085 123.595 -46.755 123.925 ;
        RECT -47.085 122.235 -46.755 122.565 ;
        RECT -47.085 120.875 -46.755 121.205 ;
        RECT -47.085 119.515 -46.755 119.845 ;
        RECT -47.085 118.155 -46.755 118.485 ;
        RECT -47.085 116.795 -46.755 117.125 ;
        RECT -47.085 115.435 -46.755 115.765 ;
        RECT -47.085 114.075 -46.755 114.405 ;
        RECT -47.085 112.715 -46.755 113.045 ;
        RECT -47.085 111.355 -46.755 111.685 ;
        RECT -47.085 109.995 -46.755 110.325 ;
        RECT -47.085 108.635 -46.755 108.965 ;
        RECT -47.085 107.275 -46.755 107.605 ;
        RECT -47.085 105.915 -46.755 106.245 ;
        RECT -47.085 104.555 -46.755 104.885 ;
        RECT -47.085 103.195 -46.755 103.525 ;
        RECT -47.085 101.835 -46.755 102.165 ;
        RECT -47.085 100.475 -46.755 100.805 ;
        RECT -47.085 99.115 -46.755 99.445 ;
        RECT -47.085 97.755 -46.755 98.085 ;
        RECT -47.085 96.395 -46.755 96.725 ;
        RECT -47.085 95.035 -46.755 95.365 ;
        RECT -47.085 93.675 -46.755 94.005 ;
        RECT -47.085 92.315 -46.755 92.645 ;
        RECT -47.085 90.955 -46.755 91.285 ;
        RECT -47.085 89.595 -46.755 89.925 ;
        RECT -47.085 88.235 -46.755 88.565 ;
        RECT -47.085 86.875 -46.755 87.205 ;
        RECT -47.085 85.515 -46.755 85.845 ;
        RECT -47.085 84.155 -46.755 84.485 ;
        RECT -47.085 82.795 -46.755 83.125 ;
        RECT -47.085 81.435 -46.755 81.765 ;
        RECT -47.085 80.075 -46.755 80.405 ;
        RECT -47.085 78.715 -46.755 79.045 ;
        RECT -47.085 77.355 -46.755 77.685 ;
        RECT -47.085 75.995 -46.755 76.325 ;
        RECT -47.085 74.635 -46.755 74.965 ;
        RECT -47.085 73.275 -46.755 73.605 ;
        RECT -47.085 71.915 -46.755 72.245 ;
        RECT -47.085 70.555 -46.755 70.885 ;
        RECT -47.085 69.195 -46.755 69.525 ;
        RECT -47.085 67.835 -46.755 68.165 ;
        RECT -47.085 66.475 -46.755 66.805 ;
        RECT -47.085 65.115 -46.755 65.445 ;
        RECT -47.085 63.755 -46.755 64.085 ;
        RECT -47.085 62.395 -46.755 62.725 ;
        RECT -47.085 61.035 -46.755 61.365 ;
        RECT -47.085 59.675 -46.755 60.005 ;
        RECT -47.085 58.315 -46.755 58.645 ;
        RECT -47.085 56.955 -46.755 57.285 ;
        RECT -47.085 55.595 -46.755 55.925 ;
        RECT -47.085 54.235 -46.755 54.565 ;
        RECT -47.085 52.875 -46.755 53.205 ;
        RECT -47.085 51.515 -46.755 51.845 ;
        RECT -47.085 50.155 -46.755 50.485 ;
        RECT -47.085 48.795 -46.755 49.125 ;
        RECT -47.085 47.435 -46.755 47.765 ;
        RECT -47.085 46.075 -46.755 46.405 ;
        RECT -47.085 44.715 -46.755 45.045 ;
        RECT -47.085 43.355 -46.755 43.685 ;
        RECT -47.085 41.995 -46.755 42.325 ;
        RECT -47.085 40.635 -46.755 40.965 ;
        RECT -47.085 39.275 -46.755 39.605 ;
        RECT -47.085 37.915 -46.755 38.245 ;
        RECT -47.085 36.555 -46.755 36.885 ;
        RECT -47.085 35.195 -46.755 35.525 ;
        RECT -47.085 33.835 -46.755 34.165 ;
        RECT -47.085 32.475 -46.755 32.805 ;
        RECT -47.085 31.115 -46.755 31.445 ;
        RECT -47.085 29.755 -46.755 30.085 ;
        RECT -47.085 28.395 -46.755 28.725 ;
        RECT -47.085 27.035 -46.755 27.365 ;
        RECT -47.085 25.675 -46.755 26.005 ;
        RECT -47.085 24.315 -46.755 24.645 ;
        RECT -47.085 22.955 -46.755 23.285 ;
        RECT -47.085 21.595 -46.755 21.925 ;
        RECT -47.085 20.235 -46.755 20.565 ;
        RECT -47.085 18.875 -46.755 19.205 ;
        RECT -47.085 17.515 -46.755 17.845 ;
        RECT -47.085 16.155 -46.755 16.485 ;
        RECT -47.085 14.795 -46.755 15.125 ;
        RECT -47.085 13.435 -46.755 13.765 ;
        RECT -47.085 12.075 -46.755 12.405 ;
        RECT -47.085 10.715 -46.755 11.045 ;
        RECT -47.085 9.355 -46.755 9.685 ;
        RECT -47.085 7.995 -46.755 8.325 ;
        RECT -47.085 6.635 -46.755 6.965 ;
        RECT -47.085 5.275 -46.755 5.605 ;
        RECT -47.085 3.915 -46.755 4.245 ;
        RECT -47.085 2.555 -46.755 2.885 ;
        RECT -47.085 1.195 -46.755 1.525 ;
        RECT -47.085 -0.165 -46.755 0.165 ;
        RECT -47.08 -1.52 -46.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -47.085 -32.805 -46.755 -32.475 ;
        RECT -47.085 -35.525 -46.755 -35.195 ;
        RECT -47.085 -36.885 -46.755 -36.555 ;
        RECT -47.085 -37.93 -46.755 -37.6 ;
        RECT -47.085 -40.965 -46.755 -40.635 ;
        RECT -47.085 -42.77 -46.755 -42.44 ;
        RECT -47.085 -43.685 -46.755 -43.355 ;
        RECT -47.085 -50.485 -46.755 -50.155 ;
        RECT -47.085 -51.845 -46.755 -51.515 ;
        RECT -47.085 -54.565 -46.755 -54.235 ;
        RECT -47.085 -55.925 -46.755 -55.595 ;
        RECT -47.085 -60.005 -46.755 -59.675 ;
        RECT -47.085 -62.725 -46.755 -62.395 ;
        RECT -47.085 -69.525 -46.755 -69.195 ;
        RECT -47.085 -70.885 -46.755 -70.555 ;
        RECT -47.085 -72.245 -46.755 -71.915 ;
        RECT -47.085 -73.605 -46.755 -73.275 ;
        RECT -47.085 -74.965 -46.755 -74.635 ;
        RECT -47.085 -76.325 -46.755 -75.995 ;
        RECT -47.085 -77.685 -46.755 -77.355 ;
        RECT -47.085 -79.045 -46.755 -78.715 ;
        RECT -47.085 -80.405 -46.755 -80.075 ;
        RECT -47.085 -81.765 -46.755 -81.435 ;
        RECT -47.085 -83.125 -46.755 -82.795 ;
        RECT -47.085 -84.485 -46.755 -84.155 ;
        RECT -47.085 -85.845 -46.755 -85.515 ;
        RECT -47.085 -87.205 -46.755 -86.875 ;
        RECT -47.085 -88.565 -46.755 -88.235 ;
        RECT -47.085 -89.925 -46.755 -89.595 ;
        RECT -47.085 -92.645 -46.755 -92.315 ;
        RECT -47.085 -94.005 -46.755 -93.675 ;
        RECT -47.085 -95.365 -46.755 -95.035 ;
        RECT -47.085 -96.725 -46.755 -96.395 ;
        RECT -47.085 -98.085 -46.755 -97.755 ;
        RECT -47.085 -99.69 -46.755 -99.36 ;
        RECT -47.085 -100.805 -46.755 -100.475 ;
        RECT -47.085 -103.525 -46.755 -103.195 ;
        RECT -47.085 -104.885 -46.755 -104.555 ;
        RECT -47.085 -106.245 -46.755 -105.915 ;
        RECT -47.085 -107.83 -46.755 -107.5 ;
        RECT -47.085 -108.965 -46.755 -108.635 ;
        RECT -47.085 -110.325 -46.755 -109.995 ;
        RECT -47.085 -111.685 -46.755 -111.355 ;
        RECT -47.085 -114.405 -46.755 -114.075 ;
        RECT -47.085 -115.765 -46.755 -115.435 ;
        RECT -47.085 -117.125 -46.755 -116.795 ;
        RECT -47.085 -118.485 -46.755 -118.155 ;
        RECT -47.085 -121.205 -46.755 -120.875 ;
        RECT -47.085 -123.925 -46.755 -123.595 ;
        RECT -47.085 -125.285 -46.755 -124.955 ;
        RECT -47.085 -126.645 -46.755 -126.315 ;
        RECT -47.085 -128.005 -46.755 -127.675 ;
        RECT -47.085 -129.365 -46.755 -129.035 ;
        RECT -47.085 -130.725 -46.755 -130.395 ;
        RECT -47.085 -132.085 -46.755 -131.755 ;
        RECT -47.085 -133.445 -46.755 -133.115 ;
        RECT -47.085 -134.805 -46.755 -134.475 ;
        RECT -47.085 -136.165 -46.755 -135.835 ;
        RECT -47.085 -137.525 -46.755 -137.195 ;
        RECT -47.085 -138.885 -46.755 -138.555 ;
        RECT -47.085 -140.245 -46.755 -139.915 ;
        RECT -47.085 -141.605 -46.755 -141.275 ;
        RECT -47.085 -142.965 -46.755 -142.635 ;
        RECT -47.085 -144.325 -46.755 -143.995 ;
        RECT -47.085 -145.685 -46.755 -145.355 ;
        RECT -47.085 -147.045 -46.755 -146.715 ;
        RECT -47.085 -148.405 -46.755 -148.075 ;
        RECT -47.085 -149.765 -46.755 -149.435 ;
        RECT -47.085 -151.125 -46.755 -150.795 ;
        RECT -47.085 -152.485 -46.755 -152.155 ;
        RECT -47.085 -153.845 -46.755 -153.515 ;
        RECT -47.085 -155.205 -46.755 -154.875 ;
        RECT -47.085 -156.565 -46.755 -156.235 ;
        RECT -47.085 -157.925 -46.755 -157.595 ;
        RECT -47.085 -159.285 -46.755 -158.955 ;
        RECT -47.085 -160.645 -46.755 -160.315 ;
        RECT -47.085 -162.005 -46.755 -161.675 ;
        RECT -47.085 -163.365 -46.755 -163.035 ;
        RECT -47.085 -164.725 -46.755 -164.395 ;
        RECT -47.085 -166.085 -46.755 -165.755 ;
        RECT -47.085 -167.445 -46.755 -167.115 ;
        RECT -47.085 -168.805 -46.755 -168.475 ;
        RECT -47.085 -171.525 -46.755 -171.195 ;
        RECT -47.085 -172.885 -46.755 -172.555 ;
        RECT -47.085 -175.605 -46.755 -175.275 ;
        RECT -47.085 -178.325 -46.755 -177.995 ;
        RECT -47.085 -179.685 -46.755 -179.355 ;
        RECT -47.085 -181.93 -46.755 -180.8 ;
        RECT -47.08 -182.045 -46.76 -31.12 ;
    END
    PORT
      LAYER met3 ;
        RECT -45.725 33.835 -45.395 34.165 ;
        RECT -45.725 32.475 -45.395 32.805 ;
        RECT -45.725 31.115 -45.395 31.445 ;
        RECT -45.725 29.755 -45.395 30.085 ;
        RECT -45.725 28.395 -45.395 28.725 ;
        RECT -45.725 27.035 -45.395 27.365 ;
        RECT -45.725 25.675 -45.395 26.005 ;
        RECT -45.725 24.315 -45.395 24.645 ;
        RECT -45.725 22.955 -45.395 23.285 ;
        RECT -45.725 21.595 -45.395 21.925 ;
        RECT -45.725 20.235 -45.395 20.565 ;
        RECT -45.725 18.875 -45.395 19.205 ;
        RECT -45.725 17.515 -45.395 17.845 ;
        RECT -45.725 16.155 -45.395 16.485 ;
        RECT -45.725 14.795 -45.395 15.125 ;
        RECT -45.725 13.435 -45.395 13.765 ;
        RECT -45.725 12.075 -45.395 12.405 ;
        RECT -45.725 10.715 -45.395 11.045 ;
        RECT -45.725 9.355 -45.395 9.685 ;
        RECT -45.725 7.995 -45.395 8.325 ;
        RECT -45.725 6.635 -45.395 6.965 ;
        RECT -45.725 5.275 -45.395 5.605 ;
        RECT -45.725 3.915 -45.395 4.245 ;
        RECT -45.725 2.555 -45.395 2.885 ;
        RECT -45.725 1.195 -45.395 1.525 ;
        RECT -45.725 -0.165 -45.395 0.165 ;
        RECT -45.725 -4.245 -45.395 -3.915 ;
        RECT -45.725 -5.605 -45.395 -5.275 ;
        RECT -45.725 -6.965 -45.395 -6.635 ;
        RECT -45.725 -8.325 -45.395 -7.995 ;
        RECT -45.725 -11.045 -45.395 -10.715 ;
        RECT -45.725 -15.125 -45.395 -14.795 ;
        RECT -45.725 -16.485 -45.395 -16.155 ;
        RECT -45.725 -17.845 -45.395 -17.515 ;
        RECT -45.725 -19.205 -45.395 -18.875 ;
        RECT -45.725 -20.565 -45.395 -20.235 ;
        RECT -45.725 -21.925 -45.395 -21.595 ;
        RECT -45.725 -23.285 -45.395 -22.955 ;
        RECT -45.725 -24.645 -45.395 -24.315 ;
        RECT -45.725 -32.805 -45.395 -32.475 ;
        RECT -45.725 -35.525 -45.395 -35.195 ;
        RECT -45.725 -36.885 -45.395 -36.555 ;
        RECT -45.725 -37.93 -45.395 -37.6 ;
        RECT -45.725 -40.965 -45.395 -40.635 ;
        RECT -45.725 -42.77 -45.395 -42.44 ;
        RECT -45.725 -43.685 -45.395 -43.355 ;
        RECT -45.725 -50.485 -45.395 -50.155 ;
        RECT -45.725 -51.845 -45.395 -51.515 ;
        RECT -45.725 -54.565 -45.395 -54.235 ;
        RECT -45.725 -55.925 -45.395 -55.595 ;
        RECT -45.725 -60.005 -45.395 -59.675 ;
        RECT -45.725 -62.725 -45.395 -62.395 ;
        RECT -45.725 -69.525 -45.395 -69.195 ;
        RECT -45.725 -70.885 -45.395 -70.555 ;
        RECT -45.725 -72.245 -45.395 -71.915 ;
        RECT -45.725 -73.605 -45.395 -73.275 ;
        RECT -45.725 -74.965 -45.395 -74.635 ;
        RECT -45.725 -76.325 -45.395 -75.995 ;
        RECT -45.725 -77.685 -45.395 -77.355 ;
        RECT -45.725 -79.045 -45.395 -78.715 ;
        RECT -45.725 -80.405 -45.395 -80.075 ;
        RECT -45.725 -81.765 -45.395 -81.435 ;
        RECT -45.725 -83.125 -45.395 -82.795 ;
        RECT -45.725 -84.485 -45.395 -84.155 ;
        RECT -45.725 -85.845 -45.395 -85.515 ;
        RECT -45.725 -87.205 -45.395 -86.875 ;
        RECT -45.725 -88.565 -45.395 -88.235 ;
        RECT -45.725 -89.925 -45.395 -89.595 ;
        RECT -45.725 -92.645 -45.395 -92.315 ;
        RECT -45.725 -94.005 -45.395 -93.675 ;
        RECT -45.725 -95.365 -45.395 -95.035 ;
        RECT -45.725 -96.725 -45.395 -96.395 ;
        RECT -45.725 -98.085 -45.395 -97.755 ;
        RECT -45.725 -99.69 -45.395 -99.36 ;
        RECT -45.725 -100.805 -45.395 -100.475 ;
        RECT -45.725 -103.525 -45.395 -103.195 ;
        RECT -45.725 -104.885 -45.395 -104.555 ;
        RECT -45.725 -106.245 -45.395 -105.915 ;
        RECT -45.725 -107.83 -45.395 -107.5 ;
        RECT -45.725 -108.965 -45.395 -108.635 ;
        RECT -45.725 -110.325 -45.395 -109.995 ;
        RECT -45.725 -111.685 -45.395 -111.355 ;
        RECT -45.725 -114.405 -45.395 -114.075 ;
        RECT -45.725 -115.765 -45.395 -115.435 ;
        RECT -45.725 -117.125 -45.395 -116.795 ;
        RECT -45.725 -118.485 -45.395 -118.155 ;
        RECT -45.725 -121.205 -45.395 -120.875 ;
        RECT -45.725 -123.925 -45.395 -123.595 ;
        RECT -45.725 -125.285 -45.395 -124.955 ;
        RECT -45.725 -126.645 -45.395 -126.315 ;
        RECT -45.725 -128.005 -45.395 -127.675 ;
        RECT -45.725 -129.365 -45.395 -129.035 ;
        RECT -45.725 -130.725 -45.395 -130.395 ;
        RECT -45.725 -132.085 -45.395 -131.755 ;
        RECT -45.725 -133.445 -45.395 -133.115 ;
        RECT -45.725 -134.805 -45.395 -134.475 ;
        RECT -45.725 -136.165 -45.395 -135.835 ;
        RECT -45.725 -137.525 -45.395 -137.195 ;
        RECT -45.725 -138.885 -45.395 -138.555 ;
        RECT -45.725 -140.245 -45.395 -139.915 ;
        RECT -45.725 -141.605 -45.395 -141.275 ;
        RECT -45.725 -142.965 -45.395 -142.635 ;
        RECT -45.725 -144.325 -45.395 -143.995 ;
        RECT -45.725 -145.685 -45.395 -145.355 ;
        RECT -45.725 -147.045 -45.395 -146.715 ;
        RECT -45.725 -148.405 -45.395 -148.075 ;
        RECT -45.725 -149.765 -45.395 -149.435 ;
        RECT -45.725 -151.125 -45.395 -150.795 ;
        RECT -45.725 -152.485 -45.395 -152.155 ;
        RECT -45.725 -153.845 -45.395 -153.515 ;
        RECT -45.725 -155.205 -45.395 -154.875 ;
        RECT -45.725 -156.565 -45.395 -156.235 ;
        RECT -45.725 -157.925 -45.395 -157.595 ;
        RECT -45.725 -159.285 -45.395 -158.955 ;
        RECT -45.725 -160.645 -45.395 -160.315 ;
        RECT -45.725 -162.005 -45.395 -161.675 ;
        RECT -45.725 -163.365 -45.395 -163.035 ;
        RECT -45.725 -164.725 -45.395 -164.395 ;
        RECT -45.725 -166.085 -45.395 -165.755 ;
        RECT -45.725 -167.445 -45.395 -167.115 ;
        RECT -45.725 -168.805 -45.395 -168.475 ;
        RECT -45.725 -171.525 -45.395 -171.195 ;
        RECT -45.725 -175.605 -45.395 -175.275 ;
        RECT -45.725 -176.685 -45.395 -176.355 ;
        RECT -45.725 -178.325 -45.395 -177.995 ;
        RECT -45.725 -179.685 -45.395 -179.355 ;
        RECT -45.725 -181.93 -45.395 -180.8 ;
        RECT -45.72 -182.045 -45.4 242.565 ;
        RECT -45.725 241.32 -45.395 242.45 ;
        RECT -45.725 239.195 -45.395 239.525 ;
        RECT -45.725 237.835 -45.395 238.165 ;
        RECT -45.725 236.475 -45.395 236.805 ;
        RECT -45.725 235.115 -45.395 235.445 ;
        RECT -45.725 233.755 -45.395 234.085 ;
        RECT -45.725 232.395 -45.395 232.725 ;
        RECT -45.725 231.035 -45.395 231.365 ;
        RECT -45.725 229.675 -45.395 230.005 ;
        RECT -45.725 228.315 -45.395 228.645 ;
        RECT -45.725 226.955 -45.395 227.285 ;
        RECT -45.725 225.595 -45.395 225.925 ;
        RECT -45.725 224.235 -45.395 224.565 ;
        RECT -45.725 222.875 -45.395 223.205 ;
        RECT -45.725 221.515 -45.395 221.845 ;
        RECT -45.725 220.155 -45.395 220.485 ;
        RECT -45.725 218.795 -45.395 219.125 ;
        RECT -45.725 217.435 -45.395 217.765 ;
        RECT -45.725 216.075 -45.395 216.405 ;
        RECT -45.725 214.715 -45.395 215.045 ;
        RECT -45.725 213.355 -45.395 213.685 ;
        RECT -45.725 211.995 -45.395 212.325 ;
        RECT -45.725 210.635 -45.395 210.965 ;
        RECT -45.725 209.275 -45.395 209.605 ;
        RECT -45.725 207.915 -45.395 208.245 ;
        RECT -45.725 206.555 -45.395 206.885 ;
        RECT -45.725 205.195 -45.395 205.525 ;
        RECT -45.725 203.835 -45.395 204.165 ;
        RECT -45.725 202.475 -45.395 202.805 ;
        RECT -45.725 201.115 -45.395 201.445 ;
        RECT -45.725 199.755 -45.395 200.085 ;
        RECT -45.725 198.395 -45.395 198.725 ;
        RECT -45.725 197.035 -45.395 197.365 ;
        RECT -45.725 195.675 -45.395 196.005 ;
        RECT -45.725 194.315 -45.395 194.645 ;
        RECT -45.725 192.955 -45.395 193.285 ;
        RECT -45.725 191.595 -45.395 191.925 ;
        RECT -45.725 190.235 -45.395 190.565 ;
        RECT -45.725 188.875 -45.395 189.205 ;
        RECT -45.725 187.515 -45.395 187.845 ;
        RECT -45.725 186.155 -45.395 186.485 ;
        RECT -45.725 184.795 -45.395 185.125 ;
        RECT -45.725 183.435 -45.395 183.765 ;
        RECT -45.725 182.075 -45.395 182.405 ;
        RECT -45.725 180.715 -45.395 181.045 ;
        RECT -45.725 179.355 -45.395 179.685 ;
        RECT -45.725 177.995 -45.395 178.325 ;
        RECT -45.725 176.635 -45.395 176.965 ;
        RECT -45.725 175.275 -45.395 175.605 ;
        RECT -45.725 173.915 -45.395 174.245 ;
        RECT -45.725 172.555 -45.395 172.885 ;
        RECT -45.725 171.195 -45.395 171.525 ;
        RECT -45.725 169.835 -45.395 170.165 ;
        RECT -45.725 168.475 -45.395 168.805 ;
        RECT -45.725 167.115 -45.395 167.445 ;
        RECT -45.725 165.755 -45.395 166.085 ;
        RECT -45.725 164.395 -45.395 164.725 ;
        RECT -45.725 163.035 -45.395 163.365 ;
        RECT -45.725 161.675 -45.395 162.005 ;
        RECT -45.725 160.315 -45.395 160.645 ;
        RECT -45.725 158.955 -45.395 159.285 ;
        RECT -45.725 157.595 -45.395 157.925 ;
        RECT -45.725 156.235 -45.395 156.565 ;
        RECT -45.725 154.875 -45.395 155.205 ;
        RECT -45.725 153.515 -45.395 153.845 ;
        RECT -45.725 152.155 -45.395 152.485 ;
        RECT -45.725 150.795 -45.395 151.125 ;
        RECT -45.725 149.435 -45.395 149.765 ;
        RECT -45.725 148.075 -45.395 148.405 ;
        RECT -45.725 146.715 -45.395 147.045 ;
        RECT -45.725 145.355 -45.395 145.685 ;
        RECT -45.725 143.995 -45.395 144.325 ;
        RECT -45.725 142.635 -45.395 142.965 ;
        RECT -45.725 141.275 -45.395 141.605 ;
        RECT -45.725 139.915 -45.395 140.245 ;
        RECT -45.725 138.555 -45.395 138.885 ;
        RECT -45.725 137.195 -45.395 137.525 ;
        RECT -45.725 135.835 -45.395 136.165 ;
        RECT -45.725 134.475 -45.395 134.805 ;
        RECT -45.725 133.115 -45.395 133.445 ;
        RECT -45.725 131.755 -45.395 132.085 ;
        RECT -45.725 130.395 -45.395 130.725 ;
        RECT -45.725 129.035 -45.395 129.365 ;
        RECT -45.725 127.675 -45.395 128.005 ;
        RECT -45.725 126.315 -45.395 126.645 ;
        RECT -45.725 124.955 -45.395 125.285 ;
        RECT -45.725 123.595 -45.395 123.925 ;
        RECT -45.725 122.235 -45.395 122.565 ;
        RECT -45.725 120.875 -45.395 121.205 ;
        RECT -45.725 119.515 -45.395 119.845 ;
        RECT -45.725 118.155 -45.395 118.485 ;
        RECT -45.725 116.795 -45.395 117.125 ;
        RECT -45.725 115.435 -45.395 115.765 ;
        RECT -45.725 114.075 -45.395 114.405 ;
        RECT -45.725 112.715 -45.395 113.045 ;
        RECT -45.725 111.355 -45.395 111.685 ;
        RECT -45.725 109.995 -45.395 110.325 ;
        RECT -45.725 108.635 -45.395 108.965 ;
        RECT -45.725 107.275 -45.395 107.605 ;
        RECT -45.725 105.915 -45.395 106.245 ;
        RECT -45.725 104.555 -45.395 104.885 ;
        RECT -45.725 103.195 -45.395 103.525 ;
        RECT -45.725 101.835 -45.395 102.165 ;
        RECT -45.725 100.475 -45.395 100.805 ;
        RECT -45.725 99.115 -45.395 99.445 ;
        RECT -45.725 97.755 -45.395 98.085 ;
        RECT -45.725 96.395 -45.395 96.725 ;
        RECT -45.725 95.035 -45.395 95.365 ;
        RECT -45.725 93.675 -45.395 94.005 ;
        RECT -45.725 92.315 -45.395 92.645 ;
        RECT -45.725 90.955 -45.395 91.285 ;
        RECT -45.725 89.595 -45.395 89.925 ;
        RECT -45.725 88.235 -45.395 88.565 ;
        RECT -45.725 86.875 -45.395 87.205 ;
        RECT -45.725 85.515 -45.395 85.845 ;
        RECT -45.725 84.155 -45.395 84.485 ;
        RECT -45.725 82.795 -45.395 83.125 ;
        RECT -45.725 81.435 -45.395 81.765 ;
        RECT -45.725 80.075 -45.395 80.405 ;
        RECT -45.725 78.715 -45.395 79.045 ;
        RECT -45.725 77.355 -45.395 77.685 ;
        RECT -45.725 75.995 -45.395 76.325 ;
        RECT -45.725 74.635 -45.395 74.965 ;
        RECT -45.725 73.275 -45.395 73.605 ;
        RECT -45.725 71.915 -45.395 72.245 ;
        RECT -45.725 70.555 -45.395 70.885 ;
        RECT -45.725 69.195 -45.395 69.525 ;
        RECT -45.725 67.835 -45.395 68.165 ;
        RECT -45.725 66.475 -45.395 66.805 ;
        RECT -45.725 65.115 -45.395 65.445 ;
        RECT -45.725 63.755 -45.395 64.085 ;
        RECT -45.725 62.395 -45.395 62.725 ;
        RECT -45.725 61.035 -45.395 61.365 ;
        RECT -45.725 59.675 -45.395 60.005 ;
        RECT -45.725 58.315 -45.395 58.645 ;
        RECT -45.725 56.955 -45.395 57.285 ;
        RECT -45.725 55.595 -45.395 55.925 ;
        RECT -45.725 54.235 -45.395 54.565 ;
        RECT -45.725 52.875 -45.395 53.205 ;
        RECT -45.725 51.515 -45.395 51.845 ;
        RECT -45.725 50.155 -45.395 50.485 ;
        RECT -45.725 48.795 -45.395 49.125 ;
        RECT -45.725 47.435 -45.395 47.765 ;
        RECT -45.725 46.075 -45.395 46.405 ;
        RECT -45.725 44.715 -45.395 45.045 ;
        RECT -45.725 43.355 -45.395 43.685 ;
        RECT -45.725 41.995 -45.395 42.325 ;
        RECT -45.725 40.635 -45.395 40.965 ;
        RECT -45.725 39.275 -45.395 39.605 ;
        RECT -45.725 37.915 -45.395 38.245 ;
        RECT -45.725 36.555 -45.395 36.885 ;
        RECT -45.725 35.195 -45.395 35.525 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.245 241.32 -54.915 242.45 ;
        RECT -55.245 239.195 -54.915 239.525 ;
        RECT -55.245 237.835 -54.915 238.165 ;
        RECT -55.245 236.475 -54.915 236.805 ;
        RECT -55.245 235.115 -54.915 235.445 ;
        RECT -55.245 233.755 -54.915 234.085 ;
        RECT -55.245 232.395 -54.915 232.725 ;
        RECT -55.245 231.035 -54.915 231.365 ;
        RECT -55.245 229.675 -54.915 230.005 ;
        RECT -55.245 228.315 -54.915 228.645 ;
        RECT -55.245 226.955 -54.915 227.285 ;
        RECT -55.245 225.595 -54.915 225.925 ;
        RECT -55.245 224.235 -54.915 224.565 ;
        RECT -55.245 222.875 -54.915 223.205 ;
        RECT -55.245 221.515 -54.915 221.845 ;
        RECT -55.245 220.155 -54.915 220.485 ;
        RECT -55.245 218.795 -54.915 219.125 ;
        RECT -55.245 217.435 -54.915 217.765 ;
        RECT -55.245 216.075 -54.915 216.405 ;
        RECT -55.245 214.715 -54.915 215.045 ;
        RECT -55.245 213.355 -54.915 213.685 ;
        RECT -55.245 211.995 -54.915 212.325 ;
        RECT -55.245 210.635 -54.915 210.965 ;
        RECT -55.245 209.275 -54.915 209.605 ;
        RECT -55.245 207.915 -54.915 208.245 ;
        RECT -55.245 206.555 -54.915 206.885 ;
        RECT -55.245 205.195 -54.915 205.525 ;
        RECT -55.245 203.835 -54.915 204.165 ;
        RECT -55.245 202.475 -54.915 202.805 ;
        RECT -55.245 201.115 -54.915 201.445 ;
        RECT -55.245 199.755 -54.915 200.085 ;
        RECT -55.245 198.395 -54.915 198.725 ;
        RECT -55.245 197.035 -54.915 197.365 ;
        RECT -55.245 195.675 -54.915 196.005 ;
        RECT -55.245 194.315 -54.915 194.645 ;
        RECT -55.245 192.955 -54.915 193.285 ;
        RECT -55.245 191.595 -54.915 191.925 ;
        RECT -55.245 190.235 -54.915 190.565 ;
        RECT -55.245 188.875 -54.915 189.205 ;
        RECT -55.245 187.515 -54.915 187.845 ;
        RECT -55.245 186.155 -54.915 186.485 ;
        RECT -55.245 184.795 -54.915 185.125 ;
        RECT -55.245 183.435 -54.915 183.765 ;
        RECT -55.245 182.075 -54.915 182.405 ;
        RECT -55.245 180.715 -54.915 181.045 ;
        RECT -55.245 179.355 -54.915 179.685 ;
        RECT -55.245 177.995 -54.915 178.325 ;
        RECT -55.245 176.635 -54.915 176.965 ;
        RECT -55.245 175.275 -54.915 175.605 ;
        RECT -55.245 173.915 -54.915 174.245 ;
        RECT -55.245 172.555 -54.915 172.885 ;
        RECT -55.245 171.195 -54.915 171.525 ;
        RECT -55.245 169.835 -54.915 170.165 ;
        RECT -55.245 168.475 -54.915 168.805 ;
        RECT -55.245 167.115 -54.915 167.445 ;
        RECT -55.245 165.755 -54.915 166.085 ;
        RECT -55.245 164.395 -54.915 164.725 ;
        RECT -55.245 163.035 -54.915 163.365 ;
        RECT -55.245 161.675 -54.915 162.005 ;
        RECT -55.245 160.315 -54.915 160.645 ;
        RECT -55.245 158.955 -54.915 159.285 ;
        RECT -55.245 157.595 -54.915 157.925 ;
        RECT -55.245 156.235 -54.915 156.565 ;
        RECT -55.245 154.875 -54.915 155.205 ;
        RECT -55.245 153.515 -54.915 153.845 ;
        RECT -55.245 152.155 -54.915 152.485 ;
        RECT -55.245 150.795 -54.915 151.125 ;
        RECT -55.245 149.435 -54.915 149.765 ;
        RECT -55.245 148.075 -54.915 148.405 ;
        RECT -55.245 146.715 -54.915 147.045 ;
        RECT -55.245 145.355 -54.915 145.685 ;
        RECT -55.245 143.995 -54.915 144.325 ;
        RECT -55.245 142.635 -54.915 142.965 ;
        RECT -55.245 141.275 -54.915 141.605 ;
        RECT -55.245 139.915 -54.915 140.245 ;
        RECT -55.245 138.555 -54.915 138.885 ;
        RECT -55.24 138.555 -54.92 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -55.245 97.755 -54.915 98.085 ;
        RECT -55.245 96.395 -54.915 96.725 ;
        RECT -55.245 95.035 -54.915 95.365 ;
        RECT -55.245 93.675 -54.915 94.005 ;
        RECT -55.245 92.315 -54.915 92.645 ;
        RECT -55.245 89.595 -54.915 89.925 ;
        RECT -55.245 88.235 -54.915 88.565 ;
        RECT -55.245 84.155 -54.915 84.485 ;
        RECT -55.245 82.795 -54.915 83.125 ;
        RECT -55.245 81.435 -54.915 81.765 ;
        RECT -55.245 80.075 -54.915 80.405 ;
        RECT -55.245 78.715 -54.915 79.045 ;
        RECT -55.245 77.355 -54.915 77.685 ;
        RECT -55.245 75.995 -54.915 76.325 ;
        RECT -55.245 74.635 -54.915 74.965 ;
        RECT -55.245 73.275 -54.915 73.605 ;
        RECT -55.245 71.915 -54.915 72.245 ;
        RECT -55.245 70.555 -54.915 70.885 ;
        RECT -55.245 69.195 -54.915 69.525 ;
        RECT -55.245 67.835 -54.915 68.165 ;
        RECT -55.245 66.475 -54.915 66.805 ;
        RECT -55.245 65.115 -54.915 65.445 ;
        RECT -55.245 63.755 -54.915 64.085 ;
        RECT -55.245 62.395 -54.915 62.725 ;
        RECT -55.245 61.035 -54.915 61.365 ;
        RECT -55.245 59.675 -54.915 60.005 ;
        RECT -55.245 58.315 -54.915 58.645 ;
        RECT -55.245 56.955 -54.915 57.285 ;
        RECT -55.245 55.595 -54.915 55.925 ;
        RECT -55.245 54.235 -54.915 54.565 ;
        RECT -55.245 52.875 -54.915 53.205 ;
        RECT -55.245 51.515 -54.915 51.845 ;
        RECT -55.245 50.155 -54.915 50.485 ;
        RECT -55.245 48.795 -54.915 49.125 ;
        RECT -55.245 47.435 -54.915 47.765 ;
        RECT -55.245 46.075 -54.915 46.405 ;
        RECT -55.245 44.715 -54.915 45.045 ;
        RECT -55.245 43.355 -54.915 43.685 ;
        RECT -55.245 41.995 -54.915 42.325 ;
        RECT -55.245 40.635 -54.915 40.965 ;
        RECT -55.245 39.275 -54.915 39.605 ;
        RECT -55.245 37.915 -54.915 38.245 ;
        RECT -55.245 36.555 -54.915 36.885 ;
        RECT -55.245 35.195 -54.915 35.525 ;
        RECT -55.245 33.835 -54.915 34.165 ;
        RECT -55.245 32.475 -54.915 32.805 ;
        RECT -55.245 31.115 -54.915 31.445 ;
        RECT -55.245 29.755 -54.915 30.085 ;
        RECT -55.245 28.395 -54.915 28.725 ;
        RECT -55.245 27.035 -54.915 27.365 ;
        RECT -55.245 25.675 -54.915 26.005 ;
        RECT -55.245 24.315 -54.915 24.645 ;
        RECT -55.245 22.955 -54.915 23.285 ;
        RECT -55.245 21.595 -54.915 21.925 ;
        RECT -55.245 20.235 -54.915 20.565 ;
        RECT -55.245 18.875 -54.915 19.205 ;
        RECT -55.245 17.515 -54.915 17.845 ;
        RECT -55.245 16.155 -54.915 16.485 ;
        RECT -55.245 14.795 -54.915 15.125 ;
        RECT -55.245 13.435 -54.915 13.765 ;
        RECT -55.245 12.075 -54.915 12.405 ;
        RECT -55.245 10.715 -54.915 11.045 ;
        RECT -55.245 9.355 -54.915 9.685 ;
        RECT -55.245 7.995 -54.915 8.325 ;
        RECT -55.245 6.635 -54.915 6.965 ;
        RECT -55.245 5.275 -54.915 5.605 ;
        RECT -55.245 3.915 -54.915 4.245 ;
        RECT -55.245 2.555 -54.915 2.885 ;
        RECT -55.245 1.195 -54.915 1.525 ;
        RECT -55.245 -0.165 -54.915 0.165 ;
        RECT -55.245 -2.885 -54.915 -2.555 ;
        RECT -55.245 -4.245 -54.915 -3.915 ;
        RECT -55.245 -5.605 -54.915 -5.275 ;
        RECT -55.245 -6.965 -54.915 -6.635 ;
        RECT -55.245 -8.325 -54.915 -7.995 ;
        RECT -55.245 -9.685 -54.915 -9.355 ;
        RECT -55.245 -11.045 -54.915 -10.715 ;
        RECT -55.245 -12.405 -54.915 -12.075 ;
        RECT -55.245 -13.765 -54.915 -13.435 ;
        RECT -55.245 -15.125 -54.915 -14.795 ;
        RECT -55.245 -16.485 -54.915 -16.155 ;
        RECT -55.245 -17.845 -54.915 -17.515 ;
        RECT -55.245 -19.205 -54.915 -18.875 ;
        RECT -55.245 -20.565 -54.915 -20.235 ;
        RECT -55.245 -21.925 -54.915 -21.595 ;
        RECT -55.245 -23.285 -54.915 -22.955 ;
        RECT -55.245 -24.645 -54.915 -24.315 ;
        RECT -55.245 -30.085 -54.915 -29.755 ;
        RECT -55.245 -31.445 -54.915 -31.115 ;
        RECT -55.245 -32.805 -54.915 -32.475 ;
        RECT -55.245 -34.165 -54.915 -33.835 ;
        RECT -55.245 -35.525 -54.915 -35.195 ;
        RECT -55.245 -36.885 -54.915 -36.555 ;
        RECT -55.245 -38.245 -54.915 -37.915 ;
        RECT -55.245 -39.605 -54.915 -39.275 ;
        RECT -55.245 -40.965 -54.915 -40.635 ;
        RECT -55.245 -42.325 -54.915 -41.995 ;
        RECT -55.245 -43.685 -54.915 -43.355 ;
        RECT -55.245 -45.045 -54.915 -44.715 ;
        RECT -55.245 -46.405 -54.915 -46.075 ;
        RECT -55.245 -47.765 -54.915 -47.435 ;
        RECT -55.245 -49.125 -54.915 -48.795 ;
        RECT -55.245 -50.485 -54.915 -50.155 ;
        RECT -55.245 -51.845 -54.915 -51.515 ;
        RECT -55.245 -53.205 -54.915 -52.875 ;
        RECT -55.245 -54.565 -54.915 -54.235 ;
        RECT -55.245 -55.925 -54.915 -55.595 ;
        RECT -55.245 -57.285 -54.915 -56.955 ;
        RECT -55.245 -58.645 -54.915 -58.315 ;
        RECT -55.245 -60.005 -54.915 -59.675 ;
        RECT -55.245 -61.365 -54.915 -61.035 ;
        RECT -55.245 -62.725 -54.915 -62.395 ;
        RECT -55.245 -64.085 -54.915 -63.755 ;
        RECT -55.245 -65.445 -54.915 -65.115 ;
        RECT -55.245 -66.805 -54.915 -66.475 ;
        RECT -55.245 -68.165 -54.915 -67.835 ;
        RECT -55.245 -69.525 -54.915 -69.195 ;
        RECT -55.245 -70.885 -54.915 -70.555 ;
        RECT -55.245 -72.245 -54.915 -71.915 ;
        RECT -55.245 -73.605 -54.915 -73.275 ;
        RECT -55.245 -74.965 -54.915 -74.635 ;
        RECT -55.245 -76.325 -54.915 -75.995 ;
        RECT -55.245 -77.685 -54.915 -77.355 ;
        RECT -55.245 -79.045 -54.915 -78.715 ;
        RECT -55.245 -80.405 -54.915 -80.075 ;
        RECT -55.245 -81.765 -54.915 -81.435 ;
        RECT -55.245 -83.125 -54.915 -82.795 ;
        RECT -55.245 -84.485 -54.915 -84.155 ;
        RECT -55.245 -85.845 -54.915 -85.515 ;
        RECT -55.245 -87.205 -54.915 -86.875 ;
        RECT -55.245 -88.565 -54.915 -88.235 ;
        RECT -55.245 -89.925 -54.915 -89.595 ;
        RECT -55.245 -92.645 -54.915 -92.315 ;
        RECT -55.245 -94.005 -54.915 -93.675 ;
        RECT -55.245 -95.365 -54.915 -95.035 ;
        RECT -55.245 -96.725 -54.915 -96.395 ;
        RECT -55.245 -98.085 -54.915 -97.755 ;
        RECT -55.245 -99.69 -54.915 -99.36 ;
        RECT -55.245 -100.805 -54.915 -100.475 ;
        RECT -55.245 -103.525 -54.915 -103.195 ;
        RECT -55.245 -104.885 -54.915 -104.555 ;
        RECT -55.245 -106.245 -54.915 -105.915 ;
        RECT -55.245 -107.83 -54.915 -107.5 ;
        RECT -55.245 -108.965 -54.915 -108.635 ;
        RECT -55.245 -110.325 -54.915 -109.995 ;
        RECT -55.245 -111.685 -54.915 -111.355 ;
        RECT -55.245 -114.405 -54.915 -114.075 ;
        RECT -55.245 -115.765 -54.915 -115.435 ;
        RECT -55.245 -117.125 -54.915 -116.795 ;
        RECT -55.245 -118.485 -54.915 -118.155 ;
        RECT -55.245 -119.845 -54.915 -119.515 ;
        RECT -55.245 -121.205 -54.915 -120.875 ;
        RECT -55.245 -123.925 -54.915 -123.595 ;
        RECT -55.245 -125.285 -54.915 -124.955 ;
        RECT -55.245 -126.645 -54.915 -126.315 ;
        RECT -55.245 -128.005 -54.915 -127.675 ;
        RECT -55.245 -129.365 -54.915 -129.035 ;
        RECT -55.245 -130.725 -54.915 -130.395 ;
        RECT -55.245 -132.085 -54.915 -131.755 ;
        RECT -55.245 -133.445 -54.915 -133.115 ;
        RECT -55.245 -134.805 -54.915 -134.475 ;
        RECT -55.245 -136.165 -54.915 -135.835 ;
        RECT -55.245 -137.525 -54.915 -137.195 ;
        RECT -55.245 -138.885 -54.915 -138.555 ;
        RECT -55.245 -140.245 -54.915 -139.915 ;
        RECT -55.245 -141.605 -54.915 -141.275 ;
        RECT -55.245 -142.965 -54.915 -142.635 ;
        RECT -55.245 -144.325 -54.915 -143.995 ;
        RECT -55.245 -145.685 -54.915 -145.355 ;
        RECT -55.245 -147.045 -54.915 -146.715 ;
        RECT -55.245 -148.405 -54.915 -148.075 ;
        RECT -55.245 -149.765 -54.915 -149.435 ;
        RECT -55.245 -151.125 -54.915 -150.795 ;
        RECT -55.245 -152.485 -54.915 -152.155 ;
        RECT -55.245 -153.845 -54.915 -153.515 ;
        RECT -55.245 -155.205 -54.915 -154.875 ;
        RECT -55.245 -156.565 -54.915 -156.235 ;
        RECT -55.245 -157.925 -54.915 -157.595 ;
        RECT -55.245 -159.285 -54.915 -158.955 ;
        RECT -55.245 -160.645 -54.915 -160.315 ;
        RECT -55.245 -162.005 -54.915 -161.675 ;
        RECT -55.245 -163.365 -54.915 -163.035 ;
        RECT -55.245 -164.725 -54.915 -164.395 ;
        RECT -55.245 -166.085 -54.915 -165.755 ;
        RECT -55.245 -167.445 -54.915 -167.115 ;
        RECT -55.245 -168.805 -54.915 -168.475 ;
        RECT -55.245 -171.525 -54.915 -171.195 ;
        RECT -55.245 -172.885 -54.915 -172.555 ;
        RECT -55.245 -174.245 -54.915 -173.915 ;
        RECT -55.245 -175.605 -54.915 -175.275 ;
        RECT -55.245 -176.685 -54.915 -176.355 ;
        RECT -55.245 -178.325 -54.915 -177.995 ;
        RECT -55.245 -179.685 -54.915 -179.355 ;
        RECT -55.245 -181.93 -54.915 -180.8 ;
        RECT -55.24 -182.045 -54.92 98.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.885 241.32 -53.555 242.45 ;
        RECT -53.885 239.195 -53.555 239.525 ;
        RECT -53.885 237.835 -53.555 238.165 ;
        RECT -53.885 236.475 -53.555 236.805 ;
        RECT -53.885 235.115 -53.555 235.445 ;
        RECT -53.885 233.755 -53.555 234.085 ;
        RECT -53.885 232.395 -53.555 232.725 ;
        RECT -53.885 231.035 -53.555 231.365 ;
        RECT -53.885 229.675 -53.555 230.005 ;
        RECT -53.885 228.315 -53.555 228.645 ;
        RECT -53.885 226.955 -53.555 227.285 ;
        RECT -53.885 225.595 -53.555 225.925 ;
        RECT -53.885 224.235 -53.555 224.565 ;
        RECT -53.885 222.875 -53.555 223.205 ;
        RECT -53.885 221.515 -53.555 221.845 ;
        RECT -53.885 220.155 -53.555 220.485 ;
        RECT -53.885 218.795 -53.555 219.125 ;
        RECT -53.885 217.435 -53.555 217.765 ;
        RECT -53.885 216.075 -53.555 216.405 ;
        RECT -53.885 214.715 -53.555 215.045 ;
        RECT -53.885 213.355 -53.555 213.685 ;
        RECT -53.885 211.995 -53.555 212.325 ;
        RECT -53.885 210.635 -53.555 210.965 ;
        RECT -53.885 209.275 -53.555 209.605 ;
        RECT -53.885 207.915 -53.555 208.245 ;
        RECT -53.885 206.555 -53.555 206.885 ;
        RECT -53.885 205.195 -53.555 205.525 ;
        RECT -53.885 203.835 -53.555 204.165 ;
        RECT -53.885 202.475 -53.555 202.805 ;
        RECT -53.885 201.115 -53.555 201.445 ;
        RECT -53.885 199.755 -53.555 200.085 ;
        RECT -53.885 198.395 -53.555 198.725 ;
        RECT -53.885 197.035 -53.555 197.365 ;
        RECT -53.885 195.675 -53.555 196.005 ;
        RECT -53.885 194.315 -53.555 194.645 ;
        RECT -53.885 192.955 -53.555 193.285 ;
        RECT -53.885 191.595 -53.555 191.925 ;
        RECT -53.885 190.235 -53.555 190.565 ;
        RECT -53.885 188.875 -53.555 189.205 ;
        RECT -53.885 187.515 -53.555 187.845 ;
        RECT -53.885 186.155 -53.555 186.485 ;
        RECT -53.885 184.795 -53.555 185.125 ;
        RECT -53.885 183.435 -53.555 183.765 ;
        RECT -53.885 182.075 -53.555 182.405 ;
        RECT -53.885 180.715 -53.555 181.045 ;
        RECT -53.885 179.355 -53.555 179.685 ;
        RECT -53.885 177.995 -53.555 178.325 ;
        RECT -53.885 176.635 -53.555 176.965 ;
        RECT -53.885 175.275 -53.555 175.605 ;
        RECT -53.885 173.915 -53.555 174.245 ;
        RECT -53.885 172.555 -53.555 172.885 ;
        RECT -53.885 171.195 -53.555 171.525 ;
        RECT -53.885 169.835 -53.555 170.165 ;
        RECT -53.885 168.475 -53.555 168.805 ;
        RECT -53.885 167.115 -53.555 167.445 ;
        RECT -53.885 165.755 -53.555 166.085 ;
        RECT -53.885 164.395 -53.555 164.725 ;
        RECT -53.885 163.035 -53.555 163.365 ;
        RECT -53.885 161.675 -53.555 162.005 ;
        RECT -53.885 160.315 -53.555 160.645 ;
        RECT -53.885 158.955 -53.555 159.285 ;
        RECT -53.885 157.595 -53.555 157.925 ;
        RECT -53.885 156.235 -53.555 156.565 ;
        RECT -53.885 154.875 -53.555 155.205 ;
        RECT -53.885 153.515 -53.555 153.845 ;
        RECT -53.885 152.155 -53.555 152.485 ;
        RECT -53.885 150.795 -53.555 151.125 ;
        RECT -53.885 149.435 -53.555 149.765 ;
        RECT -53.885 148.075 -53.555 148.405 ;
        RECT -53.885 146.715 -53.555 147.045 ;
        RECT -53.885 145.355 -53.555 145.685 ;
        RECT -53.885 143.995 -53.555 144.325 ;
        RECT -53.885 142.635 -53.555 142.965 ;
        RECT -53.885 141.275 -53.555 141.605 ;
        RECT -53.885 139.915 -53.555 140.245 ;
        RECT -53.885 138.555 -53.555 138.885 ;
        RECT -53.88 138.555 -53.56 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.885 97.755 -53.555 98.085 ;
        RECT -53.885 96.395 -53.555 96.725 ;
        RECT -53.885 95.035 -53.555 95.365 ;
        RECT -53.885 93.675 -53.555 94.005 ;
        RECT -53.885 92.315 -53.555 92.645 ;
        RECT -53.885 89.595 -53.555 89.925 ;
        RECT -53.885 88.235 -53.555 88.565 ;
        RECT -53.885 84.155 -53.555 84.485 ;
        RECT -53.885 82.795 -53.555 83.125 ;
        RECT -53.885 81.435 -53.555 81.765 ;
        RECT -53.885 80.075 -53.555 80.405 ;
        RECT -53.885 78.715 -53.555 79.045 ;
        RECT -53.885 77.355 -53.555 77.685 ;
        RECT -53.885 75.995 -53.555 76.325 ;
        RECT -53.885 74.635 -53.555 74.965 ;
        RECT -53.885 73.275 -53.555 73.605 ;
        RECT -53.885 71.915 -53.555 72.245 ;
        RECT -53.885 70.555 -53.555 70.885 ;
        RECT -53.885 69.195 -53.555 69.525 ;
        RECT -53.885 67.835 -53.555 68.165 ;
        RECT -53.885 66.475 -53.555 66.805 ;
        RECT -53.885 65.115 -53.555 65.445 ;
        RECT -53.885 63.755 -53.555 64.085 ;
        RECT -53.885 62.395 -53.555 62.725 ;
        RECT -53.885 61.035 -53.555 61.365 ;
        RECT -53.885 59.675 -53.555 60.005 ;
        RECT -53.885 58.315 -53.555 58.645 ;
        RECT -53.885 56.955 -53.555 57.285 ;
        RECT -53.885 55.595 -53.555 55.925 ;
        RECT -53.885 54.235 -53.555 54.565 ;
        RECT -53.885 52.875 -53.555 53.205 ;
        RECT -53.885 51.515 -53.555 51.845 ;
        RECT -53.885 50.155 -53.555 50.485 ;
        RECT -53.885 48.795 -53.555 49.125 ;
        RECT -53.885 47.435 -53.555 47.765 ;
        RECT -53.885 46.075 -53.555 46.405 ;
        RECT -53.885 44.715 -53.555 45.045 ;
        RECT -53.885 43.355 -53.555 43.685 ;
        RECT -53.885 41.995 -53.555 42.325 ;
        RECT -53.885 40.635 -53.555 40.965 ;
        RECT -53.885 39.275 -53.555 39.605 ;
        RECT -53.885 37.915 -53.555 38.245 ;
        RECT -53.885 36.555 -53.555 36.885 ;
        RECT -53.885 35.195 -53.555 35.525 ;
        RECT -53.885 33.835 -53.555 34.165 ;
        RECT -53.885 32.475 -53.555 32.805 ;
        RECT -53.885 31.115 -53.555 31.445 ;
        RECT -53.885 29.755 -53.555 30.085 ;
        RECT -53.885 28.395 -53.555 28.725 ;
        RECT -53.885 27.035 -53.555 27.365 ;
        RECT -53.885 25.675 -53.555 26.005 ;
        RECT -53.885 24.315 -53.555 24.645 ;
        RECT -53.885 22.955 -53.555 23.285 ;
        RECT -53.885 21.595 -53.555 21.925 ;
        RECT -53.885 20.235 -53.555 20.565 ;
        RECT -53.885 18.875 -53.555 19.205 ;
        RECT -53.885 17.515 -53.555 17.845 ;
        RECT -53.885 16.155 -53.555 16.485 ;
        RECT -53.885 14.795 -53.555 15.125 ;
        RECT -53.885 13.435 -53.555 13.765 ;
        RECT -53.885 12.075 -53.555 12.405 ;
        RECT -53.885 10.715 -53.555 11.045 ;
        RECT -53.885 9.355 -53.555 9.685 ;
        RECT -53.885 7.995 -53.555 8.325 ;
        RECT -53.885 6.635 -53.555 6.965 ;
        RECT -53.885 5.275 -53.555 5.605 ;
        RECT -53.885 3.915 -53.555 4.245 ;
        RECT -53.885 2.555 -53.555 2.885 ;
        RECT -53.885 1.195 -53.555 1.525 ;
        RECT -53.885 -0.165 -53.555 0.165 ;
        RECT -53.885 -2.885 -53.555 -2.555 ;
        RECT -53.885 -4.245 -53.555 -3.915 ;
        RECT -53.885 -5.605 -53.555 -5.275 ;
        RECT -53.885 -6.965 -53.555 -6.635 ;
        RECT -53.885 -8.325 -53.555 -7.995 ;
        RECT -53.885 -9.685 -53.555 -9.355 ;
        RECT -53.885 -11.045 -53.555 -10.715 ;
        RECT -53.885 -12.405 -53.555 -12.075 ;
        RECT -53.885 -13.765 -53.555 -13.435 ;
        RECT -53.885 -15.125 -53.555 -14.795 ;
        RECT -53.885 -16.485 -53.555 -16.155 ;
        RECT -53.885 -17.845 -53.555 -17.515 ;
        RECT -53.885 -19.205 -53.555 -18.875 ;
        RECT -53.885 -20.565 -53.555 -20.235 ;
        RECT -53.885 -21.925 -53.555 -21.595 ;
        RECT -53.885 -23.285 -53.555 -22.955 ;
        RECT -53.885 -24.645 -53.555 -24.315 ;
        RECT -53.885 -30.085 -53.555 -29.755 ;
        RECT -53.885 -31.445 -53.555 -31.115 ;
        RECT -53.885 -32.805 -53.555 -32.475 ;
        RECT -53.885 -34.165 -53.555 -33.835 ;
        RECT -53.885 -35.525 -53.555 -35.195 ;
        RECT -53.885 -36.885 -53.555 -36.555 ;
        RECT -53.885 -38.245 -53.555 -37.915 ;
        RECT -53.885 -39.605 -53.555 -39.275 ;
        RECT -53.885 -40.965 -53.555 -40.635 ;
        RECT -53.885 -42.325 -53.555 -41.995 ;
        RECT -53.885 -43.685 -53.555 -43.355 ;
        RECT -53.885 -45.045 -53.555 -44.715 ;
        RECT -53.885 -46.405 -53.555 -46.075 ;
        RECT -53.885 -47.765 -53.555 -47.435 ;
        RECT -53.885 -49.125 -53.555 -48.795 ;
        RECT -53.885 -50.485 -53.555 -50.155 ;
        RECT -53.885 -51.845 -53.555 -51.515 ;
        RECT -53.885 -53.205 -53.555 -52.875 ;
        RECT -53.885 -54.565 -53.555 -54.235 ;
        RECT -53.885 -55.925 -53.555 -55.595 ;
        RECT -53.885 -57.285 -53.555 -56.955 ;
        RECT -53.885 -58.645 -53.555 -58.315 ;
        RECT -53.885 -60.005 -53.555 -59.675 ;
        RECT -53.885 -61.365 -53.555 -61.035 ;
        RECT -53.885 -62.725 -53.555 -62.395 ;
        RECT -53.885 -64.085 -53.555 -63.755 ;
        RECT -53.885 -65.445 -53.555 -65.115 ;
        RECT -53.885 -68.165 -53.555 -67.835 ;
        RECT -53.885 -69.525 -53.555 -69.195 ;
        RECT -53.885 -70.885 -53.555 -70.555 ;
        RECT -53.885 -72.245 -53.555 -71.915 ;
        RECT -53.885 -73.605 -53.555 -73.275 ;
        RECT -53.885 -74.965 -53.555 -74.635 ;
        RECT -53.885 -76.325 -53.555 -75.995 ;
        RECT -53.885 -77.685 -53.555 -77.355 ;
        RECT -53.885 -79.045 -53.555 -78.715 ;
        RECT -53.885 -80.405 -53.555 -80.075 ;
        RECT -53.885 -81.765 -53.555 -81.435 ;
        RECT -53.885 -83.125 -53.555 -82.795 ;
        RECT -53.885 -84.485 -53.555 -84.155 ;
        RECT -53.885 -85.845 -53.555 -85.515 ;
        RECT -53.885 -87.205 -53.555 -86.875 ;
        RECT -53.885 -88.565 -53.555 -88.235 ;
        RECT -53.885 -89.925 -53.555 -89.595 ;
        RECT -53.885 -92.645 -53.555 -92.315 ;
        RECT -53.885 -94.005 -53.555 -93.675 ;
        RECT -53.885 -95.365 -53.555 -95.035 ;
        RECT -53.885 -96.725 -53.555 -96.395 ;
        RECT -53.885 -98.085 -53.555 -97.755 ;
        RECT -53.885 -99.69 -53.555 -99.36 ;
        RECT -53.885 -100.805 -53.555 -100.475 ;
        RECT -53.885 -103.525 -53.555 -103.195 ;
        RECT -53.885 -104.885 -53.555 -104.555 ;
        RECT -53.885 -106.245 -53.555 -105.915 ;
        RECT -53.885 -107.83 -53.555 -107.5 ;
        RECT -53.885 -108.965 -53.555 -108.635 ;
        RECT -53.885 -110.325 -53.555 -109.995 ;
        RECT -53.885 -111.685 -53.555 -111.355 ;
        RECT -53.88 -113.04 -53.56 98.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -53.885 -175.605 -53.555 -175.275 ;
        RECT -53.885 -178.325 -53.555 -177.995 ;
        RECT -53.885 -179.685 -53.555 -179.355 ;
        RECT -53.885 -181.93 -53.555 -180.8 ;
        RECT -53.88 -182.045 -53.56 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.525 241.32 -52.195 242.45 ;
        RECT -52.525 239.195 -52.195 239.525 ;
        RECT -52.525 237.835 -52.195 238.165 ;
        RECT -52.525 236.475 -52.195 236.805 ;
        RECT -52.525 235.115 -52.195 235.445 ;
        RECT -52.525 233.755 -52.195 234.085 ;
        RECT -52.525 232.395 -52.195 232.725 ;
        RECT -52.525 231.035 -52.195 231.365 ;
        RECT -52.525 229.675 -52.195 230.005 ;
        RECT -52.525 228.315 -52.195 228.645 ;
        RECT -52.525 226.955 -52.195 227.285 ;
        RECT -52.525 225.595 -52.195 225.925 ;
        RECT -52.525 224.235 -52.195 224.565 ;
        RECT -52.525 222.875 -52.195 223.205 ;
        RECT -52.525 221.515 -52.195 221.845 ;
        RECT -52.525 220.155 -52.195 220.485 ;
        RECT -52.525 218.795 -52.195 219.125 ;
        RECT -52.525 217.435 -52.195 217.765 ;
        RECT -52.525 216.075 -52.195 216.405 ;
        RECT -52.525 214.715 -52.195 215.045 ;
        RECT -52.525 213.355 -52.195 213.685 ;
        RECT -52.525 211.995 -52.195 212.325 ;
        RECT -52.525 210.635 -52.195 210.965 ;
        RECT -52.525 209.275 -52.195 209.605 ;
        RECT -52.525 207.915 -52.195 208.245 ;
        RECT -52.525 206.555 -52.195 206.885 ;
        RECT -52.525 205.195 -52.195 205.525 ;
        RECT -52.525 203.835 -52.195 204.165 ;
        RECT -52.525 202.475 -52.195 202.805 ;
        RECT -52.525 201.115 -52.195 201.445 ;
        RECT -52.525 199.755 -52.195 200.085 ;
        RECT -52.525 198.395 -52.195 198.725 ;
        RECT -52.525 197.035 -52.195 197.365 ;
        RECT -52.525 195.675 -52.195 196.005 ;
        RECT -52.525 194.315 -52.195 194.645 ;
        RECT -52.525 192.955 -52.195 193.285 ;
        RECT -52.525 191.595 -52.195 191.925 ;
        RECT -52.525 190.235 -52.195 190.565 ;
        RECT -52.525 188.875 -52.195 189.205 ;
        RECT -52.525 187.515 -52.195 187.845 ;
        RECT -52.525 186.155 -52.195 186.485 ;
        RECT -52.525 184.795 -52.195 185.125 ;
        RECT -52.525 183.435 -52.195 183.765 ;
        RECT -52.525 182.075 -52.195 182.405 ;
        RECT -52.525 180.715 -52.195 181.045 ;
        RECT -52.525 179.355 -52.195 179.685 ;
        RECT -52.525 177.995 -52.195 178.325 ;
        RECT -52.525 176.635 -52.195 176.965 ;
        RECT -52.525 175.275 -52.195 175.605 ;
        RECT -52.525 173.915 -52.195 174.245 ;
        RECT -52.525 172.555 -52.195 172.885 ;
        RECT -52.525 171.195 -52.195 171.525 ;
        RECT -52.525 169.835 -52.195 170.165 ;
        RECT -52.525 168.475 -52.195 168.805 ;
        RECT -52.525 167.115 -52.195 167.445 ;
        RECT -52.525 165.755 -52.195 166.085 ;
        RECT -52.525 164.395 -52.195 164.725 ;
        RECT -52.525 163.035 -52.195 163.365 ;
        RECT -52.525 161.675 -52.195 162.005 ;
        RECT -52.525 160.315 -52.195 160.645 ;
        RECT -52.525 158.955 -52.195 159.285 ;
        RECT -52.525 157.595 -52.195 157.925 ;
        RECT -52.525 156.235 -52.195 156.565 ;
        RECT -52.525 154.875 -52.195 155.205 ;
        RECT -52.525 153.515 -52.195 153.845 ;
        RECT -52.525 152.155 -52.195 152.485 ;
        RECT -52.525 150.795 -52.195 151.125 ;
        RECT -52.525 149.435 -52.195 149.765 ;
        RECT -52.525 148.075 -52.195 148.405 ;
        RECT -52.525 146.715 -52.195 147.045 ;
        RECT -52.525 145.355 -52.195 145.685 ;
        RECT -52.525 143.995 -52.195 144.325 ;
        RECT -52.525 142.635 -52.195 142.965 ;
        RECT -52.525 141.275 -52.195 141.605 ;
        RECT -52.525 139.915 -52.195 140.245 ;
        RECT -52.525 138.555 -52.195 138.885 ;
        RECT -52.525 137.225 -52.195 137.555 ;
        RECT -52.525 135.175 -52.195 135.505 ;
        RECT -52.525 132.815 -52.195 133.145 ;
        RECT -52.525 131.665 -52.195 131.995 ;
        RECT -52.525 129.655 -52.195 129.985 ;
        RECT -52.525 128.505 -52.195 128.835 ;
        RECT -52.525 126.495 -52.195 126.825 ;
        RECT -52.525 125.345 -52.195 125.675 ;
        RECT -52.525 123.335 -52.195 123.665 ;
        RECT -52.525 122.185 -52.195 122.515 ;
        RECT -52.525 120.175 -52.195 120.505 ;
        RECT -52.525 119.025 -52.195 119.355 ;
        RECT -52.52 117.48 -52.2 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -52.525 -121.205 -52.195 -120.875 ;
        RECT -52.525 -123.925 -52.195 -123.595 ;
        RECT -52.525 -125.285 -52.195 -124.955 ;
        RECT -52.525 -126.645 -52.195 -126.315 ;
        RECT -52.525 -128.005 -52.195 -127.675 ;
        RECT -52.525 -129.365 -52.195 -129.035 ;
        RECT -52.525 -130.725 -52.195 -130.395 ;
        RECT -52.525 -132.085 -52.195 -131.755 ;
        RECT -52.525 -133.445 -52.195 -133.115 ;
        RECT -52.525 -134.805 -52.195 -134.475 ;
        RECT -52.525 -136.165 -52.195 -135.835 ;
        RECT -52.525 -137.525 -52.195 -137.195 ;
        RECT -52.525 -138.885 -52.195 -138.555 ;
        RECT -52.525 -140.245 -52.195 -139.915 ;
        RECT -52.525 -141.605 -52.195 -141.275 ;
        RECT -52.525 -142.965 -52.195 -142.635 ;
        RECT -52.525 -144.325 -52.195 -143.995 ;
        RECT -52.525 -145.685 -52.195 -145.355 ;
        RECT -52.525 -147.045 -52.195 -146.715 ;
        RECT -52.525 -148.405 -52.195 -148.075 ;
        RECT -52.525 -149.765 -52.195 -149.435 ;
        RECT -52.525 -151.125 -52.195 -150.795 ;
        RECT -52.525 -152.485 -52.195 -152.155 ;
        RECT -52.525 -153.845 -52.195 -153.515 ;
        RECT -52.525 -155.205 -52.195 -154.875 ;
        RECT -52.525 -156.565 -52.195 -156.235 ;
        RECT -52.525 -157.925 -52.195 -157.595 ;
        RECT -52.525 -159.285 -52.195 -158.955 ;
        RECT -52.525 -160.645 -52.195 -160.315 ;
        RECT -52.525 -162.005 -52.195 -161.675 ;
        RECT -52.525 -163.365 -52.195 -163.035 ;
        RECT -52.525 -164.725 -52.195 -164.395 ;
        RECT -52.525 -166.085 -52.195 -165.755 ;
        RECT -52.525 -167.445 -52.195 -167.115 ;
        RECT -52.525 -168.805 -52.195 -168.475 ;
        RECT -52.525 -171.525 -52.195 -171.195 ;
        RECT -52.525 -172.885 -52.195 -172.555 ;
        RECT -52.52 -172.885 -52.2 -120.2 ;
    END
    PORT
      LAYER met3 ;
        RECT -51.165 135.175 -50.835 135.505 ;
        RECT -51.165 132.815 -50.835 133.145 ;
        RECT -51.165 131.665 -50.835 131.995 ;
        RECT -51.165 129.655 -50.835 129.985 ;
        RECT -51.165 128.505 -50.835 128.835 ;
        RECT -51.165 126.495 -50.835 126.825 ;
        RECT -51.165 125.345 -50.835 125.675 ;
        RECT -51.165 123.335 -50.835 123.665 ;
        RECT -51.165 122.185 -50.835 122.515 ;
        RECT -51.165 120.175 -50.835 120.505 ;
        RECT -51.165 119.025 -50.835 119.355 ;
        RECT -51.165 117.185 -50.835 117.515 ;
        RECT -51.165 115.865 -50.835 116.195 ;
        RECT -51.165 113.855 -50.835 114.185 ;
        RECT -51.165 112.705 -50.835 113.035 ;
        RECT -51.165 110.695 -50.835 111.025 ;
        RECT -51.165 109.545 -50.835 109.875 ;
        RECT -51.165 107.535 -50.835 107.865 ;
        RECT -51.165 106.385 -50.835 106.715 ;
        RECT -51.165 104.375 -50.835 104.705 ;
        RECT -51.165 103.225 -50.835 103.555 ;
        RECT -51.165 100.865 -50.835 101.195 ;
        RECT -51.165 98.81 -50.835 99.14 ;
        RECT -51.165 97.755 -50.835 98.085 ;
        RECT -51.165 96.395 -50.835 96.725 ;
        RECT -51.165 95.035 -50.835 95.365 ;
        RECT -51.165 93.675 -50.835 94.005 ;
        RECT -51.165 92.315 -50.835 92.645 ;
        RECT -51.165 90.955 -50.835 91.285 ;
        RECT -51.165 89.595 -50.835 89.925 ;
        RECT -51.165 88.235 -50.835 88.565 ;
        RECT -51.165 86.875 -50.835 87.205 ;
        RECT -51.165 85.515 -50.835 85.845 ;
        RECT -51.165 84.155 -50.835 84.485 ;
        RECT -51.165 82.795 -50.835 83.125 ;
        RECT -51.165 81.435 -50.835 81.765 ;
        RECT -51.165 80.075 -50.835 80.405 ;
        RECT -51.165 78.715 -50.835 79.045 ;
        RECT -51.165 77.355 -50.835 77.685 ;
        RECT -51.165 75.995 -50.835 76.325 ;
        RECT -51.165 74.635 -50.835 74.965 ;
        RECT -51.165 73.275 -50.835 73.605 ;
        RECT -51.165 71.915 -50.835 72.245 ;
        RECT -51.165 70.555 -50.835 70.885 ;
        RECT -51.165 69.195 -50.835 69.525 ;
        RECT -51.165 67.835 -50.835 68.165 ;
        RECT -51.165 66.475 -50.835 66.805 ;
        RECT -51.165 65.115 -50.835 65.445 ;
        RECT -51.165 63.755 -50.835 64.085 ;
        RECT -51.165 62.395 -50.835 62.725 ;
        RECT -51.165 61.035 -50.835 61.365 ;
        RECT -51.165 59.675 -50.835 60.005 ;
        RECT -51.165 58.315 -50.835 58.645 ;
        RECT -51.165 56.955 -50.835 57.285 ;
        RECT -51.165 55.595 -50.835 55.925 ;
        RECT -51.165 54.235 -50.835 54.565 ;
        RECT -51.165 52.875 -50.835 53.205 ;
        RECT -51.165 51.515 -50.835 51.845 ;
        RECT -51.165 50.155 -50.835 50.485 ;
        RECT -51.165 48.795 -50.835 49.125 ;
        RECT -51.165 47.435 -50.835 47.765 ;
        RECT -51.165 46.075 -50.835 46.405 ;
        RECT -51.165 44.715 -50.835 45.045 ;
        RECT -51.165 43.355 -50.835 43.685 ;
        RECT -51.165 41.995 -50.835 42.325 ;
        RECT -51.165 40.635 -50.835 40.965 ;
        RECT -51.165 39.275 -50.835 39.605 ;
        RECT -51.165 37.915 -50.835 38.245 ;
        RECT -51.165 36.555 -50.835 36.885 ;
        RECT -51.165 35.195 -50.835 35.525 ;
        RECT -51.165 33.835 -50.835 34.165 ;
        RECT -51.165 32.475 -50.835 32.805 ;
        RECT -51.165 31.115 -50.835 31.445 ;
        RECT -51.165 29.755 -50.835 30.085 ;
        RECT -51.165 28.395 -50.835 28.725 ;
        RECT -51.165 27.035 -50.835 27.365 ;
        RECT -51.165 25.675 -50.835 26.005 ;
        RECT -51.165 24.315 -50.835 24.645 ;
        RECT -51.165 22.955 -50.835 23.285 ;
        RECT -51.165 21.595 -50.835 21.925 ;
        RECT -51.165 20.235 -50.835 20.565 ;
        RECT -51.165 18.875 -50.835 19.205 ;
        RECT -51.165 17.515 -50.835 17.845 ;
        RECT -51.165 16.155 -50.835 16.485 ;
        RECT -51.165 14.795 -50.835 15.125 ;
        RECT -51.165 13.435 -50.835 13.765 ;
        RECT -51.165 12.075 -50.835 12.405 ;
        RECT -51.165 10.715 -50.835 11.045 ;
        RECT -51.165 9.355 -50.835 9.685 ;
        RECT -51.165 7.995 -50.835 8.325 ;
        RECT -51.165 6.635 -50.835 6.965 ;
        RECT -51.165 5.275 -50.835 5.605 ;
        RECT -51.165 3.915 -50.835 4.245 ;
        RECT -51.165 2.555 -50.835 2.885 ;
        RECT -51.165 1.195 -50.835 1.525 ;
        RECT -51.165 -0.165 -50.835 0.165 ;
        RECT -51.165 -2.885 -50.835 -2.555 ;
        RECT -51.165 -4.245 -50.835 -3.915 ;
        RECT -51.165 -5.605 -50.835 -5.275 ;
        RECT -51.165 -6.965 -50.835 -6.635 ;
        RECT -51.165 -8.325 -50.835 -7.995 ;
        RECT -51.165 -9.685 -50.835 -9.355 ;
        RECT -51.165 -11.045 -50.835 -10.715 ;
        RECT -51.165 -12.405 -50.835 -12.075 ;
        RECT -51.165 -13.765 -50.835 -13.435 ;
        RECT -51.165 -15.125 -50.835 -14.795 ;
        RECT -51.165 -16.485 -50.835 -16.155 ;
        RECT -51.165 -17.845 -50.835 -17.515 ;
        RECT -51.165 -19.205 -50.835 -18.875 ;
        RECT -51.165 -20.565 -50.835 -20.235 ;
        RECT -51.165 -21.925 -50.835 -21.595 ;
        RECT -51.165 -23.285 -50.835 -22.955 ;
        RECT -51.165 -24.645 -50.835 -24.315 ;
        RECT -51.165 -30.085 -50.835 -29.755 ;
        RECT -51.165 -31.445 -50.835 -31.115 ;
        RECT -51.165 -32.805 -50.835 -32.475 ;
        RECT -51.165 -34.165 -50.835 -33.835 ;
        RECT -51.165 -35.525 -50.835 -35.195 ;
        RECT -51.165 -36.885 -50.835 -36.555 ;
        RECT -51.165 -38.245 -50.835 -37.915 ;
        RECT -51.165 -39.605 -50.835 -39.275 ;
        RECT -51.165 -40.965 -50.835 -40.635 ;
        RECT -51.165 -42.325 -50.835 -41.995 ;
        RECT -51.165 -43.685 -50.835 -43.355 ;
        RECT -51.165 -45.045 -50.835 -44.715 ;
        RECT -51.165 -46.405 -50.835 -46.075 ;
        RECT -51.165 -47.765 -50.835 -47.435 ;
        RECT -51.165 -49.125 -50.835 -48.795 ;
        RECT -51.165 -50.485 -50.835 -50.155 ;
        RECT -51.165 -51.845 -50.835 -51.515 ;
        RECT -51.165 -53.205 -50.835 -52.875 ;
        RECT -51.165 -54.565 -50.835 -54.235 ;
        RECT -51.165 -55.925 -50.835 -55.595 ;
        RECT -51.165 -57.285 -50.835 -56.955 ;
        RECT -51.165 -58.645 -50.835 -58.315 ;
        RECT -51.165 -60.005 -50.835 -59.675 ;
        RECT -51.165 -61.365 -50.835 -61.035 ;
        RECT -51.165 -62.725 -50.835 -62.395 ;
        RECT -51.165 -64.085 -50.835 -63.755 ;
        RECT -51.165 -65.445 -50.835 -65.115 ;
        RECT -51.165 -68.165 -50.835 -67.835 ;
        RECT -51.165 -69.525 -50.835 -69.195 ;
        RECT -51.165 -70.885 -50.835 -70.555 ;
        RECT -51.165 -72.245 -50.835 -71.915 ;
        RECT -51.165 -73.605 -50.835 -73.275 ;
        RECT -51.165 -74.965 -50.835 -74.635 ;
        RECT -51.165 -76.325 -50.835 -75.995 ;
        RECT -51.165 -77.685 -50.835 -77.355 ;
        RECT -51.165 -79.045 -50.835 -78.715 ;
        RECT -51.165 -80.405 -50.835 -80.075 ;
        RECT -51.165 -81.765 -50.835 -81.435 ;
        RECT -51.165 -83.125 -50.835 -82.795 ;
        RECT -51.165 -84.485 -50.835 -84.155 ;
        RECT -51.165 -85.845 -50.835 -85.515 ;
        RECT -51.165 -87.205 -50.835 -86.875 ;
        RECT -51.165 -88.565 -50.835 -88.235 ;
        RECT -51.165 -89.925 -50.835 -89.595 ;
        RECT -51.165 -92.645 -50.835 -92.315 ;
        RECT -51.165 -94.005 -50.835 -93.675 ;
        RECT -51.165 -95.365 -50.835 -95.035 ;
        RECT -51.165 -96.725 -50.835 -96.395 ;
        RECT -51.165 -98.085 -50.835 -97.755 ;
        RECT -51.165 -99.69 -50.835 -99.36 ;
        RECT -51.165 -100.805 -50.835 -100.475 ;
        RECT -51.165 -103.525 -50.835 -103.195 ;
        RECT -51.165 -104.885 -50.835 -104.555 ;
        RECT -51.165 -106.245 -50.835 -105.915 ;
        RECT -51.165 -107.83 -50.835 -107.5 ;
        RECT -51.165 -108.965 -50.835 -108.635 ;
        RECT -51.165 -110.325 -50.835 -109.995 ;
        RECT -51.165 -111.685 -50.835 -111.355 ;
        RECT -51.165 -114.405 -50.835 -114.075 ;
        RECT -51.165 -115.765 -50.835 -115.435 ;
        RECT -51.165 -117.125 -50.835 -116.795 ;
        RECT -51.165 -118.485 -50.835 -118.155 ;
        RECT -51.165 -121.205 -50.835 -120.875 ;
        RECT -51.165 -123.925 -50.835 -123.595 ;
        RECT -51.165 -125.285 -50.835 -124.955 ;
        RECT -51.165 -126.645 -50.835 -126.315 ;
        RECT -51.165 -128.005 -50.835 -127.675 ;
        RECT -51.165 -129.365 -50.835 -129.035 ;
        RECT -51.165 -130.725 -50.835 -130.395 ;
        RECT -51.165 -132.085 -50.835 -131.755 ;
        RECT -51.165 -133.445 -50.835 -133.115 ;
        RECT -51.165 -134.805 -50.835 -134.475 ;
        RECT -51.165 -136.165 -50.835 -135.835 ;
        RECT -51.165 -137.525 -50.835 -137.195 ;
        RECT -51.165 -138.885 -50.835 -138.555 ;
        RECT -51.165 -140.245 -50.835 -139.915 ;
        RECT -51.165 -141.605 -50.835 -141.275 ;
        RECT -51.165 -142.965 -50.835 -142.635 ;
        RECT -51.165 -144.325 -50.835 -143.995 ;
        RECT -51.165 -145.685 -50.835 -145.355 ;
        RECT -51.165 -147.045 -50.835 -146.715 ;
        RECT -51.165 -148.405 -50.835 -148.075 ;
        RECT -51.165 -149.765 -50.835 -149.435 ;
        RECT -51.165 -151.125 -50.835 -150.795 ;
        RECT -51.165 -152.485 -50.835 -152.155 ;
        RECT -51.165 -153.845 -50.835 -153.515 ;
        RECT -51.165 -155.205 -50.835 -154.875 ;
        RECT -51.165 -156.565 -50.835 -156.235 ;
        RECT -51.165 -157.925 -50.835 -157.595 ;
        RECT -51.165 -159.285 -50.835 -158.955 ;
        RECT -51.165 -160.645 -50.835 -160.315 ;
        RECT -51.165 -162.005 -50.835 -161.675 ;
        RECT -51.165 -163.365 -50.835 -163.035 ;
        RECT -51.165 -164.725 -50.835 -164.395 ;
        RECT -51.165 -166.085 -50.835 -165.755 ;
        RECT -51.165 -167.445 -50.835 -167.115 ;
        RECT -51.16 -167.445 -50.84 242.565 ;
        RECT -51.165 241.32 -50.835 242.45 ;
        RECT -51.165 239.195 -50.835 239.525 ;
        RECT -51.165 237.835 -50.835 238.165 ;
        RECT -51.165 236.475 -50.835 236.805 ;
        RECT -51.165 235.115 -50.835 235.445 ;
        RECT -51.165 233.755 -50.835 234.085 ;
        RECT -51.165 232.395 -50.835 232.725 ;
        RECT -51.165 231.035 -50.835 231.365 ;
        RECT -51.165 229.675 -50.835 230.005 ;
        RECT -51.165 228.315 -50.835 228.645 ;
        RECT -51.165 226.955 -50.835 227.285 ;
        RECT -51.165 225.595 -50.835 225.925 ;
        RECT -51.165 224.235 -50.835 224.565 ;
        RECT -51.165 222.875 -50.835 223.205 ;
        RECT -51.165 221.515 -50.835 221.845 ;
        RECT -51.165 220.155 -50.835 220.485 ;
        RECT -51.165 218.795 -50.835 219.125 ;
        RECT -51.165 217.435 -50.835 217.765 ;
        RECT -51.165 216.075 -50.835 216.405 ;
        RECT -51.165 214.715 -50.835 215.045 ;
        RECT -51.165 213.355 -50.835 213.685 ;
        RECT -51.165 211.995 -50.835 212.325 ;
        RECT -51.165 210.635 -50.835 210.965 ;
        RECT -51.165 209.275 -50.835 209.605 ;
        RECT -51.165 207.915 -50.835 208.245 ;
        RECT -51.165 206.555 -50.835 206.885 ;
        RECT -51.165 205.195 -50.835 205.525 ;
        RECT -51.165 203.835 -50.835 204.165 ;
        RECT -51.165 202.475 -50.835 202.805 ;
        RECT -51.165 201.115 -50.835 201.445 ;
        RECT -51.165 199.755 -50.835 200.085 ;
        RECT -51.165 198.395 -50.835 198.725 ;
        RECT -51.165 197.035 -50.835 197.365 ;
        RECT -51.165 195.675 -50.835 196.005 ;
        RECT -51.165 194.315 -50.835 194.645 ;
        RECT -51.165 192.955 -50.835 193.285 ;
        RECT -51.165 191.595 -50.835 191.925 ;
        RECT -51.165 190.235 -50.835 190.565 ;
        RECT -51.165 188.875 -50.835 189.205 ;
        RECT -51.165 187.515 -50.835 187.845 ;
        RECT -51.165 186.155 -50.835 186.485 ;
        RECT -51.165 184.795 -50.835 185.125 ;
        RECT -51.165 183.435 -50.835 183.765 ;
        RECT -51.165 182.075 -50.835 182.405 ;
        RECT -51.165 180.715 -50.835 181.045 ;
        RECT -51.165 179.355 -50.835 179.685 ;
        RECT -51.165 177.995 -50.835 178.325 ;
        RECT -51.165 176.635 -50.835 176.965 ;
        RECT -51.165 175.275 -50.835 175.605 ;
        RECT -51.165 173.915 -50.835 174.245 ;
        RECT -51.165 172.555 -50.835 172.885 ;
        RECT -51.165 171.195 -50.835 171.525 ;
        RECT -51.165 169.835 -50.835 170.165 ;
        RECT -51.165 168.475 -50.835 168.805 ;
        RECT -51.165 167.115 -50.835 167.445 ;
        RECT -51.165 165.755 -50.835 166.085 ;
        RECT -51.165 164.395 -50.835 164.725 ;
        RECT -51.165 163.035 -50.835 163.365 ;
        RECT -51.165 161.675 -50.835 162.005 ;
        RECT -51.165 160.315 -50.835 160.645 ;
        RECT -51.165 158.955 -50.835 159.285 ;
        RECT -51.165 157.595 -50.835 157.925 ;
        RECT -51.165 156.235 -50.835 156.565 ;
        RECT -51.165 154.875 -50.835 155.205 ;
        RECT -51.165 153.515 -50.835 153.845 ;
        RECT -51.165 152.155 -50.835 152.485 ;
        RECT -51.165 150.795 -50.835 151.125 ;
        RECT -51.165 149.435 -50.835 149.765 ;
        RECT -51.165 148.075 -50.835 148.405 ;
        RECT -51.165 146.715 -50.835 147.045 ;
        RECT -51.165 145.355 -50.835 145.685 ;
        RECT -51.165 143.995 -50.835 144.325 ;
        RECT -51.165 142.635 -50.835 142.965 ;
        RECT -51.165 141.275 -50.835 141.605 ;
        RECT -51.165 139.915 -50.835 140.245 ;
        RECT -51.165 138.555 -50.835 138.885 ;
        RECT -51.165 137.225 -50.835 137.555 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.685 241.32 -60.355 242.45 ;
        RECT -60.685 239.195 -60.355 239.525 ;
        RECT -60.685 237.835 -60.355 238.165 ;
        RECT -60.685 236.475 -60.355 236.805 ;
        RECT -60.685 235.115 -60.355 235.445 ;
        RECT -60.685 233.755 -60.355 234.085 ;
        RECT -60.685 232.395 -60.355 232.725 ;
        RECT -60.685 231.035 -60.355 231.365 ;
        RECT -60.685 229.675 -60.355 230.005 ;
        RECT -60.685 228.315 -60.355 228.645 ;
        RECT -60.685 226.955 -60.355 227.285 ;
        RECT -60.685 225.595 -60.355 225.925 ;
        RECT -60.685 224.235 -60.355 224.565 ;
        RECT -60.685 222.875 -60.355 223.205 ;
        RECT -60.685 221.515 -60.355 221.845 ;
        RECT -60.685 220.155 -60.355 220.485 ;
        RECT -60.685 218.795 -60.355 219.125 ;
        RECT -60.685 217.435 -60.355 217.765 ;
        RECT -60.685 216.075 -60.355 216.405 ;
        RECT -60.685 214.715 -60.355 215.045 ;
        RECT -60.685 213.355 -60.355 213.685 ;
        RECT -60.685 211.995 -60.355 212.325 ;
        RECT -60.685 210.635 -60.355 210.965 ;
        RECT -60.685 209.275 -60.355 209.605 ;
        RECT -60.685 207.915 -60.355 208.245 ;
        RECT -60.685 206.555 -60.355 206.885 ;
        RECT -60.685 205.195 -60.355 205.525 ;
        RECT -60.685 203.835 -60.355 204.165 ;
        RECT -60.685 202.475 -60.355 202.805 ;
        RECT -60.685 201.115 -60.355 201.445 ;
        RECT -60.685 199.755 -60.355 200.085 ;
        RECT -60.685 198.395 -60.355 198.725 ;
        RECT -60.685 197.035 -60.355 197.365 ;
        RECT -60.685 195.675 -60.355 196.005 ;
        RECT -60.685 194.315 -60.355 194.645 ;
        RECT -60.685 192.955 -60.355 193.285 ;
        RECT -60.685 191.595 -60.355 191.925 ;
        RECT -60.685 190.235 -60.355 190.565 ;
        RECT -60.685 188.875 -60.355 189.205 ;
        RECT -60.685 187.515 -60.355 187.845 ;
        RECT -60.685 186.155 -60.355 186.485 ;
        RECT -60.685 184.795 -60.355 185.125 ;
        RECT -60.685 183.435 -60.355 183.765 ;
        RECT -60.685 182.075 -60.355 182.405 ;
        RECT -60.685 180.715 -60.355 181.045 ;
        RECT -60.685 179.355 -60.355 179.685 ;
        RECT -60.685 177.995 -60.355 178.325 ;
        RECT -60.685 176.635 -60.355 176.965 ;
        RECT -60.685 175.275 -60.355 175.605 ;
        RECT -60.685 173.915 -60.355 174.245 ;
        RECT -60.685 172.555 -60.355 172.885 ;
        RECT -60.685 171.195 -60.355 171.525 ;
        RECT -60.685 169.835 -60.355 170.165 ;
        RECT -60.685 168.475 -60.355 168.805 ;
        RECT -60.685 167.115 -60.355 167.445 ;
        RECT -60.685 165.755 -60.355 166.085 ;
        RECT -60.685 164.395 -60.355 164.725 ;
        RECT -60.685 163.035 -60.355 163.365 ;
        RECT -60.685 161.675 -60.355 162.005 ;
        RECT -60.685 160.315 -60.355 160.645 ;
        RECT -60.685 158.955 -60.355 159.285 ;
        RECT -60.685 157.595 -60.355 157.925 ;
        RECT -60.685 156.235 -60.355 156.565 ;
        RECT -60.685 154.875 -60.355 155.205 ;
        RECT -60.685 153.515 -60.355 153.845 ;
        RECT -60.685 152.155 -60.355 152.485 ;
        RECT -60.685 150.795 -60.355 151.125 ;
        RECT -60.685 149.435 -60.355 149.765 ;
        RECT -60.685 148.075 -60.355 148.405 ;
        RECT -60.685 146.715 -60.355 147.045 ;
        RECT -60.685 145.355 -60.355 145.685 ;
        RECT -60.685 143.995 -60.355 144.325 ;
        RECT -60.685 142.635 -60.355 142.965 ;
        RECT -60.685 141.275 -60.355 141.605 ;
        RECT -60.685 139.915 -60.355 140.245 ;
        RECT -60.685 138.555 -60.355 138.885 ;
        RECT -60.685 137.225 -60.355 137.555 ;
        RECT -60.685 135.175 -60.355 135.505 ;
        RECT -60.685 132.815 -60.355 133.145 ;
        RECT -60.685 131.665 -60.355 131.995 ;
        RECT -60.685 129.655 -60.355 129.985 ;
        RECT -60.685 128.505 -60.355 128.835 ;
        RECT -60.685 126.495 -60.355 126.825 ;
        RECT -60.685 125.345 -60.355 125.675 ;
        RECT -60.685 123.335 -60.355 123.665 ;
        RECT -60.685 122.185 -60.355 122.515 ;
        RECT -60.685 120.175 -60.355 120.505 ;
        RECT -60.685 119.025 -60.355 119.355 ;
        RECT -60.685 117.185 -60.355 117.515 ;
        RECT -60.685 115.865 -60.355 116.195 ;
        RECT -60.685 113.855 -60.355 114.185 ;
        RECT -60.685 112.705 -60.355 113.035 ;
        RECT -60.685 110.695 -60.355 111.025 ;
        RECT -60.685 109.545 -60.355 109.875 ;
        RECT -60.685 107.535 -60.355 107.865 ;
        RECT -60.685 106.385 -60.355 106.715 ;
        RECT -60.685 104.375 -60.355 104.705 ;
        RECT -60.685 103.225 -60.355 103.555 ;
        RECT -60.685 100.865 -60.355 101.195 ;
        RECT -60.685 98.81 -60.355 99.14 ;
        RECT -60.685 97.755 -60.355 98.085 ;
        RECT -60.685 96.395 -60.355 96.725 ;
        RECT -60.685 95.035 -60.355 95.365 ;
        RECT -60.685 93.675 -60.355 94.005 ;
        RECT -60.685 92.315 -60.355 92.645 ;
        RECT -60.685 90.955 -60.355 91.285 ;
        RECT -60.685 89.595 -60.355 89.925 ;
        RECT -60.685 88.235 -60.355 88.565 ;
        RECT -60.685 86.875 -60.355 87.205 ;
        RECT -60.685 85.515 -60.355 85.845 ;
        RECT -60.685 84.155 -60.355 84.485 ;
        RECT -60.685 82.795 -60.355 83.125 ;
        RECT -60.685 81.435 -60.355 81.765 ;
        RECT -60.685 80.075 -60.355 80.405 ;
        RECT -60.685 78.715 -60.355 79.045 ;
        RECT -60.685 77.355 -60.355 77.685 ;
        RECT -60.685 75.995 -60.355 76.325 ;
        RECT -60.685 74.635 -60.355 74.965 ;
        RECT -60.685 73.275 -60.355 73.605 ;
        RECT -60.685 71.915 -60.355 72.245 ;
        RECT -60.685 70.555 -60.355 70.885 ;
        RECT -60.685 69.195 -60.355 69.525 ;
        RECT -60.685 67.835 -60.355 68.165 ;
        RECT -60.685 66.475 -60.355 66.805 ;
        RECT -60.685 65.115 -60.355 65.445 ;
        RECT -60.685 63.755 -60.355 64.085 ;
        RECT -60.685 62.395 -60.355 62.725 ;
        RECT -60.685 61.035 -60.355 61.365 ;
        RECT -60.685 59.675 -60.355 60.005 ;
        RECT -60.685 58.315 -60.355 58.645 ;
        RECT -60.685 56.955 -60.355 57.285 ;
        RECT -60.685 55.595 -60.355 55.925 ;
        RECT -60.685 54.235 -60.355 54.565 ;
        RECT -60.685 52.875 -60.355 53.205 ;
        RECT -60.685 51.515 -60.355 51.845 ;
        RECT -60.685 50.155 -60.355 50.485 ;
        RECT -60.685 48.795 -60.355 49.125 ;
        RECT -60.685 47.435 -60.355 47.765 ;
        RECT -60.685 46.075 -60.355 46.405 ;
        RECT -60.685 44.715 -60.355 45.045 ;
        RECT -60.685 43.355 -60.355 43.685 ;
        RECT -60.685 41.995 -60.355 42.325 ;
        RECT -60.685 40.635 -60.355 40.965 ;
        RECT -60.685 39.275 -60.355 39.605 ;
        RECT -60.685 37.915 -60.355 38.245 ;
        RECT -60.685 36.555 -60.355 36.885 ;
        RECT -60.685 35.195 -60.355 35.525 ;
        RECT -60.685 33.835 -60.355 34.165 ;
        RECT -60.685 32.475 -60.355 32.805 ;
        RECT -60.685 31.115 -60.355 31.445 ;
        RECT -60.685 29.755 -60.355 30.085 ;
        RECT -60.685 28.395 -60.355 28.725 ;
        RECT -60.685 27.035 -60.355 27.365 ;
        RECT -60.685 25.675 -60.355 26.005 ;
        RECT -60.685 24.315 -60.355 24.645 ;
        RECT -60.685 22.955 -60.355 23.285 ;
        RECT -60.685 21.595 -60.355 21.925 ;
        RECT -60.685 20.235 -60.355 20.565 ;
        RECT -60.685 18.875 -60.355 19.205 ;
        RECT -60.685 17.515 -60.355 17.845 ;
        RECT -60.685 16.155 -60.355 16.485 ;
        RECT -60.685 14.795 -60.355 15.125 ;
        RECT -60.685 13.435 -60.355 13.765 ;
        RECT -60.685 12.075 -60.355 12.405 ;
        RECT -60.685 10.715 -60.355 11.045 ;
        RECT -60.685 9.355 -60.355 9.685 ;
        RECT -60.685 7.995 -60.355 8.325 ;
        RECT -60.685 6.635 -60.355 6.965 ;
        RECT -60.685 5.275 -60.355 5.605 ;
        RECT -60.685 3.915 -60.355 4.245 ;
        RECT -60.685 2.555 -60.355 2.885 ;
        RECT -60.685 1.195 -60.355 1.525 ;
        RECT -60.685 -0.165 -60.355 0.165 ;
        RECT -60.685 -1.525 -60.355 -1.195 ;
        RECT -60.685 -2.885 -60.355 -2.555 ;
        RECT -60.685 -4.245 -60.355 -3.915 ;
        RECT -60.685 -5.605 -60.355 -5.275 ;
        RECT -60.685 -6.965 -60.355 -6.635 ;
        RECT -60.685 -8.325 -60.355 -7.995 ;
        RECT -60.685 -9.685 -60.355 -9.355 ;
        RECT -60.685 -11.045 -60.355 -10.715 ;
        RECT -60.685 -12.405 -60.355 -12.075 ;
        RECT -60.685 -13.765 -60.355 -13.435 ;
        RECT -60.685 -15.125 -60.355 -14.795 ;
        RECT -60.685 -16.485 -60.355 -16.155 ;
        RECT -60.685 -17.845 -60.355 -17.515 ;
        RECT -60.685 -19.205 -60.355 -18.875 ;
        RECT -60.685 -20.565 -60.355 -20.235 ;
        RECT -60.685 -21.925 -60.355 -21.595 ;
        RECT -60.685 -23.285 -60.355 -22.955 ;
        RECT -60.685 -24.645 -60.355 -24.315 ;
        RECT -60.685 -28.725 -60.355 -28.395 ;
        RECT -60.685 -30.085 -60.355 -29.755 ;
        RECT -60.685 -31.445 -60.355 -31.115 ;
        RECT -60.685 -32.805 -60.355 -32.475 ;
        RECT -60.685 -34.165 -60.355 -33.835 ;
        RECT -60.685 -35.525 -60.355 -35.195 ;
        RECT -60.685 -36.885 -60.355 -36.555 ;
        RECT -60.685 -38.245 -60.355 -37.915 ;
        RECT -60.685 -39.605 -60.355 -39.275 ;
        RECT -60.685 -40.965 -60.355 -40.635 ;
        RECT -60.685 -42.325 -60.355 -41.995 ;
        RECT -60.685 -43.685 -60.355 -43.355 ;
        RECT -60.685 -45.045 -60.355 -44.715 ;
        RECT -60.685 -46.405 -60.355 -46.075 ;
        RECT -60.685 -47.765 -60.355 -47.435 ;
        RECT -60.685 -49.125 -60.355 -48.795 ;
        RECT -60.685 -50.485 -60.355 -50.155 ;
        RECT -60.685 -51.845 -60.355 -51.515 ;
        RECT -60.685 -53.205 -60.355 -52.875 ;
        RECT -60.685 -54.565 -60.355 -54.235 ;
        RECT -60.685 -55.925 -60.355 -55.595 ;
        RECT -60.685 -57.285 -60.355 -56.955 ;
        RECT -60.685 -58.645 -60.355 -58.315 ;
        RECT -60.685 -60.005 -60.355 -59.675 ;
        RECT -60.685 -61.365 -60.355 -61.035 ;
        RECT -60.685 -62.725 -60.355 -62.395 ;
        RECT -60.685 -64.085 -60.355 -63.755 ;
        RECT -60.685 -65.445 -60.355 -65.115 ;
        RECT -60.685 -66.805 -60.355 -66.475 ;
        RECT -60.685 -68.165 -60.355 -67.835 ;
        RECT -60.685 -69.525 -60.355 -69.195 ;
        RECT -60.685 -70.885 -60.355 -70.555 ;
        RECT -60.685 -72.245 -60.355 -71.915 ;
        RECT -60.685 -73.605 -60.355 -73.275 ;
        RECT -60.685 -74.965 -60.355 -74.635 ;
        RECT -60.685 -76.325 -60.355 -75.995 ;
        RECT -60.685 -77.685 -60.355 -77.355 ;
        RECT -60.685 -79.045 -60.355 -78.715 ;
        RECT -60.685 -80.405 -60.355 -80.075 ;
        RECT -60.685 -81.765 -60.355 -81.435 ;
        RECT -60.685 -83.125 -60.355 -82.795 ;
        RECT -60.685 -84.485 -60.355 -84.155 ;
        RECT -60.685 -85.845 -60.355 -85.515 ;
        RECT -60.685 -87.205 -60.355 -86.875 ;
        RECT -60.685 -88.565 -60.355 -88.235 ;
        RECT -60.685 -89.925 -60.355 -89.595 ;
        RECT -60.685 -92.645 -60.355 -92.315 ;
        RECT -60.685 -94.005 -60.355 -93.675 ;
        RECT -60.685 -95.365 -60.355 -95.035 ;
        RECT -60.685 -96.725 -60.355 -96.395 ;
        RECT -60.685 -98.085 -60.355 -97.755 ;
        RECT -60.685 -99.69 -60.355 -99.36 ;
        RECT -60.685 -100.805 -60.355 -100.475 ;
        RECT -60.685 -103.525 -60.355 -103.195 ;
        RECT -60.685 -104.885 -60.355 -104.555 ;
        RECT -60.685 -106.245 -60.355 -105.915 ;
        RECT -60.685 -107.83 -60.355 -107.5 ;
        RECT -60.685 -108.965 -60.355 -108.635 ;
        RECT -60.685 -110.325 -60.355 -109.995 ;
        RECT -60.685 -111.685 -60.355 -111.355 ;
        RECT -60.68 -113.72 -60.36 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -60.685 -175.605 -60.355 -175.275 ;
        RECT -60.685 -176.685 -60.355 -176.355 ;
        RECT -60.685 -178.325 -60.355 -177.995 ;
        RECT -60.685 -179.685 -60.355 -179.355 ;
        RECT -60.685 -181.93 -60.355 -180.8 ;
        RECT -60.68 -182.045 -60.36 -175.275 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.325 241.32 -58.995 242.45 ;
        RECT -59.325 239.195 -58.995 239.525 ;
        RECT -59.325 237.835 -58.995 238.165 ;
        RECT -59.325 236.475 -58.995 236.805 ;
        RECT -59.325 235.115 -58.995 235.445 ;
        RECT -59.325 233.755 -58.995 234.085 ;
        RECT -59.325 232.395 -58.995 232.725 ;
        RECT -59.325 231.035 -58.995 231.365 ;
        RECT -59.325 229.675 -58.995 230.005 ;
        RECT -59.325 228.315 -58.995 228.645 ;
        RECT -59.325 226.955 -58.995 227.285 ;
        RECT -59.325 225.595 -58.995 225.925 ;
        RECT -59.325 224.235 -58.995 224.565 ;
        RECT -59.325 222.875 -58.995 223.205 ;
        RECT -59.325 221.515 -58.995 221.845 ;
        RECT -59.325 220.155 -58.995 220.485 ;
        RECT -59.325 218.795 -58.995 219.125 ;
        RECT -59.325 217.435 -58.995 217.765 ;
        RECT -59.325 216.075 -58.995 216.405 ;
        RECT -59.325 214.715 -58.995 215.045 ;
        RECT -59.325 213.355 -58.995 213.685 ;
        RECT -59.325 211.995 -58.995 212.325 ;
        RECT -59.325 210.635 -58.995 210.965 ;
        RECT -59.325 209.275 -58.995 209.605 ;
        RECT -59.325 207.915 -58.995 208.245 ;
        RECT -59.325 206.555 -58.995 206.885 ;
        RECT -59.325 205.195 -58.995 205.525 ;
        RECT -59.325 203.835 -58.995 204.165 ;
        RECT -59.325 202.475 -58.995 202.805 ;
        RECT -59.325 201.115 -58.995 201.445 ;
        RECT -59.325 199.755 -58.995 200.085 ;
        RECT -59.325 198.395 -58.995 198.725 ;
        RECT -59.325 197.035 -58.995 197.365 ;
        RECT -59.325 195.675 -58.995 196.005 ;
        RECT -59.325 194.315 -58.995 194.645 ;
        RECT -59.325 192.955 -58.995 193.285 ;
        RECT -59.325 191.595 -58.995 191.925 ;
        RECT -59.325 190.235 -58.995 190.565 ;
        RECT -59.325 188.875 -58.995 189.205 ;
        RECT -59.325 187.515 -58.995 187.845 ;
        RECT -59.325 186.155 -58.995 186.485 ;
        RECT -59.325 184.795 -58.995 185.125 ;
        RECT -59.325 183.435 -58.995 183.765 ;
        RECT -59.325 182.075 -58.995 182.405 ;
        RECT -59.325 180.715 -58.995 181.045 ;
        RECT -59.325 179.355 -58.995 179.685 ;
        RECT -59.325 177.995 -58.995 178.325 ;
        RECT -59.325 176.635 -58.995 176.965 ;
        RECT -59.325 175.275 -58.995 175.605 ;
        RECT -59.325 173.915 -58.995 174.245 ;
        RECT -59.325 172.555 -58.995 172.885 ;
        RECT -59.325 171.195 -58.995 171.525 ;
        RECT -59.325 169.835 -58.995 170.165 ;
        RECT -59.325 168.475 -58.995 168.805 ;
        RECT -59.325 167.115 -58.995 167.445 ;
        RECT -59.325 165.755 -58.995 166.085 ;
        RECT -59.325 164.395 -58.995 164.725 ;
        RECT -59.325 163.035 -58.995 163.365 ;
        RECT -59.325 161.675 -58.995 162.005 ;
        RECT -59.325 160.315 -58.995 160.645 ;
        RECT -59.325 158.955 -58.995 159.285 ;
        RECT -59.325 157.595 -58.995 157.925 ;
        RECT -59.325 156.235 -58.995 156.565 ;
        RECT -59.325 154.875 -58.995 155.205 ;
        RECT -59.325 153.515 -58.995 153.845 ;
        RECT -59.325 152.155 -58.995 152.485 ;
        RECT -59.325 150.795 -58.995 151.125 ;
        RECT -59.325 149.435 -58.995 149.765 ;
        RECT -59.325 148.075 -58.995 148.405 ;
        RECT -59.325 146.715 -58.995 147.045 ;
        RECT -59.325 145.355 -58.995 145.685 ;
        RECT -59.325 143.995 -58.995 144.325 ;
        RECT -59.325 142.635 -58.995 142.965 ;
        RECT -59.325 141.275 -58.995 141.605 ;
        RECT -59.325 139.915 -58.995 140.245 ;
        RECT -59.325 138.555 -58.995 138.885 ;
        RECT -59.325 137.225 -58.995 137.555 ;
        RECT -59.325 135.175 -58.995 135.505 ;
        RECT -59.325 132.815 -58.995 133.145 ;
        RECT -59.325 131.665 -58.995 131.995 ;
        RECT -59.325 129.655 -58.995 129.985 ;
        RECT -59.325 128.505 -58.995 128.835 ;
        RECT -59.325 126.495 -58.995 126.825 ;
        RECT -59.325 125.345 -58.995 125.675 ;
        RECT -59.325 123.335 -58.995 123.665 ;
        RECT -59.325 122.185 -58.995 122.515 ;
        RECT -59.325 120.175 -58.995 120.505 ;
        RECT -59.325 119.025 -58.995 119.355 ;
        RECT -59.325 117.185 -58.995 117.515 ;
        RECT -59.325 115.865 -58.995 116.195 ;
        RECT -59.325 113.855 -58.995 114.185 ;
        RECT -59.325 112.705 -58.995 113.035 ;
        RECT -59.325 110.695 -58.995 111.025 ;
        RECT -59.325 109.545 -58.995 109.875 ;
        RECT -59.325 107.535 -58.995 107.865 ;
        RECT -59.325 106.385 -58.995 106.715 ;
        RECT -59.325 104.375 -58.995 104.705 ;
        RECT -59.325 103.225 -58.995 103.555 ;
        RECT -59.325 100.865 -58.995 101.195 ;
        RECT -59.325 98.81 -58.995 99.14 ;
        RECT -59.325 97.755 -58.995 98.085 ;
        RECT -59.325 96.395 -58.995 96.725 ;
        RECT -59.325 95.035 -58.995 95.365 ;
        RECT -59.325 93.675 -58.995 94.005 ;
        RECT -59.325 92.315 -58.995 92.645 ;
        RECT -59.325 90.955 -58.995 91.285 ;
        RECT -59.325 89.595 -58.995 89.925 ;
        RECT -59.325 88.235 -58.995 88.565 ;
        RECT -59.32 87.56 -59 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -59.325 -2.885 -58.995 -2.555 ;
        RECT -59.325 -4.245 -58.995 -3.915 ;
        RECT -59.325 -5.605 -58.995 -5.275 ;
        RECT -59.325 -6.965 -58.995 -6.635 ;
        RECT -59.325 -8.325 -58.995 -7.995 ;
        RECT -59.325 -9.685 -58.995 -9.355 ;
        RECT -59.325 -11.045 -58.995 -10.715 ;
        RECT -59.325 -12.405 -58.995 -12.075 ;
        RECT -59.325 -13.765 -58.995 -13.435 ;
        RECT -59.325 -15.125 -58.995 -14.795 ;
        RECT -59.325 -16.485 -58.995 -16.155 ;
        RECT -59.325 -17.845 -58.995 -17.515 ;
        RECT -59.325 -19.205 -58.995 -18.875 ;
        RECT -59.325 -20.565 -58.995 -20.235 ;
        RECT -59.325 -21.925 -58.995 -21.595 ;
        RECT -59.325 -23.285 -58.995 -22.955 ;
        RECT -59.325 -24.645 -58.995 -24.315 ;
        RECT -59.325 -28.725 -58.995 -28.395 ;
        RECT -59.325 -30.085 -58.995 -29.755 ;
        RECT -59.325 -31.445 -58.995 -31.115 ;
        RECT -59.325 -32.805 -58.995 -32.475 ;
        RECT -59.325 -34.165 -58.995 -33.835 ;
        RECT -59.325 -35.525 -58.995 -35.195 ;
        RECT -59.325 -36.885 -58.995 -36.555 ;
        RECT -59.325 -38.245 -58.995 -37.915 ;
        RECT -59.325 -39.605 -58.995 -39.275 ;
        RECT -59.325 -40.965 -58.995 -40.635 ;
        RECT -59.325 -42.325 -58.995 -41.995 ;
        RECT -59.325 -43.685 -58.995 -43.355 ;
        RECT -59.325 -45.045 -58.995 -44.715 ;
        RECT -59.325 -46.405 -58.995 -46.075 ;
        RECT -59.325 -47.765 -58.995 -47.435 ;
        RECT -59.325 -49.125 -58.995 -48.795 ;
        RECT -59.325 -50.485 -58.995 -50.155 ;
        RECT -59.325 -51.845 -58.995 -51.515 ;
        RECT -59.325 -53.205 -58.995 -52.875 ;
        RECT -59.325 -54.565 -58.995 -54.235 ;
        RECT -59.325 -55.925 -58.995 -55.595 ;
        RECT -59.325 -57.285 -58.995 -56.955 ;
        RECT -59.325 -58.645 -58.995 -58.315 ;
        RECT -59.325 -60.005 -58.995 -59.675 ;
        RECT -59.325 -61.365 -58.995 -61.035 ;
        RECT -59.325 -62.725 -58.995 -62.395 ;
        RECT -59.325 -64.085 -58.995 -63.755 ;
        RECT -59.325 -65.445 -58.995 -65.115 ;
        RECT -59.325 -66.805 -58.995 -66.475 ;
        RECT -59.325 -68.165 -58.995 -67.835 ;
        RECT -59.325 -69.525 -58.995 -69.195 ;
        RECT -59.325 -70.885 -58.995 -70.555 ;
        RECT -59.325 -72.245 -58.995 -71.915 ;
        RECT -59.325 -73.605 -58.995 -73.275 ;
        RECT -59.325 -74.965 -58.995 -74.635 ;
        RECT -59.325 -76.325 -58.995 -75.995 ;
        RECT -59.325 -77.685 -58.995 -77.355 ;
        RECT -59.325 -79.045 -58.995 -78.715 ;
        RECT -59.325 -80.405 -58.995 -80.075 ;
        RECT -59.325 -81.765 -58.995 -81.435 ;
        RECT -59.325 -83.125 -58.995 -82.795 ;
        RECT -59.325 -84.485 -58.995 -84.155 ;
        RECT -59.325 -85.845 -58.995 -85.515 ;
        RECT -59.325 -87.205 -58.995 -86.875 ;
        RECT -59.325 -88.565 -58.995 -88.235 ;
        RECT -59.325 -89.925 -58.995 -89.595 ;
        RECT -59.325 -92.645 -58.995 -92.315 ;
        RECT -59.325 -94.005 -58.995 -93.675 ;
        RECT -59.325 -95.365 -58.995 -95.035 ;
        RECT -59.325 -96.725 -58.995 -96.395 ;
        RECT -59.325 -98.085 -58.995 -97.755 ;
        RECT -59.325 -99.69 -58.995 -99.36 ;
        RECT -59.325 -100.805 -58.995 -100.475 ;
        RECT -59.325 -103.525 -58.995 -103.195 ;
        RECT -59.325 -104.885 -58.995 -104.555 ;
        RECT -59.325 -106.245 -58.995 -105.915 ;
        RECT -59.325 -107.83 -58.995 -107.5 ;
        RECT -59.325 -108.965 -58.995 -108.635 ;
        RECT -59.325 -110.325 -58.995 -109.995 ;
        RECT -59.325 -111.685 -58.995 -111.355 ;
        RECT -59.325 -115.765 -58.995 -115.435 ;
        RECT -59.325 -117.125 -58.995 -116.795 ;
        RECT -59.325 -118.485 -58.995 -118.155 ;
        RECT -59.325 -119.845 -58.995 -119.515 ;
        RECT -59.325 -121.205 -58.995 -120.875 ;
        RECT -59.325 -123.925 -58.995 -123.595 ;
        RECT -59.325 -125.285 -58.995 -124.955 ;
        RECT -59.325 -126.645 -58.995 -126.315 ;
        RECT -59.325 -128.005 -58.995 -127.675 ;
        RECT -59.325 -129.365 -58.995 -129.035 ;
        RECT -59.325 -130.725 -58.995 -130.395 ;
        RECT -59.325 -132.085 -58.995 -131.755 ;
        RECT -59.325 -133.445 -58.995 -133.115 ;
        RECT -59.325 -134.805 -58.995 -134.475 ;
        RECT -59.325 -136.165 -58.995 -135.835 ;
        RECT -59.325 -137.525 -58.995 -137.195 ;
        RECT -59.325 -138.885 -58.995 -138.555 ;
        RECT -59.325 -140.245 -58.995 -139.915 ;
        RECT -59.325 -141.605 -58.995 -141.275 ;
        RECT -59.325 -142.965 -58.995 -142.635 ;
        RECT -59.325 -144.325 -58.995 -143.995 ;
        RECT -59.325 -145.685 -58.995 -145.355 ;
        RECT -59.325 -147.045 -58.995 -146.715 ;
        RECT -59.325 -148.405 -58.995 -148.075 ;
        RECT -59.325 -149.765 -58.995 -149.435 ;
        RECT -59.325 -151.125 -58.995 -150.795 ;
        RECT -59.325 -152.485 -58.995 -152.155 ;
        RECT -59.325 -153.845 -58.995 -153.515 ;
        RECT -59.325 -155.205 -58.995 -154.875 ;
        RECT -59.325 -156.565 -58.995 -156.235 ;
        RECT -59.325 -157.925 -58.995 -157.595 ;
        RECT -59.325 -159.285 -58.995 -158.955 ;
        RECT -59.325 -160.645 -58.995 -160.315 ;
        RECT -59.325 -162.005 -58.995 -161.675 ;
        RECT -59.325 -163.365 -58.995 -163.035 ;
        RECT -59.325 -164.725 -58.995 -164.395 ;
        RECT -59.325 -166.085 -58.995 -165.755 ;
        RECT -59.325 -167.445 -58.995 -167.115 ;
        RECT -59.325 -168.805 -58.995 -168.475 ;
        RECT -59.325 -171.525 -58.995 -171.195 ;
        RECT -59.325 -175.605 -58.995 -175.275 ;
        RECT -59.325 -176.685 -58.995 -176.355 ;
        RECT -59.325 -178.325 -58.995 -177.995 ;
        RECT -59.325 -179.685 -58.995 -179.355 ;
        RECT -59.325 -181.93 -58.995 -180.8 ;
        RECT -59.32 -182.045 -59 -1.88 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.965 241.32 -57.635 242.45 ;
        RECT -57.965 239.195 -57.635 239.525 ;
        RECT -57.965 237.835 -57.635 238.165 ;
        RECT -57.965 236.475 -57.635 236.805 ;
        RECT -57.965 235.115 -57.635 235.445 ;
        RECT -57.965 233.755 -57.635 234.085 ;
        RECT -57.965 232.395 -57.635 232.725 ;
        RECT -57.965 231.035 -57.635 231.365 ;
        RECT -57.965 229.675 -57.635 230.005 ;
        RECT -57.965 228.315 -57.635 228.645 ;
        RECT -57.965 226.955 -57.635 227.285 ;
        RECT -57.965 225.595 -57.635 225.925 ;
        RECT -57.965 224.235 -57.635 224.565 ;
        RECT -57.965 222.875 -57.635 223.205 ;
        RECT -57.965 221.515 -57.635 221.845 ;
        RECT -57.965 220.155 -57.635 220.485 ;
        RECT -57.965 218.795 -57.635 219.125 ;
        RECT -57.965 217.435 -57.635 217.765 ;
        RECT -57.965 216.075 -57.635 216.405 ;
        RECT -57.965 214.715 -57.635 215.045 ;
        RECT -57.965 213.355 -57.635 213.685 ;
        RECT -57.965 211.995 -57.635 212.325 ;
        RECT -57.965 210.635 -57.635 210.965 ;
        RECT -57.965 209.275 -57.635 209.605 ;
        RECT -57.965 207.915 -57.635 208.245 ;
        RECT -57.965 206.555 -57.635 206.885 ;
        RECT -57.965 205.195 -57.635 205.525 ;
        RECT -57.965 203.835 -57.635 204.165 ;
        RECT -57.965 202.475 -57.635 202.805 ;
        RECT -57.965 201.115 -57.635 201.445 ;
        RECT -57.965 199.755 -57.635 200.085 ;
        RECT -57.965 198.395 -57.635 198.725 ;
        RECT -57.965 197.035 -57.635 197.365 ;
        RECT -57.965 195.675 -57.635 196.005 ;
        RECT -57.965 194.315 -57.635 194.645 ;
        RECT -57.965 192.955 -57.635 193.285 ;
        RECT -57.965 191.595 -57.635 191.925 ;
        RECT -57.965 190.235 -57.635 190.565 ;
        RECT -57.965 188.875 -57.635 189.205 ;
        RECT -57.965 187.515 -57.635 187.845 ;
        RECT -57.965 186.155 -57.635 186.485 ;
        RECT -57.965 184.795 -57.635 185.125 ;
        RECT -57.965 183.435 -57.635 183.765 ;
        RECT -57.965 182.075 -57.635 182.405 ;
        RECT -57.965 180.715 -57.635 181.045 ;
        RECT -57.965 179.355 -57.635 179.685 ;
        RECT -57.965 177.995 -57.635 178.325 ;
        RECT -57.965 176.635 -57.635 176.965 ;
        RECT -57.965 175.275 -57.635 175.605 ;
        RECT -57.965 173.915 -57.635 174.245 ;
        RECT -57.965 172.555 -57.635 172.885 ;
        RECT -57.965 171.195 -57.635 171.525 ;
        RECT -57.965 169.835 -57.635 170.165 ;
        RECT -57.965 168.475 -57.635 168.805 ;
        RECT -57.965 167.115 -57.635 167.445 ;
        RECT -57.965 165.755 -57.635 166.085 ;
        RECT -57.965 164.395 -57.635 164.725 ;
        RECT -57.965 163.035 -57.635 163.365 ;
        RECT -57.965 161.675 -57.635 162.005 ;
        RECT -57.965 160.315 -57.635 160.645 ;
        RECT -57.965 158.955 -57.635 159.285 ;
        RECT -57.965 157.595 -57.635 157.925 ;
        RECT -57.965 156.235 -57.635 156.565 ;
        RECT -57.965 154.875 -57.635 155.205 ;
        RECT -57.965 153.515 -57.635 153.845 ;
        RECT -57.965 152.155 -57.635 152.485 ;
        RECT -57.965 150.795 -57.635 151.125 ;
        RECT -57.965 149.435 -57.635 149.765 ;
        RECT -57.965 148.075 -57.635 148.405 ;
        RECT -57.965 146.715 -57.635 147.045 ;
        RECT -57.965 145.355 -57.635 145.685 ;
        RECT -57.965 143.995 -57.635 144.325 ;
        RECT -57.965 142.635 -57.635 142.965 ;
        RECT -57.965 141.275 -57.635 141.605 ;
        RECT -57.965 139.915 -57.635 140.245 ;
        RECT -57.965 138.555 -57.635 138.885 ;
        RECT -57.96 138.555 -57.64 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -57.965 97.755 -57.635 98.085 ;
        RECT -57.965 96.395 -57.635 96.725 ;
        RECT -57.965 95.035 -57.635 95.365 ;
        RECT -57.965 93.675 -57.635 94.005 ;
        RECT -57.965 92.315 -57.635 92.645 ;
        RECT -57.965 89.595 -57.635 89.925 ;
        RECT -57.965 88.235 -57.635 88.565 ;
        RECT -57.965 84.155 -57.635 84.485 ;
        RECT -57.965 82.795 -57.635 83.125 ;
        RECT -57.965 81.435 -57.635 81.765 ;
        RECT -57.965 80.075 -57.635 80.405 ;
        RECT -57.965 78.715 -57.635 79.045 ;
        RECT -57.965 77.355 -57.635 77.685 ;
        RECT -57.965 75.995 -57.635 76.325 ;
        RECT -57.965 74.635 -57.635 74.965 ;
        RECT -57.965 73.275 -57.635 73.605 ;
        RECT -57.965 71.915 -57.635 72.245 ;
        RECT -57.965 70.555 -57.635 70.885 ;
        RECT -57.965 69.195 -57.635 69.525 ;
        RECT -57.965 67.835 -57.635 68.165 ;
        RECT -57.965 66.475 -57.635 66.805 ;
        RECT -57.965 65.115 -57.635 65.445 ;
        RECT -57.965 63.755 -57.635 64.085 ;
        RECT -57.965 62.395 -57.635 62.725 ;
        RECT -57.965 61.035 -57.635 61.365 ;
        RECT -57.965 59.675 -57.635 60.005 ;
        RECT -57.965 58.315 -57.635 58.645 ;
        RECT -57.965 56.955 -57.635 57.285 ;
        RECT -57.965 55.595 -57.635 55.925 ;
        RECT -57.965 54.235 -57.635 54.565 ;
        RECT -57.965 52.875 -57.635 53.205 ;
        RECT -57.965 51.515 -57.635 51.845 ;
        RECT -57.965 50.155 -57.635 50.485 ;
        RECT -57.965 48.795 -57.635 49.125 ;
        RECT -57.965 47.435 -57.635 47.765 ;
        RECT -57.965 46.075 -57.635 46.405 ;
        RECT -57.965 44.715 -57.635 45.045 ;
        RECT -57.965 43.355 -57.635 43.685 ;
        RECT -57.965 41.995 -57.635 42.325 ;
        RECT -57.965 40.635 -57.635 40.965 ;
        RECT -57.965 39.275 -57.635 39.605 ;
        RECT -57.965 37.915 -57.635 38.245 ;
        RECT -57.965 36.555 -57.635 36.885 ;
        RECT -57.965 35.195 -57.635 35.525 ;
        RECT -57.965 33.835 -57.635 34.165 ;
        RECT -57.965 32.475 -57.635 32.805 ;
        RECT -57.965 31.115 -57.635 31.445 ;
        RECT -57.965 29.755 -57.635 30.085 ;
        RECT -57.965 28.395 -57.635 28.725 ;
        RECT -57.965 27.035 -57.635 27.365 ;
        RECT -57.965 25.675 -57.635 26.005 ;
        RECT -57.965 24.315 -57.635 24.645 ;
        RECT -57.965 22.955 -57.635 23.285 ;
        RECT -57.965 21.595 -57.635 21.925 ;
        RECT -57.965 20.235 -57.635 20.565 ;
        RECT -57.965 18.875 -57.635 19.205 ;
        RECT -57.965 17.515 -57.635 17.845 ;
        RECT -57.965 16.155 -57.635 16.485 ;
        RECT -57.965 14.795 -57.635 15.125 ;
        RECT -57.965 13.435 -57.635 13.765 ;
        RECT -57.965 12.075 -57.635 12.405 ;
        RECT -57.965 10.715 -57.635 11.045 ;
        RECT -57.965 9.355 -57.635 9.685 ;
        RECT -57.965 7.995 -57.635 8.325 ;
        RECT -57.965 6.635 -57.635 6.965 ;
        RECT -57.965 5.275 -57.635 5.605 ;
        RECT -57.965 3.915 -57.635 4.245 ;
        RECT -57.965 2.555 -57.635 2.885 ;
        RECT -57.965 1.195 -57.635 1.525 ;
        RECT -57.965 -0.165 -57.635 0.165 ;
        RECT -57.965 -2.885 -57.635 -2.555 ;
        RECT -57.965 -4.245 -57.635 -3.915 ;
        RECT -57.965 -5.605 -57.635 -5.275 ;
        RECT -57.965 -6.965 -57.635 -6.635 ;
        RECT -57.965 -8.325 -57.635 -7.995 ;
        RECT -57.965 -9.685 -57.635 -9.355 ;
        RECT -57.965 -11.045 -57.635 -10.715 ;
        RECT -57.965 -12.405 -57.635 -12.075 ;
        RECT -57.965 -13.765 -57.635 -13.435 ;
        RECT -57.965 -15.125 -57.635 -14.795 ;
        RECT -57.965 -16.485 -57.635 -16.155 ;
        RECT -57.965 -17.845 -57.635 -17.515 ;
        RECT -57.965 -19.205 -57.635 -18.875 ;
        RECT -57.965 -20.565 -57.635 -20.235 ;
        RECT -57.965 -21.925 -57.635 -21.595 ;
        RECT -57.965 -23.285 -57.635 -22.955 ;
        RECT -57.965 -24.645 -57.635 -24.315 ;
        RECT -57.965 -30.085 -57.635 -29.755 ;
        RECT -57.965 -31.445 -57.635 -31.115 ;
        RECT -57.965 -32.805 -57.635 -32.475 ;
        RECT -57.965 -34.165 -57.635 -33.835 ;
        RECT -57.965 -35.525 -57.635 -35.195 ;
        RECT -57.965 -36.885 -57.635 -36.555 ;
        RECT -57.965 -38.245 -57.635 -37.915 ;
        RECT -57.965 -39.605 -57.635 -39.275 ;
        RECT -57.965 -40.965 -57.635 -40.635 ;
        RECT -57.965 -42.325 -57.635 -41.995 ;
        RECT -57.965 -43.685 -57.635 -43.355 ;
        RECT -57.965 -45.045 -57.635 -44.715 ;
        RECT -57.965 -46.405 -57.635 -46.075 ;
        RECT -57.965 -47.765 -57.635 -47.435 ;
        RECT -57.965 -49.125 -57.635 -48.795 ;
        RECT -57.965 -50.485 -57.635 -50.155 ;
        RECT -57.965 -51.845 -57.635 -51.515 ;
        RECT -57.965 -53.205 -57.635 -52.875 ;
        RECT -57.965 -54.565 -57.635 -54.235 ;
        RECT -57.965 -55.925 -57.635 -55.595 ;
        RECT -57.965 -57.285 -57.635 -56.955 ;
        RECT -57.965 -58.645 -57.635 -58.315 ;
        RECT -57.965 -60.005 -57.635 -59.675 ;
        RECT -57.965 -61.365 -57.635 -61.035 ;
        RECT -57.965 -62.725 -57.635 -62.395 ;
        RECT -57.965 -64.085 -57.635 -63.755 ;
        RECT -57.965 -65.445 -57.635 -65.115 ;
        RECT -57.965 -66.805 -57.635 -66.475 ;
        RECT -57.965 -68.165 -57.635 -67.835 ;
        RECT -57.965 -69.525 -57.635 -69.195 ;
        RECT -57.965 -70.885 -57.635 -70.555 ;
        RECT -57.965 -72.245 -57.635 -71.915 ;
        RECT -57.965 -73.605 -57.635 -73.275 ;
        RECT -57.965 -74.965 -57.635 -74.635 ;
        RECT -57.965 -76.325 -57.635 -75.995 ;
        RECT -57.965 -77.685 -57.635 -77.355 ;
        RECT -57.965 -79.045 -57.635 -78.715 ;
        RECT -57.965 -80.405 -57.635 -80.075 ;
        RECT -57.965 -81.765 -57.635 -81.435 ;
        RECT -57.965 -83.125 -57.635 -82.795 ;
        RECT -57.965 -84.485 -57.635 -84.155 ;
        RECT -57.965 -85.845 -57.635 -85.515 ;
        RECT -57.965 -87.205 -57.635 -86.875 ;
        RECT -57.965 -88.565 -57.635 -88.235 ;
        RECT -57.965 -89.925 -57.635 -89.595 ;
        RECT -57.965 -92.645 -57.635 -92.315 ;
        RECT -57.965 -94.005 -57.635 -93.675 ;
        RECT -57.965 -95.365 -57.635 -95.035 ;
        RECT -57.965 -96.725 -57.635 -96.395 ;
        RECT -57.965 -98.085 -57.635 -97.755 ;
        RECT -57.965 -99.69 -57.635 -99.36 ;
        RECT -57.965 -100.805 -57.635 -100.475 ;
        RECT -57.965 -103.525 -57.635 -103.195 ;
        RECT -57.965 -104.885 -57.635 -104.555 ;
        RECT -57.965 -106.245 -57.635 -105.915 ;
        RECT -57.965 -107.83 -57.635 -107.5 ;
        RECT -57.965 -108.965 -57.635 -108.635 ;
        RECT -57.965 -110.325 -57.635 -109.995 ;
        RECT -57.965 -111.685 -57.635 -111.355 ;
        RECT -57.965 -115.765 -57.635 -115.435 ;
        RECT -57.965 -117.125 -57.635 -116.795 ;
        RECT -57.965 -118.485 -57.635 -118.155 ;
        RECT -57.965 -119.845 -57.635 -119.515 ;
        RECT -57.965 -121.205 -57.635 -120.875 ;
        RECT -57.965 -123.925 -57.635 -123.595 ;
        RECT -57.965 -125.285 -57.635 -124.955 ;
        RECT -57.965 -126.645 -57.635 -126.315 ;
        RECT -57.965 -128.005 -57.635 -127.675 ;
        RECT -57.965 -129.365 -57.635 -129.035 ;
        RECT -57.965 -130.725 -57.635 -130.395 ;
        RECT -57.965 -132.085 -57.635 -131.755 ;
        RECT -57.965 -133.445 -57.635 -133.115 ;
        RECT -57.965 -134.805 -57.635 -134.475 ;
        RECT -57.965 -136.165 -57.635 -135.835 ;
        RECT -57.965 -137.525 -57.635 -137.195 ;
        RECT -57.965 -138.885 -57.635 -138.555 ;
        RECT -57.965 -140.245 -57.635 -139.915 ;
        RECT -57.965 -141.605 -57.635 -141.275 ;
        RECT -57.965 -142.965 -57.635 -142.635 ;
        RECT -57.965 -144.325 -57.635 -143.995 ;
        RECT -57.965 -145.685 -57.635 -145.355 ;
        RECT -57.965 -147.045 -57.635 -146.715 ;
        RECT -57.965 -148.405 -57.635 -148.075 ;
        RECT -57.965 -149.765 -57.635 -149.435 ;
        RECT -57.965 -151.125 -57.635 -150.795 ;
        RECT -57.965 -152.485 -57.635 -152.155 ;
        RECT -57.965 -153.845 -57.635 -153.515 ;
        RECT -57.965 -155.205 -57.635 -154.875 ;
        RECT -57.965 -156.565 -57.635 -156.235 ;
        RECT -57.965 -157.925 -57.635 -157.595 ;
        RECT -57.965 -159.285 -57.635 -158.955 ;
        RECT -57.965 -160.645 -57.635 -160.315 ;
        RECT -57.965 -162.005 -57.635 -161.675 ;
        RECT -57.965 -163.365 -57.635 -163.035 ;
        RECT -57.965 -164.725 -57.635 -164.395 ;
        RECT -57.965 -166.085 -57.635 -165.755 ;
        RECT -57.965 -167.445 -57.635 -167.115 ;
        RECT -57.965 -168.805 -57.635 -168.475 ;
        RECT -57.965 -171.525 -57.635 -171.195 ;
        RECT -57.965 -174.245 -57.635 -173.915 ;
        RECT -57.965 -175.605 -57.635 -175.275 ;
        RECT -57.965 -176.685 -57.635 -176.355 ;
        RECT -57.965 -178.325 -57.635 -177.995 ;
        RECT -57.965 -179.685 -57.635 -179.355 ;
        RECT -57.965 -181.93 -57.635 -180.8 ;
        RECT -57.96 -182.045 -57.64 98.085 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.605 241.32 -56.275 242.45 ;
        RECT -56.605 239.195 -56.275 239.525 ;
        RECT -56.605 237.835 -56.275 238.165 ;
        RECT -56.605 236.475 -56.275 236.805 ;
        RECT -56.605 235.115 -56.275 235.445 ;
        RECT -56.605 233.755 -56.275 234.085 ;
        RECT -56.605 232.395 -56.275 232.725 ;
        RECT -56.605 231.035 -56.275 231.365 ;
        RECT -56.605 229.675 -56.275 230.005 ;
        RECT -56.605 228.315 -56.275 228.645 ;
        RECT -56.605 226.955 -56.275 227.285 ;
        RECT -56.605 225.595 -56.275 225.925 ;
        RECT -56.605 224.235 -56.275 224.565 ;
        RECT -56.605 222.875 -56.275 223.205 ;
        RECT -56.605 221.515 -56.275 221.845 ;
        RECT -56.605 220.155 -56.275 220.485 ;
        RECT -56.605 218.795 -56.275 219.125 ;
        RECT -56.605 217.435 -56.275 217.765 ;
        RECT -56.605 216.075 -56.275 216.405 ;
        RECT -56.605 214.715 -56.275 215.045 ;
        RECT -56.605 213.355 -56.275 213.685 ;
        RECT -56.605 211.995 -56.275 212.325 ;
        RECT -56.605 210.635 -56.275 210.965 ;
        RECT -56.605 209.275 -56.275 209.605 ;
        RECT -56.605 207.915 -56.275 208.245 ;
        RECT -56.605 206.555 -56.275 206.885 ;
        RECT -56.605 205.195 -56.275 205.525 ;
        RECT -56.605 203.835 -56.275 204.165 ;
        RECT -56.605 202.475 -56.275 202.805 ;
        RECT -56.605 201.115 -56.275 201.445 ;
        RECT -56.605 199.755 -56.275 200.085 ;
        RECT -56.605 198.395 -56.275 198.725 ;
        RECT -56.605 197.035 -56.275 197.365 ;
        RECT -56.605 195.675 -56.275 196.005 ;
        RECT -56.605 194.315 -56.275 194.645 ;
        RECT -56.605 192.955 -56.275 193.285 ;
        RECT -56.605 191.595 -56.275 191.925 ;
        RECT -56.605 190.235 -56.275 190.565 ;
        RECT -56.605 188.875 -56.275 189.205 ;
        RECT -56.605 187.515 -56.275 187.845 ;
        RECT -56.605 186.155 -56.275 186.485 ;
        RECT -56.605 184.795 -56.275 185.125 ;
        RECT -56.605 183.435 -56.275 183.765 ;
        RECT -56.605 182.075 -56.275 182.405 ;
        RECT -56.605 180.715 -56.275 181.045 ;
        RECT -56.605 179.355 -56.275 179.685 ;
        RECT -56.605 177.995 -56.275 178.325 ;
        RECT -56.605 176.635 -56.275 176.965 ;
        RECT -56.605 175.275 -56.275 175.605 ;
        RECT -56.605 173.915 -56.275 174.245 ;
        RECT -56.605 172.555 -56.275 172.885 ;
        RECT -56.605 171.195 -56.275 171.525 ;
        RECT -56.605 169.835 -56.275 170.165 ;
        RECT -56.605 168.475 -56.275 168.805 ;
        RECT -56.605 167.115 -56.275 167.445 ;
        RECT -56.605 165.755 -56.275 166.085 ;
        RECT -56.605 164.395 -56.275 164.725 ;
        RECT -56.605 163.035 -56.275 163.365 ;
        RECT -56.605 161.675 -56.275 162.005 ;
        RECT -56.605 160.315 -56.275 160.645 ;
        RECT -56.605 158.955 -56.275 159.285 ;
        RECT -56.605 157.595 -56.275 157.925 ;
        RECT -56.605 156.235 -56.275 156.565 ;
        RECT -56.605 154.875 -56.275 155.205 ;
        RECT -56.605 153.515 -56.275 153.845 ;
        RECT -56.605 152.155 -56.275 152.485 ;
        RECT -56.605 150.795 -56.275 151.125 ;
        RECT -56.605 149.435 -56.275 149.765 ;
        RECT -56.605 148.075 -56.275 148.405 ;
        RECT -56.605 146.715 -56.275 147.045 ;
        RECT -56.605 145.355 -56.275 145.685 ;
        RECT -56.605 143.995 -56.275 144.325 ;
        RECT -56.605 142.635 -56.275 142.965 ;
        RECT -56.605 141.275 -56.275 141.605 ;
        RECT -56.605 139.915 -56.275 140.245 ;
        RECT -56.605 138.555 -56.275 138.885 ;
        RECT -56.6 138.555 -56.28 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -56.605 -138.885 -56.275 -138.555 ;
        RECT -56.605 -140.245 -56.275 -139.915 ;
        RECT -56.605 -141.605 -56.275 -141.275 ;
        RECT -56.605 -142.965 -56.275 -142.635 ;
        RECT -56.605 -144.325 -56.275 -143.995 ;
        RECT -56.605 -145.685 -56.275 -145.355 ;
        RECT -56.605 -147.045 -56.275 -146.715 ;
        RECT -56.605 -148.405 -56.275 -148.075 ;
        RECT -56.605 -149.765 -56.275 -149.435 ;
        RECT -56.605 -151.125 -56.275 -150.795 ;
        RECT -56.605 -152.485 -56.275 -152.155 ;
        RECT -56.605 -153.845 -56.275 -153.515 ;
        RECT -56.605 -155.205 -56.275 -154.875 ;
        RECT -56.605 -156.565 -56.275 -156.235 ;
        RECT -56.605 -157.925 -56.275 -157.595 ;
        RECT -56.605 -159.285 -56.275 -158.955 ;
        RECT -56.605 -160.645 -56.275 -160.315 ;
        RECT -56.605 -162.005 -56.275 -161.675 ;
        RECT -56.605 -163.365 -56.275 -163.035 ;
        RECT -56.605 -164.725 -56.275 -164.395 ;
        RECT -56.605 -166.085 -56.275 -165.755 ;
        RECT -56.605 -167.445 -56.275 -167.115 ;
        RECT -56.605 -168.805 -56.275 -168.475 ;
        RECT -56.605 -171.525 -56.275 -171.195 ;
        RECT -56.605 -172.885 -56.275 -172.555 ;
        RECT -56.605 -174.245 -56.275 -173.915 ;
        RECT -56.605 -175.605 -56.275 -175.275 ;
        RECT -56.605 -176.685 -56.275 -176.355 ;
        RECT -56.605 -178.325 -56.275 -177.995 ;
        RECT -56.605 -179.685 -56.275 -179.355 ;
        RECT -56.605 -181.93 -56.275 -180.8 ;
        RECT -56.6 -182.045 -56.28 98.085 ;
        RECT -56.605 97.755 -56.275 98.085 ;
        RECT -56.605 96.395 -56.275 96.725 ;
        RECT -56.605 95.035 -56.275 95.365 ;
        RECT -56.605 93.675 -56.275 94.005 ;
        RECT -56.605 92.315 -56.275 92.645 ;
        RECT -56.605 89.595 -56.275 89.925 ;
        RECT -56.605 88.235 -56.275 88.565 ;
        RECT -56.605 84.155 -56.275 84.485 ;
        RECT -56.605 82.795 -56.275 83.125 ;
        RECT -56.605 81.435 -56.275 81.765 ;
        RECT -56.605 80.075 -56.275 80.405 ;
        RECT -56.605 78.715 -56.275 79.045 ;
        RECT -56.605 77.355 -56.275 77.685 ;
        RECT -56.605 75.995 -56.275 76.325 ;
        RECT -56.605 74.635 -56.275 74.965 ;
        RECT -56.605 73.275 -56.275 73.605 ;
        RECT -56.605 71.915 -56.275 72.245 ;
        RECT -56.605 70.555 -56.275 70.885 ;
        RECT -56.605 69.195 -56.275 69.525 ;
        RECT -56.605 67.835 -56.275 68.165 ;
        RECT -56.605 66.475 -56.275 66.805 ;
        RECT -56.605 65.115 -56.275 65.445 ;
        RECT -56.605 63.755 -56.275 64.085 ;
        RECT -56.605 62.395 -56.275 62.725 ;
        RECT -56.605 61.035 -56.275 61.365 ;
        RECT -56.605 59.675 -56.275 60.005 ;
        RECT -56.605 58.315 -56.275 58.645 ;
        RECT -56.605 56.955 -56.275 57.285 ;
        RECT -56.605 55.595 -56.275 55.925 ;
        RECT -56.605 54.235 -56.275 54.565 ;
        RECT -56.605 52.875 -56.275 53.205 ;
        RECT -56.605 51.515 -56.275 51.845 ;
        RECT -56.605 50.155 -56.275 50.485 ;
        RECT -56.605 48.795 -56.275 49.125 ;
        RECT -56.605 47.435 -56.275 47.765 ;
        RECT -56.605 46.075 -56.275 46.405 ;
        RECT -56.605 44.715 -56.275 45.045 ;
        RECT -56.605 43.355 -56.275 43.685 ;
        RECT -56.605 41.995 -56.275 42.325 ;
        RECT -56.605 40.635 -56.275 40.965 ;
        RECT -56.605 39.275 -56.275 39.605 ;
        RECT -56.605 37.915 -56.275 38.245 ;
        RECT -56.605 36.555 -56.275 36.885 ;
        RECT -56.605 35.195 -56.275 35.525 ;
        RECT -56.605 33.835 -56.275 34.165 ;
        RECT -56.605 32.475 -56.275 32.805 ;
        RECT -56.605 31.115 -56.275 31.445 ;
        RECT -56.605 29.755 -56.275 30.085 ;
        RECT -56.605 28.395 -56.275 28.725 ;
        RECT -56.605 27.035 -56.275 27.365 ;
        RECT -56.605 25.675 -56.275 26.005 ;
        RECT -56.605 24.315 -56.275 24.645 ;
        RECT -56.605 22.955 -56.275 23.285 ;
        RECT -56.605 21.595 -56.275 21.925 ;
        RECT -56.605 20.235 -56.275 20.565 ;
        RECT -56.605 18.875 -56.275 19.205 ;
        RECT -56.605 17.515 -56.275 17.845 ;
        RECT -56.605 16.155 -56.275 16.485 ;
        RECT -56.605 14.795 -56.275 15.125 ;
        RECT -56.605 13.435 -56.275 13.765 ;
        RECT -56.605 12.075 -56.275 12.405 ;
        RECT -56.605 10.715 -56.275 11.045 ;
        RECT -56.605 9.355 -56.275 9.685 ;
        RECT -56.605 7.995 -56.275 8.325 ;
        RECT -56.605 6.635 -56.275 6.965 ;
        RECT -56.605 5.275 -56.275 5.605 ;
        RECT -56.605 3.915 -56.275 4.245 ;
        RECT -56.605 2.555 -56.275 2.885 ;
        RECT -56.605 1.195 -56.275 1.525 ;
        RECT -56.605 -0.165 -56.275 0.165 ;
        RECT -56.605 -2.885 -56.275 -2.555 ;
        RECT -56.605 -4.245 -56.275 -3.915 ;
        RECT -56.605 -5.605 -56.275 -5.275 ;
        RECT -56.605 -6.965 -56.275 -6.635 ;
        RECT -56.605 -8.325 -56.275 -7.995 ;
        RECT -56.605 -9.685 -56.275 -9.355 ;
        RECT -56.605 -11.045 -56.275 -10.715 ;
        RECT -56.605 -12.405 -56.275 -12.075 ;
        RECT -56.605 -13.765 -56.275 -13.435 ;
        RECT -56.605 -15.125 -56.275 -14.795 ;
        RECT -56.605 -16.485 -56.275 -16.155 ;
        RECT -56.605 -17.845 -56.275 -17.515 ;
        RECT -56.605 -19.205 -56.275 -18.875 ;
        RECT -56.605 -20.565 -56.275 -20.235 ;
        RECT -56.605 -21.925 -56.275 -21.595 ;
        RECT -56.605 -23.285 -56.275 -22.955 ;
        RECT -56.605 -24.645 -56.275 -24.315 ;
        RECT -56.605 -30.085 -56.275 -29.755 ;
        RECT -56.605 -31.445 -56.275 -31.115 ;
        RECT -56.605 -32.805 -56.275 -32.475 ;
        RECT -56.605 -34.165 -56.275 -33.835 ;
        RECT -56.605 -35.525 -56.275 -35.195 ;
        RECT -56.605 -36.885 -56.275 -36.555 ;
        RECT -56.605 -38.245 -56.275 -37.915 ;
        RECT -56.605 -39.605 -56.275 -39.275 ;
        RECT -56.605 -40.965 -56.275 -40.635 ;
        RECT -56.605 -42.325 -56.275 -41.995 ;
        RECT -56.605 -43.685 -56.275 -43.355 ;
        RECT -56.605 -45.045 -56.275 -44.715 ;
        RECT -56.605 -46.405 -56.275 -46.075 ;
        RECT -56.605 -47.765 -56.275 -47.435 ;
        RECT -56.605 -49.125 -56.275 -48.795 ;
        RECT -56.605 -50.485 -56.275 -50.155 ;
        RECT -56.605 -51.845 -56.275 -51.515 ;
        RECT -56.605 -53.205 -56.275 -52.875 ;
        RECT -56.605 -54.565 -56.275 -54.235 ;
        RECT -56.605 -55.925 -56.275 -55.595 ;
        RECT -56.605 -57.285 -56.275 -56.955 ;
        RECT -56.605 -58.645 -56.275 -58.315 ;
        RECT -56.605 -60.005 -56.275 -59.675 ;
        RECT -56.605 -61.365 -56.275 -61.035 ;
        RECT -56.605 -62.725 -56.275 -62.395 ;
        RECT -56.605 -64.085 -56.275 -63.755 ;
        RECT -56.605 -65.445 -56.275 -65.115 ;
        RECT -56.605 -66.805 -56.275 -66.475 ;
        RECT -56.605 -68.165 -56.275 -67.835 ;
        RECT -56.605 -69.525 -56.275 -69.195 ;
        RECT -56.605 -70.885 -56.275 -70.555 ;
        RECT -56.605 -72.245 -56.275 -71.915 ;
        RECT -56.605 -73.605 -56.275 -73.275 ;
        RECT -56.605 -74.965 -56.275 -74.635 ;
        RECT -56.605 -76.325 -56.275 -75.995 ;
        RECT -56.605 -77.685 -56.275 -77.355 ;
        RECT -56.605 -79.045 -56.275 -78.715 ;
        RECT -56.605 -80.405 -56.275 -80.075 ;
        RECT -56.605 -81.765 -56.275 -81.435 ;
        RECT -56.605 -83.125 -56.275 -82.795 ;
        RECT -56.605 -84.485 -56.275 -84.155 ;
        RECT -56.605 -85.845 -56.275 -85.515 ;
        RECT -56.605 -87.205 -56.275 -86.875 ;
        RECT -56.605 -88.565 -56.275 -88.235 ;
        RECT -56.605 -89.925 -56.275 -89.595 ;
        RECT -56.605 -92.645 -56.275 -92.315 ;
        RECT -56.605 -94.005 -56.275 -93.675 ;
        RECT -56.605 -95.365 -56.275 -95.035 ;
        RECT -56.605 -96.725 -56.275 -96.395 ;
        RECT -56.605 -98.085 -56.275 -97.755 ;
        RECT -56.605 -99.69 -56.275 -99.36 ;
        RECT -56.605 -100.805 -56.275 -100.475 ;
        RECT -56.605 -103.525 -56.275 -103.195 ;
        RECT -56.605 -104.885 -56.275 -104.555 ;
        RECT -56.605 -106.245 -56.275 -105.915 ;
        RECT -56.605 -107.83 -56.275 -107.5 ;
        RECT -56.605 -108.965 -56.275 -108.635 ;
        RECT -56.605 -110.325 -56.275 -109.995 ;
        RECT -56.605 -111.685 -56.275 -111.355 ;
        RECT -56.605 -114.405 -56.275 -114.075 ;
        RECT -56.605 -115.765 -56.275 -115.435 ;
        RECT -56.605 -117.125 -56.275 -116.795 ;
        RECT -56.605 -118.485 -56.275 -118.155 ;
        RECT -56.605 -119.845 -56.275 -119.515 ;
        RECT -56.605 -121.205 -56.275 -120.875 ;
        RECT -56.605 -123.925 -56.275 -123.595 ;
        RECT -56.605 -125.285 -56.275 -124.955 ;
        RECT -56.605 -126.645 -56.275 -126.315 ;
        RECT -56.605 -128.005 -56.275 -127.675 ;
        RECT -56.605 -129.365 -56.275 -129.035 ;
        RECT -56.605 -130.725 -56.275 -130.395 ;
        RECT -56.605 -132.085 -56.275 -131.755 ;
        RECT -56.605 -133.445 -56.275 -133.115 ;
        RECT -56.605 -134.805 -56.275 -134.475 ;
        RECT -56.605 -136.165 -56.275 -135.835 ;
        RECT -56.605 -137.525 -56.275 -137.195 ;
    END
    PORT
      LAYER met3 ;
        RECT -64.765 241.32 -64.435 242.45 ;
        RECT -64.765 239.195 -64.435 239.525 ;
        RECT -64.765 237.835 -64.435 238.165 ;
        RECT -64.765 236.475 -64.435 236.805 ;
        RECT -64.765 235.115 -64.435 235.445 ;
        RECT -64.765 233.755 -64.435 234.085 ;
        RECT -64.765 232.395 -64.435 232.725 ;
        RECT -64.765 231.035 -64.435 231.365 ;
        RECT -64.765 229.675 -64.435 230.005 ;
        RECT -64.765 228.315 -64.435 228.645 ;
        RECT -64.765 226.955 -64.435 227.285 ;
        RECT -64.765 225.595 -64.435 225.925 ;
        RECT -64.765 224.235 -64.435 224.565 ;
        RECT -64.765 222.875 -64.435 223.205 ;
        RECT -64.765 221.515 -64.435 221.845 ;
        RECT -64.765 220.155 -64.435 220.485 ;
        RECT -64.765 218.795 -64.435 219.125 ;
        RECT -64.765 217.435 -64.435 217.765 ;
        RECT -64.765 216.075 -64.435 216.405 ;
        RECT -64.765 214.715 -64.435 215.045 ;
        RECT -64.765 213.355 -64.435 213.685 ;
        RECT -64.765 211.995 -64.435 212.325 ;
        RECT -64.765 210.635 -64.435 210.965 ;
        RECT -64.765 209.275 -64.435 209.605 ;
        RECT -64.765 207.915 -64.435 208.245 ;
        RECT -64.765 206.555 -64.435 206.885 ;
        RECT -64.765 205.195 -64.435 205.525 ;
        RECT -64.765 203.835 -64.435 204.165 ;
        RECT -64.765 202.475 -64.435 202.805 ;
        RECT -64.765 201.115 -64.435 201.445 ;
        RECT -64.765 199.755 -64.435 200.085 ;
        RECT -64.765 198.395 -64.435 198.725 ;
        RECT -64.765 197.035 -64.435 197.365 ;
        RECT -64.765 195.675 -64.435 196.005 ;
        RECT -64.765 194.315 -64.435 194.645 ;
        RECT -64.765 192.955 -64.435 193.285 ;
        RECT -64.765 191.595 -64.435 191.925 ;
        RECT -64.765 190.235 -64.435 190.565 ;
        RECT -64.765 188.875 -64.435 189.205 ;
        RECT -64.765 187.515 -64.435 187.845 ;
        RECT -64.765 186.155 -64.435 186.485 ;
        RECT -64.765 184.795 -64.435 185.125 ;
        RECT -64.765 183.435 -64.435 183.765 ;
        RECT -64.765 182.075 -64.435 182.405 ;
        RECT -64.765 180.715 -64.435 181.045 ;
        RECT -64.765 179.355 -64.435 179.685 ;
        RECT -64.765 177.995 -64.435 178.325 ;
        RECT -64.765 176.635 -64.435 176.965 ;
        RECT -64.765 175.275 -64.435 175.605 ;
        RECT -64.765 173.915 -64.435 174.245 ;
        RECT -64.765 172.555 -64.435 172.885 ;
        RECT -64.765 171.195 -64.435 171.525 ;
        RECT -64.765 169.835 -64.435 170.165 ;
        RECT -64.765 168.475 -64.435 168.805 ;
        RECT -64.765 167.115 -64.435 167.445 ;
        RECT -64.765 165.755 -64.435 166.085 ;
        RECT -64.765 164.395 -64.435 164.725 ;
        RECT -64.765 163.035 -64.435 163.365 ;
        RECT -64.765 161.675 -64.435 162.005 ;
        RECT -64.765 160.315 -64.435 160.645 ;
        RECT -64.765 158.955 -64.435 159.285 ;
        RECT -64.765 157.595 -64.435 157.925 ;
        RECT -64.765 156.235 -64.435 156.565 ;
        RECT -64.765 154.875 -64.435 155.205 ;
        RECT -64.765 153.515 -64.435 153.845 ;
        RECT -64.765 152.155 -64.435 152.485 ;
        RECT -64.765 150.795 -64.435 151.125 ;
        RECT -64.765 149.435 -64.435 149.765 ;
        RECT -64.765 148.075 -64.435 148.405 ;
        RECT -64.765 146.715 -64.435 147.045 ;
        RECT -64.765 145.355 -64.435 145.685 ;
        RECT -64.765 143.995 -64.435 144.325 ;
        RECT -64.765 142.635 -64.435 142.965 ;
        RECT -64.765 141.275 -64.435 141.605 ;
        RECT -64.765 139.915 -64.435 140.245 ;
        RECT -64.765 138.555 -64.435 138.885 ;
        RECT -64.765 97.755 -64.435 98.085 ;
        RECT -64.765 96.395 -64.435 96.725 ;
        RECT -64.765 95.035 -64.435 95.365 ;
        RECT -64.765 93.675 -64.435 94.005 ;
        RECT -64.765 92.315 -64.435 92.645 ;
        RECT -64.765 90.955 -64.435 91.285 ;
        RECT -64.765 89.595 -64.435 89.925 ;
        RECT -64.765 88.235 -64.435 88.565 ;
        RECT -64.765 86.875 -64.435 87.205 ;
        RECT -64.765 85.515 -64.435 85.845 ;
        RECT -64.765 84.155 -64.435 84.485 ;
        RECT -64.765 82.795 -64.435 83.125 ;
        RECT -64.765 81.435 -64.435 81.765 ;
        RECT -64.765 80.075 -64.435 80.405 ;
        RECT -64.765 78.715 -64.435 79.045 ;
        RECT -64.765 77.355 -64.435 77.685 ;
        RECT -64.765 75.995 -64.435 76.325 ;
        RECT -64.765 74.635 -64.435 74.965 ;
        RECT -64.765 73.275 -64.435 73.605 ;
        RECT -64.765 71.915 -64.435 72.245 ;
        RECT -64.765 70.555 -64.435 70.885 ;
        RECT -64.765 69.195 -64.435 69.525 ;
        RECT -64.765 67.835 -64.435 68.165 ;
        RECT -64.765 66.475 -64.435 66.805 ;
        RECT -64.765 65.115 -64.435 65.445 ;
        RECT -64.765 63.755 -64.435 64.085 ;
        RECT -64.765 62.395 -64.435 62.725 ;
        RECT -64.765 61.035 -64.435 61.365 ;
        RECT -64.765 59.675 -64.435 60.005 ;
        RECT -64.765 58.315 -64.435 58.645 ;
        RECT -64.765 56.955 -64.435 57.285 ;
        RECT -64.765 55.595 -64.435 55.925 ;
        RECT -64.765 54.235 -64.435 54.565 ;
        RECT -64.765 52.875 -64.435 53.205 ;
        RECT -64.765 51.515 -64.435 51.845 ;
        RECT -64.765 50.155 -64.435 50.485 ;
        RECT -64.765 48.795 -64.435 49.125 ;
        RECT -64.765 47.435 -64.435 47.765 ;
        RECT -64.765 46.075 -64.435 46.405 ;
        RECT -64.765 44.715 -64.435 45.045 ;
        RECT -64.765 43.355 -64.435 43.685 ;
        RECT -64.765 41.995 -64.435 42.325 ;
        RECT -64.765 40.635 -64.435 40.965 ;
        RECT -64.765 39.275 -64.435 39.605 ;
        RECT -64.765 37.915 -64.435 38.245 ;
        RECT -64.765 36.555 -64.435 36.885 ;
        RECT -64.765 35.195 -64.435 35.525 ;
        RECT -64.765 33.835 -64.435 34.165 ;
        RECT -64.765 32.475 -64.435 32.805 ;
        RECT -64.765 31.115 -64.435 31.445 ;
        RECT -64.765 29.755 -64.435 30.085 ;
        RECT -64.765 28.395 -64.435 28.725 ;
        RECT -64.765 27.035 -64.435 27.365 ;
        RECT -64.765 25.675 -64.435 26.005 ;
        RECT -64.765 24.315 -64.435 24.645 ;
        RECT -64.765 22.955 -64.435 23.285 ;
        RECT -64.765 21.595 -64.435 21.925 ;
        RECT -64.765 20.235 -64.435 20.565 ;
        RECT -64.765 18.875 -64.435 19.205 ;
        RECT -64.765 17.515 -64.435 17.845 ;
        RECT -64.765 16.155 -64.435 16.485 ;
        RECT -64.765 14.795 -64.435 15.125 ;
        RECT -64.765 13.435 -64.435 13.765 ;
        RECT -64.765 12.075 -64.435 12.405 ;
        RECT -64.765 10.715 -64.435 11.045 ;
        RECT -64.765 9.355 -64.435 9.685 ;
        RECT -64.765 7.995 -64.435 8.325 ;
        RECT -64.765 6.635 -64.435 6.965 ;
        RECT -64.765 5.275 -64.435 5.605 ;
        RECT -64.765 3.915 -64.435 4.245 ;
        RECT -64.765 2.555 -64.435 2.885 ;
        RECT -64.765 1.195 -64.435 1.525 ;
        RECT -64.765 -0.165 -64.435 0.165 ;
        RECT -64.765 -1.525 -64.435 -1.195 ;
        RECT -64.765 -2.885 -64.435 -2.555 ;
        RECT -64.765 -4.245 -64.435 -3.915 ;
        RECT -64.765 -5.605 -64.435 -5.275 ;
        RECT -64.765 -6.965 -64.435 -6.635 ;
        RECT -64.765 -8.325 -64.435 -7.995 ;
        RECT -64.765 -9.685 -64.435 -9.355 ;
        RECT -64.765 -11.045 -64.435 -10.715 ;
        RECT -64.765 -12.405 -64.435 -12.075 ;
        RECT -64.765 -13.765 -64.435 -13.435 ;
        RECT -64.765 -15.125 -64.435 -14.795 ;
        RECT -64.765 -16.485 -64.435 -16.155 ;
        RECT -64.765 -17.845 -64.435 -17.515 ;
        RECT -64.765 -19.205 -64.435 -18.875 ;
        RECT -64.765 -20.565 -64.435 -20.235 ;
        RECT -64.765 -21.925 -64.435 -21.595 ;
        RECT -64.765 -23.285 -64.435 -22.955 ;
        RECT -64.765 -24.645 -64.435 -24.315 ;
        RECT -64.765 -27.365 -64.435 -27.035 ;
        RECT -64.765 -28.725 -64.435 -28.395 ;
        RECT -64.765 -30.085 -64.435 -29.755 ;
        RECT -64.765 -31.445 -64.435 -31.115 ;
        RECT -64.765 -32.805 -64.435 -32.475 ;
        RECT -64.765 -34.165 -64.435 -33.835 ;
        RECT -64.765 -35.525 -64.435 -35.195 ;
        RECT -64.765 -36.885 -64.435 -36.555 ;
        RECT -64.765 -38.245 -64.435 -37.915 ;
        RECT -64.765 -39.605 -64.435 -39.275 ;
        RECT -64.765 -40.965 -64.435 -40.635 ;
        RECT -64.765 -42.325 -64.435 -41.995 ;
        RECT -64.765 -43.685 -64.435 -43.355 ;
        RECT -64.765 -45.045 -64.435 -44.715 ;
        RECT -64.765 -46.405 -64.435 -46.075 ;
        RECT -64.765 -47.765 -64.435 -47.435 ;
        RECT -64.765 -49.125 -64.435 -48.795 ;
        RECT -64.765 -50.485 -64.435 -50.155 ;
        RECT -64.765 -51.845 -64.435 -51.515 ;
        RECT -64.765 -53.205 -64.435 -52.875 ;
        RECT -64.765 -54.565 -64.435 -54.235 ;
        RECT -64.765 -55.925 -64.435 -55.595 ;
        RECT -64.765 -57.285 -64.435 -56.955 ;
        RECT -64.765 -58.645 -64.435 -58.315 ;
        RECT -64.765 -60.005 -64.435 -59.675 ;
        RECT -64.765 -61.365 -64.435 -61.035 ;
        RECT -64.765 -62.725 -64.435 -62.395 ;
        RECT -64.765 -64.085 -64.435 -63.755 ;
        RECT -64.765 -65.445 -64.435 -65.115 ;
        RECT -64.765 -66.805 -64.435 -66.475 ;
        RECT -64.765 -68.165 -64.435 -67.835 ;
        RECT -64.765 -69.525 -64.435 -69.195 ;
        RECT -64.765 -70.885 -64.435 -70.555 ;
        RECT -64.765 -72.245 -64.435 -71.915 ;
        RECT -64.765 -73.605 -64.435 -73.275 ;
        RECT -64.765 -74.965 -64.435 -74.635 ;
        RECT -64.765 -76.325 -64.435 -75.995 ;
        RECT -64.765 -77.685 -64.435 -77.355 ;
        RECT -64.765 -79.045 -64.435 -78.715 ;
        RECT -64.765 -80.405 -64.435 -80.075 ;
        RECT -64.765 -81.765 -64.435 -81.435 ;
        RECT -64.765 -83.125 -64.435 -82.795 ;
        RECT -64.765 -84.485 -64.435 -84.155 ;
        RECT -64.765 -85.845 -64.435 -85.515 ;
        RECT -64.765 -87.205 -64.435 -86.875 ;
        RECT -64.765 -88.565 -64.435 -88.235 ;
        RECT -64.765 -89.925 -64.435 -89.595 ;
        RECT -64.765 -92.645 -64.435 -92.315 ;
        RECT -64.765 -94.005 -64.435 -93.675 ;
        RECT -64.765 -95.365 -64.435 -95.035 ;
        RECT -64.765 -96.725 -64.435 -96.395 ;
        RECT -64.765 -98.085 -64.435 -97.755 ;
        RECT -64.765 -99.69 -64.435 -99.36 ;
        RECT -64.765 -100.805 -64.435 -100.475 ;
        RECT -64.765 -103.525 -64.435 -103.195 ;
        RECT -64.765 -104.885 -64.435 -104.555 ;
        RECT -64.765 -106.245 -64.435 -105.915 ;
        RECT -64.765 -107.83 -64.435 -107.5 ;
        RECT -64.765 -108.965 -64.435 -108.635 ;
        RECT -64.765 -110.325 -64.435 -109.995 ;
        RECT -64.765 -111.685 -64.435 -111.355 ;
        RECT -64.76 -113.04 -64.44 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -63.405 241.32 -63.075 242.45 ;
        RECT -63.405 239.195 -63.075 239.525 ;
        RECT -63.405 237.835 -63.075 238.165 ;
        RECT -63.405 236.475 -63.075 236.805 ;
        RECT -63.405 235.115 -63.075 235.445 ;
        RECT -63.405 233.755 -63.075 234.085 ;
        RECT -63.405 232.395 -63.075 232.725 ;
        RECT -63.405 231.035 -63.075 231.365 ;
        RECT -63.405 229.675 -63.075 230.005 ;
        RECT -63.405 228.315 -63.075 228.645 ;
        RECT -63.405 226.955 -63.075 227.285 ;
        RECT -63.405 225.595 -63.075 225.925 ;
        RECT -63.405 224.235 -63.075 224.565 ;
        RECT -63.405 222.875 -63.075 223.205 ;
        RECT -63.405 221.515 -63.075 221.845 ;
        RECT -63.405 220.155 -63.075 220.485 ;
        RECT -63.405 218.795 -63.075 219.125 ;
        RECT -63.405 217.435 -63.075 217.765 ;
        RECT -63.405 216.075 -63.075 216.405 ;
        RECT -63.405 214.715 -63.075 215.045 ;
        RECT -63.405 213.355 -63.075 213.685 ;
        RECT -63.405 211.995 -63.075 212.325 ;
        RECT -63.405 210.635 -63.075 210.965 ;
        RECT -63.405 209.275 -63.075 209.605 ;
        RECT -63.405 207.915 -63.075 208.245 ;
        RECT -63.405 206.555 -63.075 206.885 ;
        RECT -63.405 205.195 -63.075 205.525 ;
        RECT -63.405 203.835 -63.075 204.165 ;
        RECT -63.405 202.475 -63.075 202.805 ;
        RECT -63.405 201.115 -63.075 201.445 ;
        RECT -63.405 199.755 -63.075 200.085 ;
        RECT -63.405 198.395 -63.075 198.725 ;
        RECT -63.405 197.035 -63.075 197.365 ;
        RECT -63.405 195.675 -63.075 196.005 ;
        RECT -63.405 194.315 -63.075 194.645 ;
        RECT -63.405 192.955 -63.075 193.285 ;
        RECT -63.405 191.595 -63.075 191.925 ;
        RECT -63.405 190.235 -63.075 190.565 ;
        RECT -63.405 188.875 -63.075 189.205 ;
        RECT -63.405 187.515 -63.075 187.845 ;
        RECT -63.405 186.155 -63.075 186.485 ;
        RECT -63.405 184.795 -63.075 185.125 ;
        RECT -63.405 183.435 -63.075 183.765 ;
        RECT -63.405 182.075 -63.075 182.405 ;
        RECT -63.405 180.715 -63.075 181.045 ;
        RECT -63.405 179.355 -63.075 179.685 ;
        RECT -63.405 177.995 -63.075 178.325 ;
        RECT -63.405 176.635 -63.075 176.965 ;
        RECT -63.405 175.275 -63.075 175.605 ;
        RECT -63.405 173.915 -63.075 174.245 ;
        RECT -63.405 172.555 -63.075 172.885 ;
        RECT -63.405 171.195 -63.075 171.525 ;
        RECT -63.405 169.835 -63.075 170.165 ;
        RECT -63.405 168.475 -63.075 168.805 ;
        RECT -63.405 167.115 -63.075 167.445 ;
        RECT -63.405 165.755 -63.075 166.085 ;
        RECT -63.405 164.395 -63.075 164.725 ;
        RECT -63.405 163.035 -63.075 163.365 ;
        RECT -63.405 161.675 -63.075 162.005 ;
        RECT -63.405 160.315 -63.075 160.645 ;
        RECT -63.405 158.955 -63.075 159.285 ;
        RECT -63.405 157.595 -63.075 157.925 ;
        RECT -63.405 156.235 -63.075 156.565 ;
        RECT -63.405 154.875 -63.075 155.205 ;
        RECT -63.405 153.515 -63.075 153.845 ;
        RECT -63.405 152.155 -63.075 152.485 ;
        RECT -63.405 150.795 -63.075 151.125 ;
        RECT -63.405 149.435 -63.075 149.765 ;
        RECT -63.405 148.075 -63.075 148.405 ;
        RECT -63.405 146.715 -63.075 147.045 ;
        RECT -63.405 145.355 -63.075 145.685 ;
        RECT -63.405 143.995 -63.075 144.325 ;
        RECT -63.405 142.635 -63.075 142.965 ;
        RECT -63.405 141.275 -63.075 141.605 ;
        RECT -63.405 139.915 -63.075 140.245 ;
        RECT -63.405 138.555 -63.075 138.885 ;
        RECT -63.405 137.225 -63.075 137.555 ;
        RECT -63.405 135.175 -63.075 135.505 ;
        RECT -63.405 132.815 -63.075 133.145 ;
        RECT -63.405 131.665 -63.075 131.995 ;
        RECT -63.405 129.655 -63.075 129.985 ;
        RECT -63.405 128.505 -63.075 128.835 ;
        RECT -63.405 126.495 -63.075 126.825 ;
        RECT -63.405 125.345 -63.075 125.675 ;
        RECT -63.405 123.335 -63.075 123.665 ;
        RECT -63.405 122.185 -63.075 122.515 ;
        RECT -63.405 120.175 -63.075 120.505 ;
        RECT -63.405 119.025 -63.075 119.355 ;
        RECT -63.405 117.185 -63.075 117.515 ;
        RECT -63.405 115.865 -63.075 116.195 ;
        RECT -63.405 113.855 -63.075 114.185 ;
        RECT -63.405 112.705 -63.075 113.035 ;
        RECT -63.405 110.695 -63.075 111.025 ;
        RECT -63.405 109.545 -63.075 109.875 ;
        RECT -63.405 107.535 -63.075 107.865 ;
        RECT -63.405 106.385 -63.075 106.715 ;
        RECT -63.405 104.375 -63.075 104.705 ;
        RECT -63.405 103.225 -63.075 103.555 ;
        RECT -63.405 100.865 -63.075 101.195 ;
        RECT -63.405 98.81 -63.075 99.14 ;
        RECT -63.405 97.755 -63.075 98.085 ;
        RECT -63.405 96.395 -63.075 96.725 ;
        RECT -63.405 95.035 -63.075 95.365 ;
        RECT -63.405 93.675 -63.075 94.005 ;
        RECT -63.405 92.315 -63.075 92.645 ;
        RECT -63.405 90.955 -63.075 91.285 ;
        RECT -63.405 89.595 -63.075 89.925 ;
        RECT -63.405 88.235 -63.075 88.565 ;
        RECT -63.405 86.875 -63.075 87.205 ;
        RECT -63.405 85.515 -63.075 85.845 ;
        RECT -63.405 84.155 -63.075 84.485 ;
        RECT -63.405 82.795 -63.075 83.125 ;
        RECT -63.405 81.435 -63.075 81.765 ;
        RECT -63.405 80.075 -63.075 80.405 ;
        RECT -63.405 78.715 -63.075 79.045 ;
        RECT -63.405 77.355 -63.075 77.685 ;
        RECT -63.405 75.995 -63.075 76.325 ;
        RECT -63.405 74.635 -63.075 74.965 ;
        RECT -63.405 73.275 -63.075 73.605 ;
        RECT -63.405 71.915 -63.075 72.245 ;
        RECT -63.405 70.555 -63.075 70.885 ;
        RECT -63.405 69.195 -63.075 69.525 ;
        RECT -63.405 67.835 -63.075 68.165 ;
        RECT -63.405 66.475 -63.075 66.805 ;
        RECT -63.405 65.115 -63.075 65.445 ;
        RECT -63.405 63.755 -63.075 64.085 ;
        RECT -63.405 62.395 -63.075 62.725 ;
        RECT -63.405 61.035 -63.075 61.365 ;
        RECT -63.405 59.675 -63.075 60.005 ;
        RECT -63.405 58.315 -63.075 58.645 ;
        RECT -63.405 56.955 -63.075 57.285 ;
        RECT -63.405 55.595 -63.075 55.925 ;
        RECT -63.405 54.235 -63.075 54.565 ;
        RECT -63.405 52.875 -63.075 53.205 ;
        RECT -63.405 51.515 -63.075 51.845 ;
        RECT -63.405 50.155 -63.075 50.485 ;
        RECT -63.405 48.795 -63.075 49.125 ;
        RECT -63.405 47.435 -63.075 47.765 ;
        RECT -63.405 46.075 -63.075 46.405 ;
        RECT -63.405 44.715 -63.075 45.045 ;
        RECT -63.405 43.355 -63.075 43.685 ;
        RECT -63.405 41.995 -63.075 42.325 ;
        RECT -63.405 40.635 -63.075 40.965 ;
        RECT -63.405 39.275 -63.075 39.605 ;
        RECT -63.405 37.915 -63.075 38.245 ;
        RECT -63.405 36.555 -63.075 36.885 ;
        RECT -63.405 35.195 -63.075 35.525 ;
        RECT -63.405 33.835 -63.075 34.165 ;
        RECT -63.405 32.475 -63.075 32.805 ;
        RECT -63.405 31.115 -63.075 31.445 ;
        RECT -63.405 29.755 -63.075 30.085 ;
        RECT -63.405 28.395 -63.075 28.725 ;
        RECT -63.405 27.035 -63.075 27.365 ;
        RECT -63.405 25.675 -63.075 26.005 ;
        RECT -63.405 24.315 -63.075 24.645 ;
        RECT -63.405 22.955 -63.075 23.285 ;
        RECT -63.405 21.595 -63.075 21.925 ;
        RECT -63.405 20.235 -63.075 20.565 ;
        RECT -63.405 18.875 -63.075 19.205 ;
        RECT -63.405 17.515 -63.075 17.845 ;
        RECT -63.405 16.155 -63.075 16.485 ;
        RECT -63.405 14.795 -63.075 15.125 ;
        RECT -63.405 13.435 -63.075 13.765 ;
        RECT -63.405 12.075 -63.075 12.405 ;
        RECT -63.405 10.715 -63.075 11.045 ;
        RECT -63.405 9.355 -63.075 9.685 ;
        RECT -63.405 7.995 -63.075 8.325 ;
        RECT -63.405 6.635 -63.075 6.965 ;
        RECT -63.405 5.275 -63.075 5.605 ;
        RECT -63.405 3.915 -63.075 4.245 ;
        RECT -63.405 2.555 -63.075 2.885 ;
        RECT -63.405 1.195 -63.075 1.525 ;
        RECT -63.405 -0.165 -63.075 0.165 ;
        RECT -63.405 -1.525 -63.075 -1.195 ;
        RECT -63.405 -2.885 -63.075 -2.555 ;
        RECT -63.405 -4.245 -63.075 -3.915 ;
        RECT -63.405 -5.605 -63.075 -5.275 ;
        RECT -63.405 -6.965 -63.075 -6.635 ;
        RECT -63.405 -8.325 -63.075 -7.995 ;
        RECT -63.405 -9.685 -63.075 -9.355 ;
        RECT -63.405 -11.045 -63.075 -10.715 ;
        RECT -63.405 -12.405 -63.075 -12.075 ;
        RECT -63.405 -13.765 -63.075 -13.435 ;
        RECT -63.405 -15.125 -63.075 -14.795 ;
        RECT -63.405 -16.485 -63.075 -16.155 ;
        RECT -63.405 -17.845 -63.075 -17.515 ;
        RECT -63.405 -19.205 -63.075 -18.875 ;
        RECT -63.405 -20.565 -63.075 -20.235 ;
        RECT -63.405 -21.925 -63.075 -21.595 ;
        RECT -63.405 -23.285 -63.075 -22.955 ;
        RECT -63.405 -24.645 -63.075 -24.315 ;
        RECT -63.405 -28.725 -63.075 -28.395 ;
        RECT -63.405 -30.085 -63.075 -29.755 ;
        RECT -63.405 -31.445 -63.075 -31.115 ;
        RECT -63.405 -32.805 -63.075 -32.475 ;
        RECT -63.405 -34.165 -63.075 -33.835 ;
        RECT -63.405 -35.525 -63.075 -35.195 ;
        RECT -63.405 -36.885 -63.075 -36.555 ;
        RECT -63.405 -38.245 -63.075 -37.915 ;
        RECT -63.405 -39.605 -63.075 -39.275 ;
        RECT -63.405 -40.965 -63.075 -40.635 ;
        RECT -63.405 -42.325 -63.075 -41.995 ;
        RECT -63.405 -43.685 -63.075 -43.355 ;
        RECT -63.405 -45.045 -63.075 -44.715 ;
        RECT -63.405 -46.405 -63.075 -46.075 ;
        RECT -63.405 -47.765 -63.075 -47.435 ;
        RECT -63.405 -49.125 -63.075 -48.795 ;
        RECT -63.405 -50.485 -63.075 -50.155 ;
        RECT -63.405 -51.845 -63.075 -51.515 ;
        RECT -63.405 -53.205 -63.075 -52.875 ;
        RECT -63.405 -54.565 -63.075 -54.235 ;
        RECT -63.405 -55.925 -63.075 -55.595 ;
        RECT -63.405 -57.285 -63.075 -56.955 ;
        RECT -63.405 -58.645 -63.075 -58.315 ;
        RECT -63.405 -60.005 -63.075 -59.675 ;
        RECT -63.405 -61.365 -63.075 -61.035 ;
        RECT -63.405 -62.725 -63.075 -62.395 ;
        RECT -63.405 -64.085 -63.075 -63.755 ;
        RECT -63.405 -65.445 -63.075 -65.115 ;
        RECT -63.405 -66.805 -63.075 -66.475 ;
        RECT -63.405 -68.165 -63.075 -67.835 ;
        RECT -63.405 -69.525 -63.075 -69.195 ;
        RECT -63.405 -70.885 -63.075 -70.555 ;
        RECT -63.405 -72.245 -63.075 -71.915 ;
        RECT -63.405 -73.605 -63.075 -73.275 ;
        RECT -63.405 -74.965 -63.075 -74.635 ;
        RECT -63.405 -76.325 -63.075 -75.995 ;
        RECT -63.405 -77.685 -63.075 -77.355 ;
        RECT -63.405 -79.045 -63.075 -78.715 ;
        RECT -63.405 -80.405 -63.075 -80.075 ;
        RECT -63.405 -81.765 -63.075 -81.435 ;
        RECT -63.405 -83.125 -63.075 -82.795 ;
        RECT -63.405 -84.485 -63.075 -84.155 ;
        RECT -63.405 -85.845 -63.075 -85.515 ;
        RECT -63.405 -87.205 -63.075 -86.875 ;
        RECT -63.405 -88.565 -63.075 -88.235 ;
        RECT -63.405 -89.925 -63.075 -89.595 ;
        RECT -63.405 -92.645 -63.075 -92.315 ;
        RECT -63.405 -94.005 -63.075 -93.675 ;
        RECT -63.405 -95.365 -63.075 -95.035 ;
        RECT -63.405 -96.725 -63.075 -96.395 ;
        RECT -63.405 -98.085 -63.075 -97.755 ;
        RECT -63.405 -99.69 -63.075 -99.36 ;
        RECT -63.405 -100.805 -63.075 -100.475 ;
        RECT -63.405 -103.525 -63.075 -103.195 ;
        RECT -63.405 -104.885 -63.075 -104.555 ;
        RECT -63.405 -106.245 -63.075 -105.915 ;
        RECT -63.405 -107.83 -63.075 -107.5 ;
        RECT -63.405 -108.965 -63.075 -108.635 ;
        RECT -63.405 -110.325 -63.075 -109.995 ;
        RECT -63.405 -111.685 -63.075 -111.355 ;
        RECT -63.405 -114.405 -63.075 -114.075 ;
        RECT -63.405 -115.765 -63.075 -115.435 ;
        RECT -63.405 -117.125 -63.075 -116.795 ;
        RECT -63.405 -118.485 -63.075 -118.155 ;
        RECT -63.405 -119.845 -63.075 -119.515 ;
        RECT -63.405 -121.205 -63.075 -120.875 ;
        RECT -63.405 -122.565 -63.075 -122.235 ;
        RECT -63.405 -123.925 -63.075 -123.595 ;
        RECT -63.405 -125.285 -63.075 -124.955 ;
        RECT -63.405 -126.645 -63.075 -126.315 ;
        RECT -63.405 -128.005 -63.075 -127.675 ;
        RECT -63.405 -129.365 -63.075 -129.035 ;
        RECT -63.405 -130.725 -63.075 -130.395 ;
        RECT -63.405 -132.085 -63.075 -131.755 ;
        RECT -63.405 -133.445 -63.075 -133.115 ;
        RECT -63.405 -134.805 -63.075 -134.475 ;
        RECT -63.405 -136.165 -63.075 -135.835 ;
        RECT -63.405 -137.525 -63.075 -137.195 ;
        RECT -63.405 -138.885 -63.075 -138.555 ;
        RECT -63.405 -140.245 -63.075 -139.915 ;
        RECT -63.405 -141.605 -63.075 -141.275 ;
        RECT -63.405 -142.965 -63.075 -142.635 ;
        RECT -63.405 -144.325 -63.075 -143.995 ;
        RECT -63.405 -145.685 -63.075 -145.355 ;
        RECT -63.405 -147.045 -63.075 -146.715 ;
        RECT -63.405 -148.405 -63.075 -148.075 ;
        RECT -63.405 -149.765 -63.075 -149.435 ;
        RECT -63.405 -151.125 -63.075 -150.795 ;
        RECT -63.405 -152.485 -63.075 -152.155 ;
        RECT -63.405 -153.845 -63.075 -153.515 ;
        RECT -63.405 -155.205 -63.075 -154.875 ;
        RECT -63.405 -156.565 -63.075 -156.235 ;
        RECT -63.405 -157.925 -63.075 -157.595 ;
        RECT -63.405 -159.285 -63.075 -158.955 ;
        RECT -63.405 -160.645 -63.075 -160.315 ;
        RECT -63.405 -162.005 -63.075 -161.675 ;
        RECT -63.405 -163.365 -63.075 -163.035 ;
        RECT -63.405 -164.725 -63.075 -164.395 ;
        RECT -63.405 -166.085 -63.075 -165.755 ;
        RECT -63.405 -167.445 -63.075 -167.115 ;
        RECT -63.405 -168.805 -63.075 -168.475 ;
        RECT -63.405 -171.525 -63.075 -171.195 ;
        RECT -63.405 -174.245 -63.075 -173.915 ;
        RECT -63.405 -175.605 -63.075 -175.275 ;
        RECT -63.405 -176.685 -63.075 -176.355 ;
        RECT -63.405 -178.325 -63.075 -177.995 ;
        RECT -63.405 -179.685 -63.075 -179.355 ;
        RECT -63.405 -181.93 -63.075 -180.8 ;
        RECT -63.4 -182.045 -63.08 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -62.045 55.595 -61.715 55.925 ;
        RECT -62.045 54.235 -61.715 54.565 ;
        RECT -62.045 52.875 -61.715 53.205 ;
        RECT -62.045 51.515 -61.715 51.845 ;
        RECT -62.045 50.155 -61.715 50.485 ;
        RECT -62.045 48.795 -61.715 49.125 ;
        RECT -62.045 47.435 -61.715 47.765 ;
        RECT -62.045 46.075 -61.715 46.405 ;
        RECT -62.045 44.715 -61.715 45.045 ;
        RECT -62.045 43.355 -61.715 43.685 ;
        RECT -62.045 41.995 -61.715 42.325 ;
        RECT -62.045 40.635 -61.715 40.965 ;
        RECT -62.045 39.275 -61.715 39.605 ;
        RECT -62.045 37.915 -61.715 38.245 ;
        RECT -62.045 36.555 -61.715 36.885 ;
        RECT -62.045 35.195 -61.715 35.525 ;
        RECT -62.045 33.835 -61.715 34.165 ;
        RECT -62.045 32.475 -61.715 32.805 ;
        RECT -62.045 31.115 -61.715 31.445 ;
        RECT -62.045 29.755 -61.715 30.085 ;
        RECT -62.045 28.395 -61.715 28.725 ;
        RECT -62.045 27.035 -61.715 27.365 ;
        RECT -62.045 25.675 -61.715 26.005 ;
        RECT -62.045 24.315 -61.715 24.645 ;
        RECT -62.045 22.955 -61.715 23.285 ;
        RECT -62.045 21.595 -61.715 21.925 ;
        RECT -62.045 20.235 -61.715 20.565 ;
        RECT -62.045 18.875 -61.715 19.205 ;
        RECT -62.045 17.515 -61.715 17.845 ;
        RECT -62.045 16.155 -61.715 16.485 ;
        RECT -62.045 14.795 -61.715 15.125 ;
        RECT -62.045 13.435 -61.715 13.765 ;
        RECT -62.045 12.075 -61.715 12.405 ;
        RECT -62.045 10.715 -61.715 11.045 ;
        RECT -62.045 9.355 -61.715 9.685 ;
        RECT -62.045 7.995 -61.715 8.325 ;
        RECT -62.045 6.635 -61.715 6.965 ;
        RECT -62.045 5.275 -61.715 5.605 ;
        RECT -62.045 3.915 -61.715 4.245 ;
        RECT -62.045 2.555 -61.715 2.885 ;
        RECT -62.045 1.195 -61.715 1.525 ;
        RECT -62.045 -0.165 -61.715 0.165 ;
        RECT -62.045 -1.525 -61.715 -1.195 ;
        RECT -62.045 -2.885 -61.715 -2.555 ;
        RECT -62.045 -4.245 -61.715 -3.915 ;
        RECT -62.045 -5.605 -61.715 -5.275 ;
        RECT -62.045 -6.965 -61.715 -6.635 ;
        RECT -62.045 -8.325 -61.715 -7.995 ;
        RECT -62.045 -9.685 -61.715 -9.355 ;
        RECT -62.045 -11.045 -61.715 -10.715 ;
        RECT -62.045 -12.405 -61.715 -12.075 ;
        RECT -62.045 -13.765 -61.715 -13.435 ;
        RECT -62.045 -15.125 -61.715 -14.795 ;
        RECT -62.045 -16.485 -61.715 -16.155 ;
        RECT -62.045 -17.845 -61.715 -17.515 ;
        RECT -62.045 -19.205 -61.715 -18.875 ;
        RECT -62.045 -20.565 -61.715 -20.235 ;
        RECT -62.045 -21.925 -61.715 -21.595 ;
        RECT -62.045 -23.285 -61.715 -22.955 ;
        RECT -62.045 -24.645 -61.715 -24.315 ;
        RECT -62.045 -28.725 -61.715 -28.395 ;
        RECT -62.045 -30.085 -61.715 -29.755 ;
        RECT -62.045 -31.445 -61.715 -31.115 ;
        RECT -62.045 -32.805 -61.715 -32.475 ;
        RECT -62.045 -34.165 -61.715 -33.835 ;
        RECT -62.045 -35.525 -61.715 -35.195 ;
        RECT -62.045 -36.885 -61.715 -36.555 ;
        RECT -62.045 -38.245 -61.715 -37.915 ;
        RECT -62.045 -39.605 -61.715 -39.275 ;
        RECT -62.045 -40.965 -61.715 -40.635 ;
        RECT -62.045 -42.325 -61.715 -41.995 ;
        RECT -62.045 -43.685 -61.715 -43.355 ;
        RECT -62.045 -45.045 -61.715 -44.715 ;
        RECT -62.045 -46.405 -61.715 -46.075 ;
        RECT -62.045 -47.765 -61.715 -47.435 ;
        RECT -62.045 -49.125 -61.715 -48.795 ;
        RECT -62.045 -50.485 -61.715 -50.155 ;
        RECT -62.045 -51.845 -61.715 -51.515 ;
        RECT -62.045 -53.205 -61.715 -52.875 ;
        RECT -62.045 -54.565 -61.715 -54.235 ;
        RECT -62.045 -55.925 -61.715 -55.595 ;
        RECT -62.045 -57.285 -61.715 -56.955 ;
        RECT -62.045 -58.645 -61.715 -58.315 ;
        RECT -62.045 -60.005 -61.715 -59.675 ;
        RECT -62.045 -61.365 -61.715 -61.035 ;
        RECT -62.045 -62.725 -61.715 -62.395 ;
        RECT -62.045 -64.085 -61.715 -63.755 ;
        RECT -62.045 -65.445 -61.715 -65.115 ;
        RECT -62.045 -66.805 -61.715 -66.475 ;
        RECT -62.045 -68.165 -61.715 -67.835 ;
        RECT -62.045 -69.525 -61.715 -69.195 ;
        RECT -62.045 -70.885 -61.715 -70.555 ;
        RECT -62.045 -72.245 -61.715 -71.915 ;
        RECT -62.045 -73.605 -61.715 -73.275 ;
        RECT -62.045 -74.965 -61.715 -74.635 ;
        RECT -62.045 -76.325 -61.715 -75.995 ;
        RECT -62.045 -77.685 -61.715 -77.355 ;
        RECT -62.045 -79.045 -61.715 -78.715 ;
        RECT -62.045 -80.405 -61.715 -80.075 ;
        RECT -62.045 -81.765 -61.715 -81.435 ;
        RECT -62.045 -83.125 -61.715 -82.795 ;
        RECT -62.045 -84.485 -61.715 -84.155 ;
        RECT -62.045 -85.845 -61.715 -85.515 ;
        RECT -62.045 -87.205 -61.715 -86.875 ;
        RECT -62.045 -88.565 -61.715 -88.235 ;
        RECT -62.045 -89.925 -61.715 -89.595 ;
        RECT -62.045 -92.645 -61.715 -92.315 ;
        RECT -62.045 -94.005 -61.715 -93.675 ;
        RECT -62.045 -95.365 -61.715 -95.035 ;
        RECT -62.045 -96.725 -61.715 -96.395 ;
        RECT -62.045 -98.085 -61.715 -97.755 ;
        RECT -62.045 -99.69 -61.715 -99.36 ;
        RECT -62.045 -100.805 -61.715 -100.475 ;
        RECT -62.045 -103.525 -61.715 -103.195 ;
        RECT -62.045 -104.885 -61.715 -104.555 ;
        RECT -62.045 -106.245 -61.715 -105.915 ;
        RECT -62.045 -107.83 -61.715 -107.5 ;
        RECT -62.045 -108.965 -61.715 -108.635 ;
        RECT -62.045 -110.325 -61.715 -109.995 ;
        RECT -62.045 -111.685 -61.715 -111.355 ;
        RECT -62.045 -114.405 -61.715 -114.075 ;
        RECT -62.045 -115.765 -61.715 -115.435 ;
        RECT -62.045 -117.125 -61.715 -116.795 ;
        RECT -62.045 -118.485 -61.715 -118.155 ;
        RECT -62.045 -119.845 -61.715 -119.515 ;
        RECT -62.045 -121.205 -61.715 -120.875 ;
        RECT -62.045 -122.565 -61.715 -122.235 ;
        RECT -62.045 -123.925 -61.715 -123.595 ;
        RECT -62.045 -125.285 -61.715 -124.955 ;
        RECT -62.045 -126.645 -61.715 -126.315 ;
        RECT -62.045 -128.005 -61.715 -127.675 ;
        RECT -62.045 -129.365 -61.715 -129.035 ;
        RECT -62.045 -130.725 -61.715 -130.395 ;
        RECT -62.045 -132.085 -61.715 -131.755 ;
        RECT -62.045 -133.445 -61.715 -133.115 ;
        RECT -62.045 -134.805 -61.715 -134.475 ;
        RECT -62.045 -136.165 -61.715 -135.835 ;
        RECT -62.045 -137.525 -61.715 -137.195 ;
        RECT -62.045 -138.885 -61.715 -138.555 ;
        RECT -62.045 -140.245 -61.715 -139.915 ;
        RECT -62.045 -141.605 -61.715 -141.275 ;
        RECT -62.045 -142.965 -61.715 -142.635 ;
        RECT -62.045 -144.325 -61.715 -143.995 ;
        RECT -62.045 -145.685 -61.715 -145.355 ;
        RECT -62.045 -147.045 -61.715 -146.715 ;
        RECT -62.045 -148.405 -61.715 -148.075 ;
        RECT -62.045 -149.765 -61.715 -149.435 ;
        RECT -62.045 -151.125 -61.715 -150.795 ;
        RECT -62.045 -152.485 -61.715 -152.155 ;
        RECT -62.045 -153.845 -61.715 -153.515 ;
        RECT -62.045 -155.205 -61.715 -154.875 ;
        RECT -62.045 -156.565 -61.715 -156.235 ;
        RECT -62.045 -157.925 -61.715 -157.595 ;
        RECT -62.045 -159.285 -61.715 -158.955 ;
        RECT -62.045 -160.645 -61.715 -160.315 ;
        RECT -62.045 -162.005 -61.715 -161.675 ;
        RECT -62.045 -163.365 -61.715 -163.035 ;
        RECT -62.045 -164.725 -61.715 -164.395 ;
        RECT -62.045 -166.085 -61.715 -165.755 ;
        RECT -62.045 -167.445 -61.715 -167.115 ;
        RECT -62.045 -168.805 -61.715 -168.475 ;
        RECT -62.045 -171.525 -61.715 -171.195 ;
        RECT -62.045 -172.885 -61.715 -172.555 ;
        RECT -62.045 -174.245 -61.715 -173.915 ;
        RECT -62.045 -175.605 -61.715 -175.275 ;
        RECT -62.045 -176.685 -61.715 -176.355 ;
        RECT -62.045 -178.325 -61.715 -177.995 ;
        RECT -62.045 -179.685 -61.715 -179.355 ;
        RECT -62.045 -181.93 -61.715 -180.8 ;
        RECT -62.04 -182.045 -61.72 242.565 ;
        RECT -62.045 241.32 -61.715 242.45 ;
        RECT -62.045 239.195 -61.715 239.525 ;
        RECT -62.045 237.835 -61.715 238.165 ;
        RECT -62.045 236.475 -61.715 236.805 ;
        RECT -62.045 235.115 -61.715 235.445 ;
        RECT -62.045 233.755 -61.715 234.085 ;
        RECT -62.045 232.395 -61.715 232.725 ;
        RECT -62.045 231.035 -61.715 231.365 ;
        RECT -62.045 229.675 -61.715 230.005 ;
        RECT -62.045 228.315 -61.715 228.645 ;
        RECT -62.045 226.955 -61.715 227.285 ;
        RECT -62.045 225.595 -61.715 225.925 ;
        RECT -62.045 224.235 -61.715 224.565 ;
        RECT -62.045 222.875 -61.715 223.205 ;
        RECT -62.045 221.515 -61.715 221.845 ;
        RECT -62.045 220.155 -61.715 220.485 ;
        RECT -62.045 218.795 -61.715 219.125 ;
        RECT -62.045 217.435 -61.715 217.765 ;
        RECT -62.045 216.075 -61.715 216.405 ;
        RECT -62.045 214.715 -61.715 215.045 ;
        RECT -62.045 213.355 -61.715 213.685 ;
        RECT -62.045 211.995 -61.715 212.325 ;
        RECT -62.045 210.635 -61.715 210.965 ;
        RECT -62.045 209.275 -61.715 209.605 ;
        RECT -62.045 207.915 -61.715 208.245 ;
        RECT -62.045 206.555 -61.715 206.885 ;
        RECT -62.045 205.195 -61.715 205.525 ;
        RECT -62.045 203.835 -61.715 204.165 ;
        RECT -62.045 202.475 -61.715 202.805 ;
        RECT -62.045 201.115 -61.715 201.445 ;
        RECT -62.045 199.755 -61.715 200.085 ;
        RECT -62.045 198.395 -61.715 198.725 ;
        RECT -62.045 197.035 -61.715 197.365 ;
        RECT -62.045 195.675 -61.715 196.005 ;
        RECT -62.045 194.315 -61.715 194.645 ;
        RECT -62.045 192.955 -61.715 193.285 ;
        RECT -62.045 191.595 -61.715 191.925 ;
        RECT -62.045 190.235 -61.715 190.565 ;
        RECT -62.045 188.875 -61.715 189.205 ;
        RECT -62.045 187.515 -61.715 187.845 ;
        RECT -62.045 186.155 -61.715 186.485 ;
        RECT -62.045 184.795 -61.715 185.125 ;
        RECT -62.045 183.435 -61.715 183.765 ;
        RECT -62.045 182.075 -61.715 182.405 ;
        RECT -62.045 180.715 -61.715 181.045 ;
        RECT -62.045 179.355 -61.715 179.685 ;
        RECT -62.045 177.995 -61.715 178.325 ;
        RECT -62.045 176.635 -61.715 176.965 ;
        RECT -62.045 175.275 -61.715 175.605 ;
        RECT -62.045 173.915 -61.715 174.245 ;
        RECT -62.045 172.555 -61.715 172.885 ;
        RECT -62.045 171.195 -61.715 171.525 ;
        RECT -62.045 169.835 -61.715 170.165 ;
        RECT -62.045 168.475 -61.715 168.805 ;
        RECT -62.045 167.115 -61.715 167.445 ;
        RECT -62.045 165.755 -61.715 166.085 ;
        RECT -62.045 164.395 -61.715 164.725 ;
        RECT -62.045 163.035 -61.715 163.365 ;
        RECT -62.045 161.675 -61.715 162.005 ;
        RECT -62.045 160.315 -61.715 160.645 ;
        RECT -62.045 158.955 -61.715 159.285 ;
        RECT -62.045 157.595 -61.715 157.925 ;
        RECT -62.045 156.235 -61.715 156.565 ;
        RECT -62.045 154.875 -61.715 155.205 ;
        RECT -62.045 153.515 -61.715 153.845 ;
        RECT -62.045 152.155 -61.715 152.485 ;
        RECT -62.045 150.795 -61.715 151.125 ;
        RECT -62.045 149.435 -61.715 149.765 ;
        RECT -62.045 148.075 -61.715 148.405 ;
        RECT -62.045 146.715 -61.715 147.045 ;
        RECT -62.045 145.355 -61.715 145.685 ;
        RECT -62.045 143.995 -61.715 144.325 ;
        RECT -62.045 142.635 -61.715 142.965 ;
        RECT -62.045 141.275 -61.715 141.605 ;
        RECT -62.045 139.915 -61.715 140.245 ;
        RECT -62.045 138.555 -61.715 138.885 ;
        RECT -62.045 137.225 -61.715 137.555 ;
        RECT -62.045 135.175 -61.715 135.505 ;
        RECT -62.045 132.815 -61.715 133.145 ;
        RECT -62.045 131.665 -61.715 131.995 ;
        RECT -62.045 129.655 -61.715 129.985 ;
        RECT -62.045 128.505 -61.715 128.835 ;
        RECT -62.045 126.495 -61.715 126.825 ;
        RECT -62.045 125.345 -61.715 125.675 ;
        RECT -62.045 123.335 -61.715 123.665 ;
        RECT -62.045 122.185 -61.715 122.515 ;
        RECT -62.045 120.175 -61.715 120.505 ;
        RECT -62.045 119.025 -61.715 119.355 ;
        RECT -62.045 117.185 -61.715 117.515 ;
        RECT -62.045 115.865 -61.715 116.195 ;
        RECT -62.045 113.855 -61.715 114.185 ;
        RECT -62.045 112.705 -61.715 113.035 ;
        RECT -62.045 110.695 -61.715 111.025 ;
        RECT -62.045 109.545 -61.715 109.875 ;
        RECT -62.045 107.535 -61.715 107.865 ;
        RECT -62.045 106.385 -61.715 106.715 ;
        RECT -62.045 104.375 -61.715 104.705 ;
        RECT -62.045 103.225 -61.715 103.555 ;
        RECT -62.045 100.865 -61.715 101.195 ;
        RECT -62.045 98.81 -61.715 99.14 ;
        RECT -62.045 97.755 -61.715 98.085 ;
        RECT -62.045 96.395 -61.715 96.725 ;
        RECT -62.045 95.035 -61.715 95.365 ;
        RECT -62.045 93.675 -61.715 94.005 ;
        RECT -62.045 92.315 -61.715 92.645 ;
        RECT -62.045 90.955 -61.715 91.285 ;
        RECT -62.045 89.595 -61.715 89.925 ;
        RECT -62.045 88.235 -61.715 88.565 ;
        RECT -62.045 86.875 -61.715 87.205 ;
        RECT -62.045 85.515 -61.715 85.845 ;
        RECT -62.045 84.155 -61.715 84.485 ;
        RECT -62.045 82.795 -61.715 83.125 ;
        RECT -62.045 81.435 -61.715 81.765 ;
        RECT -62.045 80.075 -61.715 80.405 ;
        RECT -62.045 78.715 -61.715 79.045 ;
        RECT -62.045 77.355 -61.715 77.685 ;
        RECT -62.045 75.995 -61.715 76.325 ;
        RECT -62.045 74.635 -61.715 74.965 ;
        RECT -62.045 73.275 -61.715 73.605 ;
        RECT -62.045 71.915 -61.715 72.245 ;
        RECT -62.045 70.555 -61.715 70.885 ;
        RECT -62.045 69.195 -61.715 69.525 ;
        RECT -62.045 67.835 -61.715 68.165 ;
        RECT -62.045 66.475 -61.715 66.805 ;
        RECT -62.045 65.115 -61.715 65.445 ;
        RECT -62.045 63.755 -61.715 64.085 ;
        RECT -62.045 62.395 -61.715 62.725 ;
        RECT -62.045 61.035 -61.715 61.365 ;
        RECT -62.045 59.675 -61.715 60.005 ;
        RECT -62.045 58.315 -61.715 58.645 ;
        RECT -62.045 56.955 -61.715 57.285 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.565 -122.565 -71.235 -122.235 ;
        RECT -71.565 -123.925 -71.235 -123.595 ;
        RECT -71.565 -125.285 -71.235 -124.955 ;
        RECT -71.565 -126.645 -71.235 -126.315 ;
        RECT -71.565 -128.005 -71.235 -127.675 ;
        RECT -71.565 -129.365 -71.235 -129.035 ;
        RECT -71.565 -130.725 -71.235 -130.395 ;
        RECT -71.565 -132.085 -71.235 -131.755 ;
        RECT -71.565 -133.445 -71.235 -133.115 ;
        RECT -71.565 -134.805 -71.235 -134.475 ;
        RECT -71.565 -136.165 -71.235 -135.835 ;
        RECT -71.565 -137.525 -71.235 -137.195 ;
        RECT -71.565 -138.885 -71.235 -138.555 ;
        RECT -71.565 -140.245 -71.235 -139.915 ;
        RECT -71.565 -141.605 -71.235 -141.275 ;
        RECT -71.565 -142.965 -71.235 -142.635 ;
        RECT -71.565 -144.325 -71.235 -143.995 ;
        RECT -71.565 -145.685 -71.235 -145.355 ;
        RECT -71.565 -147.045 -71.235 -146.715 ;
        RECT -71.565 -148.405 -71.235 -148.075 ;
        RECT -71.565 -149.765 -71.235 -149.435 ;
        RECT -71.565 -151.125 -71.235 -150.795 ;
        RECT -71.565 -152.485 -71.235 -152.155 ;
        RECT -71.565 -153.845 -71.235 -153.515 ;
        RECT -71.565 -155.205 -71.235 -154.875 ;
        RECT -71.565 -156.565 -71.235 -156.235 ;
        RECT -71.565 -157.925 -71.235 -157.595 ;
        RECT -71.565 -159.285 -71.235 -158.955 ;
        RECT -71.565 -160.645 -71.235 -160.315 ;
        RECT -71.565 -162.005 -71.235 -161.675 ;
        RECT -71.565 -163.365 -71.235 -163.035 ;
        RECT -71.565 -164.725 -71.235 -164.395 ;
        RECT -71.565 -166.085 -71.235 -165.755 ;
        RECT -71.565 -167.445 -71.235 -167.115 ;
        RECT -71.565 -168.805 -71.235 -168.475 ;
        RECT -71.565 -171.525 -71.235 -171.195 ;
        RECT -71.56 -171.525 -71.24 -122.235 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.565 -175.605 -71.235 -175.275 ;
        RECT -71.565 -176.685 -71.235 -176.355 ;
        RECT -71.565 -178.325 -71.235 -177.995 ;
        RECT -71.565 -179.685 -71.235 -179.355 ;
        RECT -71.565 -181.93 -71.235 -180.8 ;
        RECT -71.56 -182.045 -71.24 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -70.205 241.32 -69.875 242.45 ;
        RECT -70.205 239.195 -69.875 239.525 ;
        RECT -70.205 237.835 -69.875 238.165 ;
        RECT -70.205 236.475 -69.875 236.805 ;
        RECT -70.205 235.115 -69.875 235.445 ;
        RECT -70.205 233.755 -69.875 234.085 ;
        RECT -70.205 232.395 -69.875 232.725 ;
        RECT -70.205 231.035 -69.875 231.365 ;
        RECT -70.205 229.675 -69.875 230.005 ;
        RECT -70.205 228.315 -69.875 228.645 ;
        RECT -70.205 226.955 -69.875 227.285 ;
        RECT -70.205 225.595 -69.875 225.925 ;
        RECT -70.205 224.235 -69.875 224.565 ;
        RECT -70.205 222.875 -69.875 223.205 ;
        RECT -70.205 221.515 -69.875 221.845 ;
        RECT -70.205 220.155 -69.875 220.485 ;
        RECT -70.205 218.795 -69.875 219.125 ;
        RECT -70.205 217.435 -69.875 217.765 ;
        RECT -70.205 216.075 -69.875 216.405 ;
        RECT -70.205 214.715 -69.875 215.045 ;
        RECT -70.205 213.355 -69.875 213.685 ;
        RECT -70.205 211.995 -69.875 212.325 ;
        RECT -70.205 210.635 -69.875 210.965 ;
        RECT -70.205 209.275 -69.875 209.605 ;
        RECT -70.205 207.915 -69.875 208.245 ;
        RECT -70.205 206.555 -69.875 206.885 ;
        RECT -70.205 205.195 -69.875 205.525 ;
        RECT -70.205 203.835 -69.875 204.165 ;
        RECT -70.205 202.475 -69.875 202.805 ;
        RECT -70.205 201.115 -69.875 201.445 ;
        RECT -70.205 199.755 -69.875 200.085 ;
        RECT -70.205 198.395 -69.875 198.725 ;
        RECT -70.205 197.035 -69.875 197.365 ;
        RECT -70.205 195.675 -69.875 196.005 ;
        RECT -70.205 194.315 -69.875 194.645 ;
        RECT -70.205 192.955 -69.875 193.285 ;
        RECT -70.205 191.595 -69.875 191.925 ;
        RECT -70.205 190.235 -69.875 190.565 ;
        RECT -70.205 188.875 -69.875 189.205 ;
        RECT -70.205 187.515 -69.875 187.845 ;
        RECT -70.205 186.155 -69.875 186.485 ;
        RECT -70.205 184.795 -69.875 185.125 ;
        RECT -70.205 183.435 -69.875 183.765 ;
        RECT -70.205 182.075 -69.875 182.405 ;
        RECT -70.205 180.715 -69.875 181.045 ;
        RECT -70.205 179.355 -69.875 179.685 ;
        RECT -70.205 177.995 -69.875 178.325 ;
        RECT -70.205 176.635 -69.875 176.965 ;
        RECT -70.205 175.275 -69.875 175.605 ;
        RECT -70.205 173.915 -69.875 174.245 ;
        RECT -70.205 172.555 -69.875 172.885 ;
        RECT -70.205 171.195 -69.875 171.525 ;
        RECT -70.205 169.835 -69.875 170.165 ;
        RECT -70.205 168.475 -69.875 168.805 ;
        RECT -70.205 167.115 -69.875 167.445 ;
        RECT -70.205 165.755 -69.875 166.085 ;
        RECT -70.205 164.395 -69.875 164.725 ;
        RECT -70.205 163.035 -69.875 163.365 ;
        RECT -70.205 161.675 -69.875 162.005 ;
        RECT -70.205 160.315 -69.875 160.645 ;
        RECT -70.205 158.955 -69.875 159.285 ;
        RECT -70.205 157.595 -69.875 157.925 ;
        RECT -70.205 156.235 -69.875 156.565 ;
        RECT -70.205 154.875 -69.875 155.205 ;
        RECT -70.205 153.515 -69.875 153.845 ;
        RECT -70.205 152.155 -69.875 152.485 ;
        RECT -70.205 150.795 -69.875 151.125 ;
        RECT -70.205 149.435 -69.875 149.765 ;
        RECT -70.205 148.075 -69.875 148.405 ;
        RECT -70.205 146.715 -69.875 147.045 ;
        RECT -70.205 145.355 -69.875 145.685 ;
        RECT -70.205 143.995 -69.875 144.325 ;
        RECT -70.205 142.635 -69.875 142.965 ;
        RECT -70.205 141.275 -69.875 141.605 ;
        RECT -70.205 139.915 -69.875 140.245 ;
        RECT -70.205 138.555 -69.875 138.885 ;
        RECT -70.205 137.195 -69.875 137.525 ;
        RECT -70.205 135.835 -69.875 136.165 ;
        RECT -70.205 134.475 -69.875 134.805 ;
        RECT -70.205 133.115 -69.875 133.445 ;
        RECT -70.205 131.755 -69.875 132.085 ;
        RECT -70.205 130.395 -69.875 130.725 ;
        RECT -70.205 129.035 -69.875 129.365 ;
        RECT -70.205 127.675 -69.875 128.005 ;
        RECT -70.205 126.315 -69.875 126.645 ;
        RECT -70.205 124.955 -69.875 125.285 ;
        RECT -70.205 123.595 -69.875 123.925 ;
        RECT -70.205 122.235 -69.875 122.565 ;
        RECT -70.205 120.875 -69.875 121.205 ;
        RECT -70.205 119.515 -69.875 119.845 ;
        RECT -70.205 118.155 -69.875 118.485 ;
        RECT -70.205 116.795 -69.875 117.125 ;
        RECT -70.205 115.435 -69.875 115.765 ;
        RECT -70.205 114.075 -69.875 114.405 ;
        RECT -70.205 112.715 -69.875 113.045 ;
        RECT -70.205 111.355 -69.875 111.685 ;
        RECT -70.205 109.995 -69.875 110.325 ;
        RECT -70.205 108.635 -69.875 108.965 ;
        RECT -70.205 107.275 -69.875 107.605 ;
        RECT -70.205 105.915 -69.875 106.245 ;
        RECT -70.205 104.555 -69.875 104.885 ;
        RECT -70.205 103.195 -69.875 103.525 ;
        RECT -70.205 101.835 -69.875 102.165 ;
        RECT -70.205 100.475 -69.875 100.805 ;
        RECT -70.205 99.115 -69.875 99.445 ;
        RECT -70.205 97.755 -69.875 98.085 ;
        RECT -70.205 96.395 -69.875 96.725 ;
        RECT -70.205 95.035 -69.875 95.365 ;
        RECT -70.205 93.675 -69.875 94.005 ;
        RECT -70.205 92.315 -69.875 92.645 ;
        RECT -70.205 90.955 -69.875 91.285 ;
        RECT -70.205 89.595 -69.875 89.925 ;
        RECT -70.205 88.235 -69.875 88.565 ;
        RECT -70.205 86.875 -69.875 87.205 ;
        RECT -70.205 85.515 -69.875 85.845 ;
        RECT -70.205 84.155 -69.875 84.485 ;
        RECT -70.205 82.795 -69.875 83.125 ;
        RECT -70.205 81.435 -69.875 81.765 ;
        RECT -70.205 80.075 -69.875 80.405 ;
        RECT -70.205 78.715 -69.875 79.045 ;
        RECT -70.205 77.355 -69.875 77.685 ;
        RECT -70.205 75.995 -69.875 76.325 ;
        RECT -70.205 74.635 -69.875 74.965 ;
        RECT -70.205 73.275 -69.875 73.605 ;
        RECT -70.205 71.915 -69.875 72.245 ;
        RECT -70.205 70.555 -69.875 70.885 ;
        RECT -70.205 69.195 -69.875 69.525 ;
        RECT -70.205 67.835 -69.875 68.165 ;
        RECT -70.205 66.475 -69.875 66.805 ;
        RECT -70.205 65.115 -69.875 65.445 ;
        RECT -70.205 63.755 -69.875 64.085 ;
        RECT -70.205 62.395 -69.875 62.725 ;
        RECT -70.205 61.035 -69.875 61.365 ;
        RECT -70.205 59.675 -69.875 60.005 ;
        RECT -70.205 58.315 -69.875 58.645 ;
        RECT -70.205 56.955 -69.875 57.285 ;
        RECT -70.205 55.595 -69.875 55.925 ;
        RECT -70.205 54.235 -69.875 54.565 ;
        RECT -70.205 52.875 -69.875 53.205 ;
        RECT -70.205 51.515 -69.875 51.845 ;
        RECT -70.205 50.155 -69.875 50.485 ;
        RECT -70.205 48.795 -69.875 49.125 ;
        RECT -70.205 47.435 -69.875 47.765 ;
        RECT -70.205 46.075 -69.875 46.405 ;
        RECT -70.205 44.715 -69.875 45.045 ;
        RECT -70.205 43.355 -69.875 43.685 ;
        RECT -70.205 41.995 -69.875 42.325 ;
        RECT -70.205 40.635 -69.875 40.965 ;
        RECT -70.205 39.275 -69.875 39.605 ;
        RECT -70.205 37.915 -69.875 38.245 ;
        RECT -70.205 36.555 -69.875 36.885 ;
        RECT -70.205 35.195 -69.875 35.525 ;
        RECT -70.205 33.835 -69.875 34.165 ;
        RECT -70.205 32.475 -69.875 32.805 ;
        RECT -70.205 31.115 -69.875 31.445 ;
        RECT -70.205 29.755 -69.875 30.085 ;
        RECT -70.205 28.395 -69.875 28.725 ;
        RECT -70.205 27.035 -69.875 27.365 ;
        RECT -70.205 25.675 -69.875 26.005 ;
        RECT -70.205 24.315 -69.875 24.645 ;
        RECT -70.205 22.955 -69.875 23.285 ;
        RECT -70.205 21.595 -69.875 21.925 ;
        RECT -70.205 20.235 -69.875 20.565 ;
        RECT -70.205 18.875 -69.875 19.205 ;
        RECT -70.205 17.515 -69.875 17.845 ;
        RECT -70.205 16.155 -69.875 16.485 ;
        RECT -70.205 14.795 -69.875 15.125 ;
        RECT -70.205 13.435 -69.875 13.765 ;
        RECT -70.205 12.075 -69.875 12.405 ;
        RECT -70.205 10.715 -69.875 11.045 ;
        RECT -70.205 9.355 -69.875 9.685 ;
        RECT -70.205 7.995 -69.875 8.325 ;
        RECT -70.205 6.635 -69.875 6.965 ;
        RECT -70.205 5.275 -69.875 5.605 ;
        RECT -70.205 3.915 -69.875 4.245 ;
        RECT -70.205 2.555 -69.875 2.885 ;
        RECT -70.205 1.195 -69.875 1.525 ;
        RECT -70.205 -0.165 -69.875 0.165 ;
        RECT -70.205 -1.525 -69.875 -1.195 ;
        RECT -70.205 -2.885 -69.875 -2.555 ;
        RECT -70.205 -4.245 -69.875 -3.915 ;
        RECT -70.205 -5.605 -69.875 -5.275 ;
        RECT -70.205 -6.965 -69.875 -6.635 ;
        RECT -70.205 -8.325 -69.875 -7.995 ;
        RECT -70.205 -9.685 -69.875 -9.355 ;
        RECT -70.205 -11.045 -69.875 -10.715 ;
        RECT -70.205 -12.405 -69.875 -12.075 ;
        RECT -70.205 -13.765 -69.875 -13.435 ;
        RECT -70.205 -15.125 -69.875 -14.795 ;
        RECT -70.205 -16.485 -69.875 -16.155 ;
        RECT -70.205 -17.845 -69.875 -17.515 ;
        RECT -70.205 -19.205 -69.875 -18.875 ;
        RECT -70.205 -20.565 -69.875 -20.235 ;
        RECT -70.205 -21.925 -69.875 -21.595 ;
        RECT -70.205 -23.285 -69.875 -22.955 ;
        RECT -70.205 -24.645 -69.875 -24.315 ;
        RECT -70.205 -26.005 -69.875 -25.675 ;
        RECT -70.205 -27.365 -69.875 -27.035 ;
        RECT -70.205 -28.725 -69.875 -28.395 ;
        RECT -70.205 -30.085 -69.875 -29.755 ;
        RECT -70.205 -31.445 -69.875 -31.115 ;
        RECT -70.205 -32.805 -69.875 -32.475 ;
        RECT -70.205 -34.165 -69.875 -33.835 ;
        RECT -70.205 -35.525 -69.875 -35.195 ;
        RECT -70.205 -36.885 -69.875 -36.555 ;
        RECT -70.205 -38.245 -69.875 -37.915 ;
        RECT -70.205 -39.605 -69.875 -39.275 ;
        RECT -70.205 -40.965 -69.875 -40.635 ;
        RECT -70.205 -42.325 -69.875 -41.995 ;
        RECT -70.205 -43.685 -69.875 -43.355 ;
        RECT -70.205 -45.045 -69.875 -44.715 ;
        RECT -70.205 -46.405 -69.875 -46.075 ;
        RECT -70.205 -47.765 -69.875 -47.435 ;
        RECT -70.205 -49.125 -69.875 -48.795 ;
        RECT -70.205 -50.485 -69.875 -50.155 ;
        RECT -70.205 -51.845 -69.875 -51.515 ;
        RECT -70.205 -53.205 -69.875 -52.875 ;
        RECT -70.205 -54.565 -69.875 -54.235 ;
        RECT -70.205 -55.925 -69.875 -55.595 ;
        RECT -70.205 -57.285 -69.875 -56.955 ;
        RECT -70.205 -58.645 -69.875 -58.315 ;
        RECT -70.205 -60.005 -69.875 -59.675 ;
        RECT -70.205 -61.365 -69.875 -61.035 ;
        RECT -70.205 -62.725 -69.875 -62.395 ;
        RECT -70.205 -64.085 -69.875 -63.755 ;
        RECT -70.205 -65.445 -69.875 -65.115 ;
        RECT -70.205 -66.805 -69.875 -66.475 ;
        RECT -70.205 -68.165 -69.875 -67.835 ;
        RECT -70.205 -69.525 -69.875 -69.195 ;
        RECT -70.205 -70.885 -69.875 -70.555 ;
        RECT -70.205 -72.245 -69.875 -71.915 ;
        RECT -70.205 -73.605 -69.875 -73.275 ;
        RECT -70.205 -74.965 -69.875 -74.635 ;
        RECT -70.205 -76.325 -69.875 -75.995 ;
        RECT -70.205 -77.685 -69.875 -77.355 ;
        RECT -70.205 -79.045 -69.875 -78.715 ;
        RECT -70.205 -80.405 -69.875 -80.075 ;
        RECT -70.205 -81.765 -69.875 -81.435 ;
        RECT -70.205 -83.125 -69.875 -82.795 ;
        RECT -70.205 -84.485 -69.875 -84.155 ;
        RECT -70.205 -85.845 -69.875 -85.515 ;
        RECT -70.205 -87.205 -69.875 -86.875 ;
        RECT -70.205 -88.565 -69.875 -88.235 ;
        RECT -70.205 -89.925 -69.875 -89.595 ;
        RECT -70.205 -92.645 -69.875 -92.315 ;
        RECT -70.205 -94.005 -69.875 -93.675 ;
        RECT -70.205 -95.365 -69.875 -95.035 ;
        RECT -70.205 -96.725 -69.875 -96.395 ;
        RECT -70.205 -98.085 -69.875 -97.755 ;
        RECT -70.205 -99.69 -69.875 -99.36 ;
        RECT -70.205 -100.805 -69.875 -100.475 ;
        RECT -70.205 -103.525 -69.875 -103.195 ;
        RECT -70.205 -104.885 -69.875 -104.555 ;
        RECT -70.205 -106.245 -69.875 -105.915 ;
        RECT -70.205 -107.83 -69.875 -107.5 ;
        RECT -70.205 -108.965 -69.875 -108.635 ;
        RECT -70.205 -110.325 -69.875 -109.995 ;
        RECT -70.205 -111.685 -69.875 -111.355 ;
        RECT -70.205 -114.405 -69.875 -114.075 ;
        RECT -70.205 -115.765 -69.875 -115.435 ;
        RECT -70.205 -117.125 -69.875 -116.795 ;
        RECT -70.205 -118.485 -69.875 -118.155 ;
        RECT -70.205 -119.845 -69.875 -119.515 ;
        RECT -70.205 -121.205 -69.875 -120.875 ;
        RECT -70.205 -122.565 -69.875 -122.235 ;
        RECT -70.205 -123.925 -69.875 -123.595 ;
        RECT -70.205 -125.285 -69.875 -124.955 ;
        RECT -70.205 -126.645 -69.875 -126.315 ;
        RECT -70.205 -128.005 -69.875 -127.675 ;
        RECT -70.205 -129.365 -69.875 -129.035 ;
        RECT -70.205 -130.725 -69.875 -130.395 ;
        RECT -70.205 -132.085 -69.875 -131.755 ;
        RECT -70.205 -133.445 -69.875 -133.115 ;
        RECT -70.205 -134.805 -69.875 -134.475 ;
        RECT -70.205 -136.165 -69.875 -135.835 ;
        RECT -70.205 -137.525 -69.875 -137.195 ;
        RECT -70.205 -138.885 -69.875 -138.555 ;
        RECT -70.205 -140.245 -69.875 -139.915 ;
        RECT -70.205 -141.605 -69.875 -141.275 ;
        RECT -70.205 -142.965 -69.875 -142.635 ;
        RECT -70.205 -144.325 -69.875 -143.995 ;
        RECT -70.205 -145.685 -69.875 -145.355 ;
        RECT -70.205 -147.045 -69.875 -146.715 ;
        RECT -70.205 -148.405 -69.875 -148.075 ;
        RECT -70.205 -149.765 -69.875 -149.435 ;
        RECT -70.205 -151.125 -69.875 -150.795 ;
        RECT -70.205 -152.485 -69.875 -152.155 ;
        RECT -70.205 -153.845 -69.875 -153.515 ;
        RECT -70.205 -155.205 -69.875 -154.875 ;
        RECT -70.205 -156.565 -69.875 -156.235 ;
        RECT -70.205 -157.925 -69.875 -157.595 ;
        RECT -70.205 -159.285 -69.875 -158.955 ;
        RECT -70.205 -160.645 -69.875 -160.315 ;
        RECT -70.205 -162.005 -69.875 -161.675 ;
        RECT -70.205 -163.365 -69.875 -163.035 ;
        RECT -70.205 -164.725 -69.875 -164.395 ;
        RECT -70.205 -166.085 -69.875 -165.755 ;
        RECT -70.205 -167.445 -69.875 -167.115 ;
        RECT -70.205 -168.805 -69.875 -168.475 ;
        RECT -70.205 -171.525 -69.875 -171.195 ;
        RECT -70.205 -174.245 -69.875 -173.915 ;
        RECT -70.205 -175.605 -69.875 -175.275 ;
        RECT -70.205 -176.685 -69.875 -176.355 ;
        RECT -70.205 -178.325 -69.875 -177.995 ;
        RECT -70.205 -179.685 -69.875 -179.355 ;
        RECT -70.205 -181.93 -69.875 -180.8 ;
        RECT -70.2 -182.045 -69.88 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -68.845 241.32 -68.515 242.45 ;
        RECT -68.845 239.195 -68.515 239.525 ;
        RECT -68.845 237.835 -68.515 238.165 ;
        RECT -68.845 236.475 -68.515 236.805 ;
        RECT -68.845 235.115 -68.515 235.445 ;
        RECT -68.845 233.755 -68.515 234.085 ;
        RECT -68.845 232.395 -68.515 232.725 ;
        RECT -68.845 231.035 -68.515 231.365 ;
        RECT -68.845 229.675 -68.515 230.005 ;
        RECT -68.845 228.315 -68.515 228.645 ;
        RECT -68.845 226.955 -68.515 227.285 ;
        RECT -68.845 225.595 -68.515 225.925 ;
        RECT -68.845 224.235 -68.515 224.565 ;
        RECT -68.845 222.875 -68.515 223.205 ;
        RECT -68.845 221.515 -68.515 221.845 ;
        RECT -68.845 220.155 -68.515 220.485 ;
        RECT -68.845 218.795 -68.515 219.125 ;
        RECT -68.845 217.435 -68.515 217.765 ;
        RECT -68.845 216.075 -68.515 216.405 ;
        RECT -68.845 214.715 -68.515 215.045 ;
        RECT -68.845 213.355 -68.515 213.685 ;
        RECT -68.845 211.995 -68.515 212.325 ;
        RECT -68.845 210.635 -68.515 210.965 ;
        RECT -68.845 209.275 -68.515 209.605 ;
        RECT -68.845 207.915 -68.515 208.245 ;
        RECT -68.845 206.555 -68.515 206.885 ;
        RECT -68.845 205.195 -68.515 205.525 ;
        RECT -68.845 203.835 -68.515 204.165 ;
        RECT -68.845 202.475 -68.515 202.805 ;
        RECT -68.845 201.115 -68.515 201.445 ;
        RECT -68.845 199.755 -68.515 200.085 ;
        RECT -68.845 198.395 -68.515 198.725 ;
        RECT -68.845 197.035 -68.515 197.365 ;
        RECT -68.845 195.675 -68.515 196.005 ;
        RECT -68.845 194.315 -68.515 194.645 ;
        RECT -68.845 192.955 -68.515 193.285 ;
        RECT -68.845 191.595 -68.515 191.925 ;
        RECT -68.845 190.235 -68.515 190.565 ;
        RECT -68.845 188.875 -68.515 189.205 ;
        RECT -68.845 187.515 -68.515 187.845 ;
        RECT -68.845 186.155 -68.515 186.485 ;
        RECT -68.845 184.795 -68.515 185.125 ;
        RECT -68.845 183.435 -68.515 183.765 ;
        RECT -68.845 182.075 -68.515 182.405 ;
        RECT -68.845 180.715 -68.515 181.045 ;
        RECT -68.845 179.355 -68.515 179.685 ;
        RECT -68.845 177.995 -68.515 178.325 ;
        RECT -68.845 176.635 -68.515 176.965 ;
        RECT -68.845 175.275 -68.515 175.605 ;
        RECT -68.845 173.915 -68.515 174.245 ;
        RECT -68.845 172.555 -68.515 172.885 ;
        RECT -68.845 171.195 -68.515 171.525 ;
        RECT -68.845 169.835 -68.515 170.165 ;
        RECT -68.845 168.475 -68.515 168.805 ;
        RECT -68.845 167.115 -68.515 167.445 ;
        RECT -68.845 165.755 -68.515 166.085 ;
        RECT -68.845 164.395 -68.515 164.725 ;
        RECT -68.845 163.035 -68.515 163.365 ;
        RECT -68.845 161.675 -68.515 162.005 ;
        RECT -68.845 160.315 -68.515 160.645 ;
        RECT -68.845 158.955 -68.515 159.285 ;
        RECT -68.845 157.595 -68.515 157.925 ;
        RECT -68.845 156.235 -68.515 156.565 ;
        RECT -68.845 154.875 -68.515 155.205 ;
        RECT -68.845 153.515 -68.515 153.845 ;
        RECT -68.845 152.155 -68.515 152.485 ;
        RECT -68.845 150.795 -68.515 151.125 ;
        RECT -68.845 149.435 -68.515 149.765 ;
        RECT -68.845 148.075 -68.515 148.405 ;
        RECT -68.845 146.715 -68.515 147.045 ;
        RECT -68.845 145.355 -68.515 145.685 ;
        RECT -68.845 143.995 -68.515 144.325 ;
        RECT -68.845 142.635 -68.515 142.965 ;
        RECT -68.845 141.275 -68.515 141.605 ;
        RECT -68.845 139.915 -68.515 140.245 ;
        RECT -68.845 138.555 -68.515 138.885 ;
        RECT -68.845 137.195 -68.515 137.525 ;
        RECT -68.845 135.835 -68.515 136.165 ;
        RECT -68.845 134.475 -68.515 134.805 ;
        RECT -68.845 133.115 -68.515 133.445 ;
        RECT -68.845 131.755 -68.515 132.085 ;
        RECT -68.845 130.395 -68.515 130.725 ;
        RECT -68.845 129.035 -68.515 129.365 ;
        RECT -68.845 127.675 -68.515 128.005 ;
        RECT -68.845 126.315 -68.515 126.645 ;
        RECT -68.845 124.955 -68.515 125.285 ;
        RECT -68.845 123.595 -68.515 123.925 ;
        RECT -68.845 122.235 -68.515 122.565 ;
        RECT -68.845 120.875 -68.515 121.205 ;
        RECT -68.845 119.515 -68.515 119.845 ;
        RECT -68.845 118.155 -68.515 118.485 ;
        RECT -68.845 116.795 -68.515 117.125 ;
        RECT -68.845 115.435 -68.515 115.765 ;
        RECT -68.845 114.075 -68.515 114.405 ;
        RECT -68.845 112.715 -68.515 113.045 ;
        RECT -68.845 111.355 -68.515 111.685 ;
        RECT -68.845 109.995 -68.515 110.325 ;
        RECT -68.845 108.635 -68.515 108.965 ;
        RECT -68.845 107.275 -68.515 107.605 ;
        RECT -68.845 105.915 -68.515 106.245 ;
        RECT -68.845 104.555 -68.515 104.885 ;
        RECT -68.845 103.195 -68.515 103.525 ;
        RECT -68.845 101.835 -68.515 102.165 ;
        RECT -68.845 100.475 -68.515 100.805 ;
        RECT -68.845 99.115 -68.515 99.445 ;
        RECT -68.845 97.755 -68.515 98.085 ;
        RECT -68.845 96.395 -68.515 96.725 ;
        RECT -68.845 95.035 -68.515 95.365 ;
        RECT -68.845 93.675 -68.515 94.005 ;
        RECT -68.845 92.315 -68.515 92.645 ;
        RECT -68.845 90.955 -68.515 91.285 ;
        RECT -68.845 89.595 -68.515 89.925 ;
        RECT -68.845 88.235 -68.515 88.565 ;
        RECT -68.845 86.875 -68.515 87.205 ;
        RECT -68.845 85.515 -68.515 85.845 ;
        RECT -68.845 84.155 -68.515 84.485 ;
        RECT -68.845 82.795 -68.515 83.125 ;
        RECT -68.845 81.435 -68.515 81.765 ;
        RECT -68.845 80.075 -68.515 80.405 ;
        RECT -68.845 78.715 -68.515 79.045 ;
        RECT -68.845 77.355 -68.515 77.685 ;
        RECT -68.845 75.995 -68.515 76.325 ;
        RECT -68.845 74.635 -68.515 74.965 ;
        RECT -68.845 73.275 -68.515 73.605 ;
        RECT -68.845 71.915 -68.515 72.245 ;
        RECT -68.845 70.555 -68.515 70.885 ;
        RECT -68.845 69.195 -68.515 69.525 ;
        RECT -68.845 67.835 -68.515 68.165 ;
        RECT -68.845 66.475 -68.515 66.805 ;
        RECT -68.845 65.115 -68.515 65.445 ;
        RECT -68.845 63.755 -68.515 64.085 ;
        RECT -68.845 62.395 -68.515 62.725 ;
        RECT -68.845 61.035 -68.515 61.365 ;
        RECT -68.845 59.675 -68.515 60.005 ;
        RECT -68.845 58.315 -68.515 58.645 ;
        RECT -68.845 56.955 -68.515 57.285 ;
        RECT -68.845 55.595 -68.515 55.925 ;
        RECT -68.845 54.235 -68.515 54.565 ;
        RECT -68.845 52.875 -68.515 53.205 ;
        RECT -68.845 51.515 -68.515 51.845 ;
        RECT -68.845 50.155 -68.515 50.485 ;
        RECT -68.845 48.795 -68.515 49.125 ;
        RECT -68.845 47.435 -68.515 47.765 ;
        RECT -68.845 46.075 -68.515 46.405 ;
        RECT -68.845 44.715 -68.515 45.045 ;
        RECT -68.845 43.355 -68.515 43.685 ;
        RECT -68.845 41.995 -68.515 42.325 ;
        RECT -68.845 40.635 -68.515 40.965 ;
        RECT -68.845 39.275 -68.515 39.605 ;
        RECT -68.845 37.915 -68.515 38.245 ;
        RECT -68.845 36.555 -68.515 36.885 ;
        RECT -68.845 35.195 -68.515 35.525 ;
        RECT -68.845 33.835 -68.515 34.165 ;
        RECT -68.845 32.475 -68.515 32.805 ;
        RECT -68.845 31.115 -68.515 31.445 ;
        RECT -68.845 29.755 -68.515 30.085 ;
        RECT -68.845 28.395 -68.515 28.725 ;
        RECT -68.845 27.035 -68.515 27.365 ;
        RECT -68.845 25.675 -68.515 26.005 ;
        RECT -68.845 24.315 -68.515 24.645 ;
        RECT -68.845 22.955 -68.515 23.285 ;
        RECT -68.845 21.595 -68.515 21.925 ;
        RECT -68.845 20.235 -68.515 20.565 ;
        RECT -68.845 18.875 -68.515 19.205 ;
        RECT -68.845 17.515 -68.515 17.845 ;
        RECT -68.845 16.155 -68.515 16.485 ;
        RECT -68.845 14.795 -68.515 15.125 ;
        RECT -68.845 13.435 -68.515 13.765 ;
        RECT -68.845 12.075 -68.515 12.405 ;
        RECT -68.845 10.715 -68.515 11.045 ;
        RECT -68.845 9.355 -68.515 9.685 ;
        RECT -68.845 7.995 -68.515 8.325 ;
        RECT -68.845 6.635 -68.515 6.965 ;
        RECT -68.845 5.275 -68.515 5.605 ;
        RECT -68.845 3.915 -68.515 4.245 ;
        RECT -68.845 2.555 -68.515 2.885 ;
        RECT -68.845 1.195 -68.515 1.525 ;
        RECT -68.845 -0.165 -68.515 0.165 ;
        RECT -68.845 -1.525 -68.515 -1.195 ;
        RECT -68.845 -2.885 -68.515 -2.555 ;
        RECT -68.845 -4.245 -68.515 -3.915 ;
        RECT -68.845 -5.605 -68.515 -5.275 ;
        RECT -68.845 -6.965 -68.515 -6.635 ;
        RECT -68.845 -8.325 -68.515 -7.995 ;
        RECT -68.845 -9.685 -68.515 -9.355 ;
        RECT -68.845 -11.045 -68.515 -10.715 ;
        RECT -68.845 -12.405 -68.515 -12.075 ;
        RECT -68.845 -13.765 -68.515 -13.435 ;
        RECT -68.845 -15.125 -68.515 -14.795 ;
        RECT -68.845 -16.485 -68.515 -16.155 ;
        RECT -68.845 -17.845 -68.515 -17.515 ;
        RECT -68.845 -19.205 -68.515 -18.875 ;
        RECT -68.845 -20.565 -68.515 -20.235 ;
        RECT -68.845 -21.925 -68.515 -21.595 ;
        RECT -68.845 -23.285 -68.515 -22.955 ;
        RECT -68.845 -24.645 -68.515 -24.315 ;
        RECT -68.845 -26.005 -68.515 -25.675 ;
        RECT -68.845 -27.365 -68.515 -27.035 ;
        RECT -68.845 -28.725 -68.515 -28.395 ;
        RECT -68.845 -30.085 -68.515 -29.755 ;
        RECT -68.845 -31.445 -68.515 -31.115 ;
        RECT -68.845 -32.805 -68.515 -32.475 ;
        RECT -68.845 -34.165 -68.515 -33.835 ;
        RECT -68.845 -35.525 -68.515 -35.195 ;
        RECT -68.845 -36.885 -68.515 -36.555 ;
        RECT -68.845 -38.245 -68.515 -37.915 ;
        RECT -68.845 -39.605 -68.515 -39.275 ;
        RECT -68.845 -40.965 -68.515 -40.635 ;
        RECT -68.845 -42.325 -68.515 -41.995 ;
        RECT -68.845 -43.685 -68.515 -43.355 ;
        RECT -68.845 -45.045 -68.515 -44.715 ;
        RECT -68.845 -46.405 -68.515 -46.075 ;
        RECT -68.845 -47.765 -68.515 -47.435 ;
        RECT -68.845 -49.125 -68.515 -48.795 ;
        RECT -68.845 -50.485 -68.515 -50.155 ;
        RECT -68.845 -51.845 -68.515 -51.515 ;
        RECT -68.845 -53.205 -68.515 -52.875 ;
        RECT -68.845 -54.565 -68.515 -54.235 ;
        RECT -68.845 -55.925 -68.515 -55.595 ;
        RECT -68.845 -57.285 -68.515 -56.955 ;
        RECT -68.845 -58.645 -68.515 -58.315 ;
        RECT -68.845 -60.005 -68.515 -59.675 ;
        RECT -68.845 -61.365 -68.515 -61.035 ;
        RECT -68.845 -62.725 -68.515 -62.395 ;
        RECT -68.845 -64.085 -68.515 -63.755 ;
        RECT -68.845 -65.445 -68.515 -65.115 ;
        RECT -68.845 -66.805 -68.515 -66.475 ;
        RECT -68.845 -68.165 -68.515 -67.835 ;
        RECT -68.845 -69.525 -68.515 -69.195 ;
        RECT -68.845 -70.885 -68.515 -70.555 ;
        RECT -68.845 -72.245 -68.515 -71.915 ;
        RECT -68.845 -73.605 -68.515 -73.275 ;
        RECT -68.845 -74.965 -68.515 -74.635 ;
        RECT -68.845 -76.325 -68.515 -75.995 ;
        RECT -68.845 -77.685 -68.515 -77.355 ;
        RECT -68.845 -79.045 -68.515 -78.715 ;
        RECT -68.845 -80.405 -68.515 -80.075 ;
        RECT -68.845 -81.765 -68.515 -81.435 ;
        RECT -68.845 -83.125 -68.515 -82.795 ;
        RECT -68.845 -84.485 -68.515 -84.155 ;
        RECT -68.845 -85.845 -68.515 -85.515 ;
        RECT -68.845 -87.205 -68.515 -86.875 ;
        RECT -68.845 -88.565 -68.515 -88.235 ;
        RECT -68.845 -89.925 -68.515 -89.595 ;
        RECT -68.845 -92.645 -68.515 -92.315 ;
        RECT -68.845 -94.005 -68.515 -93.675 ;
        RECT -68.845 -95.365 -68.515 -95.035 ;
        RECT -68.845 -96.725 -68.515 -96.395 ;
        RECT -68.845 -98.085 -68.515 -97.755 ;
        RECT -68.845 -99.69 -68.515 -99.36 ;
        RECT -68.845 -100.805 -68.515 -100.475 ;
        RECT -68.845 -103.525 -68.515 -103.195 ;
        RECT -68.845 -104.885 -68.515 -104.555 ;
        RECT -68.845 -106.245 -68.515 -105.915 ;
        RECT -68.845 -107.83 -68.515 -107.5 ;
        RECT -68.845 -108.965 -68.515 -108.635 ;
        RECT -68.845 -110.325 -68.515 -109.995 ;
        RECT -68.845 -111.685 -68.515 -111.355 ;
        RECT -68.845 -114.405 -68.515 -114.075 ;
        RECT -68.845 -115.765 -68.515 -115.435 ;
        RECT -68.845 -117.125 -68.515 -116.795 ;
        RECT -68.845 -118.485 -68.515 -118.155 ;
        RECT -68.845 -119.845 -68.515 -119.515 ;
        RECT -68.845 -121.205 -68.515 -120.875 ;
        RECT -68.845 -122.565 -68.515 -122.235 ;
        RECT -68.845 -123.925 -68.515 -123.595 ;
        RECT -68.845 -125.285 -68.515 -124.955 ;
        RECT -68.845 -126.645 -68.515 -126.315 ;
        RECT -68.845 -128.005 -68.515 -127.675 ;
        RECT -68.845 -129.365 -68.515 -129.035 ;
        RECT -68.845 -130.725 -68.515 -130.395 ;
        RECT -68.845 -132.085 -68.515 -131.755 ;
        RECT -68.845 -133.445 -68.515 -133.115 ;
        RECT -68.845 -134.805 -68.515 -134.475 ;
        RECT -68.845 -136.165 -68.515 -135.835 ;
        RECT -68.845 -137.525 -68.515 -137.195 ;
        RECT -68.845 -138.885 -68.515 -138.555 ;
        RECT -68.845 -140.245 -68.515 -139.915 ;
        RECT -68.845 -141.605 -68.515 -141.275 ;
        RECT -68.845 -142.965 -68.515 -142.635 ;
        RECT -68.845 -144.325 -68.515 -143.995 ;
        RECT -68.845 -145.685 -68.515 -145.355 ;
        RECT -68.845 -147.045 -68.515 -146.715 ;
        RECT -68.845 -148.405 -68.515 -148.075 ;
        RECT -68.845 -149.765 -68.515 -149.435 ;
        RECT -68.845 -151.125 -68.515 -150.795 ;
        RECT -68.845 -152.485 -68.515 -152.155 ;
        RECT -68.845 -153.845 -68.515 -153.515 ;
        RECT -68.845 -155.205 -68.515 -154.875 ;
        RECT -68.845 -156.565 -68.515 -156.235 ;
        RECT -68.845 -157.925 -68.515 -157.595 ;
        RECT -68.845 -159.285 -68.515 -158.955 ;
        RECT -68.845 -160.645 -68.515 -160.315 ;
        RECT -68.845 -162.005 -68.515 -161.675 ;
        RECT -68.845 -163.365 -68.515 -163.035 ;
        RECT -68.845 -164.725 -68.515 -164.395 ;
        RECT -68.845 -166.085 -68.515 -165.755 ;
        RECT -68.845 -167.445 -68.515 -167.115 ;
        RECT -68.845 -168.805 -68.515 -168.475 ;
        RECT -68.845 -171.525 -68.515 -171.195 ;
        RECT -68.845 -172.885 -68.515 -172.555 ;
        RECT -68.845 -174.245 -68.515 -173.915 ;
        RECT -68.845 -175.605 -68.515 -175.275 ;
        RECT -68.845 -176.685 -68.515 -176.355 ;
        RECT -68.845 -178.325 -68.515 -177.995 ;
        RECT -68.845 -179.685 -68.515 -179.355 ;
        RECT -68.845 -181.93 -68.515 -180.8 ;
        RECT -68.84 -182.045 -68.52 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -67.485 241.32 -67.155 242.45 ;
        RECT -67.485 239.195 -67.155 239.525 ;
        RECT -67.485 237.835 -67.155 238.165 ;
        RECT -67.485 236.475 -67.155 236.805 ;
        RECT -67.485 235.115 -67.155 235.445 ;
        RECT -67.485 233.755 -67.155 234.085 ;
        RECT -67.485 232.395 -67.155 232.725 ;
        RECT -67.485 231.035 -67.155 231.365 ;
        RECT -67.485 229.675 -67.155 230.005 ;
        RECT -67.485 228.315 -67.155 228.645 ;
        RECT -67.485 226.955 -67.155 227.285 ;
        RECT -67.485 225.595 -67.155 225.925 ;
        RECT -67.485 224.235 -67.155 224.565 ;
        RECT -67.485 222.875 -67.155 223.205 ;
        RECT -67.485 221.515 -67.155 221.845 ;
        RECT -67.485 220.155 -67.155 220.485 ;
        RECT -67.485 218.795 -67.155 219.125 ;
        RECT -67.485 217.435 -67.155 217.765 ;
        RECT -67.485 216.075 -67.155 216.405 ;
        RECT -67.485 214.715 -67.155 215.045 ;
        RECT -67.485 213.355 -67.155 213.685 ;
        RECT -67.485 211.995 -67.155 212.325 ;
        RECT -67.485 210.635 -67.155 210.965 ;
        RECT -67.485 209.275 -67.155 209.605 ;
        RECT -67.485 207.915 -67.155 208.245 ;
        RECT -67.485 206.555 -67.155 206.885 ;
        RECT -67.485 205.195 -67.155 205.525 ;
        RECT -67.485 203.835 -67.155 204.165 ;
        RECT -67.485 202.475 -67.155 202.805 ;
        RECT -67.485 201.115 -67.155 201.445 ;
        RECT -67.485 199.755 -67.155 200.085 ;
        RECT -67.485 198.395 -67.155 198.725 ;
        RECT -67.485 197.035 -67.155 197.365 ;
        RECT -67.485 195.675 -67.155 196.005 ;
        RECT -67.485 194.315 -67.155 194.645 ;
        RECT -67.485 192.955 -67.155 193.285 ;
        RECT -67.485 191.595 -67.155 191.925 ;
        RECT -67.485 190.235 -67.155 190.565 ;
        RECT -67.485 188.875 -67.155 189.205 ;
        RECT -67.485 187.515 -67.155 187.845 ;
        RECT -67.485 186.155 -67.155 186.485 ;
        RECT -67.485 184.795 -67.155 185.125 ;
        RECT -67.485 183.435 -67.155 183.765 ;
        RECT -67.485 182.075 -67.155 182.405 ;
        RECT -67.485 180.715 -67.155 181.045 ;
        RECT -67.485 179.355 -67.155 179.685 ;
        RECT -67.485 177.995 -67.155 178.325 ;
        RECT -67.485 176.635 -67.155 176.965 ;
        RECT -67.485 175.275 -67.155 175.605 ;
        RECT -67.485 173.915 -67.155 174.245 ;
        RECT -67.485 172.555 -67.155 172.885 ;
        RECT -67.485 171.195 -67.155 171.525 ;
        RECT -67.485 169.835 -67.155 170.165 ;
        RECT -67.485 168.475 -67.155 168.805 ;
        RECT -67.485 167.115 -67.155 167.445 ;
        RECT -67.485 165.755 -67.155 166.085 ;
        RECT -67.485 164.395 -67.155 164.725 ;
        RECT -67.485 163.035 -67.155 163.365 ;
        RECT -67.485 161.675 -67.155 162.005 ;
        RECT -67.485 160.315 -67.155 160.645 ;
        RECT -67.485 158.955 -67.155 159.285 ;
        RECT -67.485 157.595 -67.155 157.925 ;
        RECT -67.485 156.235 -67.155 156.565 ;
        RECT -67.485 154.875 -67.155 155.205 ;
        RECT -67.485 153.515 -67.155 153.845 ;
        RECT -67.485 152.155 -67.155 152.485 ;
        RECT -67.485 150.795 -67.155 151.125 ;
        RECT -67.485 149.435 -67.155 149.765 ;
        RECT -67.485 148.075 -67.155 148.405 ;
        RECT -67.485 146.715 -67.155 147.045 ;
        RECT -67.485 145.355 -67.155 145.685 ;
        RECT -67.485 143.995 -67.155 144.325 ;
        RECT -67.485 142.635 -67.155 142.965 ;
        RECT -67.485 141.275 -67.155 141.605 ;
        RECT -67.485 139.915 -67.155 140.245 ;
        RECT -67.485 138.555 -67.155 138.885 ;
        RECT -67.485 137.195 -67.155 137.525 ;
        RECT -67.485 135.835 -67.155 136.165 ;
        RECT -67.485 134.475 -67.155 134.805 ;
        RECT -67.485 133.115 -67.155 133.445 ;
        RECT -67.485 131.755 -67.155 132.085 ;
        RECT -67.485 130.395 -67.155 130.725 ;
        RECT -67.485 129.035 -67.155 129.365 ;
        RECT -67.485 127.675 -67.155 128.005 ;
        RECT -67.485 126.315 -67.155 126.645 ;
        RECT -67.485 124.955 -67.155 125.285 ;
        RECT -67.485 123.595 -67.155 123.925 ;
        RECT -67.485 122.235 -67.155 122.565 ;
        RECT -67.485 120.875 -67.155 121.205 ;
        RECT -67.485 119.515 -67.155 119.845 ;
        RECT -67.485 118.155 -67.155 118.485 ;
        RECT -67.485 116.795 -67.155 117.125 ;
        RECT -67.485 115.435 -67.155 115.765 ;
        RECT -67.485 114.075 -67.155 114.405 ;
        RECT -67.485 112.715 -67.155 113.045 ;
        RECT -67.485 111.355 -67.155 111.685 ;
        RECT -67.485 109.995 -67.155 110.325 ;
        RECT -67.485 108.635 -67.155 108.965 ;
        RECT -67.485 107.275 -67.155 107.605 ;
        RECT -67.485 105.915 -67.155 106.245 ;
        RECT -67.485 104.555 -67.155 104.885 ;
        RECT -67.485 103.195 -67.155 103.525 ;
        RECT -67.485 101.835 -67.155 102.165 ;
        RECT -67.485 100.475 -67.155 100.805 ;
        RECT -67.485 99.115 -67.155 99.445 ;
        RECT -67.485 97.755 -67.155 98.085 ;
        RECT -67.485 96.395 -67.155 96.725 ;
        RECT -67.485 95.035 -67.155 95.365 ;
        RECT -67.485 93.675 -67.155 94.005 ;
        RECT -67.485 92.315 -67.155 92.645 ;
        RECT -67.485 90.955 -67.155 91.285 ;
        RECT -67.485 89.595 -67.155 89.925 ;
        RECT -67.485 88.235 -67.155 88.565 ;
        RECT -67.485 86.875 -67.155 87.205 ;
        RECT -67.485 85.515 -67.155 85.845 ;
        RECT -67.485 84.155 -67.155 84.485 ;
        RECT -67.485 82.795 -67.155 83.125 ;
        RECT -67.485 81.435 -67.155 81.765 ;
        RECT -67.485 80.075 -67.155 80.405 ;
        RECT -67.485 78.715 -67.155 79.045 ;
        RECT -67.485 77.355 -67.155 77.685 ;
        RECT -67.485 75.995 -67.155 76.325 ;
        RECT -67.485 74.635 -67.155 74.965 ;
        RECT -67.485 73.275 -67.155 73.605 ;
        RECT -67.485 71.915 -67.155 72.245 ;
        RECT -67.485 70.555 -67.155 70.885 ;
        RECT -67.485 69.195 -67.155 69.525 ;
        RECT -67.485 67.835 -67.155 68.165 ;
        RECT -67.485 66.475 -67.155 66.805 ;
        RECT -67.485 65.115 -67.155 65.445 ;
        RECT -67.485 63.755 -67.155 64.085 ;
        RECT -67.485 62.395 -67.155 62.725 ;
        RECT -67.485 61.035 -67.155 61.365 ;
        RECT -67.485 59.675 -67.155 60.005 ;
        RECT -67.485 58.315 -67.155 58.645 ;
        RECT -67.485 56.955 -67.155 57.285 ;
        RECT -67.485 55.595 -67.155 55.925 ;
        RECT -67.485 54.235 -67.155 54.565 ;
        RECT -67.485 52.875 -67.155 53.205 ;
        RECT -67.485 51.515 -67.155 51.845 ;
        RECT -67.485 50.155 -67.155 50.485 ;
        RECT -67.485 48.795 -67.155 49.125 ;
        RECT -67.485 47.435 -67.155 47.765 ;
        RECT -67.485 46.075 -67.155 46.405 ;
        RECT -67.485 44.715 -67.155 45.045 ;
        RECT -67.485 43.355 -67.155 43.685 ;
        RECT -67.485 41.995 -67.155 42.325 ;
        RECT -67.485 40.635 -67.155 40.965 ;
        RECT -67.485 39.275 -67.155 39.605 ;
        RECT -67.485 37.915 -67.155 38.245 ;
        RECT -67.485 36.555 -67.155 36.885 ;
        RECT -67.485 35.195 -67.155 35.525 ;
        RECT -67.485 33.835 -67.155 34.165 ;
        RECT -67.485 32.475 -67.155 32.805 ;
        RECT -67.485 31.115 -67.155 31.445 ;
        RECT -67.485 29.755 -67.155 30.085 ;
        RECT -67.485 28.395 -67.155 28.725 ;
        RECT -67.485 27.035 -67.155 27.365 ;
        RECT -67.485 25.675 -67.155 26.005 ;
        RECT -67.485 24.315 -67.155 24.645 ;
        RECT -67.485 22.955 -67.155 23.285 ;
        RECT -67.485 21.595 -67.155 21.925 ;
        RECT -67.485 20.235 -67.155 20.565 ;
        RECT -67.485 18.875 -67.155 19.205 ;
        RECT -67.485 17.515 -67.155 17.845 ;
        RECT -67.485 16.155 -67.155 16.485 ;
        RECT -67.485 14.795 -67.155 15.125 ;
        RECT -67.485 13.435 -67.155 13.765 ;
        RECT -67.485 12.075 -67.155 12.405 ;
        RECT -67.485 10.715 -67.155 11.045 ;
        RECT -67.485 9.355 -67.155 9.685 ;
        RECT -67.485 7.995 -67.155 8.325 ;
        RECT -67.485 6.635 -67.155 6.965 ;
        RECT -67.485 5.275 -67.155 5.605 ;
        RECT -67.485 3.915 -67.155 4.245 ;
        RECT -67.485 2.555 -67.155 2.885 ;
        RECT -67.485 1.195 -67.155 1.525 ;
        RECT -67.485 -0.165 -67.155 0.165 ;
        RECT -67.485 -1.525 -67.155 -1.195 ;
        RECT -67.485 -2.885 -67.155 -2.555 ;
        RECT -67.485 -4.245 -67.155 -3.915 ;
        RECT -67.485 -5.605 -67.155 -5.275 ;
        RECT -67.485 -6.965 -67.155 -6.635 ;
        RECT -67.485 -8.325 -67.155 -7.995 ;
        RECT -67.485 -9.685 -67.155 -9.355 ;
        RECT -67.485 -11.045 -67.155 -10.715 ;
        RECT -67.485 -12.405 -67.155 -12.075 ;
        RECT -67.485 -13.765 -67.155 -13.435 ;
        RECT -67.485 -15.125 -67.155 -14.795 ;
        RECT -67.485 -16.485 -67.155 -16.155 ;
        RECT -67.485 -17.845 -67.155 -17.515 ;
        RECT -67.485 -19.205 -67.155 -18.875 ;
        RECT -67.485 -20.565 -67.155 -20.235 ;
        RECT -67.485 -21.925 -67.155 -21.595 ;
        RECT -67.485 -23.285 -67.155 -22.955 ;
        RECT -67.485 -24.645 -67.155 -24.315 ;
        RECT -67.485 -27.365 -67.155 -27.035 ;
        RECT -67.485 -28.725 -67.155 -28.395 ;
        RECT -67.485 -30.085 -67.155 -29.755 ;
        RECT -67.485 -31.445 -67.155 -31.115 ;
        RECT -67.485 -32.805 -67.155 -32.475 ;
        RECT -67.485 -34.165 -67.155 -33.835 ;
        RECT -67.485 -35.525 -67.155 -35.195 ;
        RECT -67.485 -36.885 -67.155 -36.555 ;
        RECT -67.485 -38.245 -67.155 -37.915 ;
        RECT -67.485 -39.605 -67.155 -39.275 ;
        RECT -67.485 -40.965 -67.155 -40.635 ;
        RECT -67.485 -42.325 -67.155 -41.995 ;
        RECT -67.485 -43.685 -67.155 -43.355 ;
        RECT -67.485 -45.045 -67.155 -44.715 ;
        RECT -67.485 -46.405 -67.155 -46.075 ;
        RECT -67.485 -47.765 -67.155 -47.435 ;
        RECT -67.485 -49.125 -67.155 -48.795 ;
        RECT -67.485 -50.485 -67.155 -50.155 ;
        RECT -67.485 -51.845 -67.155 -51.515 ;
        RECT -67.485 -53.205 -67.155 -52.875 ;
        RECT -67.485 -54.565 -67.155 -54.235 ;
        RECT -67.485 -55.925 -67.155 -55.595 ;
        RECT -67.485 -57.285 -67.155 -56.955 ;
        RECT -67.485 -58.645 -67.155 -58.315 ;
        RECT -67.485 -60.005 -67.155 -59.675 ;
        RECT -67.485 -61.365 -67.155 -61.035 ;
        RECT -67.485 -62.725 -67.155 -62.395 ;
        RECT -67.485 -64.085 -67.155 -63.755 ;
        RECT -67.485 -65.445 -67.155 -65.115 ;
        RECT -67.485 -66.805 -67.155 -66.475 ;
        RECT -67.485 -68.165 -67.155 -67.835 ;
        RECT -67.485 -69.525 -67.155 -69.195 ;
        RECT -67.485 -70.885 -67.155 -70.555 ;
        RECT -67.485 -72.245 -67.155 -71.915 ;
        RECT -67.485 -73.605 -67.155 -73.275 ;
        RECT -67.485 -74.965 -67.155 -74.635 ;
        RECT -67.485 -76.325 -67.155 -75.995 ;
        RECT -67.485 -77.685 -67.155 -77.355 ;
        RECT -67.485 -79.045 -67.155 -78.715 ;
        RECT -67.485 -80.405 -67.155 -80.075 ;
        RECT -67.485 -81.765 -67.155 -81.435 ;
        RECT -67.485 -83.125 -67.155 -82.795 ;
        RECT -67.485 -84.485 -67.155 -84.155 ;
        RECT -67.485 -85.845 -67.155 -85.515 ;
        RECT -67.485 -87.205 -67.155 -86.875 ;
        RECT -67.485 -88.565 -67.155 -88.235 ;
        RECT -67.485 -89.925 -67.155 -89.595 ;
        RECT -67.485 -92.645 -67.155 -92.315 ;
        RECT -67.485 -94.005 -67.155 -93.675 ;
        RECT -67.485 -95.365 -67.155 -95.035 ;
        RECT -67.485 -96.725 -67.155 -96.395 ;
        RECT -67.485 -98.085 -67.155 -97.755 ;
        RECT -67.485 -99.69 -67.155 -99.36 ;
        RECT -67.485 -100.805 -67.155 -100.475 ;
        RECT -67.485 -103.525 -67.155 -103.195 ;
        RECT -67.485 -104.885 -67.155 -104.555 ;
        RECT -67.485 -106.245 -67.155 -105.915 ;
        RECT -67.485 -107.83 -67.155 -107.5 ;
        RECT -67.485 -108.965 -67.155 -108.635 ;
        RECT -67.485 -110.325 -67.155 -109.995 ;
        RECT -67.485 -111.685 -67.155 -111.355 ;
        RECT -67.485 -115.765 -67.155 -115.435 ;
        RECT -67.485 -117.125 -67.155 -116.795 ;
        RECT -67.485 -118.485 -67.155 -118.155 ;
        RECT -67.485 -119.845 -67.155 -119.515 ;
        RECT -67.485 -121.205 -67.155 -120.875 ;
        RECT -67.485 -122.565 -67.155 -122.235 ;
        RECT -67.485 -123.925 -67.155 -123.595 ;
        RECT -67.485 -125.285 -67.155 -124.955 ;
        RECT -67.485 -126.645 -67.155 -126.315 ;
        RECT -67.485 -128.005 -67.155 -127.675 ;
        RECT -67.485 -129.365 -67.155 -129.035 ;
        RECT -67.485 -130.725 -67.155 -130.395 ;
        RECT -67.485 -132.085 -67.155 -131.755 ;
        RECT -67.485 -133.445 -67.155 -133.115 ;
        RECT -67.485 -134.805 -67.155 -134.475 ;
        RECT -67.485 -136.165 -67.155 -135.835 ;
        RECT -67.485 -137.525 -67.155 -137.195 ;
        RECT -67.485 -138.885 -67.155 -138.555 ;
        RECT -67.485 -140.245 -67.155 -139.915 ;
        RECT -67.485 -141.605 -67.155 -141.275 ;
        RECT -67.485 -142.965 -67.155 -142.635 ;
        RECT -67.485 -144.325 -67.155 -143.995 ;
        RECT -67.485 -145.685 -67.155 -145.355 ;
        RECT -67.485 -147.045 -67.155 -146.715 ;
        RECT -67.485 -148.405 -67.155 -148.075 ;
        RECT -67.485 -149.765 -67.155 -149.435 ;
        RECT -67.485 -151.125 -67.155 -150.795 ;
        RECT -67.485 -152.485 -67.155 -152.155 ;
        RECT -67.485 -153.845 -67.155 -153.515 ;
        RECT -67.485 -155.205 -67.155 -154.875 ;
        RECT -67.485 -156.565 -67.155 -156.235 ;
        RECT -67.485 -157.925 -67.155 -157.595 ;
        RECT -67.485 -159.285 -67.155 -158.955 ;
        RECT -67.485 -160.645 -67.155 -160.315 ;
        RECT -67.485 -162.005 -67.155 -161.675 ;
        RECT -67.485 -163.365 -67.155 -163.035 ;
        RECT -67.485 -164.725 -67.155 -164.395 ;
        RECT -67.485 -166.085 -67.155 -165.755 ;
        RECT -67.485 -167.445 -67.155 -167.115 ;
        RECT -67.485 -168.805 -67.155 -168.475 ;
        RECT -67.485 -171.525 -67.155 -171.195 ;
        RECT -67.485 -172.885 -67.155 -172.555 ;
        RECT -67.485 -175.605 -67.155 -175.275 ;
        RECT -67.485 -176.685 -67.155 -176.355 ;
        RECT -67.485 -178.325 -67.155 -177.995 ;
        RECT -67.485 -179.685 -67.155 -179.355 ;
        RECT -67.485 -181.93 -67.155 -180.8 ;
        RECT -67.48 -182.045 -67.16 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -66.125 -179.685 -65.795 -179.355 ;
        RECT -66.125 -181.93 -65.795 -180.8 ;
        RECT -66.12 -182.045 -65.8 242.565 ;
        RECT -66.125 241.32 -65.795 242.45 ;
        RECT -66.125 239.195 -65.795 239.525 ;
        RECT -66.125 237.835 -65.795 238.165 ;
        RECT -66.125 236.475 -65.795 236.805 ;
        RECT -66.125 235.115 -65.795 235.445 ;
        RECT -66.125 233.755 -65.795 234.085 ;
        RECT -66.125 232.395 -65.795 232.725 ;
        RECT -66.125 231.035 -65.795 231.365 ;
        RECT -66.125 229.675 -65.795 230.005 ;
        RECT -66.125 228.315 -65.795 228.645 ;
        RECT -66.125 226.955 -65.795 227.285 ;
        RECT -66.125 225.595 -65.795 225.925 ;
        RECT -66.125 224.235 -65.795 224.565 ;
        RECT -66.125 222.875 -65.795 223.205 ;
        RECT -66.125 221.515 -65.795 221.845 ;
        RECT -66.125 220.155 -65.795 220.485 ;
        RECT -66.125 218.795 -65.795 219.125 ;
        RECT -66.125 217.435 -65.795 217.765 ;
        RECT -66.125 216.075 -65.795 216.405 ;
        RECT -66.125 214.715 -65.795 215.045 ;
        RECT -66.125 213.355 -65.795 213.685 ;
        RECT -66.125 211.995 -65.795 212.325 ;
        RECT -66.125 210.635 -65.795 210.965 ;
        RECT -66.125 209.275 -65.795 209.605 ;
        RECT -66.125 207.915 -65.795 208.245 ;
        RECT -66.125 206.555 -65.795 206.885 ;
        RECT -66.125 205.195 -65.795 205.525 ;
        RECT -66.125 203.835 -65.795 204.165 ;
        RECT -66.125 202.475 -65.795 202.805 ;
        RECT -66.125 201.115 -65.795 201.445 ;
        RECT -66.125 199.755 -65.795 200.085 ;
        RECT -66.125 198.395 -65.795 198.725 ;
        RECT -66.125 197.035 -65.795 197.365 ;
        RECT -66.125 195.675 -65.795 196.005 ;
        RECT -66.125 194.315 -65.795 194.645 ;
        RECT -66.125 192.955 -65.795 193.285 ;
        RECT -66.125 191.595 -65.795 191.925 ;
        RECT -66.125 190.235 -65.795 190.565 ;
        RECT -66.125 188.875 -65.795 189.205 ;
        RECT -66.125 187.515 -65.795 187.845 ;
        RECT -66.125 186.155 -65.795 186.485 ;
        RECT -66.125 184.795 -65.795 185.125 ;
        RECT -66.125 183.435 -65.795 183.765 ;
        RECT -66.125 182.075 -65.795 182.405 ;
        RECT -66.125 180.715 -65.795 181.045 ;
        RECT -66.125 179.355 -65.795 179.685 ;
        RECT -66.125 177.995 -65.795 178.325 ;
        RECT -66.125 176.635 -65.795 176.965 ;
        RECT -66.125 175.275 -65.795 175.605 ;
        RECT -66.125 173.915 -65.795 174.245 ;
        RECT -66.125 172.555 -65.795 172.885 ;
        RECT -66.125 171.195 -65.795 171.525 ;
        RECT -66.125 169.835 -65.795 170.165 ;
        RECT -66.125 168.475 -65.795 168.805 ;
        RECT -66.125 167.115 -65.795 167.445 ;
        RECT -66.125 165.755 -65.795 166.085 ;
        RECT -66.125 164.395 -65.795 164.725 ;
        RECT -66.125 163.035 -65.795 163.365 ;
        RECT -66.125 161.675 -65.795 162.005 ;
        RECT -66.125 160.315 -65.795 160.645 ;
        RECT -66.125 158.955 -65.795 159.285 ;
        RECT -66.125 157.595 -65.795 157.925 ;
        RECT -66.125 156.235 -65.795 156.565 ;
        RECT -66.125 154.875 -65.795 155.205 ;
        RECT -66.125 153.515 -65.795 153.845 ;
        RECT -66.125 152.155 -65.795 152.485 ;
        RECT -66.125 150.795 -65.795 151.125 ;
        RECT -66.125 149.435 -65.795 149.765 ;
        RECT -66.125 148.075 -65.795 148.405 ;
        RECT -66.125 146.715 -65.795 147.045 ;
        RECT -66.125 145.355 -65.795 145.685 ;
        RECT -66.125 143.995 -65.795 144.325 ;
        RECT -66.125 142.635 -65.795 142.965 ;
        RECT -66.125 141.275 -65.795 141.605 ;
        RECT -66.125 139.915 -65.795 140.245 ;
        RECT -66.125 138.555 -65.795 138.885 ;
        RECT -66.125 137.195 -65.795 137.525 ;
        RECT -66.125 135.835 -65.795 136.165 ;
        RECT -66.125 134.475 -65.795 134.805 ;
        RECT -66.125 133.115 -65.795 133.445 ;
        RECT -66.125 131.755 -65.795 132.085 ;
        RECT -66.125 130.395 -65.795 130.725 ;
        RECT -66.125 129.035 -65.795 129.365 ;
        RECT -66.125 127.675 -65.795 128.005 ;
        RECT -66.125 126.315 -65.795 126.645 ;
        RECT -66.125 124.955 -65.795 125.285 ;
        RECT -66.125 123.595 -65.795 123.925 ;
        RECT -66.125 122.235 -65.795 122.565 ;
        RECT -66.125 120.875 -65.795 121.205 ;
        RECT -66.125 119.515 -65.795 119.845 ;
        RECT -66.125 118.155 -65.795 118.485 ;
        RECT -66.125 116.795 -65.795 117.125 ;
        RECT -66.125 115.435 -65.795 115.765 ;
        RECT -66.125 114.075 -65.795 114.405 ;
        RECT -66.125 112.715 -65.795 113.045 ;
        RECT -66.125 111.355 -65.795 111.685 ;
        RECT -66.125 109.995 -65.795 110.325 ;
        RECT -66.125 108.635 -65.795 108.965 ;
        RECT -66.125 107.275 -65.795 107.605 ;
        RECT -66.125 105.915 -65.795 106.245 ;
        RECT -66.125 104.555 -65.795 104.885 ;
        RECT -66.125 103.195 -65.795 103.525 ;
        RECT -66.125 101.835 -65.795 102.165 ;
        RECT -66.125 100.475 -65.795 100.805 ;
        RECT -66.125 99.115 -65.795 99.445 ;
        RECT -66.125 97.755 -65.795 98.085 ;
        RECT -66.125 96.395 -65.795 96.725 ;
        RECT -66.125 95.035 -65.795 95.365 ;
        RECT -66.125 93.675 -65.795 94.005 ;
        RECT -66.125 92.315 -65.795 92.645 ;
        RECT -66.125 90.955 -65.795 91.285 ;
        RECT -66.125 89.595 -65.795 89.925 ;
        RECT -66.125 88.235 -65.795 88.565 ;
        RECT -66.125 86.875 -65.795 87.205 ;
        RECT -66.125 85.515 -65.795 85.845 ;
        RECT -66.125 84.155 -65.795 84.485 ;
        RECT -66.125 82.795 -65.795 83.125 ;
        RECT -66.125 81.435 -65.795 81.765 ;
        RECT -66.125 80.075 -65.795 80.405 ;
        RECT -66.125 78.715 -65.795 79.045 ;
        RECT -66.125 77.355 -65.795 77.685 ;
        RECT -66.125 75.995 -65.795 76.325 ;
        RECT -66.125 74.635 -65.795 74.965 ;
        RECT -66.125 73.275 -65.795 73.605 ;
        RECT -66.125 71.915 -65.795 72.245 ;
        RECT -66.125 70.555 -65.795 70.885 ;
        RECT -66.125 69.195 -65.795 69.525 ;
        RECT -66.125 67.835 -65.795 68.165 ;
        RECT -66.125 66.475 -65.795 66.805 ;
        RECT -66.125 65.115 -65.795 65.445 ;
        RECT -66.125 63.755 -65.795 64.085 ;
        RECT -66.125 62.395 -65.795 62.725 ;
        RECT -66.125 61.035 -65.795 61.365 ;
        RECT -66.125 59.675 -65.795 60.005 ;
        RECT -66.125 58.315 -65.795 58.645 ;
        RECT -66.125 56.955 -65.795 57.285 ;
        RECT -66.125 55.595 -65.795 55.925 ;
        RECT -66.125 54.235 -65.795 54.565 ;
        RECT -66.125 52.875 -65.795 53.205 ;
        RECT -66.125 51.515 -65.795 51.845 ;
        RECT -66.125 50.155 -65.795 50.485 ;
        RECT -66.125 48.795 -65.795 49.125 ;
        RECT -66.125 47.435 -65.795 47.765 ;
        RECT -66.125 46.075 -65.795 46.405 ;
        RECT -66.125 44.715 -65.795 45.045 ;
        RECT -66.125 43.355 -65.795 43.685 ;
        RECT -66.125 41.995 -65.795 42.325 ;
        RECT -66.125 40.635 -65.795 40.965 ;
        RECT -66.125 39.275 -65.795 39.605 ;
        RECT -66.125 37.915 -65.795 38.245 ;
        RECT -66.125 36.555 -65.795 36.885 ;
        RECT -66.125 35.195 -65.795 35.525 ;
        RECT -66.125 33.835 -65.795 34.165 ;
        RECT -66.125 32.475 -65.795 32.805 ;
        RECT -66.125 31.115 -65.795 31.445 ;
        RECT -66.125 29.755 -65.795 30.085 ;
        RECT -66.125 28.395 -65.795 28.725 ;
        RECT -66.125 27.035 -65.795 27.365 ;
        RECT -66.125 25.675 -65.795 26.005 ;
        RECT -66.125 24.315 -65.795 24.645 ;
        RECT -66.125 22.955 -65.795 23.285 ;
        RECT -66.125 21.595 -65.795 21.925 ;
        RECT -66.125 20.235 -65.795 20.565 ;
        RECT -66.125 18.875 -65.795 19.205 ;
        RECT -66.125 17.515 -65.795 17.845 ;
        RECT -66.125 16.155 -65.795 16.485 ;
        RECT -66.125 14.795 -65.795 15.125 ;
        RECT -66.125 13.435 -65.795 13.765 ;
        RECT -66.125 12.075 -65.795 12.405 ;
        RECT -66.125 10.715 -65.795 11.045 ;
        RECT -66.125 9.355 -65.795 9.685 ;
        RECT -66.125 7.995 -65.795 8.325 ;
        RECT -66.125 6.635 -65.795 6.965 ;
        RECT -66.125 5.275 -65.795 5.605 ;
        RECT -66.125 3.915 -65.795 4.245 ;
        RECT -66.125 2.555 -65.795 2.885 ;
        RECT -66.125 1.195 -65.795 1.525 ;
        RECT -66.125 -0.165 -65.795 0.165 ;
        RECT -66.125 -1.525 -65.795 -1.195 ;
        RECT -66.125 -2.885 -65.795 -2.555 ;
        RECT -66.125 -4.245 -65.795 -3.915 ;
        RECT -66.125 -5.605 -65.795 -5.275 ;
        RECT -66.125 -6.965 -65.795 -6.635 ;
        RECT -66.125 -8.325 -65.795 -7.995 ;
        RECT -66.125 -9.685 -65.795 -9.355 ;
        RECT -66.125 -11.045 -65.795 -10.715 ;
        RECT -66.125 -12.405 -65.795 -12.075 ;
        RECT -66.125 -13.765 -65.795 -13.435 ;
        RECT -66.125 -15.125 -65.795 -14.795 ;
        RECT -66.125 -16.485 -65.795 -16.155 ;
        RECT -66.125 -17.845 -65.795 -17.515 ;
        RECT -66.125 -19.205 -65.795 -18.875 ;
        RECT -66.125 -20.565 -65.795 -20.235 ;
        RECT -66.125 -21.925 -65.795 -21.595 ;
        RECT -66.125 -23.285 -65.795 -22.955 ;
        RECT -66.125 -24.645 -65.795 -24.315 ;
        RECT -66.125 -27.365 -65.795 -27.035 ;
        RECT -66.125 -28.725 -65.795 -28.395 ;
        RECT -66.125 -30.085 -65.795 -29.755 ;
        RECT -66.125 -31.445 -65.795 -31.115 ;
        RECT -66.125 -32.805 -65.795 -32.475 ;
        RECT -66.125 -34.165 -65.795 -33.835 ;
        RECT -66.125 -35.525 -65.795 -35.195 ;
        RECT -66.125 -36.885 -65.795 -36.555 ;
        RECT -66.125 -38.245 -65.795 -37.915 ;
        RECT -66.125 -39.605 -65.795 -39.275 ;
        RECT -66.125 -40.965 -65.795 -40.635 ;
        RECT -66.125 -42.325 -65.795 -41.995 ;
        RECT -66.125 -43.685 -65.795 -43.355 ;
        RECT -66.125 -45.045 -65.795 -44.715 ;
        RECT -66.125 -46.405 -65.795 -46.075 ;
        RECT -66.125 -47.765 -65.795 -47.435 ;
        RECT -66.125 -49.125 -65.795 -48.795 ;
        RECT -66.125 -50.485 -65.795 -50.155 ;
        RECT -66.125 -51.845 -65.795 -51.515 ;
        RECT -66.125 -53.205 -65.795 -52.875 ;
        RECT -66.125 -54.565 -65.795 -54.235 ;
        RECT -66.125 -55.925 -65.795 -55.595 ;
        RECT -66.125 -57.285 -65.795 -56.955 ;
        RECT -66.125 -58.645 -65.795 -58.315 ;
        RECT -66.125 -60.005 -65.795 -59.675 ;
        RECT -66.125 -61.365 -65.795 -61.035 ;
        RECT -66.125 -62.725 -65.795 -62.395 ;
        RECT -66.125 -64.085 -65.795 -63.755 ;
        RECT -66.125 -65.445 -65.795 -65.115 ;
        RECT -66.125 -66.805 -65.795 -66.475 ;
        RECT -66.125 -68.165 -65.795 -67.835 ;
        RECT -66.125 -69.525 -65.795 -69.195 ;
        RECT -66.125 -70.885 -65.795 -70.555 ;
        RECT -66.125 -72.245 -65.795 -71.915 ;
        RECT -66.125 -73.605 -65.795 -73.275 ;
        RECT -66.125 -74.965 -65.795 -74.635 ;
        RECT -66.125 -76.325 -65.795 -75.995 ;
        RECT -66.125 -77.685 -65.795 -77.355 ;
        RECT -66.125 -79.045 -65.795 -78.715 ;
        RECT -66.125 -80.405 -65.795 -80.075 ;
        RECT -66.125 -81.765 -65.795 -81.435 ;
        RECT -66.125 -83.125 -65.795 -82.795 ;
        RECT -66.125 -84.485 -65.795 -84.155 ;
        RECT -66.125 -85.845 -65.795 -85.515 ;
        RECT -66.125 -87.205 -65.795 -86.875 ;
        RECT -66.125 -88.565 -65.795 -88.235 ;
        RECT -66.125 -89.925 -65.795 -89.595 ;
        RECT -66.125 -92.645 -65.795 -92.315 ;
        RECT -66.125 -94.005 -65.795 -93.675 ;
        RECT -66.125 -95.365 -65.795 -95.035 ;
        RECT -66.125 -96.725 -65.795 -96.395 ;
        RECT -66.125 -98.085 -65.795 -97.755 ;
        RECT -66.125 -99.69 -65.795 -99.36 ;
        RECT -66.125 -100.805 -65.795 -100.475 ;
        RECT -66.125 -103.525 -65.795 -103.195 ;
        RECT -66.125 -104.885 -65.795 -104.555 ;
        RECT -66.125 -106.245 -65.795 -105.915 ;
        RECT -66.125 -107.83 -65.795 -107.5 ;
        RECT -66.125 -108.965 -65.795 -108.635 ;
        RECT -66.125 -110.325 -65.795 -109.995 ;
        RECT -66.125 -111.685 -65.795 -111.355 ;
        RECT -66.125 -114.405 -65.795 -114.075 ;
        RECT -66.125 -115.765 -65.795 -115.435 ;
        RECT -66.125 -117.125 -65.795 -116.795 ;
        RECT -66.125 -118.485 -65.795 -118.155 ;
        RECT -66.125 -119.845 -65.795 -119.515 ;
        RECT -66.125 -121.205 -65.795 -120.875 ;
        RECT -66.125 -122.565 -65.795 -122.235 ;
        RECT -66.125 -123.925 -65.795 -123.595 ;
        RECT -66.125 -125.285 -65.795 -124.955 ;
        RECT -66.125 -126.645 -65.795 -126.315 ;
        RECT -66.125 -128.005 -65.795 -127.675 ;
        RECT -66.125 -129.365 -65.795 -129.035 ;
        RECT -66.125 -130.725 -65.795 -130.395 ;
        RECT -66.125 -132.085 -65.795 -131.755 ;
        RECT -66.125 -133.445 -65.795 -133.115 ;
        RECT -66.125 -134.805 -65.795 -134.475 ;
        RECT -66.125 -136.165 -65.795 -135.835 ;
        RECT -66.125 -137.525 -65.795 -137.195 ;
        RECT -66.125 -138.885 -65.795 -138.555 ;
        RECT -66.125 -140.245 -65.795 -139.915 ;
        RECT -66.125 -141.605 -65.795 -141.275 ;
        RECT -66.125 -142.965 -65.795 -142.635 ;
        RECT -66.125 -144.325 -65.795 -143.995 ;
        RECT -66.125 -145.685 -65.795 -145.355 ;
        RECT -66.125 -147.045 -65.795 -146.715 ;
        RECT -66.125 -148.405 -65.795 -148.075 ;
        RECT -66.125 -149.765 -65.795 -149.435 ;
        RECT -66.125 -151.125 -65.795 -150.795 ;
        RECT -66.125 -152.485 -65.795 -152.155 ;
        RECT -66.125 -153.845 -65.795 -153.515 ;
        RECT -66.125 -155.205 -65.795 -154.875 ;
        RECT -66.125 -156.565 -65.795 -156.235 ;
        RECT -66.125 -157.925 -65.795 -157.595 ;
        RECT -66.125 -159.285 -65.795 -158.955 ;
        RECT -66.125 -160.645 -65.795 -160.315 ;
        RECT -66.125 -162.005 -65.795 -161.675 ;
        RECT -66.125 -163.365 -65.795 -163.035 ;
        RECT -66.125 -164.725 -65.795 -164.395 ;
        RECT -66.125 -166.085 -65.795 -165.755 ;
        RECT -66.125 -167.445 -65.795 -167.115 ;
        RECT -66.125 -168.805 -65.795 -168.475 ;
        RECT -66.125 -171.525 -65.795 -171.195 ;
        RECT -66.125 -175.605 -65.795 -175.275 ;
        RECT -66.125 -178.325 -65.795 -177.995 ;
    END
    PORT
      LAYER met3 ;
        RECT -74.285 241.32 -73.955 242.45 ;
        RECT -74.285 239.195 -73.955 239.525 ;
        RECT -74.285 237.835 -73.955 238.165 ;
        RECT -74.285 236.475 -73.955 236.805 ;
        RECT -74.285 235.115 -73.955 235.445 ;
        RECT -74.285 233.755 -73.955 234.085 ;
        RECT -74.285 232.395 -73.955 232.725 ;
        RECT -74.285 231.035 -73.955 231.365 ;
        RECT -74.285 229.675 -73.955 230.005 ;
        RECT -74.285 228.315 -73.955 228.645 ;
        RECT -74.285 226.955 -73.955 227.285 ;
        RECT -74.285 225.595 -73.955 225.925 ;
        RECT -74.285 224.235 -73.955 224.565 ;
        RECT -74.285 222.875 -73.955 223.205 ;
        RECT -74.285 221.515 -73.955 221.845 ;
        RECT -74.285 220.155 -73.955 220.485 ;
        RECT -74.285 218.795 -73.955 219.125 ;
        RECT -74.285 217.435 -73.955 217.765 ;
        RECT -74.285 216.075 -73.955 216.405 ;
        RECT -74.285 214.715 -73.955 215.045 ;
        RECT -74.285 213.355 -73.955 213.685 ;
        RECT -74.285 211.995 -73.955 212.325 ;
        RECT -74.285 210.635 -73.955 210.965 ;
        RECT -74.285 209.275 -73.955 209.605 ;
        RECT -74.285 207.915 -73.955 208.245 ;
        RECT -74.285 206.555 -73.955 206.885 ;
        RECT -74.285 205.195 -73.955 205.525 ;
        RECT -74.285 203.835 -73.955 204.165 ;
        RECT -74.285 202.475 -73.955 202.805 ;
        RECT -74.285 201.115 -73.955 201.445 ;
        RECT -74.285 199.755 -73.955 200.085 ;
        RECT -74.285 198.395 -73.955 198.725 ;
        RECT -74.285 197.035 -73.955 197.365 ;
        RECT -74.285 195.675 -73.955 196.005 ;
        RECT -74.285 194.315 -73.955 194.645 ;
        RECT -74.285 192.955 -73.955 193.285 ;
        RECT -74.285 191.595 -73.955 191.925 ;
        RECT -74.285 190.235 -73.955 190.565 ;
        RECT -74.285 188.875 -73.955 189.205 ;
        RECT -74.285 187.515 -73.955 187.845 ;
        RECT -74.285 186.155 -73.955 186.485 ;
        RECT -74.285 184.795 -73.955 185.125 ;
        RECT -74.285 183.435 -73.955 183.765 ;
        RECT -74.285 182.075 -73.955 182.405 ;
        RECT -74.285 180.715 -73.955 181.045 ;
        RECT -74.285 179.355 -73.955 179.685 ;
        RECT -74.285 177.995 -73.955 178.325 ;
        RECT -74.285 176.635 -73.955 176.965 ;
        RECT -74.285 175.275 -73.955 175.605 ;
        RECT -74.285 173.915 -73.955 174.245 ;
        RECT -74.285 172.555 -73.955 172.885 ;
        RECT -74.285 171.195 -73.955 171.525 ;
        RECT -74.285 169.835 -73.955 170.165 ;
        RECT -74.285 168.475 -73.955 168.805 ;
        RECT -74.285 167.115 -73.955 167.445 ;
        RECT -74.285 165.755 -73.955 166.085 ;
        RECT -74.285 164.395 -73.955 164.725 ;
        RECT -74.285 163.035 -73.955 163.365 ;
        RECT -74.285 161.675 -73.955 162.005 ;
        RECT -74.285 160.315 -73.955 160.645 ;
        RECT -74.285 158.955 -73.955 159.285 ;
        RECT -74.285 157.595 -73.955 157.925 ;
        RECT -74.285 156.235 -73.955 156.565 ;
        RECT -74.285 154.875 -73.955 155.205 ;
        RECT -74.285 153.515 -73.955 153.845 ;
        RECT -74.285 152.155 -73.955 152.485 ;
        RECT -74.285 150.795 -73.955 151.125 ;
        RECT -74.285 149.435 -73.955 149.765 ;
        RECT -74.285 148.075 -73.955 148.405 ;
        RECT -74.285 146.715 -73.955 147.045 ;
        RECT -74.285 145.355 -73.955 145.685 ;
        RECT -74.285 143.995 -73.955 144.325 ;
        RECT -74.285 142.635 -73.955 142.965 ;
        RECT -74.285 141.275 -73.955 141.605 ;
        RECT -74.285 139.915 -73.955 140.245 ;
        RECT -74.285 138.555 -73.955 138.885 ;
        RECT -74.285 137.195 -73.955 137.525 ;
        RECT -74.285 135.835 -73.955 136.165 ;
        RECT -74.285 134.475 -73.955 134.805 ;
        RECT -74.285 133.115 -73.955 133.445 ;
        RECT -74.285 131.755 -73.955 132.085 ;
        RECT -74.285 130.395 -73.955 130.725 ;
        RECT -74.285 129.035 -73.955 129.365 ;
        RECT -74.285 127.675 -73.955 128.005 ;
        RECT -74.285 126.315 -73.955 126.645 ;
        RECT -74.285 124.955 -73.955 125.285 ;
        RECT -74.285 123.595 -73.955 123.925 ;
        RECT -74.285 122.235 -73.955 122.565 ;
        RECT -74.285 120.875 -73.955 121.205 ;
        RECT -74.285 119.515 -73.955 119.845 ;
        RECT -74.285 118.155 -73.955 118.485 ;
        RECT -74.285 116.795 -73.955 117.125 ;
        RECT -74.285 115.435 -73.955 115.765 ;
        RECT -74.285 114.075 -73.955 114.405 ;
        RECT -74.285 112.715 -73.955 113.045 ;
        RECT -74.285 111.355 -73.955 111.685 ;
        RECT -74.285 109.995 -73.955 110.325 ;
        RECT -74.285 108.635 -73.955 108.965 ;
        RECT -74.285 107.275 -73.955 107.605 ;
        RECT -74.285 105.915 -73.955 106.245 ;
        RECT -74.285 104.555 -73.955 104.885 ;
        RECT -74.285 103.195 -73.955 103.525 ;
        RECT -74.285 101.835 -73.955 102.165 ;
        RECT -74.285 100.475 -73.955 100.805 ;
        RECT -74.285 99.115 -73.955 99.445 ;
        RECT -74.285 97.755 -73.955 98.085 ;
        RECT -74.285 96.395 -73.955 96.725 ;
        RECT -74.285 95.035 -73.955 95.365 ;
        RECT -74.285 93.675 -73.955 94.005 ;
        RECT -74.285 92.315 -73.955 92.645 ;
        RECT -74.285 90.955 -73.955 91.285 ;
        RECT -74.285 89.595 -73.955 89.925 ;
        RECT -74.285 88.235 -73.955 88.565 ;
        RECT -74.285 86.875 -73.955 87.205 ;
        RECT -74.285 85.515 -73.955 85.845 ;
        RECT -74.285 84.155 -73.955 84.485 ;
        RECT -74.285 82.795 -73.955 83.125 ;
        RECT -74.285 81.435 -73.955 81.765 ;
        RECT -74.285 80.075 -73.955 80.405 ;
        RECT -74.285 78.715 -73.955 79.045 ;
        RECT -74.285 77.355 -73.955 77.685 ;
        RECT -74.285 75.995 -73.955 76.325 ;
        RECT -74.285 74.635 -73.955 74.965 ;
        RECT -74.285 73.275 -73.955 73.605 ;
        RECT -74.285 71.915 -73.955 72.245 ;
        RECT -74.285 70.555 -73.955 70.885 ;
        RECT -74.285 69.195 -73.955 69.525 ;
        RECT -74.285 67.835 -73.955 68.165 ;
        RECT -74.285 66.475 -73.955 66.805 ;
        RECT -74.285 65.115 -73.955 65.445 ;
        RECT -74.285 63.755 -73.955 64.085 ;
        RECT -74.285 62.395 -73.955 62.725 ;
        RECT -74.285 61.035 -73.955 61.365 ;
        RECT -74.285 59.675 -73.955 60.005 ;
        RECT -74.285 58.315 -73.955 58.645 ;
        RECT -74.285 56.955 -73.955 57.285 ;
        RECT -74.285 55.595 -73.955 55.925 ;
        RECT -74.285 54.235 -73.955 54.565 ;
        RECT -74.285 52.875 -73.955 53.205 ;
        RECT -74.285 51.515 -73.955 51.845 ;
        RECT -74.285 50.155 -73.955 50.485 ;
        RECT -74.285 48.795 -73.955 49.125 ;
        RECT -74.285 47.435 -73.955 47.765 ;
        RECT -74.285 46.075 -73.955 46.405 ;
        RECT -74.285 44.715 -73.955 45.045 ;
        RECT -74.285 43.355 -73.955 43.685 ;
        RECT -74.285 41.995 -73.955 42.325 ;
        RECT -74.285 40.635 -73.955 40.965 ;
        RECT -74.285 39.275 -73.955 39.605 ;
        RECT -74.285 37.915 -73.955 38.245 ;
        RECT -74.285 36.555 -73.955 36.885 ;
        RECT -74.285 35.195 -73.955 35.525 ;
        RECT -74.285 33.835 -73.955 34.165 ;
        RECT -74.285 32.475 -73.955 32.805 ;
        RECT -74.285 31.115 -73.955 31.445 ;
        RECT -74.285 29.755 -73.955 30.085 ;
        RECT -74.285 28.395 -73.955 28.725 ;
        RECT -74.285 27.035 -73.955 27.365 ;
        RECT -74.285 25.675 -73.955 26.005 ;
        RECT -74.285 24.315 -73.955 24.645 ;
        RECT -74.285 22.955 -73.955 23.285 ;
        RECT -74.285 21.595 -73.955 21.925 ;
        RECT -74.285 20.235 -73.955 20.565 ;
        RECT -74.285 18.875 -73.955 19.205 ;
        RECT -74.285 17.515 -73.955 17.845 ;
        RECT -74.285 16.155 -73.955 16.485 ;
        RECT -74.285 14.795 -73.955 15.125 ;
        RECT -74.285 13.435 -73.955 13.765 ;
        RECT -74.285 12.075 -73.955 12.405 ;
        RECT -74.285 10.715 -73.955 11.045 ;
        RECT -74.285 9.355 -73.955 9.685 ;
        RECT -74.285 7.995 -73.955 8.325 ;
        RECT -74.285 6.635 -73.955 6.965 ;
        RECT -74.285 5.275 -73.955 5.605 ;
        RECT -74.285 3.915 -73.955 4.245 ;
        RECT -74.285 2.555 -73.955 2.885 ;
        RECT -74.285 1.195 -73.955 1.525 ;
        RECT -74.285 -0.165 -73.955 0.165 ;
        RECT -74.285 -1.525 -73.955 -1.195 ;
        RECT -74.285 -2.885 -73.955 -2.555 ;
        RECT -74.285 -4.245 -73.955 -3.915 ;
        RECT -74.285 -5.605 -73.955 -5.275 ;
        RECT -74.285 -6.965 -73.955 -6.635 ;
        RECT -74.285 -8.325 -73.955 -7.995 ;
        RECT -74.285 -9.685 -73.955 -9.355 ;
        RECT -74.285 -11.045 -73.955 -10.715 ;
        RECT -74.285 -12.405 -73.955 -12.075 ;
        RECT -74.285 -13.765 -73.955 -13.435 ;
        RECT -74.285 -15.125 -73.955 -14.795 ;
        RECT -74.285 -16.485 -73.955 -16.155 ;
        RECT -74.285 -17.845 -73.955 -17.515 ;
        RECT -74.285 -19.205 -73.955 -18.875 ;
        RECT -74.285 -20.565 -73.955 -20.235 ;
        RECT -74.285 -21.925 -73.955 -21.595 ;
        RECT -74.285 -23.285 -73.955 -22.955 ;
        RECT -74.285 -24.645 -73.955 -24.315 ;
        RECT -74.285 -26.005 -73.955 -25.675 ;
        RECT -74.285 -27.365 -73.955 -27.035 ;
        RECT -74.285 -28.725 -73.955 -28.395 ;
        RECT -74.285 -30.085 -73.955 -29.755 ;
        RECT -74.285 -31.445 -73.955 -31.115 ;
        RECT -74.285 -32.805 -73.955 -32.475 ;
        RECT -74.285 -34.165 -73.955 -33.835 ;
        RECT -74.285 -35.525 -73.955 -35.195 ;
        RECT -74.285 -36.885 -73.955 -36.555 ;
        RECT -74.285 -38.245 -73.955 -37.915 ;
        RECT -74.285 -39.605 -73.955 -39.275 ;
        RECT -74.285 -40.965 -73.955 -40.635 ;
        RECT -74.285 -42.325 -73.955 -41.995 ;
        RECT -74.285 -43.685 -73.955 -43.355 ;
        RECT -74.285 -45.045 -73.955 -44.715 ;
        RECT -74.285 -46.405 -73.955 -46.075 ;
        RECT -74.285 -47.765 -73.955 -47.435 ;
        RECT -74.285 -49.125 -73.955 -48.795 ;
        RECT -74.285 -50.485 -73.955 -50.155 ;
        RECT -74.285 -51.845 -73.955 -51.515 ;
        RECT -74.285 -53.205 -73.955 -52.875 ;
        RECT -74.285 -54.565 -73.955 -54.235 ;
        RECT -74.285 -55.925 -73.955 -55.595 ;
        RECT -74.285 -57.285 -73.955 -56.955 ;
        RECT -74.285 -58.645 -73.955 -58.315 ;
        RECT -74.285 -60.005 -73.955 -59.675 ;
        RECT -74.285 -61.365 -73.955 -61.035 ;
        RECT -74.285 -62.725 -73.955 -62.395 ;
        RECT -74.285 -64.085 -73.955 -63.755 ;
        RECT -74.285 -65.445 -73.955 -65.115 ;
        RECT -74.285 -66.805 -73.955 -66.475 ;
        RECT -74.285 -68.165 -73.955 -67.835 ;
        RECT -74.285 -69.525 -73.955 -69.195 ;
        RECT -74.285 -70.885 -73.955 -70.555 ;
        RECT -74.285 -72.245 -73.955 -71.915 ;
        RECT -74.285 -73.605 -73.955 -73.275 ;
        RECT -74.285 -74.965 -73.955 -74.635 ;
        RECT -74.285 -76.325 -73.955 -75.995 ;
        RECT -74.285 -77.685 -73.955 -77.355 ;
        RECT -74.285 -79.045 -73.955 -78.715 ;
        RECT -74.285 -80.405 -73.955 -80.075 ;
        RECT -74.285 -81.765 -73.955 -81.435 ;
        RECT -74.285 -83.125 -73.955 -82.795 ;
        RECT -74.285 -84.485 -73.955 -84.155 ;
        RECT -74.285 -85.845 -73.955 -85.515 ;
        RECT -74.285 -87.205 -73.955 -86.875 ;
        RECT -74.285 -88.565 -73.955 -88.235 ;
        RECT -74.285 -89.925 -73.955 -89.595 ;
        RECT -74.285 -91.285 -73.955 -90.955 ;
        RECT -74.285 -92.645 -73.955 -92.315 ;
        RECT -74.285 -94.005 -73.955 -93.675 ;
        RECT -74.285 -95.365 -73.955 -95.035 ;
        RECT -74.285 -96.725 -73.955 -96.395 ;
        RECT -74.285 -98.085 -73.955 -97.755 ;
        RECT -74.285 -99.445 -73.955 -99.115 ;
        RECT -74.285 -100.805 -73.955 -100.475 ;
        RECT -74.285 -102.165 -73.955 -101.835 ;
        RECT -74.285 -103.525 -73.955 -103.195 ;
        RECT -74.285 -104.885 -73.955 -104.555 ;
        RECT -74.285 -106.245 -73.955 -105.915 ;
        RECT -74.285 -107.605 -73.955 -107.275 ;
        RECT -74.285 -108.965 -73.955 -108.635 ;
        RECT -74.285 -110.325 -73.955 -109.995 ;
        RECT -74.285 -111.685 -73.955 -111.355 ;
        RECT -74.285 -113.045 -73.955 -112.715 ;
        RECT -74.285 -114.405 -73.955 -114.075 ;
        RECT -74.285 -115.765 -73.955 -115.435 ;
        RECT -74.285 -117.125 -73.955 -116.795 ;
        RECT -74.285 -118.485 -73.955 -118.155 ;
        RECT -74.285 -119.845 -73.955 -119.515 ;
        RECT -74.285 -121.205 -73.955 -120.875 ;
        RECT -74.285 -122.565 -73.955 -122.235 ;
        RECT -74.285 -123.925 -73.955 -123.595 ;
        RECT -74.285 -125.285 -73.955 -124.955 ;
        RECT -74.285 -126.645 -73.955 -126.315 ;
        RECT -74.285 -128.005 -73.955 -127.675 ;
        RECT -74.285 -129.365 -73.955 -129.035 ;
        RECT -74.285 -130.725 -73.955 -130.395 ;
        RECT -74.285 -132.085 -73.955 -131.755 ;
        RECT -74.285 -133.445 -73.955 -133.115 ;
        RECT -74.285 -134.805 -73.955 -134.475 ;
        RECT -74.285 -136.165 -73.955 -135.835 ;
        RECT -74.285 -137.525 -73.955 -137.195 ;
        RECT -74.285 -138.885 -73.955 -138.555 ;
        RECT -74.285 -140.245 -73.955 -139.915 ;
        RECT -74.285 -141.605 -73.955 -141.275 ;
        RECT -74.285 -142.965 -73.955 -142.635 ;
        RECT -74.285 -144.325 -73.955 -143.995 ;
        RECT -74.285 -145.685 -73.955 -145.355 ;
        RECT -74.285 -147.045 -73.955 -146.715 ;
        RECT -74.285 -148.405 -73.955 -148.075 ;
        RECT -74.285 -149.765 -73.955 -149.435 ;
        RECT -74.285 -151.125 -73.955 -150.795 ;
        RECT -74.285 -152.485 -73.955 -152.155 ;
        RECT -74.285 -153.845 -73.955 -153.515 ;
        RECT -74.285 -155.205 -73.955 -154.875 ;
        RECT -74.285 -156.565 -73.955 -156.235 ;
        RECT -74.285 -157.925 -73.955 -157.595 ;
        RECT -74.285 -159.285 -73.955 -158.955 ;
        RECT -74.285 -160.645 -73.955 -160.315 ;
        RECT -74.285 -162.005 -73.955 -161.675 ;
        RECT -74.285 -163.365 -73.955 -163.035 ;
        RECT -74.285 -164.725 -73.955 -164.395 ;
        RECT -74.285 -166.085 -73.955 -165.755 ;
        RECT -74.285 -167.445 -73.955 -167.115 ;
        RECT -74.285 -168.805 -73.955 -168.475 ;
        RECT -74.285 -171.525 -73.955 -171.195 ;
        RECT -74.285 -174.245 -73.955 -173.915 ;
        RECT -74.285 -175.605 -73.955 -175.275 ;
        RECT -74.285 -176.685 -73.955 -176.355 ;
        RECT -74.285 -178.325 -73.955 -177.995 ;
        RECT -74.285 -179.685 -73.955 -179.355 ;
        RECT -74.285 -181.93 -73.955 -180.8 ;
        RECT -74.28 -182.045 -73.96 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.925 241.32 -72.595 242.45 ;
        RECT -72.925 239.195 -72.595 239.525 ;
        RECT -72.925 237.835 -72.595 238.165 ;
        RECT -72.925 236.475 -72.595 236.805 ;
        RECT -72.925 235.115 -72.595 235.445 ;
        RECT -72.925 233.755 -72.595 234.085 ;
        RECT -72.925 232.395 -72.595 232.725 ;
        RECT -72.925 231.035 -72.595 231.365 ;
        RECT -72.925 229.675 -72.595 230.005 ;
        RECT -72.925 228.315 -72.595 228.645 ;
        RECT -72.925 226.955 -72.595 227.285 ;
        RECT -72.925 225.595 -72.595 225.925 ;
        RECT -72.925 224.235 -72.595 224.565 ;
        RECT -72.925 222.875 -72.595 223.205 ;
        RECT -72.925 221.515 -72.595 221.845 ;
        RECT -72.925 220.155 -72.595 220.485 ;
        RECT -72.925 218.795 -72.595 219.125 ;
        RECT -72.925 217.435 -72.595 217.765 ;
        RECT -72.925 216.075 -72.595 216.405 ;
        RECT -72.925 214.715 -72.595 215.045 ;
        RECT -72.925 213.355 -72.595 213.685 ;
        RECT -72.925 211.995 -72.595 212.325 ;
        RECT -72.925 210.635 -72.595 210.965 ;
        RECT -72.925 209.275 -72.595 209.605 ;
        RECT -72.925 207.915 -72.595 208.245 ;
        RECT -72.925 206.555 -72.595 206.885 ;
        RECT -72.925 205.195 -72.595 205.525 ;
        RECT -72.925 203.835 -72.595 204.165 ;
        RECT -72.925 202.475 -72.595 202.805 ;
        RECT -72.925 201.115 -72.595 201.445 ;
        RECT -72.925 199.755 -72.595 200.085 ;
        RECT -72.925 198.395 -72.595 198.725 ;
        RECT -72.925 197.035 -72.595 197.365 ;
        RECT -72.925 195.675 -72.595 196.005 ;
        RECT -72.925 194.315 -72.595 194.645 ;
        RECT -72.925 192.955 -72.595 193.285 ;
        RECT -72.925 191.595 -72.595 191.925 ;
        RECT -72.925 190.235 -72.595 190.565 ;
        RECT -72.925 188.875 -72.595 189.205 ;
        RECT -72.925 187.515 -72.595 187.845 ;
        RECT -72.925 186.155 -72.595 186.485 ;
        RECT -72.925 184.795 -72.595 185.125 ;
        RECT -72.925 183.435 -72.595 183.765 ;
        RECT -72.925 182.075 -72.595 182.405 ;
        RECT -72.925 180.715 -72.595 181.045 ;
        RECT -72.925 179.355 -72.595 179.685 ;
        RECT -72.925 177.995 -72.595 178.325 ;
        RECT -72.925 176.635 -72.595 176.965 ;
        RECT -72.925 175.275 -72.595 175.605 ;
        RECT -72.925 173.915 -72.595 174.245 ;
        RECT -72.925 172.555 -72.595 172.885 ;
        RECT -72.925 171.195 -72.595 171.525 ;
        RECT -72.925 169.835 -72.595 170.165 ;
        RECT -72.925 168.475 -72.595 168.805 ;
        RECT -72.925 167.115 -72.595 167.445 ;
        RECT -72.925 165.755 -72.595 166.085 ;
        RECT -72.925 164.395 -72.595 164.725 ;
        RECT -72.925 163.035 -72.595 163.365 ;
        RECT -72.925 161.675 -72.595 162.005 ;
        RECT -72.925 160.315 -72.595 160.645 ;
        RECT -72.925 158.955 -72.595 159.285 ;
        RECT -72.925 157.595 -72.595 157.925 ;
        RECT -72.925 156.235 -72.595 156.565 ;
        RECT -72.925 154.875 -72.595 155.205 ;
        RECT -72.925 153.515 -72.595 153.845 ;
        RECT -72.925 152.155 -72.595 152.485 ;
        RECT -72.925 150.795 -72.595 151.125 ;
        RECT -72.925 149.435 -72.595 149.765 ;
        RECT -72.925 148.075 -72.595 148.405 ;
        RECT -72.925 146.715 -72.595 147.045 ;
        RECT -72.925 145.355 -72.595 145.685 ;
        RECT -72.925 143.995 -72.595 144.325 ;
        RECT -72.925 142.635 -72.595 142.965 ;
        RECT -72.925 141.275 -72.595 141.605 ;
        RECT -72.925 139.915 -72.595 140.245 ;
        RECT -72.925 138.555 -72.595 138.885 ;
        RECT -72.925 137.195 -72.595 137.525 ;
        RECT -72.925 135.835 -72.595 136.165 ;
        RECT -72.925 134.475 -72.595 134.805 ;
        RECT -72.925 133.115 -72.595 133.445 ;
        RECT -72.925 131.755 -72.595 132.085 ;
        RECT -72.925 130.395 -72.595 130.725 ;
        RECT -72.925 129.035 -72.595 129.365 ;
        RECT -72.925 127.675 -72.595 128.005 ;
        RECT -72.925 126.315 -72.595 126.645 ;
        RECT -72.925 124.955 -72.595 125.285 ;
        RECT -72.925 123.595 -72.595 123.925 ;
        RECT -72.925 122.235 -72.595 122.565 ;
        RECT -72.925 120.875 -72.595 121.205 ;
        RECT -72.925 119.515 -72.595 119.845 ;
        RECT -72.925 118.155 -72.595 118.485 ;
        RECT -72.925 116.795 -72.595 117.125 ;
        RECT -72.925 115.435 -72.595 115.765 ;
        RECT -72.925 114.075 -72.595 114.405 ;
        RECT -72.925 112.715 -72.595 113.045 ;
        RECT -72.925 111.355 -72.595 111.685 ;
        RECT -72.925 109.995 -72.595 110.325 ;
        RECT -72.925 108.635 -72.595 108.965 ;
        RECT -72.925 107.275 -72.595 107.605 ;
        RECT -72.925 105.915 -72.595 106.245 ;
        RECT -72.925 104.555 -72.595 104.885 ;
        RECT -72.925 103.195 -72.595 103.525 ;
        RECT -72.925 101.835 -72.595 102.165 ;
        RECT -72.925 100.475 -72.595 100.805 ;
        RECT -72.925 99.115 -72.595 99.445 ;
        RECT -72.925 97.755 -72.595 98.085 ;
        RECT -72.925 96.395 -72.595 96.725 ;
        RECT -72.925 95.035 -72.595 95.365 ;
        RECT -72.925 93.675 -72.595 94.005 ;
        RECT -72.925 92.315 -72.595 92.645 ;
        RECT -72.925 90.955 -72.595 91.285 ;
        RECT -72.925 89.595 -72.595 89.925 ;
        RECT -72.925 88.235 -72.595 88.565 ;
        RECT -72.925 86.875 -72.595 87.205 ;
        RECT -72.925 85.515 -72.595 85.845 ;
        RECT -72.925 84.155 -72.595 84.485 ;
        RECT -72.925 82.795 -72.595 83.125 ;
        RECT -72.925 81.435 -72.595 81.765 ;
        RECT -72.925 80.075 -72.595 80.405 ;
        RECT -72.925 78.715 -72.595 79.045 ;
        RECT -72.925 77.355 -72.595 77.685 ;
        RECT -72.925 75.995 -72.595 76.325 ;
        RECT -72.925 74.635 -72.595 74.965 ;
        RECT -72.925 73.275 -72.595 73.605 ;
        RECT -72.925 71.915 -72.595 72.245 ;
        RECT -72.925 70.555 -72.595 70.885 ;
        RECT -72.925 69.195 -72.595 69.525 ;
        RECT -72.925 67.835 -72.595 68.165 ;
        RECT -72.925 66.475 -72.595 66.805 ;
        RECT -72.925 65.115 -72.595 65.445 ;
        RECT -72.925 63.755 -72.595 64.085 ;
        RECT -72.925 62.395 -72.595 62.725 ;
        RECT -72.925 61.035 -72.595 61.365 ;
        RECT -72.925 59.675 -72.595 60.005 ;
        RECT -72.925 58.315 -72.595 58.645 ;
        RECT -72.925 56.955 -72.595 57.285 ;
        RECT -72.925 55.595 -72.595 55.925 ;
        RECT -72.925 54.235 -72.595 54.565 ;
        RECT -72.925 52.875 -72.595 53.205 ;
        RECT -72.925 51.515 -72.595 51.845 ;
        RECT -72.925 50.155 -72.595 50.485 ;
        RECT -72.925 48.795 -72.595 49.125 ;
        RECT -72.925 47.435 -72.595 47.765 ;
        RECT -72.925 46.075 -72.595 46.405 ;
        RECT -72.925 44.715 -72.595 45.045 ;
        RECT -72.925 43.355 -72.595 43.685 ;
        RECT -72.925 41.995 -72.595 42.325 ;
        RECT -72.925 40.635 -72.595 40.965 ;
        RECT -72.925 39.275 -72.595 39.605 ;
        RECT -72.925 37.915 -72.595 38.245 ;
        RECT -72.925 36.555 -72.595 36.885 ;
        RECT -72.925 35.195 -72.595 35.525 ;
        RECT -72.925 33.835 -72.595 34.165 ;
        RECT -72.925 32.475 -72.595 32.805 ;
        RECT -72.925 31.115 -72.595 31.445 ;
        RECT -72.925 29.755 -72.595 30.085 ;
        RECT -72.925 28.395 -72.595 28.725 ;
        RECT -72.925 27.035 -72.595 27.365 ;
        RECT -72.925 25.675 -72.595 26.005 ;
        RECT -72.925 24.315 -72.595 24.645 ;
        RECT -72.925 22.955 -72.595 23.285 ;
        RECT -72.925 21.595 -72.595 21.925 ;
        RECT -72.925 20.235 -72.595 20.565 ;
        RECT -72.925 18.875 -72.595 19.205 ;
        RECT -72.925 17.515 -72.595 17.845 ;
        RECT -72.925 16.155 -72.595 16.485 ;
        RECT -72.925 14.795 -72.595 15.125 ;
        RECT -72.925 13.435 -72.595 13.765 ;
        RECT -72.925 12.075 -72.595 12.405 ;
        RECT -72.925 10.715 -72.595 11.045 ;
        RECT -72.925 9.355 -72.595 9.685 ;
        RECT -72.925 7.995 -72.595 8.325 ;
        RECT -72.925 6.635 -72.595 6.965 ;
        RECT -72.925 5.275 -72.595 5.605 ;
        RECT -72.925 3.915 -72.595 4.245 ;
        RECT -72.925 2.555 -72.595 2.885 ;
        RECT -72.925 1.195 -72.595 1.525 ;
        RECT -72.925 -0.165 -72.595 0.165 ;
        RECT -72.925 -1.525 -72.595 -1.195 ;
        RECT -72.925 -2.885 -72.595 -2.555 ;
        RECT -72.925 -4.245 -72.595 -3.915 ;
        RECT -72.925 -5.605 -72.595 -5.275 ;
        RECT -72.925 -6.965 -72.595 -6.635 ;
        RECT -72.925 -8.325 -72.595 -7.995 ;
        RECT -72.925 -9.685 -72.595 -9.355 ;
        RECT -72.925 -11.045 -72.595 -10.715 ;
        RECT -72.925 -12.405 -72.595 -12.075 ;
        RECT -72.925 -13.765 -72.595 -13.435 ;
        RECT -72.925 -15.125 -72.595 -14.795 ;
        RECT -72.925 -16.485 -72.595 -16.155 ;
        RECT -72.925 -17.845 -72.595 -17.515 ;
        RECT -72.925 -19.205 -72.595 -18.875 ;
        RECT -72.925 -20.565 -72.595 -20.235 ;
        RECT -72.925 -21.925 -72.595 -21.595 ;
        RECT -72.925 -23.285 -72.595 -22.955 ;
        RECT -72.925 -24.645 -72.595 -24.315 ;
        RECT -72.925 -26.005 -72.595 -25.675 ;
        RECT -72.925 -27.365 -72.595 -27.035 ;
        RECT -72.925 -28.725 -72.595 -28.395 ;
        RECT -72.925 -30.085 -72.595 -29.755 ;
        RECT -72.925 -31.445 -72.595 -31.115 ;
        RECT -72.925 -32.805 -72.595 -32.475 ;
        RECT -72.925 -34.165 -72.595 -33.835 ;
        RECT -72.925 -35.525 -72.595 -35.195 ;
        RECT -72.925 -36.885 -72.595 -36.555 ;
        RECT -72.925 -38.245 -72.595 -37.915 ;
        RECT -72.925 -39.605 -72.595 -39.275 ;
        RECT -72.925 -40.965 -72.595 -40.635 ;
        RECT -72.925 -42.325 -72.595 -41.995 ;
        RECT -72.925 -43.685 -72.595 -43.355 ;
        RECT -72.925 -45.045 -72.595 -44.715 ;
        RECT -72.925 -46.405 -72.595 -46.075 ;
        RECT -72.925 -47.765 -72.595 -47.435 ;
        RECT -72.925 -49.125 -72.595 -48.795 ;
        RECT -72.925 -50.485 -72.595 -50.155 ;
        RECT -72.925 -51.845 -72.595 -51.515 ;
        RECT -72.925 -53.205 -72.595 -52.875 ;
        RECT -72.925 -54.565 -72.595 -54.235 ;
        RECT -72.925 -55.925 -72.595 -55.595 ;
        RECT -72.925 -57.285 -72.595 -56.955 ;
        RECT -72.925 -58.645 -72.595 -58.315 ;
        RECT -72.925 -60.005 -72.595 -59.675 ;
        RECT -72.925 -61.365 -72.595 -61.035 ;
        RECT -72.925 -62.725 -72.595 -62.395 ;
        RECT -72.925 -64.085 -72.595 -63.755 ;
        RECT -72.925 -65.445 -72.595 -65.115 ;
        RECT -72.925 -66.805 -72.595 -66.475 ;
        RECT -72.925 -68.165 -72.595 -67.835 ;
        RECT -72.925 -69.525 -72.595 -69.195 ;
        RECT -72.925 -70.885 -72.595 -70.555 ;
        RECT -72.925 -72.245 -72.595 -71.915 ;
        RECT -72.925 -73.605 -72.595 -73.275 ;
        RECT -72.925 -74.965 -72.595 -74.635 ;
        RECT -72.925 -76.325 -72.595 -75.995 ;
        RECT -72.925 -77.685 -72.595 -77.355 ;
        RECT -72.925 -79.045 -72.595 -78.715 ;
        RECT -72.925 -80.405 -72.595 -80.075 ;
        RECT -72.925 -81.765 -72.595 -81.435 ;
        RECT -72.925 -83.125 -72.595 -82.795 ;
        RECT -72.925 -84.485 -72.595 -84.155 ;
        RECT -72.925 -85.845 -72.595 -85.515 ;
        RECT -72.925 -87.205 -72.595 -86.875 ;
        RECT -72.925 -88.565 -72.595 -88.235 ;
        RECT -72.925 -89.925 -72.595 -89.595 ;
        RECT -72.925 -91.285 -72.595 -90.955 ;
        RECT -72.925 -92.645 -72.595 -92.315 ;
        RECT -72.925 -94.005 -72.595 -93.675 ;
        RECT -72.925 -95.365 -72.595 -95.035 ;
        RECT -72.925 -96.725 -72.595 -96.395 ;
        RECT -72.925 -98.085 -72.595 -97.755 ;
        RECT -72.925 -99.445 -72.595 -99.115 ;
        RECT -72.925 -100.805 -72.595 -100.475 ;
        RECT -72.925 -102.165 -72.595 -101.835 ;
        RECT -72.925 -103.525 -72.595 -103.195 ;
        RECT -72.925 -104.885 -72.595 -104.555 ;
        RECT -72.925 -106.245 -72.595 -105.915 ;
        RECT -72.925 -107.605 -72.595 -107.275 ;
        RECT -72.925 -108.965 -72.595 -108.635 ;
        RECT -72.925 -110.325 -72.595 -109.995 ;
        RECT -72.925 -111.685 -72.595 -111.355 ;
        RECT -72.925 -113.045 -72.595 -112.715 ;
        RECT -72.92 -113.045 -72.6 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -72.925 -175.605 -72.595 -175.275 ;
        RECT -72.925 -176.685 -72.595 -176.355 ;
        RECT -72.925 -178.325 -72.595 -177.995 ;
        RECT -72.925 -179.685 -72.595 -179.355 ;
        RECT -72.925 -181.93 -72.595 -180.8 ;
        RECT -72.92 -182.045 -72.6 -173.24 ;
    END
    PORT
      LAYER met3 ;
        RECT -71.565 194.315 -71.235 194.645 ;
        RECT -71.565 192.955 -71.235 193.285 ;
        RECT -71.565 191.595 -71.235 191.925 ;
        RECT -71.565 190.235 -71.235 190.565 ;
        RECT -71.565 188.875 -71.235 189.205 ;
        RECT -71.565 187.515 -71.235 187.845 ;
        RECT -71.565 186.155 -71.235 186.485 ;
        RECT -71.565 184.795 -71.235 185.125 ;
        RECT -71.565 183.435 -71.235 183.765 ;
        RECT -71.565 182.075 -71.235 182.405 ;
        RECT -71.565 180.715 -71.235 181.045 ;
        RECT -71.565 179.355 -71.235 179.685 ;
        RECT -71.565 177.995 -71.235 178.325 ;
        RECT -71.565 176.635 -71.235 176.965 ;
        RECT -71.565 175.275 -71.235 175.605 ;
        RECT -71.565 173.915 -71.235 174.245 ;
        RECT -71.565 172.555 -71.235 172.885 ;
        RECT -71.565 171.195 -71.235 171.525 ;
        RECT -71.565 169.835 -71.235 170.165 ;
        RECT -71.565 168.475 -71.235 168.805 ;
        RECT -71.565 167.115 -71.235 167.445 ;
        RECT -71.565 165.755 -71.235 166.085 ;
        RECT -71.565 164.395 -71.235 164.725 ;
        RECT -71.565 163.035 -71.235 163.365 ;
        RECT -71.565 161.675 -71.235 162.005 ;
        RECT -71.565 160.315 -71.235 160.645 ;
        RECT -71.565 158.955 -71.235 159.285 ;
        RECT -71.565 157.595 -71.235 157.925 ;
        RECT -71.565 156.235 -71.235 156.565 ;
        RECT -71.565 154.875 -71.235 155.205 ;
        RECT -71.565 153.515 -71.235 153.845 ;
        RECT -71.565 152.155 -71.235 152.485 ;
        RECT -71.565 150.795 -71.235 151.125 ;
        RECT -71.565 149.435 -71.235 149.765 ;
        RECT -71.565 148.075 -71.235 148.405 ;
        RECT -71.565 146.715 -71.235 147.045 ;
        RECT -71.565 145.355 -71.235 145.685 ;
        RECT -71.565 143.995 -71.235 144.325 ;
        RECT -71.565 142.635 -71.235 142.965 ;
        RECT -71.565 141.275 -71.235 141.605 ;
        RECT -71.565 139.915 -71.235 140.245 ;
        RECT -71.565 138.555 -71.235 138.885 ;
        RECT -71.565 137.195 -71.235 137.525 ;
        RECT -71.565 135.835 -71.235 136.165 ;
        RECT -71.565 134.475 -71.235 134.805 ;
        RECT -71.565 133.115 -71.235 133.445 ;
        RECT -71.565 131.755 -71.235 132.085 ;
        RECT -71.565 130.395 -71.235 130.725 ;
        RECT -71.565 129.035 -71.235 129.365 ;
        RECT -71.565 127.675 -71.235 128.005 ;
        RECT -71.565 126.315 -71.235 126.645 ;
        RECT -71.565 124.955 -71.235 125.285 ;
        RECT -71.565 123.595 -71.235 123.925 ;
        RECT -71.565 122.235 -71.235 122.565 ;
        RECT -71.565 120.875 -71.235 121.205 ;
        RECT -71.565 119.515 -71.235 119.845 ;
        RECT -71.565 118.155 -71.235 118.485 ;
        RECT -71.565 116.795 -71.235 117.125 ;
        RECT -71.565 115.435 -71.235 115.765 ;
        RECT -71.565 114.075 -71.235 114.405 ;
        RECT -71.565 112.715 -71.235 113.045 ;
        RECT -71.565 111.355 -71.235 111.685 ;
        RECT -71.565 109.995 -71.235 110.325 ;
        RECT -71.565 108.635 -71.235 108.965 ;
        RECT -71.565 107.275 -71.235 107.605 ;
        RECT -71.565 105.915 -71.235 106.245 ;
        RECT -71.565 104.555 -71.235 104.885 ;
        RECT -71.565 103.195 -71.235 103.525 ;
        RECT -71.565 101.835 -71.235 102.165 ;
        RECT -71.565 100.475 -71.235 100.805 ;
        RECT -71.565 99.115 -71.235 99.445 ;
        RECT -71.565 97.755 -71.235 98.085 ;
        RECT -71.565 96.395 -71.235 96.725 ;
        RECT -71.565 95.035 -71.235 95.365 ;
        RECT -71.565 93.675 -71.235 94.005 ;
        RECT -71.565 92.315 -71.235 92.645 ;
        RECT -71.565 90.955 -71.235 91.285 ;
        RECT -71.565 89.595 -71.235 89.925 ;
        RECT -71.565 88.235 -71.235 88.565 ;
        RECT -71.565 86.875 -71.235 87.205 ;
        RECT -71.565 85.515 -71.235 85.845 ;
        RECT -71.565 84.155 -71.235 84.485 ;
        RECT -71.565 82.795 -71.235 83.125 ;
        RECT -71.565 81.435 -71.235 81.765 ;
        RECT -71.565 80.075 -71.235 80.405 ;
        RECT -71.565 78.715 -71.235 79.045 ;
        RECT -71.565 77.355 -71.235 77.685 ;
        RECT -71.565 75.995 -71.235 76.325 ;
        RECT -71.565 74.635 -71.235 74.965 ;
        RECT -71.565 73.275 -71.235 73.605 ;
        RECT -71.565 71.915 -71.235 72.245 ;
        RECT -71.565 70.555 -71.235 70.885 ;
        RECT -71.565 69.195 -71.235 69.525 ;
        RECT -71.565 67.835 -71.235 68.165 ;
        RECT -71.565 66.475 -71.235 66.805 ;
        RECT -71.565 65.115 -71.235 65.445 ;
        RECT -71.565 63.755 -71.235 64.085 ;
        RECT -71.565 62.395 -71.235 62.725 ;
        RECT -71.565 61.035 -71.235 61.365 ;
        RECT -71.565 59.675 -71.235 60.005 ;
        RECT -71.565 58.315 -71.235 58.645 ;
        RECT -71.565 56.955 -71.235 57.285 ;
        RECT -71.565 55.595 -71.235 55.925 ;
        RECT -71.565 54.235 -71.235 54.565 ;
        RECT -71.565 52.875 -71.235 53.205 ;
        RECT -71.565 51.515 -71.235 51.845 ;
        RECT -71.565 50.155 -71.235 50.485 ;
        RECT -71.565 48.795 -71.235 49.125 ;
        RECT -71.565 47.435 -71.235 47.765 ;
        RECT -71.565 46.075 -71.235 46.405 ;
        RECT -71.565 44.715 -71.235 45.045 ;
        RECT -71.565 43.355 -71.235 43.685 ;
        RECT -71.565 41.995 -71.235 42.325 ;
        RECT -71.565 40.635 -71.235 40.965 ;
        RECT -71.565 39.275 -71.235 39.605 ;
        RECT -71.565 37.915 -71.235 38.245 ;
        RECT -71.565 36.555 -71.235 36.885 ;
        RECT -71.565 35.195 -71.235 35.525 ;
        RECT -71.565 33.835 -71.235 34.165 ;
        RECT -71.565 32.475 -71.235 32.805 ;
        RECT -71.565 31.115 -71.235 31.445 ;
        RECT -71.565 29.755 -71.235 30.085 ;
        RECT -71.565 28.395 -71.235 28.725 ;
        RECT -71.565 27.035 -71.235 27.365 ;
        RECT -71.565 25.675 -71.235 26.005 ;
        RECT -71.565 24.315 -71.235 24.645 ;
        RECT -71.565 22.955 -71.235 23.285 ;
        RECT -71.565 21.595 -71.235 21.925 ;
        RECT -71.565 20.235 -71.235 20.565 ;
        RECT -71.565 18.875 -71.235 19.205 ;
        RECT -71.565 17.515 -71.235 17.845 ;
        RECT -71.565 16.155 -71.235 16.485 ;
        RECT -71.565 14.795 -71.235 15.125 ;
        RECT -71.565 13.435 -71.235 13.765 ;
        RECT -71.565 12.075 -71.235 12.405 ;
        RECT -71.565 10.715 -71.235 11.045 ;
        RECT -71.565 9.355 -71.235 9.685 ;
        RECT -71.565 7.995 -71.235 8.325 ;
        RECT -71.565 6.635 -71.235 6.965 ;
        RECT -71.565 5.275 -71.235 5.605 ;
        RECT -71.565 3.915 -71.235 4.245 ;
        RECT -71.565 2.555 -71.235 2.885 ;
        RECT -71.565 1.195 -71.235 1.525 ;
        RECT -71.565 -0.165 -71.235 0.165 ;
        RECT -71.565 -1.525 -71.235 -1.195 ;
        RECT -71.565 -2.885 -71.235 -2.555 ;
        RECT -71.565 -4.245 -71.235 -3.915 ;
        RECT -71.565 -5.605 -71.235 -5.275 ;
        RECT -71.565 -6.965 -71.235 -6.635 ;
        RECT -71.565 -8.325 -71.235 -7.995 ;
        RECT -71.565 -9.685 -71.235 -9.355 ;
        RECT -71.565 -11.045 -71.235 -10.715 ;
        RECT -71.565 -12.405 -71.235 -12.075 ;
        RECT -71.565 -13.765 -71.235 -13.435 ;
        RECT -71.565 -15.125 -71.235 -14.795 ;
        RECT -71.565 -16.485 -71.235 -16.155 ;
        RECT -71.565 -17.845 -71.235 -17.515 ;
        RECT -71.565 -19.205 -71.235 -18.875 ;
        RECT -71.565 -20.565 -71.235 -20.235 ;
        RECT -71.565 -21.925 -71.235 -21.595 ;
        RECT -71.565 -23.285 -71.235 -22.955 ;
        RECT -71.565 -24.645 -71.235 -24.315 ;
        RECT -71.565 -26.005 -71.235 -25.675 ;
        RECT -71.565 -27.365 -71.235 -27.035 ;
        RECT -71.565 -28.725 -71.235 -28.395 ;
        RECT -71.565 -30.085 -71.235 -29.755 ;
        RECT -71.565 -31.445 -71.235 -31.115 ;
        RECT -71.565 -32.805 -71.235 -32.475 ;
        RECT -71.565 -34.165 -71.235 -33.835 ;
        RECT -71.565 -35.525 -71.235 -35.195 ;
        RECT -71.565 -36.885 -71.235 -36.555 ;
        RECT -71.565 -38.245 -71.235 -37.915 ;
        RECT -71.565 -39.605 -71.235 -39.275 ;
        RECT -71.565 -40.965 -71.235 -40.635 ;
        RECT -71.565 -42.325 -71.235 -41.995 ;
        RECT -71.565 -43.685 -71.235 -43.355 ;
        RECT -71.565 -45.045 -71.235 -44.715 ;
        RECT -71.565 -46.405 -71.235 -46.075 ;
        RECT -71.565 -47.765 -71.235 -47.435 ;
        RECT -71.565 -49.125 -71.235 -48.795 ;
        RECT -71.565 -50.485 -71.235 -50.155 ;
        RECT -71.565 -51.845 -71.235 -51.515 ;
        RECT -71.565 -53.205 -71.235 -52.875 ;
        RECT -71.565 -54.565 -71.235 -54.235 ;
        RECT -71.565 -55.925 -71.235 -55.595 ;
        RECT -71.565 -57.285 -71.235 -56.955 ;
        RECT -71.565 -58.645 -71.235 -58.315 ;
        RECT -71.565 -60.005 -71.235 -59.675 ;
        RECT -71.565 -61.365 -71.235 -61.035 ;
        RECT -71.565 -62.725 -71.235 -62.395 ;
        RECT -71.565 -64.085 -71.235 -63.755 ;
        RECT -71.565 -65.445 -71.235 -65.115 ;
        RECT -71.565 -66.805 -71.235 -66.475 ;
        RECT -71.565 -68.165 -71.235 -67.835 ;
        RECT -71.565 -69.525 -71.235 -69.195 ;
        RECT -71.565 -70.885 -71.235 -70.555 ;
        RECT -71.565 -72.245 -71.235 -71.915 ;
        RECT -71.565 -73.605 -71.235 -73.275 ;
        RECT -71.565 -74.965 -71.235 -74.635 ;
        RECT -71.565 -76.325 -71.235 -75.995 ;
        RECT -71.565 -77.685 -71.235 -77.355 ;
        RECT -71.565 -79.045 -71.235 -78.715 ;
        RECT -71.565 -80.405 -71.235 -80.075 ;
        RECT -71.565 -81.765 -71.235 -81.435 ;
        RECT -71.565 -83.125 -71.235 -82.795 ;
        RECT -71.565 -84.485 -71.235 -84.155 ;
        RECT -71.565 -85.845 -71.235 -85.515 ;
        RECT -71.565 -87.205 -71.235 -86.875 ;
        RECT -71.565 -88.565 -71.235 -88.235 ;
        RECT -71.565 -89.925 -71.235 -89.595 ;
        RECT -71.565 -91.285 -71.235 -90.955 ;
        RECT -71.565 -92.645 -71.235 -92.315 ;
        RECT -71.565 -94.005 -71.235 -93.675 ;
        RECT -71.565 -95.365 -71.235 -95.035 ;
        RECT -71.565 -96.725 -71.235 -96.395 ;
        RECT -71.565 -98.085 -71.235 -97.755 ;
        RECT -71.565 -99.445 -71.235 -99.115 ;
        RECT -71.565 -100.805 -71.235 -100.475 ;
        RECT -71.565 -102.165 -71.235 -101.835 ;
        RECT -71.565 -103.525 -71.235 -103.195 ;
        RECT -71.565 -104.885 -71.235 -104.555 ;
        RECT -71.565 -106.245 -71.235 -105.915 ;
        RECT -71.565 -107.605 -71.235 -107.275 ;
        RECT -71.565 -108.965 -71.235 -108.635 ;
        RECT -71.565 -110.325 -71.235 -109.995 ;
        RECT -71.565 -111.685 -71.235 -111.355 ;
        RECT -71.56 -112.36 -71.24 242.565 ;
        RECT -71.565 241.32 -71.235 242.45 ;
        RECT -71.565 239.195 -71.235 239.525 ;
        RECT -71.565 237.835 -71.235 238.165 ;
        RECT -71.565 236.475 -71.235 236.805 ;
        RECT -71.565 235.115 -71.235 235.445 ;
        RECT -71.565 233.755 -71.235 234.085 ;
        RECT -71.565 232.395 -71.235 232.725 ;
        RECT -71.565 231.035 -71.235 231.365 ;
        RECT -71.565 229.675 -71.235 230.005 ;
        RECT -71.565 228.315 -71.235 228.645 ;
        RECT -71.565 226.955 -71.235 227.285 ;
        RECT -71.565 225.595 -71.235 225.925 ;
        RECT -71.565 224.235 -71.235 224.565 ;
        RECT -71.565 222.875 -71.235 223.205 ;
        RECT -71.565 221.515 -71.235 221.845 ;
        RECT -71.565 220.155 -71.235 220.485 ;
        RECT -71.565 218.795 -71.235 219.125 ;
        RECT -71.565 217.435 -71.235 217.765 ;
        RECT -71.565 216.075 -71.235 216.405 ;
        RECT -71.565 214.715 -71.235 215.045 ;
        RECT -71.565 213.355 -71.235 213.685 ;
        RECT -71.565 211.995 -71.235 212.325 ;
        RECT -71.565 210.635 -71.235 210.965 ;
        RECT -71.565 209.275 -71.235 209.605 ;
        RECT -71.565 207.915 -71.235 208.245 ;
        RECT -71.565 206.555 -71.235 206.885 ;
        RECT -71.565 205.195 -71.235 205.525 ;
        RECT -71.565 203.835 -71.235 204.165 ;
        RECT -71.565 202.475 -71.235 202.805 ;
        RECT -71.565 201.115 -71.235 201.445 ;
        RECT -71.565 199.755 -71.235 200.085 ;
        RECT -71.565 198.395 -71.235 198.725 ;
        RECT -71.565 197.035 -71.235 197.365 ;
        RECT -71.565 195.675 -71.235 196.005 ;
    END
    PORT
      LAYER met3 ;
        RECT -78.365 241.32 -78.035 242.45 ;
        RECT -78.365 239.195 -78.035 239.525 ;
        RECT -78.365 237.835 -78.035 238.165 ;
        RECT -78.365 236.475 -78.035 236.805 ;
        RECT -78.365 235.115 -78.035 235.445 ;
        RECT -78.365 233.755 -78.035 234.085 ;
        RECT -78.365 232.395 -78.035 232.725 ;
        RECT -78.365 231.035 -78.035 231.365 ;
        RECT -78.365 229.675 -78.035 230.005 ;
        RECT -78.365 228.315 -78.035 228.645 ;
        RECT -78.365 226.955 -78.035 227.285 ;
        RECT -78.365 225.595 -78.035 225.925 ;
        RECT -78.365 224.235 -78.035 224.565 ;
        RECT -78.365 222.875 -78.035 223.205 ;
        RECT -78.365 221.515 -78.035 221.845 ;
        RECT -78.365 220.155 -78.035 220.485 ;
        RECT -78.365 218.795 -78.035 219.125 ;
        RECT -78.365 217.435 -78.035 217.765 ;
        RECT -78.365 216.075 -78.035 216.405 ;
        RECT -78.365 214.715 -78.035 215.045 ;
        RECT -78.365 213.355 -78.035 213.685 ;
        RECT -78.365 211.995 -78.035 212.325 ;
        RECT -78.365 210.635 -78.035 210.965 ;
        RECT -78.365 209.275 -78.035 209.605 ;
        RECT -78.365 207.915 -78.035 208.245 ;
        RECT -78.365 206.555 -78.035 206.885 ;
        RECT -78.365 205.195 -78.035 205.525 ;
        RECT -78.365 203.835 -78.035 204.165 ;
        RECT -78.365 202.475 -78.035 202.805 ;
        RECT -78.365 201.115 -78.035 201.445 ;
        RECT -78.365 199.755 -78.035 200.085 ;
        RECT -78.365 198.395 -78.035 198.725 ;
        RECT -78.365 197.035 -78.035 197.365 ;
        RECT -78.365 195.675 -78.035 196.005 ;
        RECT -78.365 194.315 -78.035 194.645 ;
        RECT -78.365 192.955 -78.035 193.285 ;
        RECT -78.365 191.595 -78.035 191.925 ;
        RECT -78.365 190.235 -78.035 190.565 ;
        RECT -78.365 188.875 -78.035 189.205 ;
        RECT -78.365 187.515 -78.035 187.845 ;
        RECT -78.365 186.155 -78.035 186.485 ;
        RECT -78.365 184.795 -78.035 185.125 ;
        RECT -78.365 183.435 -78.035 183.765 ;
        RECT -78.365 182.075 -78.035 182.405 ;
        RECT -78.365 180.715 -78.035 181.045 ;
        RECT -78.365 179.355 -78.035 179.685 ;
        RECT -78.365 177.995 -78.035 178.325 ;
        RECT -78.365 176.635 -78.035 176.965 ;
        RECT -78.365 175.275 -78.035 175.605 ;
        RECT -78.365 173.915 -78.035 174.245 ;
        RECT -78.365 172.555 -78.035 172.885 ;
        RECT -78.365 171.195 -78.035 171.525 ;
        RECT -78.365 169.835 -78.035 170.165 ;
        RECT -78.365 168.475 -78.035 168.805 ;
        RECT -78.365 167.115 -78.035 167.445 ;
        RECT -78.365 165.755 -78.035 166.085 ;
        RECT -78.365 164.395 -78.035 164.725 ;
        RECT -78.365 163.035 -78.035 163.365 ;
        RECT -78.365 161.675 -78.035 162.005 ;
        RECT -78.365 160.315 -78.035 160.645 ;
        RECT -78.365 158.955 -78.035 159.285 ;
        RECT -78.365 157.595 -78.035 157.925 ;
        RECT -78.365 156.235 -78.035 156.565 ;
        RECT -78.365 154.875 -78.035 155.205 ;
        RECT -78.365 153.515 -78.035 153.845 ;
        RECT -78.365 152.155 -78.035 152.485 ;
        RECT -78.365 150.795 -78.035 151.125 ;
        RECT -78.365 149.435 -78.035 149.765 ;
        RECT -78.365 148.075 -78.035 148.405 ;
        RECT -78.365 146.715 -78.035 147.045 ;
        RECT -78.365 145.355 -78.035 145.685 ;
        RECT -78.365 143.995 -78.035 144.325 ;
        RECT -78.365 142.635 -78.035 142.965 ;
        RECT -78.365 141.275 -78.035 141.605 ;
        RECT -78.365 139.915 -78.035 140.245 ;
        RECT -78.365 138.555 -78.035 138.885 ;
        RECT -78.365 137.195 -78.035 137.525 ;
        RECT -78.365 135.835 -78.035 136.165 ;
        RECT -78.365 134.475 -78.035 134.805 ;
        RECT -78.365 133.115 -78.035 133.445 ;
        RECT -78.365 131.755 -78.035 132.085 ;
        RECT -78.365 130.395 -78.035 130.725 ;
        RECT -78.365 129.035 -78.035 129.365 ;
        RECT -78.365 127.675 -78.035 128.005 ;
        RECT -78.365 126.315 -78.035 126.645 ;
        RECT -78.365 124.955 -78.035 125.285 ;
        RECT -78.365 123.595 -78.035 123.925 ;
        RECT -78.365 122.235 -78.035 122.565 ;
        RECT -78.365 120.875 -78.035 121.205 ;
        RECT -78.365 119.515 -78.035 119.845 ;
        RECT -78.365 118.155 -78.035 118.485 ;
        RECT -78.365 116.795 -78.035 117.125 ;
        RECT -78.365 115.435 -78.035 115.765 ;
        RECT -78.365 114.075 -78.035 114.405 ;
        RECT -78.365 112.715 -78.035 113.045 ;
        RECT -78.365 111.355 -78.035 111.685 ;
        RECT -78.365 109.995 -78.035 110.325 ;
        RECT -78.365 108.635 -78.035 108.965 ;
        RECT -78.365 107.275 -78.035 107.605 ;
        RECT -78.365 105.915 -78.035 106.245 ;
        RECT -78.365 104.555 -78.035 104.885 ;
        RECT -78.365 103.195 -78.035 103.525 ;
        RECT -78.365 101.835 -78.035 102.165 ;
        RECT -78.365 100.475 -78.035 100.805 ;
        RECT -78.365 99.115 -78.035 99.445 ;
        RECT -78.365 97.755 -78.035 98.085 ;
        RECT -78.365 96.395 -78.035 96.725 ;
        RECT -78.365 95.035 -78.035 95.365 ;
        RECT -78.365 93.675 -78.035 94.005 ;
        RECT -78.365 92.315 -78.035 92.645 ;
        RECT -78.365 90.955 -78.035 91.285 ;
        RECT -78.365 89.595 -78.035 89.925 ;
        RECT -78.365 88.235 -78.035 88.565 ;
        RECT -78.365 86.875 -78.035 87.205 ;
        RECT -78.365 85.515 -78.035 85.845 ;
        RECT -78.365 84.155 -78.035 84.485 ;
        RECT -78.365 82.795 -78.035 83.125 ;
        RECT -78.365 81.435 -78.035 81.765 ;
        RECT -78.365 80.075 -78.035 80.405 ;
        RECT -78.365 78.715 -78.035 79.045 ;
        RECT -78.365 77.355 -78.035 77.685 ;
        RECT -78.365 75.995 -78.035 76.325 ;
        RECT -78.365 74.635 -78.035 74.965 ;
        RECT -78.365 73.275 -78.035 73.605 ;
        RECT -78.365 71.915 -78.035 72.245 ;
        RECT -78.365 70.555 -78.035 70.885 ;
        RECT -78.365 69.195 -78.035 69.525 ;
        RECT -78.365 67.835 -78.035 68.165 ;
        RECT -78.365 66.475 -78.035 66.805 ;
        RECT -78.365 65.115 -78.035 65.445 ;
        RECT -78.365 63.755 -78.035 64.085 ;
        RECT -78.365 62.395 -78.035 62.725 ;
        RECT -78.365 61.035 -78.035 61.365 ;
        RECT -78.365 59.675 -78.035 60.005 ;
        RECT -78.365 58.315 -78.035 58.645 ;
        RECT -78.365 56.955 -78.035 57.285 ;
        RECT -78.365 55.595 -78.035 55.925 ;
        RECT -78.365 54.235 -78.035 54.565 ;
        RECT -78.365 52.875 -78.035 53.205 ;
        RECT -78.365 51.515 -78.035 51.845 ;
        RECT -78.365 50.155 -78.035 50.485 ;
        RECT -78.365 48.795 -78.035 49.125 ;
        RECT -78.365 47.435 -78.035 47.765 ;
        RECT -78.365 46.075 -78.035 46.405 ;
        RECT -78.365 44.715 -78.035 45.045 ;
        RECT -78.365 43.355 -78.035 43.685 ;
        RECT -78.365 41.995 -78.035 42.325 ;
        RECT -78.365 40.635 -78.035 40.965 ;
        RECT -78.365 39.275 -78.035 39.605 ;
        RECT -78.365 37.915 -78.035 38.245 ;
        RECT -78.365 36.555 -78.035 36.885 ;
        RECT -78.365 35.195 -78.035 35.525 ;
        RECT -78.365 33.835 -78.035 34.165 ;
        RECT -78.365 32.475 -78.035 32.805 ;
        RECT -78.365 31.115 -78.035 31.445 ;
        RECT -78.365 29.755 -78.035 30.085 ;
        RECT -78.365 28.395 -78.035 28.725 ;
        RECT -78.365 27.035 -78.035 27.365 ;
        RECT -78.365 25.675 -78.035 26.005 ;
        RECT -78.365 24.315 -78.035 24.645 ;
        RECT -78.365 22.955 -78.035 23.285 ;
        RECT -78.365 21.595 -78.035 21.925 ;
        RECT -78.365 20.235 -78.035 20.565 ;
        RECT -78.365 18.875 -78.035 19.205 ;
        RECT -78.365 17.515 -78.035 17.845 ;
        RECT -78.365 16.155 -78.035 16.485 ;
        RECT -78.365 14.795 -78.035 15.125 ;
        RECT -78.365 13.435 -78.035 13.765 ;
        RECT -78.365 12.075 -78.035 12.405 ;
        RECT -78.365 10.715 -78.035 11.045 ;
        RECT -78.365 9.355 -78.035 9.685 ;
        RECT -78.365 7.995 -78.035 8.325 ;
        RECT -78.365 6.635 -78.035 6.965 ;
        RECT -78.365 5.275 -78.035 5.605 ;
        RECT -78.365 3.915 -78.035 4.245 ;
        RECT -78.365 2.555 -78.035 2.885 ;
        RECT -78.365 1.195 -78.035 1.525 ;
        RECT -78.365 -0.165 -78.035 0.165 ;
        RECT -78.365 -1.525 -78.035 -1.195 ;
        RECT -78.365 -2.885 -78.035 -2.555 ;
        RECT -78.365 -4.245 -78.035 -3.915 ;
        RECT -78.365 -5.605 -78.035 -5.275 ;
        RECT -78.365 -6.965 -78.035 -6.635 ;
        RECT -78.365 -8.325 -78.035 -7.995 ;
        RECT -78.365 -9.685 -78.035 -9.355 ;
        RECT -78.365 -11.045 -78.035 -10.715 ;
        RECT -78.365 -12.405 -78.035 -12.075 ;
        RECT -78.365 -13.765 -78.035 -13.435 ;
        RECT -78.365 -15.125 -78.035 -14.795 ;
        RECT -78.365 -16.485 -78.035 -16.155 ;
        RECT -78.365 -17.845 -78.035 -17.515 ;
        RECT -78.365 -19.205 -78.035 -18.875 ;
        RECT -78.365 -20.565 -78.035 -20.235 ;
        RECT -78.365 -21.925 -78.035 -21.595 ;
        RECT -78.365 -23.285 -78.035 -22.955 ;
        RECT -78.365 -24.645 -78.035 -24.315 ;
        RECT -78.365 -26.005 -78.035 -25.675 ;
        RECT -78.365 -27.365 -78.035 -27.035 ;
        RECT -78.365 -28.725 -78.035 -28.395 ;
        RECT -78.365 -30.085 -78.035 -29.755 ;
        RECT -78.365 -31.445 -78.035 -31.115 ;
        RECT -78.365 -32.805 -78.035 -32.475 ;
        RECT -78.365 -34.165 -78.035 -33.835 ;
        RECT -78.365 -35.525 -78.035 -35.195 ;
        RECT -78.365 -36.885 -78.035 -36.555 ;
        RECT -78.365 -38.245 -78.035 -37.915 ;
        RECT -78.365 -39.605 -78.035 -39.275 ;
        RECT -78.365 -40.965 -78.035 -40.635 ;
        RECT -78.365 -42.325 -78.035 -41.995 ;
        RECT -78.365 -43.685 -78.035 -43.355 ;
        RECT -78.365 -45.045 -78.035 -44.715 ;
        RECT -78.365 -46.405 -78.035 -46.075 ;
        RECT -78.365 -47.765 -78.035 -47.435 ;
        RECT -78.365 -49.125 -78.035 -48.795 ;
        RECT -78.365 -50.485 -78.035 -50.155 ;
        RECT -78.365 -51.845 -78.035 -51.515 ;
        RECT -78.365 -53.205 -78.035 -52.875 ;
        RECT -78.365 -54.565 -78.035 -54.235 ;
        RECT -78.365 -55.925 -78.035 -55.595 ;
        RECT -78.365 -57.285 -78.035 -56.955 ;
        RECT -78.365 -58.645 -78.035 -58.315 ;
        RECT -78.365 -60.005 -78.035 -59.675 ;
        RECT -78.365 -61.365 -78.035 -61.035 ;
        RECT -78.365 -62.725 -78.035 -62.395 ;
        RECT -78.365 -64.085 -78.035 -63.755 ;
        RECT -78.365 -65.445 -78.035 -65.115 ;
        RECT -78.365 -66.805 -78.035 -66.475 ;
        RECT -78.365 -68.165 -78.035 -67.835 ;
        RECT -78.365 -69.525 -78.035 -69.195 ;
        RECT -78.365 -70.885 -78.035 -70.555 ;
        RECT -78.365 -72.245 -78.035 -71.915 ;
        RECT -78.365 -73.605 -78.035 -73.275 ;
        RECT -78.365 -74.965 -78.035 -74.635 ;
        RECT -78.365 -76.325 -78.035 -75.995 ;
        RECT -78.365 -77.685 -78.035 -77.355 ;
        RECT -78.365 -79.045 -78.035 -78.715 ;
        RECT -78.365 -80.405 -78.035 -80.075 ;
        RECT -78.365 -81.765 -78.035 -81.435 ;
        RECT -78.365 -83.125 -78.035 -82.795 ;
        RECT -78.365 -84.485 -78.035 -84.155 ;
        RECT -78.365 -85.845 -78.035 -85.515 ;
        RECT -78.365 -87.205 -78.035 -86.875 ;
        RECT -78.365 -88.565 -78.035 -88.235 ;
        RECT -78.365 -89.925 -78.035 -89.595 ;
        RECT -78.365 -91.285 -78.035 -90.955 ;
        RECT -78.365 -92.645 -78.035 -92.315 ;
        RECT -78.365 -94.005 -78.035 -93.675 ;
        RECT -78.365 -95.365 -78.035 -95.035 ;
        RECT -78.365 -96.725 -78.035 -96.395 ;
        RECT -78.365 -98.085 -78.035 -97.755 ;
        RECT -78.365 -99.445 -78.035 -99.115 ;
        RECT -78.365 -100.805 -78.035 -100.475 ;
        RECT -78.365 -102.165 -78.035 -101.835 ;
        RECT -78.365 -103.525 -78.035 -103.195 ;
        RECT -78.365 -104.885 -78.035 -104.555 ;
        RECT -78.365 -106.245 -78.035 -105.915 ;
        RECT -78.365 -107.605 -78.035 -107.275 ;
        RECT -78.365 -108.965 -78.035 -108.635 ;
        RECT -78.365 -110.325 -78.035 -109.995 ;
        RECT -78.365 -111.685 -78.035 -111.355 ;
        RECT -78.365 -113.045 -78.035 -112.715 ;
        RECT -78.365 -114.405 -78.035 -114.075 ;
        RECT -78.365 -115.765 -78.035 -115.435 ;
        RECT -78.365 -117.125 -78.035 -116.795 ;
        RECT -78.365 -118.485 -78.035 -118.155 ;
        RECT -78.365 -119.845 -78.035 -119.515 ;
        RECT -78.365 -121.205 -78.035 -120.875 ;
        RECT -78.365 -122.565 -78.035 -122.235 ;
        RECT -78.365 -123.925 -78.035 -123.595 ;
        RECT -78.365 -125.285 -78.035 -124.955 ;
        RECT -78.365 -126.645 -78.035 -126.315 ;
        RECT -78.365 -128.005 -78.035 -127.675 ;
        RECT -78.365 -129.365 -78.035 -129.035 ;
        RECT -78.365 -130.725 -78.035 -130.395 ;
        RECT -78.365 -132.085 -78.035 -131.755 ;
        RECT -78.365 -133.445 -78.035 -133.115 ;
        RECT -78.365 -134.805 -78.035 -134.475 ;
        RECT -78.365 -136.165 -78.035 -135.835 ;
        RECT -78.365 -137.525 -78.035 -137.195 ;
        RECT -78.365 -138.885 -78.035 -138.555 ;
        RECT -78.365 -140.245 -78.035 -139.915 ;
        RECT -78.365 -141.605 -78.035 -141.275 ;
        RECT -78.365 -142.965 -78.035 -142.635 ;
        RECT -78.365 -144.325 -78.035 -143.995 ;
        RECT -78.365 -145.685 -78.035 -145.355 ;
        RECT -78.365 -147.045 -78.035 -146.715 ;
        RECT -78.365 -148.405 -78.035 -148.075 ;
        RECT -78.365 -149.765 -78.035 -149.435 ;
        RECT -78.365 -151.125 -78.035 -150.795 ;
        RECT -78.365 -152.485 -78.035 -152.155 ;
        RECT -78.365 -153.845 -78.035 -153.515 ;
        RECT -78.365 -155.205 -78.035 -154.875 ;
        RECT -78.365 -156.565 -78.035 -156.235 ;
        RECT -78.365 -157.925 -78.035 -157.595 ;
        RECT -78.365 -159.285 -78.035 -158.955 ;
        RECT -78.365 -160.645 -78.035 -160.315 ;
        RECT -78.365 -162.005 -78.035 -161.675 ;
        RECT -78.365 -163.365 -78.035 -163.035 ;
        RECT -78.365 -164.725 -78.035 -164.395 ;
        RECT -78.365 -166.085 -78.035 -165.755 ;
        RECT -78.365 -167.445 -78.035 -167.115 ;
        RECT -78.365 -168.805 -78.035 -168.475 ;
        RECT -78.365 -171.525 -78.035 -171.195 ;
        RECT -78.365 -172.885 -78.035 -172.555 ;
        RECT -78.365 -174.245 -78.035 -173.915 ;
        RECT -78.365 -175.605 -78.035 -175.275 ;
        RECT -78.365 -178.325 -78.035 -177.995 ;
        RECT -78.365 -179.685 -78.035 -179.355 ;
        RECT -78.365 -181.93 -78.035 -180.8 ;
        RECT -78.36 -182.045 -78.04 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -77.005 241.32 -76.675 242.45 ;
        RECT -77.005 239.195 -76.675 239.525 ;
        RECT -77.005 237.835 -76.675 238.165 ;
        RECT -77.005 236.475 -76.675 236.805 ;
        RECT -77.005 235.115 -76.675 235.445 ;
        RECT -77.005 233.755 -76.675 234.085 ;
        RECT -77.005 232.395 -76.675 232.725 ;
        RECT -77.005 231.035 -76.675 231.365 ;
        RECT -77.005 229.675 -76.675 230.005 ;
        RECT -77.005 228.315 -76.675 228.645 ;
        RECT -77.005 226.955 -76.675 227.285 ;
        RECT -77.005 225.595 -76.675 225.925 ;
        RECT -77.005 224.235 -76.675 224.565 ;
        RECT -77.005 222.875 -76.675 223.205 ;
        RECT -77.005 221.515 -76.675 221.845 ;
        RECT -77.005 220.155 -76.675 220.485 ;
        RECT -77.005 218.795 -76.675 219.125 ;
        RECT -77.005 217.435 -76.675 217.765 ;
        RECT -77.005 216.075 -76.675 216.405 ;
        RECT -77.005 214.715 -76.675 215.045 ;
        RECT -77.005 213.355 -76.675 213.685 ;
        RECT -77.005 211.995 -76.675 212.325 ;
        RECT -77.005 210.635 -76.675 210.965 ;
        RECT -77.005 209.275 -76.675 209.605 ;
        RECT -77.005 207.915 -76.675 208.245 ;
        RECT -77.005 206.555 -76.675 206.885 ;
        RECT -77.005 205.195 -76.675 205.525 ;
        RECT -77.005 203.835 -76.675 204.165 ;
        RECT -77.005 202.475 -76.675 202.805 ;
        RECT -77.005 201.115 -76.675 201.445 ;
        RECT -77.005 199.755 -76.675 200.085 ;
        RECT -77.005 198.395 -76.675 198.725 ;
        RECT -77.005 197.035 -76.675 197.365 ;
        RECT -77.005 195.675 -76.675 196.005 ;
        RECT -77.005 194.315 -76.675 194.645 ;
        RECT -77.005 192.955 -76.675 193.285 ;
        RECT -77.005 191.595 -76.675 191.925 ;
        RECT -77.005 190.235 -76.675 190.565 ;
        RECT -77.005 188.875 -76.675 189.205 ;
        RECT -77.005 187.515 -76.675 187.845 ;
        RECT -77.005 186.155 -76.675 186.485 ;
        RECT -77.005 184.795 -76.675 185.125 ;
        RECT -77.005 183.435 -76.675 183.765 ;
        RECT -77.005 182.075 -76.675 182.405 ;
        RECT -77.005 180.715 -76.675 181.045 ;
        RECT -77.005 179.355 -76.675 179.685 ;
        RECT -77.005 177.995 -76.675 178.325 ;
        RECT -77.005 176.635 -76.675 176.965 ;
        RECT -77.005 175.275 -76.675 175.605 ;
        RECT -77.005 173.915 -76.675 174.245 ;
        RECT -77.005 172.555 -76.675 172.885 ;
        RECT -77.005 171.195 -76.675 171.525 ;
        RECT -77.005 169.835 -76.675 170.165 ;
        RECT -77.005 168.475 -76.675 168.805 ;
        RECT -77.005 167.115 -76.675 167.445 ;
        RECT -77.005 165.755 -76.675 166.085 ;
        RECT -77.005 164.395 -76.675 164.725 ;
        RECT -77.005 163.035 -76.675 163.365 ;
        RECT -77.005 161.675 -76.675 162.005 ;
        RECT -77.005 160.315 -76.675 160.645 ;
        RECT -77.005 158.955 -76.675 159.285 ;
        RECT -77.005 157.595 -76.675 157.925 ;
        RECT -77.005 156.235 -76.675 156.565 ;
        RECT -77.005 154.875 -76.675 155.205 ;
        RECT -77.005 153.515 -76.675 153.845 ;
        RECT -77.005 152.155 -76.675 152.485 ;
        RECT -77.005 150.795 -76.675 151.125 ;
        RECT -77.005 149.435 -76.675 149.765 ;
        RECT -77.005 148.075 -76.675 148.405 ;
        RECT -77.005 146.715 -76.675 147.045 ;
        RECT -77.005 145.355 -76.675 145.685 ;
        RECT -77.005 143.995 -76.675 144.325 ;
        RECT -77.005 142.635 -76.675 142.965 ;
        RECT -77.005 141.275 -76.675 141.605 ;
        RECT -77.005 139.915 -76.675 140.245 ;
        RECT -77.005 138.555 -76.675 138.885 ;
        RECT -77.005 137.195 -76.675 137.525 ;
        RECT -77.005 135.835 -76.675 136.165 ;
        RECT -77.005 134.475 -76.675 134.805 ;
        RECT -77.005 133.115 -76.675 133.445 ;
        RECT -77.005 131.755 -76.675 132.085 ;
        RECT -77.005 130.395 -76.675 130.725 ;
        RECT -77.005 129.035 -76.675 129.365 ;
        RECT -77.005 127.675 -76.675 128.005 ;
        RECT -77.005 126.315 -76.675 126.645 ;
        RECT -77.005 124.955 -76.675 125.285 ;
        RECT -77.005 123.595 -76.675 123.925 ;
        RECT -77.005 122.235 -76.675 122.565 ;
        RECT -77.005 120.875 -76.675 121.205 ;
        RECT -77.005 119.515 -76.675 119.845 ;
        RECT -77.005 118.155 -76.675 118.485 ;
        RECT -77.005 116.795 -76.675 117.125 ;
        RECT -77.005 115.435 -76.675 115.765 ;
        RECT -77.005 114.075 -76.675 114.405 ;
        RECT -77.005 112.715 -76.675 113.045 ;
        RECT -77.005 111.355 -76.675 111.685 ;
        RECT -77.005 109.995 -76.675 110.325 ;
        RECT -77.005 108.635 -76.675 108.965 ;
        RECT -77.005 107.275 -76.675 107.605 ;
        RECT -77.005 105.915 -76.675 106.245 ;
        RECT -77.005 104.555 -76.675 104.885 ;
        RECT -77.005 103.195 -76.675 103.525 ;
        RECT -77.005 101.835 -76.675 102.165 ;
        RECT -77.005 100.475 -76.675 100.805 ;
        RECT -77.005 99.115 -76.675 99.445 ;
        RECT -77.005 97.755 -76.675 98.085 ;
        RECT -77.005 96.395 -76.675 96.725 ;
        RECT -77.005 95.035 -76.675 95.365 ;
        RECT -77.005 93.675 -76.675 94.005 ;
        RECT -77.005 92.315 -76.675 92.645 ;
        RECT -77.005 90.955 -76.675 91.285 ;
        RECT -77.005 89.595 -76.675 89.925 ;
        RECT -77.005 88.235 -76.675 88.565 ;
        RECT -77.005 86.875 -76.675 87.205 ;
        RECT -77.005 85.515 -76.675 85.845 ;
        RECT -77.005 84.155 -76.675 84.485 ;
        RECT -77.005 82.795 -76.675 83.125 ;
        RECT -77.005 81.435 -76.675 81.765 ;
        RECT -77.005 80.075 -76.675 80.405 ;
        RECT -77.005 78.715 -76.675 79.045 ;
        RECT -77.005 77.355 -76.675 77.685 ;
        RECT -77.005 75.995 -76.675 76.325 ;
        RECT -77.005 74.635 -76.675 74.965 ;
        RECT -77.005 73.275 -76.675 73.605 ;
        RECT -77.005 71.915 -76.675 72.245 ;
        RECT -77.005 70.555 -76.675 70.885 ;
        RECT -77.005 69.195 -76.675 69.525 ;
        RECT -77.005 67.835 -76.675 68.165 ;
        RECT -77.005 66.475 -76.675 66.805 ;
        RECT -77.005 65.115 -76.675 65.445 ;
        RECT -77.005 63.755 -76.675 64.085 ;
        RECT -77.005 62.395 -76.675 62.725 ;
        RECT -77.005 61.035 -76.675 61.365 ;
        RECT -77.005 59.675 -76.675 60.005 ;
        RECT -77.005 58.315 -76.675 58.645 ;
        RECT -77.005 56.955 -76.675 57.285 ;
        RECT -77.005 55.595 -76.675 55.925 ;
        RECT -77.005 54.235 -76.675 54.565 ;
        RECT -77.005 52.875 -76.675 53.205 ;
        RECT -77.005 51.515 -76.675 51.845 ;
        RECT -77.005 50.155 -76.675 50.485 ;
        RECT -77.005 48.795 -76.675 49.125 ;
        RECT -77.005 47.435 -76.675 47.765 ;
        RECT -77.005 46.075 -76.675 46.405 ;
        RECT -77.005 44.715 -76.675 45.045 ;
        RECT -77.005 43.355 -76.675 43.685 ;
        RECT -77.005 41.995 -76.675 42.325 ;
        RECT -77.005 40.635 -76.675 40.965 ;
        RECT -77.005 39.275 -76.675 39.605 ;
        RECT -77.005 37.915 -76.675 38.245 ;
        RECT -77.005 36.555 -76.675 36.885 ;
        RECT -77.005 35.195 -76.675 35.525 ;
        RECT -77.005 33.835 -76.675 34.165 ;
        RECT -77.005 32.475 -76.675 32.805 ;
        RECT -77.005 31.115 -76.675 31.445 ;
        RECT -77.005 29.755 -76.675 30.085 ;
        RECT -77.005 28.395 -76.675 28.725 ;
        RECT -77.005 27.035 -76.675 27.365 ;
        RECT -77.005 25.675 -76.675 26.005 ;
        RECT -77.005 24.315 -76.675 24.645 ;
        RECT -77.005 22.955 -76.675 23.285 ;
        RECT -77.005 21.595 -76.675 21.925 ;
        RECT -77.005 20.235 -76.675 20.565 ;
        RECT -77.005 18.875 -76.675 19.205 ;
        RECT -77.005 17.515 -76.675 17.845 ;
        RECT -77.005 16.155 -76.675 16.485 ;
        RECT -77.005 14.795 -76.675 15.125 ;
        RECT -77.005 13.435 -76.675 13.765 ;
        RECT -77.005 12.075 -76.675 12.405 ;
        RECT -77.005 10.715 -76.675 11.045 ;
        RECT -77.005 9.355 -76.675 9.685 ;
        RECT -77.005 7.995 -76.675 8.325 ;
        RECT -77.005 6.635 -76.675 6.965 ;
        RECT -77.005 5.275 -76.675 5.605 ;
        RECT -77.005 3.915 -76.675 4.245 ;
        RECT -77.005 2.555 -76.675 2.885 ;
        RECT -77.005 1.195 -76.675 1.525 ;
        RECT -77.005 -0.165 -76.675 0.165 ;
        RECT -77.005 -1.525 -76.675 -1.195 ;
        RECT -77.005 -2.885 -76.675 -2.555 ;
        RECT -77.005 -4.245 -76.675 -3.915 ;
        RECT -77.005 -5.605 -76.675 -5.275 ;
        RECT -77.005 -6.965 -76.675 -6.635 ;
        RECT -77.005 -8.325 -76.675 -7.995 ;
        RECT -77.005 -9.685 -76.675 -9.355 ;
        RECT -77.005 -11.045 -76.675 -10.715 ;
        RECT -77.005 -12.405 -76.675 -12.075 ;
        RECT -77.005 -13.765 -76.675 -13.435 ;
        RECT -77.005 -15.125 -76.675 -14.795 ;
        RECT -77.005 -16.485 -76.675 -16.155 ;
        RECT -77.005 -17.845 -76.675 -17.515 ;
        RECT -77.005 -19.205 -76.675 -18.875 ;
        RECT -77.005 -20.565 -76.675 -20.235 ;
        RECT -77.005 -21.925 -76.675 -21.595 ;
        RECT -77.005 -23.285 -76.675 -22.955 ;
        RECT -77.005 -24.645 -76.675 -24.315 ;
        RECT -77.005 -26.005 -76.675 -25.675 ;
        RECT -77.005 -27.365 -76.675 -27.035 ;
        RECT -77.005 -28.725 -76.675 -28.395 ;
        RECT -77.005 -30.085 -76.675 -29.755 ;
        RECT -77.005 -31.445 -76.675 -31.115 ;
        RECT -77.005 -32.805 -76.675 -32.475 ;
        RECT -77.005 -34.165 -76.675 -33.835 ;
        RECT -77.005 -35.525 -76.675 -35.195 ;
        RECT -77.005 -36.885 -76.675 -36.555 ;
        RECT -77.005 -38.245 -76.675 -37.915 ;
        RECT -77.005 -39.605 -76.675 -39.275 ;
        RECT -77.005 -40.965 -76.675 -40.635 ;
        RECT -77.005 -42.325 -76.675 -41.995 ;
        RECT -77.005 -43.685 -76.675 -43.355 ;
        RECT -77.005 -45.045 -76.675 -44.715 ;
        RECT -77.005 -46.405 -76.675 -46.075 ;
        RECT -77.005 -47.765 -76.675 -47.435 ;
        RECT -77.005 -49.125 -76.675 -48.795 ;
        RECT -77.005 -50.485 -76.675 -50.155 ;
        RECT -77.005 -51.845 -76.675 -51.515 ;
        RECT -77.005 -53.205 -76.675 -52.875 ;
        RECT -77.005 -54.565 -76.675 -54.235 ;
        RECT -77.005 -55.925 -76.675 -55.595 ;
        RECT -77.005 -57.285 -76.675 -56.955 ;
        RECT -77.005 -58.645 -76.675 -58.315 ;
        RECT -77.005 -60.005 -76.675 -59.675 ;
        RECT -77.005 -61.365 -76.675 -61.035 ;
        RECT -77.005 -62.725 -76.675 -62.395 ;
        RECT -77.005 -64.085 -76.675 -63.755 ;
        RECT -77.005 -65.445 -76.675 -65.115 ;
        RECT -77.005 -66.805 -76.675 -66.475 ;
        RECT -77.005 -68.165 -76.675 -67.835 ;
        RECT -77.005 -69.525 -76.675 -69.195 ;
        RECT -77.005 -70.885 -76.675 -70.555 ;
        RECT -77.005 -72.245 -76.675 -71.915 ;
        RECT -77.005 -73.605 -76.675 -73.275 ;
        RECT -77.005 -74.965 -76.675 -74.635 ;
        RECT -77.005 -76.325 -76.675 -75.995 ;
        RECT -77.005 -77.685 -76.675 -77.355 ;
        RECT -77.005 -79.045 -76.675 -78.715 ;
        RECT -77.005 -80.405 -76.675 -80.075 ;
        RECT -77.005 -81.765 -76.675 -81.435 ;
        RECT -77.005 -83.125 -76.675 -82.795 ;
        RECT -77.005 -84.485 -76.675 -84.155 ;
        RECT -77.005 -85.845 -76.675 -85.515 ;
        RECT -77.005 -87.205 -76.675 -86.875 ;
        RECT -77.005 -88.565 -76.675 -88.235 ;
        RECT -77.005 -89.925 -76.675 -89.595 ;
        RECT -77.005 -91.285 -76.675 -90.955 ;
        RECT -77.005 -92.645 -76.675 -92.315 ;
        RECT -77.005 -94.005 -76.675 -93.675 ;
        RECT -77.005 -95.365 -76.675 -95.035 ;
        RECT -77.005 -96.725 -76.675 -96.395 ;
        RECT -77.005 -98.085 -76.675 -97.755 ;
        RECT -77.005 -99.445 -76.675 -99.115 ;
        RECT -77.005 -100.805 -76.675 -100.475 ;
        RECT -77.005 -102.165 -76.675 -101.835 ;
        RECT -77.005 -103.525 -76.675 -103.195 ;
        RECT -77.005 -104.885 -76.675 -104.555 ;
        RECT -77.005 -106.245 -76.675 -105.915 ;
        RECT -77.005 -107.605 -76.675 -107.275 ;
        RECT -77.005 -108.965 -76.675 -108.635 ;
        RECT -77.005 -110.325 -76.675 -109.995 ;
        RECT -77.005 -111.685 -76.675 -111.355 ;
        RECT -77.005 -113.045 -76.675 -112.715 ;
        RECT -77.005 -114.405 -76.675 -114.075 ;
        RECT -77.005 -115.765 -76.675 -115.435 ;
        RECT -77.005 -117.125 -76.675 -116.795 ;
        RECT -77.005 -118.485 -76.675 -118.155 ;
        RECT -77.005 -119.845 -76.675 -119.515 ;
        RECT -77.005 -121.205 -76.675 -120.875 ;
        RECT -77.005 -122.565 -76.675 -122.235 ;
        RECT -77.005 -123.925 -76.675 -123.595 ;
        RECT -77.005 -125.285 -76.675 -124.955 ;
        RECT -77.005 -126.645 -76.675 -126.315 ;
        RECT -77.005 -128.005 -76.675 -127.675 ;
        RECT -77.005 -129.365 -76.675 -129.035 ;
        RECT -77.005 -130.725 -76.675 -130.395 ;
        RECT -77.005 -132.085 -76.675 -131.755 ;
        RECT -77.005 -133.445 -76.675 -133.115 ;
        RECT -77.005 -134.805 -76.675 -134.475 ;
        RECT -77.005 -136.165 -76.675 -135.835 ;
        RECT -77.005 -137.525 -76.675 -137.195 ;
        RECT -77.005 -138.885 -76.675 -138.555 ;
        RECT -77.005 -140.245 -76.675 -139.915 ;
        RECT -77.005 -141.605 -76.675 -141.275 ;
        RECT -77.005 -142.965 -76.675 -142.635 ;
        RECT -77.005 -144.325 -76.675 -143.995 ;
        RECT -77.005 -145.685 -76.675 -145.355 ;
        RECT -77.005 -147.045 -76.675 -146.715 ;
        RECT -77.005 -148.405 -76.675 -148.075 ;
        RECT -77.005 -149.765 -76.675 -149.435 ;
        RECT -77.005 -151.125 -76.675 -150.795 ;
        RECT -77.005 -152.485 -76.675 -152.155 ;
        RECT -77.005 -153.845 -76.675 -153.515 ;
        RECT -77.005 -155.205 -76.675 -154.875 ;
        RECT -77.005 -156.565 -76.675 -156.235 ;
        RECT -77.005 -157.925 -76.675 -157.595 ;
        RECT -77.005 -159.285 -76.675 -158.955 ;
        RECT -77.005 -160.645 -76.675 -160.315 ;
        RECT -77.005 -162.005 -76.675 -161.675 ;
        RECT -77.005 -163.365 -76.675 -163.035 ;
        RECT -77.005 -164.725 -76.675 -164.395 ;
        RECT -77.005 -166.085 -76.675 -165.755 ;
        RECT -77.005 -167.445 -76.675 -167.115 ;
        RECT -77.005 -168.805 -76.675 -168.475 ;
        RECT -77.005 -171.525 -76.675 -171.195 ;
        RECT -77.005 -172.885 -76.675 -172.555 ;
        RECT -77.005 -175.605 -76.675 -175.275 ;
        RECT -77.005 -176.685 -76.675 -176.355 ;
        RECT -77.005 -178.325 -76.675 -177.995 ;
        RECT -77.005 -179.685 -76.675 -179.355 ;
        RECT -77.005 -181.93 -76.675 -180.8 ;
        RECT -77 -182.045 -76.68 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -75.645 -24.645 -75.315 -24.315 ;
        RECT -75.645 -26.005 -75.315 -25.675 ;
        RECT -75.645 -27.365 -75.315 -27.035 ;
        RECT -75.645 -28.725 -75.315 -28.395 ;
        RECT -75.645 -30.085 -75.315 -29.755 ;
        RECT -75.645 -31.445 -75.315 -31.115 ;
        RECT -75.645 -32.805 -75.315 -32.475 ;
        RECT -75.645 -34.165 -75.315 -33.835 ;
        RECT -75.645 -35.525 -75.315 -35.195 ;
        RECT -75.645 -36.885 -75.315 -36.555 ;
        RECT -75.645 -38.245 -75.315 -37.915 ;
        RECT -75.645 -39.605 -75.315 -39.275 ;
        RECT -75.645 -40.965 -75.315 -40.635 ;
        RECT -75.645 -42.325 -75.315 -41.995 ;
        RECT -75.645 -43.685 -75.315 -43.355 ;
        RECT -75.645 -45.045 -75.315 -44.715 ;
        RECT -75.645 -46.405 -75.315 -46.075 ;
        RECT -75.645 -47.765 -75.315 -47.435 ;
        RECT -75.645 -49.125 -75.315 -48.795 ;
        RECT -75.645 -50.485 -75.315 -50.155 ;
        RECT -75.645 -51.845 -75.315 -51.515 ;
        RECT -75.645 -53.205 -75.315 -52.875 ;
        RECT -75.645 -54.565 -75.315 -54.235 ;
        RECT -75.645 -55.925 -75.315 -55.595 ;
        RECT -75.645 -57.285 -75.315 -56.955 ;
        RECT -75.645 -58.645 -75.315 -58.315 ;
        RECT -75.645 -60.005 -75.315 -59.675 ;
        RECT -75.645 -61.365 -75.315 -61.035 ;
        RECT -75.645 -62.725 -75.315 -62.395 ;
        RECT -75.645 -64.085 -75.315 -63.755 ;
        RECT -75.645 -65.445 -75.315 -65.115 ;
        RECT -75.645 -66.805 -75.315 -66.475 ;
        RECT -75.645 -68.165 -75.315 -67.835 ;
        RECT -75.645 -69.525 -75.315 -69.195 ;
        RECT -75.645 -70.885 -75.315 -70.555 ;
        RECT -75.645 -72.245 -75.315 -71.915 ;
        RECT -75.645 -73.605 -75.315 -73.275 ;
        RECT -75.645 -74.965 -75.315 -74.635 ;
        RECT -75.645 -76.325 -75.315 -75.995 ;
        RECT -75.645 -77.685 -75.315 -77.355 ;
        RECT -75.645 -79.045 -75.315 -78.715 ;
        RECT -75.645 -80.405 -75.315 -80.075 ;
        RECT -75.645 -81.765 -75.315 -81.435 ;
        RECT -75.645 -83.125 -75.315 -82.795 ;
        RECT -75.645 -84.485 -75.315 -84.155 ;
        RECT -75.645 -85.845 -75.315 -85.515 ;
        RECT -75.645 -87.205 -75.315 -86.875 ;
        RECT -75.645 -88.565 -75.315 -88.235 ;
        RECT -75.645 -89.925 -75.315 -89.595 ;
        RECT -75.645 -91.285 -75.315 -90.955 ;
        RECT -75.645 -92.645 -75.315 -92.315 ;
        RECT -75.645 -94.005 -75.315 -93.675 ;
        RECT -75.645 -95.365 -75.315 -95.035 ;
        RECT -75.645 -96.725 -75.315 -96.395 ;
        RECT -75.645 -98.085 -75.315 -97.755 ;
        RECT -75.645 -99.445 -75.315 -99.115 ;
        RECT -75.645 -100.805 -75.315 -100.475 ;
        RECT -75.645 -102.165 -75.315 -101.835 ;
        RECT -75.645 -103.525 -75.315 -103.195 ;
        RECT -75.645 -104.885 -75.315 -104.555 ;
        RECT -75.645 -106.245 -75.315 -105.915 ;
        RECT -75.645 -107.605 -75.315 -107.275 ;
        RECT -75.645 -108.965 -75.315 -108.635 ;
        RECT -75.645 -110.325 -75.315 -109.995 ;
        RECT -75.645 -111.685 -75.315 -111.355 ;
        RECT -75.645 -113.045 -75.315 -112.715 ;
        RECT -75.645 -114.405 -75.315 -114.075 ;
        RECT -75.645 -115.765 -75.315 -115.435 ;
        RECT -75.645 -117.125 -75.315 -116.795 ;
        RECT -75.645 -118.485 -75.315 -118.155 ;
        RECT -75.645 -119.845 -75.315 -119.515 ;
        RECT -75.645 -121.205 -75.315 -120.875 ;
        RECT -75.645 -122.565 -75.315 -122.235 ;
        RECT -75.645 -123.925 -75.315 -123.595 ;
        RECT -75.645 -125.285 -75.315 -124.955 ;
        RECT -75.645 -126.645 -75.315 -126.315 ;
        RECT -75.645 -128.005 -75.315 -127.675 ;
        RECT -75.645 -129.365 -75.315 -129.035 ;
        RECT -75.645 -130.725 -75.315 -130.395 ;
        RECT -75.645 -132.085 -75.315 -131.755 ;
        RECT -75.645 -133.445 -75.315 -133.115 ;
        RECT -75.645 -134.805 -75.315 -134.475 ;
        RECT -75.645 -136.165 -75.315 -135.835 ;
        RECT -75.645 -137.525 -75.315 -137.195 ;
        RECT -75.645 -138.885 -75.315 -138.555 ;
        RECT -75.645 -140.245 -75.315 -139.915 ;
        RECT -75.645 -141.605 -75.315 -141.275 ;
        RECT -75.645 -142.965 -75.315 -142.635 ;
        RECT -75.645 -144.325 -75.315 -143.995 ;
        RECT -75.645 -145.685 -75.315 -145.355 ;
        RECT -75.645 -147.045 -75.315 -146.715 ;
        RECT -75.645 -148.405 -75.315 -148.075 ;
        RECT -75.645 -149.765 -75.315 -149.435 ;
        RECT -75.645 -151.125 -75.315 -150.795 ;
        RECT -75.645 -152.485 -75.315 -152.155 ;
        RECT -75.645 -153.845 -75.315 -153.515 ;
        RECT -75.645 -155.205 -75.315 -154.875 ;
        RECT -75.645 -156.565 -75.315 -156.235 ;
        RECT -75.645 -157.925 -75.315 -157.595 ;
        RECT -75.645 -159.285 -75.315 -158.955 ;
        RECT -75.645 -160.645 -75.315 -160.315 ;
        RECT -75.645 -162.005 -75.315 -161.675 ;
        RECT -75.645 -163.365 -75.315 -163.035 ;
        RECT -75.645 -164.725 -75.315 -164.395 ;
        RECT -75.645 -166.085 -75.315 -165.755 ;
        RECT -75.645 -167.445 -75.315 -167.115 ;
        RECT -75.645 -168.805 -75.315 -168.475 ;
        RECT -75.645 -171.525 -75.315 -171.195 ;
        RECT -75.645 -174.245 -75.315 -173.915 ;
        RECT -75.645 -175.605 -75.315 -175.275 ;
        RECT -75.645 -176.685 -75.315 -176.355 ;
        RECT -75.645 -178.325 -75.315 -177.995 ;
        RECT -75.645 -179.685 -75.315 -179.355 ;
        RECT -75.645 -181.93 -75.315 -180.8 ;
        RECT -75.64 -182.045 -75.32 242.565 ;
        RECT -75.645 241.32 -75.315 242.45 ;
        RECT -75.645 239.195 -75.315 239.525 ;
        RECT -75.645 237.835 -75.315 238.165 ;
        RECT -75.645 236.475 -75.315 236.805 ;
        RECT -75.645 235.115 -75.315 235.445 ;
        RECT -75.645 233.755 -75.315 234.085 ;
        RECT -75.645 232.395 -75.315 232.725 ;
        RECT -75.645 231.035 -75.315 231.365 ;
        RECT -75.645 229.675 -75.315 230.005 ;
        RECT -75.645 228.315 -75.315 228.645 ;
        RECT -75.645 226.955 -75.315 227.285 ;
        RECT -75.645 225.595 -75.315 225.925 ;
        RECT -75.645 224.235 -75.315 224.565 ;
        RECT -75.645 222.875 -75.315 223.205 ;
        RECT -75.645 221.515 -75.315 221.845 ;
        RECT -75.645 220.155 -75.315 220.485 ;
        RECT -75.645 218.795 -75.315 219.125 ;
        RECT -75.645 217.435 -75.315 217.765 ;
        RECT -75.645 216.075 -75.315 216.405 ;
        RECT -75.645 214.715 -75.315 215.045 ;
        RECT -75.645 213.355 -75.315 213.685 ;
        RECT -75.645 211.995 -75.315 212.325 ;
        RECT -75.645 210.635 -75.315 210.965 ;
        RECT -75.645 209.275 -75.315 209.605 ;
        RECT -75.645 207.915 -75.315 208.245 ;
        RECT -75.645 206.555 -75.315 206.885 ;
        RECT -75.645 205.195 -75.315 205.525 ;
        RECT -75.645 203.835 -75.315 204.165 ;
        RECT -75.645 202.475 -75.315 202.805 ;
        RECT -75.645 201.115 -75.315 201.445 ;
        RECT -75.645 199.755 -75.315 200.085 ;
        RECT -75.645 198.395 -75.315 198.725 ;
        RECT -75.645 197.035 -75.315 197.365 ;
        RECT -75.645 195.675 -75.315 196.005 ;
        RECT -75.645 194.315 -75.315 194.645 ;
        RECT -75.645 192.955 -75.315 193.285 ;
        RECT -75.645 191.595 -75.315 191.925 ;
        RECT -75.645 190.235 -75.315 190.565 ;
        RECT -75.645 188.875 -75.315 189.205 ;
        RECT -75.645 187.515 -75.315 187.845 ;
        RECT -75.645 186.155 -75.315 186.485 ;
        RECT -75.645 184.795 -75.315 185.125 ;
        RECT -75.645 183.435 -75.315 183.765 ;
        RECT -75.645 182.075 -75.315 182.405 ;
        RECT -75.645 180.715 -75.315 181.045 ;
        RECT -75.645 179.355 -75.315 179.685 ;
        RECT -75.645 177.995 -75.315 178.325 ;
        RECT -75.645 176.635 -75.315 176.965 ;
        RECT -75.645 175.275 -75.315 175.605 ;
        RECT -75.645 173.915 -75.315 174.245 ;
        RECT -75.645 172.555 -75.315 172.885 ;
        RECT -75.645 171.195 -75.315 171.525 ;
        RECT -75.645 169.835 -75.315 170.165 ;
        RECT -75.645 168.475 -75.315 168.805 ;
        RECT -75.645 167.115 -75.315 167.445 ;
        RECT -75.645 165.755 -75.315 166.085 ;
        RECT -75.645 164.395 -75.315 164.725 ;
        RECT -75.645 163.035 -75.315 163.365 ;
        RECT -75.645 161.675 -75.315 162.005 ;
        RECT -75.645 160.315 -75.315 160.645 ;
        RECT -75.645 158.955 -75.315 159.285 ;
        RECT -75.645 157.595 -75.315 157.925 ;
        RECT -75.645 156.235 -75.315 156.565 ;
        RECT -75.645 154.875 -75.315 155.205 ;
        RECT -75.645 153.515 -75.315 153.845 ;
        RECT -75.645 152.155 -75.315 152.485 ;
        RECT -75.645 150.795 -75.315 151.125 ;
        RECT -75.645 149.435 -75.315 149.765 ;
        RECT -75.645 148.075 -75.315 148.405 ;
        RECT -75.645 146.715 -75.315 147.045 ;
        RECT -75.645 145.355 -75.315 145.685 ;
        RECT -75.645 143.995 -75.315 144.325 ;
        RECT -75.645 142.635 -75.315 142.965 ;
        RECT -75.645 141.275 -75.315 141.605 ;
        RECT -75.645 139.915 -75.315 140.245 ;
        RECT -75.645 138.555 -75.315 138.885 ;
        RECT -75.645 137.195 -75.315 137.525 ;
        RECT -75.645 135.835 -75.315 136.165 ;
        RECT -75.645 134.475 -75.315 134.805 ;
        RECT -75.645 133.115 -75.315 133.445 ;
        RECT -75.645 131.755 -75.315 132.085 ;
        RECT -75.645 130.395 -75.315 130.725 ;
        RECT -75.645 129.035 -75.315 129.365 ;
        RECT -75.645 127.675 -75.315 128.005 ;
        RECT -75.645 126.315 -75.315 126.645 ;
        RECT -75.645 124.955 -75.315 125.285 ;
        RECT -75.645 123.595 -75.315 123.925 ;
        RECT -75.645 122.235 -75.315 122.565 ;
        RECT -75.645 120.875 -75.315 121.205 ;
        RECT -75.645 119.515 -75.315 119.845 ;
        RECT -75.645 118.155 -75.315 118.485 ;
        RECT -75.645 116.795 -75.315 117.125 ;
        RECT -75.645 115.435 -75.315 115.765 ;
        RECT -75.645 114.075 -75.315 114.405 ;
        RECT -75.645 112.715 -75.315 113.045 ;
        RECT -75.645 111.355 -75.315 111.685 ;
        RECT -75.645 109.995 -75.315 110.325 ;
        RECT -75.645 108.635 -75.315 108.965 ;
        RECT -75.645 107.275 -75.315 107.605 ;
        RECT -75.645 105.915 -75.315 106.245 ;
        RECT -75.645 104.555 -75.315 104.885 ;
        RECT -75.645 103.195 -75.315 103.525 ;
        RECT -75.645 101.835 -75.315 102.165 ;
        RECT -75.645 100.475 -75.315 100.805 ;
        RECT -75.645 99.115 -75.315 99.445 ;
        RECT -75.645 97.755 -75.315 98.085 ;
        RECT -75.645 96.395 -75.315 96.725 ;
        RECT -75.645 95.035 -75.315 95.365 ;
        RECT -75.645 93.675 -75.315 94.005 ;
        RECT -75.645 92.315 -75.315 92.645 ;
        RECT -75.645 90.955 -75.315 91.285 ;
        RECT -75.645 89.595 -75.315 89.925 ;
        RECT -75.645 88.235 -75.315 88.565 ;
        RECT -75.645 86.875 -75.315 87.205 ;
        RECT -75.645 85.515 -75.315 85.845 ;
        RECT -75.645 84.155 -75.315 84.485 ;
        RECT -75.645 82.795 -75.315 83.125 ;
        RECT -75.645 81.435 -75.315 81.765 ;
        RECT -75.645 80.075 -75.315 80.405 ;
        RECT -75.645 78.715 -75.315 79.045 ;
        RECT -75.645 77.355 -75.315 77.685 ;
        RECT -75.645 75.995 -75.315 76.325 ;
        RECT -75.645 74.635 -75.315 74.965 ;
        RECT -75.645 73.275 -75.315 73.605 ;
        RECT -75.645 71.915 -75.315 72.245 ;
        RECT -75.645 70.555 -75.315 70.885 ;
        RECT -75.645 69.195 -75.315 69.525 ;
        RECT -75.645 67.835 -75.315 68.165 ;
        RECT -75.645 66.475 -75.315 66.805 ;
        RECT -75.645 65.115 -75.315 65.445 ;
        RECT -75.645 63.755 -75.315 64.085 ;
        RECT -75.645 62.395 -75.315 62.725 ;
        RECT -75.645 61.035 -75.315 61.365 ;
        RECT -75.645 59.675 -75.315 60.005 ;
        RECT -75.645 58.315 -75.315 58.645 ;
        RECT -75.645 56.955 -75.315 57.285 ;
        RECT -75.645 55.595 -75.315 55.925 ;
        RECT -75.645 54.235 -75.315 54.565 ;
        RECT -75.645 52.875 -75.315 53.205 ;
        RECT -75.645 51.515 -75.315 51.845 ;
        RECT -75.645 50.155 -75.315 50.485 ;
        RECT -75.645 48.795 -75.315 49.125 ;
        RECT -75.645 47.435 -75.315 47.765 ;
        RECT -75.645 46.075 -75.315 46.405 ;
        RECT -75.645 44.715 -75.315 45.045 ;
        RECT -75.645 43.355 -75.315 43.685 ;
        RECT -75.645 41.995 -75.315 42.325 ;
        RECT -75.645 40.635 -75.315 40.965 ;
        RECT -75.645 39.275 -75.315 39.605 ;
        RECT -75.645 37.915 -75.315 38.245 ;
        RECT -75.645 36.555 -75.315 36.885 ;
        RECT -75.645 35.195 -75.315 35.525 ;
        RECT -75.645 33.835 -75.315 34.165 ;
        RECT -75.645 32.475 -75.315 32.805 ;
        RECT -75.645 31.115 -75.315 31.445 ;
        RECT -75.645 29.755 -75.315 30.085 ;
        RECT -75.645 28.395 -75.315 28.725 ;
        RECT -75.645 27.035 -75.315 27.365 ;
        RECT -75.645 25.675 -75.315 26.005 ;
        RECT -75.645 24.315 -75.315 24.645 ;
        RECT -75.645 22.955 -75.315 23.285 ;
        RECT -75.645 21.595 -75.315 21.925 ;
        RECT -75.645 20.235 -75.315 20.565 ;
        RECT -75.645 18.875 -75.315 19.205 ;
        RECT -75.645 17.515 -75.315 17.845 ;
        RECT -75.645 16.155 -75.315 16.485 ;
        RECT -75.645 14.795 -75.315 15.125 ;
        RECT -75.645 13.435 -75.315 13.765 ;
        RECT -75.645 12.075 -75.315 12.405 ;
        RECT -75.645 10.715 -75.315 11.045 ;
        RECT -75.645 9.355 -75.315 9.685 ;
        RECT -75.645 7.995 -75.315 8.325 ;
        RECT -75.645 6.635 -75.315 6.965 ;
        RECT -75.645 5.275 -75.315 5.605 ;
        RECT -75.645 3.915 -75.315 4.245 ;
        RECT -75.645 2.555 -75.315 2.885 ;
        RECT -75.645 1.195 -75.315 1.525 ;
        RECT -75.645 -0.165 -75.315 0.165 ;
        RECT -75.645 -1.525 -75.315 -1.195 ;
        RECT -75.645 -2.885 -75.315 -2.555 ;
        RECT -75.645 -4.245 -75.315 -3.915 ;
        RECT -75.645 -5.605 -75.315 -5.275 ;
        RECT -75.645 -6.965 -75.315 -6.635 ;
        RECT -75.645 -8.325 -75.315 -7.995 ;
        RECT -75.645 -9.685 -75.315 -9.355 ;
        RECT -75.645 -11.045 -75.315 -10.715 ;
        RECT -75.645 -12.405 -75.315 -12.075 ;
        RECT -75.645 -13.765 -75.315 -13.435 ;
        RECT -75.645 -15.125 -75.315 -14.795 ;
        RECT -75.645 -16.485 -75.315 -16.155 ;
        RECT -75.645 -17.845 -75.315 -17.515 ;
        RECT -75.645 -19.205 -75.315 -18.875 ;
        RECT -75.645 -20.565 -75.315 -20.235 ;
        RECT -75.645 -21.925 -75.315 -21.595 ;
        RECT -75.645 -23.285 -75.315 -22.955 ;
    END
    PORT
      LAYER met3 ;
        RECT -81.085 241.32 -80.755 242.45 ;
        RECT -81.085 239.195 -80.755 239.525 ;
        RECT -81.085 237.835 -80.755 238.165 ;
        RECT -81.085 236.475 -80.755 236.805 ;
        RECT -81.085 235.115 -80.755 235.445 ;
        RECT -81.085 233.755 -80.755 234.085 ;
        RECT -81.085 232.395 -80.755 232.725 ;
        RECT -81.085 231.035 -80.755 231.365 ;
        RECT -81.085 229.675 -80.755 230.005 ;
        RECT -81.085 228.315 -80.755 228.645 ;
        RECT -81.085 226.955 -80.755 227.285 ;
        RECT -81.085 225.595 -80.755 225.925 ;
        RECT -81.085 224.235 -80.755 224.565 ;
        RECT -81.085 222.875 -80.755 223.205 ;
        RECT -81.085 221.515 -80.755 221.845 ;
        RECT -81.085 220.155 -80.755 220.485 ;
        RECT -81.085 218.795 -80.755 219.125 ;
        RECT -81.085 217.435 -80.755 217.765 ;
        RECT -81.085 216.075 -80.755 216.405 ;
        RECT -81.085 214.715 -80.755 215.045 ;
        RECT -81.085 213.355 -80.755 213.685 ;
        RECT -81.085 211.995 -80.755 212.325 ;
        RECT -81.085 210.635 -80.755 210.965 ;
        RECT -81.085 209.275 -80.755 209.605 ;
        RECT -81.085 207.915 -80.755 208.245 ;
        RECT -81.085 206.555 -80.755 206.885 ;
        RECT -81.085 205.195 -80.755 205.525 ;
        RECT -81.085 203.835 -80.755 204.165 ;
        RECT -81.085 202.475 -80.755 202.805 ;
        RECT -81.085 201.115 -80.755 201.445 ;
        RECT -81.085 199.755 -80.755 200.085 ;
        RECT -81.085 198.395 -80.755 198.725 ;
        RECT -81.085 197.035 -80.755 197.365 ;
        RECT -81.085 195.675 -80.755 196.005 ;
        RECT -81.085 194.315 -80.755 194.645 ;
        RECT -81.085 192.955 -80.755 193.285 ;
        RECT -81.085 191.595 -80.755 191.925 ;
        RECT -81.085 190.235 -80.755 190.565 ;
        RECT -81.085 188.875 -80.755 189.205 ;
        RECT -81.085 187.515 -80.755 187.845 ;
        RECT -81.085 186.155 -80.755 186.485 ;
        RECT -81.085 184.795 -80.755 185.125 ;
        RECT -81.085 183.435 -80.755 183.765 ;
        RECT -81.085 182.075 -80.755 182.405 ;
        RECT -81.085 180.715 -80.755 181.045 ;
        RECT -81.085 179.355 -80.755 179.685 ;
        RECT -81.085 177.995 -80.755 178.325 ;
        RECT -81.085 176.635 -80.755 176.965 ;
        RECT -81.085 175.275 -80.755 175.605 ;
        RECT -81.085 173.915 -80.755 174.245 ;
        RECT -81.085 172.555 -80.755 172.885 ;
        RECT -81.085 171.195 -80.755 171.525 ;
        RECT -81.085 169.835 -80.755 170.165 ;
        RECT -81.085 168.475 -80.755 168.805 ;
        RECT -81.085 167.115 -80.755 167.445 ;
        RECT -81.085 165.755 -80.755 166.085 ;
        RECT -81.085 164.395 -80.755 164.725 ;
        RECT -81.085 163.035 -80.755 163.365 ;
        RECT -81.085 161.675 -80.755 162.005 ;
        RECT -81.085 160.315 -80.755 160.645 ;
        RECT -81.085 158.955 -80.755 159.285 ;
        RECT -81.085 157.595 -80.755 157.925 ;
        RECT -81.085 156.235 -80.755 156.565 ;
        RECT -81.085 154.875 -80.755 155.205 ;
        RECT -81.085 153.515 -80.755 153.845 ;
        RECT -81.085 152.155 -80.755 152.485 ;
        RECT -81.085 150.795 -80.755 151.125 ;
        RECT -81.085 149.435 -80.755 149.765 ;
        RECT -81.085 148.075 -80.755 148.405 ;
        RECT -81.085 146.715 -80.755 147.045 ;
        RECT -81.085 145.355 -80.755 145.685 ;
        RECT -81.085 143.995 -80.755 144.325 ;
        RECT -81.085 142.635 -80.755 142.965 ;
        RECT -81.085 141.275 -80.755 141.605 ;
        RECT -81.085 139.915 -80.755 140.245 ;
        RECT -81.085 138.555 -80.755 138.885 ;
        RECT -81.085 137.195 -80.755 137.525 ;
        RECT -81.085 135.835 -80.755 136.165 ;
        RECT -81.085 134.475 -80.755 134.805 ;
        RECT -81.085 133.115 -80.755 133.445 ;
        RECT -81.085 131.755 -80.755 132.085 ;
        RECT -81.085 130.395 -80.755 130.725 ;
        RECT -81.085 129.035 -80.755 129.365 ;
        RECT -81.085 127.675 -80.755 128.005 ;
        RECT -81.085 126.315 -80.755 126.645 ;
        RECT -81.085 124.955 -80.755 125.285 ;
        RECT -81.085 123.595 -80.755 123.925 ;
        RECT -81.085 122.235 -80.755 122.565 ;
        RECT -81.085 120.875 -80.755 121.205 ;
        RECT -81.085 119.515 -80.755 119.845 ;
        RECT -81.085 118.155 -80.755 118.485 ;
        RECT -81.085 116.795 -80.755 117.125 ;
        RECT -81.085 115.435 -80.755 115.765 ;
        RECT -81.085 114.075 -80.755 114.405 ;
        RECT -81.085 112.715 -80.755 113.045 ;
        RECT -81.085 111.355 -80.755 111.685 ;
        RECT -81.085 109.995 -80.755 110.325 ;
        RECT -81.085 108.635 -80.755 108.965 ;
        RECT -81.085 107.275 -80.755 107.605 ;
        RECT -81.085 105.915 -80.755 106.245 ;
        RECT -81.085 104.555 -80.755 104.885 ;
        RECT -81.085 103.195 -80.755 103.525 ;
        RECT -81.085 101.835 -80.755 102.165 ;
        RECT -81.085 100.475 -80.755 100.805 ;
        RECT -81.085 99.115 -80.755 99.445 ;
        RECT -81.085 97.755 -80.755 98.085 ;
        RECT -81.085 96.395 -80.755 96.725 ;
        RECT -81.085 95.035 -80.755 95.365 ;
        RECT -81.085 93.675 -80.755 94.005 ;
        RECT -81.085 92.315 -80.755 92.645 ;
        RECT -81.085 90.955 -80.755 91.285 ;
        RECT -81.085 89.595 -80.755 89.925 ;
        RECT -81.085 88.235 -80.755 88.565 ;
        RECT -81.085 86.875 -80.755 87.205 ;
        RECT -81.085 85.515 -80.755 85.845 ;
        RECT -81.085 84.155 -80.755 84.485 ;
        RECT -81.085 82.795 -80.755 83.125 ;
        RECT -81.085 81.435 -80.755 81.765 ;
        RECT -81.085 80.075 -80.755 80.405 ;
        RECT -81.085 78.715 -80.755 79.045 ;
        RECT -81.085 77.355 -80.755 77.685 ;
        RECT -81.085 75.995 -80.755 76.325 ;
        RECT -81.085 74.635 -80.755 74.965 ;
        RECT -81.085 73.275 -80.755 73.605 ;
        RECT -81.085 71.915 -80.755 72.245 ;
        RECT -81.085 70.555 -80.755 70.885 ;
        RECT -81.085 69.195 -80.755 69.525 ;
        RECT -81.085 67.835 -80.755 68.165 ;
        RECT -81.085 66.475 -80.755 66.805 ;
        RECT -81.085 65.115 -80.755 65.445 ;
        RECT -81.085 63.755 -80.755 64.085 ;
        RECT -81.085 62.395 -80.755 62.725 ;
        RECT -81.085 61.035 -80.755 61.365 ;
        RECT -81.085 59.675 -80.755 60.005 ;
        RECT -81.085 58.315 -80.755 58.645 ;
        RECT -81.085 56.955 -80.755 57.285 ;
        RECT -81.085 55.595 -80.755 55.925 ;
        RECT -81.085 54.235 -80.755 54.565 ;
        RECT -81.085 52.875 -80.755 53.205 ;
        RECT -81.085 51.515 -80.755 51.845 ;
        RECT -81.085 50.155 -80.755 50.485 ;
        RECT -81.085 48.795 -80.755 49.125 ;
        RECT -81.085 47.435 -80.755 47.765 ;
        RECT -81.085 46.075 -80.755 46.405 ;
        RECT -81.085 44.715 -80.755 45.045 ;
        RECT -81.085 43.355 -80.755 43.685 ;
        RECT -81.085 41.995 -80.755 42.325 ;
        RECT -81.085 40.635 -80.755 40.965 ;
        RECT -81.085 39.275 -80.755 39.605 ;
        RECT -81.085 37.915 -80.755 38.245 ;
        RECT -81.085 36.555 -80.755 36.885 ;
        RECT -81.085 35.195 -80.755 35.525 ;
        RECT -81.085 33.835 -80.755 34.165 ;
        RECT -81.085 32.475 -80.755 32.805 ;
        RECT -81.085 31.115 -80.755 31.445 ;
        RECT -81.085 29.755 -80.755 30.085 ;
        RECT -81.085 28.395 -80.755 28.725 ;
        RECT -81.085 27.035 -80.755 27.365 ;
        RECT -81.085 25.675 -80.755 26.005 ;
        RECT -81.085 24.315 -80.755 24.645 ;
        RECT -81.085 22.955 -80.755 23.285 ;
        RECT -81.085 21.595 -80.755 21.925 ;
        RECT -81.085 20.235 -80.755 20.565 ;
        RECT -81.085 18.875 -80.755 19.205 ;
        RECT -81.085 17.515 -80.755 17.845 ;
        RECT -81.085 16.155 -80.755 16.485 ;
        RECT -81.085 14.795 -80.755 15.125 ;
        RECT -81.085 13.435 -80.755 13.765 ;
        RECT -81.085 12.075 -80.755 12.405 ;
        RECT -81.085 10.715 -80.755 11.045 ;
        RECT -81.085 9.355 -80.755 9.685 ;
        RECT -81.085 7.995 -80.755 8.325 ;
        RECT -81.085 6.635 -80.755 6.965 ;
        RECT -81.085 5.275 -80.755 5.605 ;
        RECT -81.085 3.915 -80.755 4.245 ;
        RECT -81.085 2.555 -80.755 2.885 ;
        RECT -81.085 1.195 -80.755 1.525 ;
        RECT -81.085 -0.165 -80.755 0.165 ;
        RECT -81.085 -1.525 -80.755 -1.195 ;
        RECT -81.085 -2.885 -80.755 -2.555 ;
        RECT -81.085 -4.245 -80.755 -3.915 ;
        RECT -81.085 -5.605 -80.755 -5.275 ;
        RECT -81.085 -6.965 -80.755 -6.635 ;
        RECT -81.085 -8.325 -80.755 -7.995 ;
        RECT -81.085 -9.685 -80.755 -9.355 ;
        RECT -81.085 -11.045 -80.755 -10.715 ;
        RECT -81.085 -12.405 -80.755 -12.075 ;
        RECT -81.085 -13.765 -80.755 -13.435 ;
        RECT -81.085 -15.125 -80.755 -14.795 ;
        RECT -81.085 -16.485 -80.755 -16.155 ;
        RECT -81.085 -17.845 -80.755 -17.515 ;
        RECT -81.085 -19.205 -80.755 -18.875 ;
        RECT -81.085 -20.565 -80.755 -20.235 ;
        RECT -81.085 -21.925 -80.755 -21.595 ;
        RECT -81.085 -23.285 -80.755 -22.955 ;
        RECT -81.085 -24.645 -80.755 -24.315 ;
        RECT -81.085 -26.005 -80.755 -25.675 ;
        RECT -81.085 -27.365 -80.755 -27.035 ;
        RECT -81.085 -28.725 -80.755 -28.395 ;
        RECT -81.085 -30.085 -80.755 -29.755 ;
        RECT -81.085 -31.445 -80.755 -31.115 ;
        RECT -81.085 -32.805 -80.755 -32.475 ;
        RECT -81.085 -34.165 -80.755 -33.835 ;
        RECT -81.085 -35.525 -80.755 -35.195 ;
        RECT -81.085 -36.885 -80.755 -36.555 ;
        RECT -81.085 -38.245 -80.755 -37.915 ;
        RECT -81.085 -39.605 -80.755 -39.275 ;
        RECT -81.085 -40.965 -80.755 -40.635 ;
        RECT -81.085 -42.325 -80.755 -41.995 ;
        RECT -81.085 -43.685 -80.755 -43.355 ;
        RECT -81.085 -45.045 -80.755 -44.715 ;
        RECT -81.085 -46.405 -80.755 -46.075 ;
        RECT -81.085 -47.765 -80.755 -47.435 ;
        RECT -81.085 -49.125 -80.755 -48.795 ;
        RECT -81.085 -50.485 -80.755 -50.155 ;
        RECT -81.085 -51.845 -80.755 -51.515 ;
        RECT -81.085 -53.205 -80.755 -52.875 ;
        RECT -81.085 -54.565 -80.755 -54.235 ;
        RECT -81.085 -55.925 -80.755 -55.595 ;
        RECT -81.085 -57.285 -80.755 -56.955 ;
        RECT -81.085 -58.645 -80.755 -58.315 ;
        RECT -81.085 -60.005 -80.755 -59.675 ;
        RECT -81.085 -61.365 -80.755 -61.035 ;
        RECT -81.085 -62.725 -80.755 -62.395 ;
        RECT -81.085 -64.085 -80.755 -63.755 ;
        RECT -81.085 -65.445 -80.755 -65.115 ;
        RECT -81.085 -66.805 -80.755 -66.475 ;
        RECT -81.085 -68.165 -80.755 -67.835 ;
        RECT -81.085 -69.525 -80.755 -69.195 ;
        RECT -81.085 -70.885 -80.755 -70.555 ;
        RECT -81.085 -72.245 -80.755 -71.915 ;
        RECT -81.085 -73.605 -80.755 -73.275 ;
        RECT -81.085 -74.965 -80.755 -74.635 ;
        RECT -81.085 -76.325 -80.755 -75.995 ;
        RECT -81.085 -77.685 -80.755 -77.355 ;
        RECT -81.085 -79.045 -80.755 -78.715 ;
        RECT -81.085 -80.405 -80.755 -80.075 ;
        RECT -81.085 -81.765 -80.755 -81.435 ;
        RECT -81.085 -83.125 -80.755 -82.795 ;
        RECT -81.085 -84.485 -80.755 -84.155 ;
        RECT -81.085 -85.845 -80.755 -85.515 ;
        RECT -81.085 -87.205 -80.755 -86.875 ;
        RECT -81.085 -88.565 -80.755 -88.235 ;
        RECT -81.085 -89.925 -80.755 -89.595 ;
        RECT -81.085 -91.285 -80.755 -90.955 ;
        RECT -81.085 -92.645 -80.755 -92.315 ;
        RECT -81.085 -94.005 -80.755 -93.675 ;
        RECT -81.085 -95.365 -80.755 -95.035 ;
        RECT -81.085 -96.725 -80.755 -96.395 ;
        RECT -81.085 -98.085 -80.755 -97.755 ;
        RECT -81.085 -99.445 -80.755 -99.115 ;
        RECT -81.085 -100.805 -80.755 -100.475 ;
        RECT -81.085 -102.165 -80.755 -101.835 ;
        RECT -81.085 -103.525 -80.755 -103.195 ;
        RECT -81.085 -104.885 -80.755 -104.555 ;
        RECT -81.085 -106.245 -80.755 -105.915 ;
        RECT -81.085 -107.605 -80.755 -107.275 ;
        RECT -81.085 -108.965 -80.755 -108.635 ;
        RECT -81.085 -110.325 -80.755 -109.995 ;
        RECT -81.085 -111.685 -80.755 -111.355 ;
        RECT -81.085 -113.045 -80.755 -112.715 ;
        RECT -81.085 -114.405 -80.755 -114.075 ;
        RECT -81.085 -115.765 -80.755 -115.435 ;
        RECT -81.085 -117.125 -80.755 -116.795 ;
        RECT -81.085 -118.485 -80.755 -118.155 ;
        RECT -81.085 -119.845 -80.755 -119.515 ;
        RECT -81.085 -121.205 -80.755 -120.875 ;
        RECT -81.085 -122.565 -80.755 -122.235 ;
        RECT -81.085 -123.925 -80.755 -123.595 ;
        RECT -81.085 -125.285 -80.755 -124.955 ;
        RECT -81.085 -126.645 -80.755 -126.315 ;
        RECT -81.085 -128.005 -80.755 -127.675 ;
        RECT -81.085 -129.365 -80.755 -129.035 ;
        RECT -81.085 -130.725 -80.755 -130.395 ;
        RECT -81.085 -132.085 -80.755 -131.755 ;
        RECT -81.085 -133.445 -80.755 -133.115 ;
        RECT -81.085 -134.805 -80.755 -134.475 ;
        RECT -81.085 -136.165 -80.755 -135.835 ;
        RECT -81.085 -137.525 -80.755 -137.195 ;
        RECT -81.085 -138.885 -80.755 -138.555 ;
        RECT -81.085 -140.245 -80.755 -139.915 ;
        RECT -81.085 -141.605 -80.755 -141.275 ;
        RECT -81.085 -142.965 -80.755 -142.635 ;
        RECT -81.085 -144.325 -80.755 -143.995 ;
        RECT -81.085 -145.685 -80.755 -145.355 ;
        RECT -81.085 -147.045 -80.755 -146.715 ;
        RECT -81.085 -148.405 -80.755 -148.075 ;
        RECT -81.085 -149.765 -80.755 -149.435 ;
        RECT -81.085 -151.125 -80.755 -150.795 ;
        RECT -81.085 -152.485 -80.755 -152.155 ;
        RECT -81.085 -153.845 -80.755 -153.515 ;
        RECT -81.085 -155.205 -80.755 -154.875 ;
        RECT -81.085 -156.565 -80.755 -156.235 ;
        RECT -81.085 -157.925 -80.755 -157.595 ;
        RECT -81.085 -159.285 -80.755 -158.955 ;
        RECT -81.085 -160.645 -80.755 -160.315 ;
        RECT -81.085 -162.005 -80.755 -161.675 ;
        RECT -81.085 -163.365 -80.755 -163.035 ;
        RECT -81.085 -164.725 -80.755 -164.395 ;
        RECT -81.085 -166.085 -80.755 -165.755 ;
        RECT -81.085 -167.445 -80.755 -167.115 ;
        RECT -81.085 -168.805 -80.755 -168.475 ;
        RECT -81.085 -170.165 -80.755 -169.835 ;
        RECT -81.085 -171.525 -80.755 -171.195 ;
        RECT -81.085 -172.885 -80.755 -172.555 ;
        RECT -81.085 -174.245 -80.755 -173.915 ;
        RECT -81.085 -175.605 -80.755 -175.275 ;
        RECT -81.085 -176.965 -80.755 -176.635 ;
        RECT -81.085 -178.325 -80.755 -177.995 ;
        RECT -81.085 -179.685 -80.755 -179.355 ;
        RECT -81.085 -181.93 -80.755 -180.8 ;
        RECT -81.08 -182.045 -80.76 242.565 ;
    END
    PORT
      LAYER met3 ;
        RECT -79.725 -119.845 -79.395 -119.515 ;
        RECT -79.725 -121.205 -79.395 -120.875 ;
        RECT -79.725 -122.565 -79.395 -122.235 ;
        RECT -79.725 -123.925 -79.395 -123.595 ;
        RECT -79.725 -125.285 -79.395 -124.955 ;
        RECT -79.725 -126.645 -79.395 -126.315 ;
        RECT -79.725 -128.005 -79.395 -127.675 ;
        RECT -79.725 -129.365 -79.395 -129.035 ;
        RECT -79.725 -130.725 -79.395 -130.395 ;
        RECT -79.725 -132.085 -79.395 -131.755 ;
        RECT -79.725 -133.445 -79.395 -133.115 ;
        RECT -79.725 -134.805 -79.395 -134.475 ;
        RECT -79.725 -136.165 -79.395 -135.835 ;
        RECT -79.725 -137.525 -79.395 -137.195 ;
        RECT -79.725 -138.885 -79.395 -138.555 ;
        RECT -79.725 -140.245 -79.395 -139.915 ;
        RECT -79.725 -141.605 -79.395 -141.275 ;
        RECT -79.725 -142.965 -79.395 -142.635 ;
        RECT -79.725 -144.325 -79.395 -143.995 ;
        RECT -79.725 -145.685 -79.395 -145.355 ;
        RECT -79.725 -147.045 -79.395 -146.715 ;
        RECT -79.725 -148.405 -79.395 -148.075 ;
        RECT -79.725 -149.765 -79.395 -149.435 ;
        RECT -79.725 -151.125 -79.395 -150.795 ;
        RECT -79.725 -152.485 -79.395 -152.155 ;
        RECT -79.725 -153.845 -79.395 -153.515 ;
        RECT -79.725 -155.205 -79.395 -154.875 ;
        RECT -79.725 -156.565 -79.395 -156.235 ;
        RECT -79.725 -157.925 -79.395 -157.595 ;
        RECT -79.725 -159.285 -79.395 -158.955 ;
        RECT -79.725 -160.645 -79.395 -160.315 ;
        RECT -79.725 -162.005 -79.395 -161.675 ;
        RECT -79.725 -163.365 -79.395 -163.035 ;
        RECT -79.725 -164.725 -79.395 -164.395 ;
        RECT -79.725 -166.085 -79.395 -165.755 ;
        RECT -79.725 -167.445 -79.395 -167.115 ;
        RECT -79.725 -168.805 -79.395 -168.475 ;
        RECT -79.725 -170.165 -79.395 -169.835 ;
        RECT -79.725 -171.525 -79.395 -171.195 ;
        RECT -79.725 -172.885 -79.395 -172.555 ;
        RECT -79.725 -174.245 -79.395 -173.915 ;
        RECT -79.725 -175.605 -79.395 -175.275 ;
        RECT -79.725 -176.965 -79.395 -176.635 ;
        RECT -79.725 -178.325 -79.395 -177.995 ;
        RECT -79.725 -179.685 -79.395 -179.355 ;
        RECT -79.725 -181.93 -79.395 -180.8 ;
        RECT -79.72 -182.045 -79.4 242.565 ;
        RECT -79.725 241.32 -79.395 242.45 ;
        RECT -79.725 239.195 -79.395 239.525 ;
        RECT -79.725 237.835 -79.395 238.165 ;
        RECT -79.725 236.475 -79.395 236.805 ;
        RECT -79.725 235.115 -79.395 235.445 ;
        RECT -79.725 233.755 -79.395 234.085 ;
        RECT -79.725 232.395 -79.395 232.725 ;
        RECT -79.725 231.035 -79.395 231.365 ;
        RECT -79.725 229.675 -79.395 230.005 ;
        RECT -79.725 228.315 -79.395 228.645 ;
        RECT -79.725 226.955 -79.395 227.285 ;
        RECT -79.725 225.595 -79.395 225.925 ;
        RECT -79.725 224.235 -79.395 224.565 ;
        RECT -79.725 222.875 -79.395 223.205 ;
        RECT -79.725 221.515 -79.395 221.845 ;
        RECT -79.725 220.155 -79.395 220.485 ;
        RECT -79.725 218.795 -79.395 219.125 ;
        RECT -79.725 217.435 -79.395 217.765 ;
        RECT -79.725 216.075 -79.395 216.405 ;
        RECT -79.725 214.715 -79.395 215.045 ;
        RECT -79.725 213.355 -79.395 213.685 ;
        RECT -79.725 211.995 -79.395 212.325 ;
        RECT -79.725 210.635 -79.395 210.965 ;
        RECT -79.725 209.275 -79.395 209.605 ;
        RECT -79.725 207.915 -79.395 208.245 ;
        RECT -79.725 206.555 -79.395 206.885 ;
        RECT -79.725 205.195 -79.395 205.525 ;
        RECT -79.725 203.835 -79.395 204.165 ;
        RECT -79.725 202.475 -79.395 202.805 ;
        RECT -79.725 201.115 -79.395 201.445 ;
        RECT -79.725 199.755 -79.395 200.085 ;
        RECT -79.725 198.395 -79.395 198.725 ;
        RECT -79.725 197.035 -79.395 197.365 ;
        RECT -79.725 195.675 -79.395 196.005 ;
        RECT -79.725 194.315 -79.395 194.645 ;
        RECT -79.725 192.955 -79.395 193.285 ;
        RECT -79.725 191.595 -79.395 191.925 ;
        RECT -79.725 190.235 -79.395 190.565 ;
        RECT -79.725 188.875 -79.395 189.205 ;
        RECT -79.725 187.515 -79.395 187.845 ;
        RECT -79.725 186.155 -79.395 186.485 ;
        RECT -79.725 184.795 -79.395 185.125 ;
        RECT -79.725 183.435 -79.395 183.765 ;
        RECT -79.725 182.075 -79.395 182.405 ;
        RECT -79.725 180.715 -79.395 181.045 ;
        RECT -79.725 179.355 -79.395 179.685 ;
        RECT -79.725 177.995 -79.395 178.325 ;
        RECT -79.725 176.635 -79.395 176.965 ;
        RECT -79.725 175.275 -79.395 175.605 ;
        RECT -79.725 173.915 -79.395 174.245 ;
        RECT -79.725 172.555 -79.395 172.885 ;
        RECT -79.725 171.195 -79.395 171.525 ;
        RECT -79.725 169.835 -79.395 170.165 ;
        RECT -79.725 168.475 -79.395 168.805 ;
        RECT -79.725 167.115 -79.395 167.445 ;
        RECT -79.725 165.755 -79.395 166.085 ;
        RECT -79.725 164.395 -79.395 164.725 ;
        RECT -79.725 163.035 -79.395 163.365 ;
        RECT -79.725 161.675 -79.395 162.005 ;
        RECT -79.725 160.315 -79.395 160.645 ;
        RECT -79.725 158.955 -79.395 159.285 ;
        RECT -79.725 157.595 -79.395 157.925 ;
        RECT -79.725 156.235 -79.395 156.565 ;
        RECT -79.725 154.875 -79.395 155.205 ;
        RECT -79.725 153.515 -79.395 153.845 ;
        RECT -79.725 152.155 -79.395 152.485 ;
        RECT -79.725 150.795 -79.395 151.125 ;
        RECT -79.725 149.435 -79.395 149.765 ;
        RECT -79.725 148.075 -79.395 148.405 ;
        RECT -79.725 146.715 -79.395 147.045 ;
        RECT -79.725 145.355 -79.395 145.685 ;
        RECT -79.725 143.995 -79.395 144.325 ;
        RECT -79.725 142.635 -79.395 142.965 ;
        RECT -79.725 141.275 -79.395 141.605 ;
        RECT -79.725 139.915 -79.395 140.245 ;
        RECT -79.725 138.555 -79.395 138.885 ;
        RECT -79.725 137.195 -79.395 137.525 ;
        RECT -79.725 135.835 -79.395 136.165 ;
        RECT -79.725 134.475 -79.395 134.805 ;
        RECT -79.725 133.115 -79.395 133.445 ;
        RECT -79.725 131.755 -79.395 132.085 ;
        RECT -79.725 130.395 -79.395 130.725 ;
        RECT -79.725 129.035 -79.395 129.365 ;
        RECT -79.725 127.675 -79.395 128.005 ;
        RECT -79.725 126.315 -79.395 126.645 ;
        RECT -79.725 124.955 -79.395 125.285 ;
        RECT -79.725 123.595 -79.395 123.925 ;
        RECT -79.725 122.235 -79.395 122.565 ;
        RECT -79.725 120.875 -79.395 121.205 ;
        RECT -79.725 119.515 -79.395 119.845 ;
        RECT -79.725 118.155 -79.395 118.485 ;
        RECT -79.725 116.795 -79.395 117.125 ;
        RECT -79.725 115.435 -79.395 115.765 ;
        RECT -79.725 114.075 -79.395 114.405 ;
        RECT -79.725 112.715 -79.395 113.045 ;
        RECT -79.725 111.355 -79.395 111.685 ;
        RECT -79.725 109.995 -79.395 110.325 ;
        RECT -79.725 108.635 -79.395 108.965 ;
        RECT -79.725 107.275 -79.395 107.605 ;
        RECT -79.725 105.915 -79.395 106.245 ;
        RECT -79.725 104.555 -79.395 104.885 ;
        RECT -79.725 103.195 -79.395 103.525 ;
        RECT -79.725 101.835 -79.395 102.165 ;
        RECT -79.725 100.475 -79.395 100.805 ;
        RECT -79.725 99.115 -79.395 99.445 ;
        RECT -79.725 97.755 -79.395 98.085 ;
        RECT -79.725 96.395 -79.395 96.725 ;
        RECT -79.725 95.035 -79.395 95.365 ;
        RECT -79.725 93.675 -79.395 94.005 ;
        RECT -79.725 92.315 -79.395 92.645 ;
        RECT -79.725 90.955 -79.395 91.285 ;
        RECT -79.725 89.595 -79.395 89.925 ;
        RECT -79.725 88.235 -79.395 88.565 ;
        RECT -79.725 86.875 -79.395 87.205 ;
        RECT -79.725 85.515 -79.395 85.845 ;
        RECT -79.725 84.155 -79.395 84.485 ;
        RECT -79.725 82.795 -79.395 83.125 ;
        RECT -79.725 81.435 -79.395 81.765 ;
        RECT -79.725 80.075 -79.395 80.405 ;
        RECT -79.725 78.715 -79.395 79.045 ;
        RECT -79.725 77.355 -79.395 77.685 ;
        RECT -79.725 75.995 -79.395 76.325 ;
        RECT -79.725 74.635 -79.395 74.965 ;
        RECT -79.725 73.275 -79.395 73.605 ;
        RECT -79.725 71.915 -79.395 72.245 ;
        RECT -79.725 70.555 -79.395 70.885 ;
        RECT -79.725 69.195 -79.395 69.525 ;
        RECT -79.725 67.835 -79.395 68.165 ;
        RECT -79.725 66.475 -79.395 66.805 ;
        RECT -79.725 65.115 -79.395 65.445 ;
        RECT -79.725 63.755 -79.395 64.085 ;
        RECT -79.725 62.395 -79.395 62.725 ;
        RECT -79.725 61.035 -79.395 61.365 ;
        RECT -79.725 59.675 -79.395 60.005 ;
        RECT -79.725 58.315 -79.395 58.645 ;
        RECT -79.725 56.955 -79.395 57.285 ;
        RECT -79.725 55.595 -79.395 55.925 ;
        RECT -79.725 54.235 -79.395 54.565 ;
        RECT -79.725 52.875 -79.395 53.205 ;
        RECT -79.725 51.515 -79.395 51.845 ;
        RECT -79.725 50.155 -79.395 50.485 ;
        RECT -79.725 48.795 -79.395 49.125 ;
        RECT -79.725 47.435 -79.395 47.765 ;
        RECT -79.725 46.075 -79.395 46.405 ;
        RECT -79.725 44.715 -79.395 45.045 ;
        RECT -79.725 43.355 -79.395 43.685 ;
        RECT -79.725 41.995 -79.395 42.325 ;
        RECT -79.725 40.635 -79.395 40.965 ;
        RECT -79.725 39.275 -79.395 39.605 ;
        RECT -79.725 37.915 -79.395 38.245 ;
        RECT -79.725 36.555 -79.395 36.885 ;
        RECT -79.725 35.195 -79.395 35.525 ;
        RECT -79.725 33.835 -79.395 34.165 ;
        RECT -79.725 32.475 -79.395 32.805 ;
        RECT -79.725 31.115 -79.395 31.445 ;
        RECT -79.725 29.755 -79.395 30.085 ;
        RECT -79.725 28.395 -79.395 28.725 ;
        RECT -79.725 27.035 -79.395 27.365 ;
        RECT -79.725 25.675 -79.395 26.005 ;
        RECT -79.725 24.315 -79.395 24.645 ;
        RECT -79.725 22.955 -79.395 23.285 ;
        RECT -79.725 21.595 -79.395 21.925 ;
        RECT -79.725 20.235 -79.395 20.565 ;
        RECT -79.725 18.875 -79.395 19.205 ;
        RECT -79.725 17.515 -79.395 17.845 ;
        RECT -79.725 16.155 -79.395 16.485 ;
        RECT -79.725 14.795 -79.395 15.125 ;
        RECT -79.725 13.435 -79.395 13.765 ;
        RECT -79.725 12.075 -79.395 12.405 ;
        RECT -79.725 10.715 -79.395 11.045 ;
        RECT -79.725 9.355 -79.395 9.685 ;
        RECT -79.725 7.995 -79.395 8.325 ;
        RECT -79.725 6.635 -79.395 6.965 ;
        RECT -79.725 5.275 -79.395 5.605 ;
        RECT -79.725 3.915 -79.395 4.245 ;
        RECT -79.725 2.555 -79.395 2.885 ;
        RECT -79.725 1.195 -79.395 1.525 ;
        RECT -79.725 -0.165 -79.395 0.165 ;
        RECT -79.725 -1.525 -79.395 -1.195 ;
        RECT -79.725 -2.885 -79.395 -2.555 ;
        RECT -79.725 -4.245 -79.395 -3.915 ;
        RECT -79.725 -5.605 -79.395 -5.275 ;
        RECT -79.725 -6.965 -79.395 -6.635 ;
        RECT -79.725 -8.325 -79.395 -7.995 ;
        RECT -79.725 -9.685 -79.395 -9.355 ;
        RECT -79.725 -11.045 -79.395 -10.715 ;
        RECT -79.725 -12.405 -79.395 -12.075 ;
        RECT -79.725 -13.765 -79.395 -13.435 ;
        RECT -79.725 -15.125 -79.395 -14.795 ;
        RECT -79.725 -16.485 -79.395 -16.155 ;
        RECT -79.725 -17.845 -79.395 -17.515 ;
        RECT -79.725 -19.205 -79.395 -18.875 ;
        RECT -79.725 -20.565 -79.395 -20.235 ;
        RECT -79.725 -21.925 -79.395 -21.595 ;
        RECT -79.725 -23.285 -79.395 -22.955 ;
        RECT -79.725 -24.645 -79.395 -24.315 ;
        RECT -79.725 -26.005 -79.395 -25.675 ;
        RECT -79.725 -27.365 -79.395 -27.035 ;
        RECT -79.725 -28.725 -79.395 -28.395 ;
        RECT -79.725 -30.085 -79.395 -29.755 ;
        RECT -79.725 -31.445 -79.395 -31.115 ;
        RECT -79.725 -32.805 -79.395 -32.475 ;
        RECT -79.725 -34.165 -79.395 -33.835 ;
        RECT -79.725 -35.525 -79.395 -35.195 ;
        RECT -79.725 -36.885 -79.395 -36.555 ;
        RECT -79.725 -38.245 -79.395 -37.915 ;
        RECT -79.725 -39.605 -79.395 -39.275 ;
        RECT -79.725 -40.965 -79.395 -40.635 ;
        RECT -79.725 -42.325 -79.395 -41.995 ;
        RECT -79.725 -43.685 -79.395 -43.355 ;
        RECT -79.725 -45.045 -79.395 -44.715 ;
        RECT -79.725 -46.405 -79.395 -46.075 ;
        RECT -79.725 -47.765 -79.395 -47.435 ;
        RECT -79.725 -49.125 -79.395 -48.795 ;
        RECT -79.725 -50.485 -79.395 -50.155 ;
        RECT -79.725 -51.845 -79.395 -51.515 ;
        RECT -79.725 -53.205 -79.395 -52.875 ;
        RECT -79.725 -54.565 -79.395 -54.235 ;
        RECT -79.725 -55.925 -79.395 -55.595 ;
        RECT -79.725 -57.285 -79.395 -56.955 ;
        RECT -79.725 -58.645 -79.395 -58.315 ;
        RECT -79.725 -60.005 -79.395 -59.675 ;
        RECT -79.725 -61.365 -79.395 -61.035 ;
        RECT -79.725 -62.725 -79.395 -62.395 ;
        RECT -79.725 -64.085 -79.395 -63.755 ;
        RECT -79.725 -65.445 -79.395 -65.115 ;
        RECT -79.725 -66.805 -79.395 -66.475 ;
        RECT -79.725 -68.165 -79.395 -67.835 ;
        RECT -79.725 -69.525 -79.395 -69.195 ;
        RECT -79.725 -70.885 -79.395 -70.555 ;
        RECT -79.725 -72.245 -79.395 -71.915 ;
        RECT -79.725 -73.605 -79.395 -73.275 ;
        RECT -79.725 -74.965 -79.395 -74.635 ;
        RECT -79.725 -76.325 -79.395 -75.995 ;
        RECT -79.725 -77.685 -79.395 -77.355 ;
        RECT -79.725 -79.045 -79.395 -78.715 ;
        RECT -79.725 -80.405 -79.395 -80.075 ;
        RECT -79.725 -81.765 -79.395 -81.435 ;
        RECT -79.725 -83.125 -79.395 -82.795 ;
        RECT -79.725 -84.485 -79.395 -84.155 ;
        RECT -79.725 -85.845 -79.395 -85.515 ;
        RECT -79.725 -87.205 -79.395 -86.875 ;
        RECT -79.725 -88.565 -79.395 -88.235 ;
        RECT -79.725 -89.925 -79.395 -89.595 ;
        RECT -79.725 -91.285 -79.395 -90.955 ;
        RECT -79.725 -92.645 -79.395 -92.315 ;
        RECT -79.725 -94.005 -79.395 -93.675 ;
        RECT -79.725 -95.365 -79.395 -95.035 ;
        RECT -79.725 -96.725 -79.395 -96.395 ;
        RECT -79.725 -98.085 -79.395 -97.755 ;
        RECT -79.725 -99.445 -79.395 -99.115 ;
        RECT -79.725 -100.805 -79.395 -100.475 ;
        RECT -79.725 -102.165 -79.395 -101.835 ;
        RECT -79.725 -103.525 -79.395 -103.195 ;
        RECT -79.725 -104.885 -79.395 -104.555 ;
        RECT -79.725 -106.245 -79.395 -105.915 ;
        RECT -79.725 -107.605 -79.395 -107.275 ;
        RECT -79.725 -108.965 -79.395 -108.635 ;
        RECT -79.725 -110.325 -79.395 -109.995 ;
        RECT -79.725 -111.685 -79.395 -111.355 ;
        RECT -79.725 -113.045 -79.395 -112.715 ;
        RECT -79.725 -114.405 -79.395 -114.075 ;
        RECT -79.725 -115.765 -79.395 -115.435 ;
        RECT -79.725 -117.125 -79.395 -116.795 ;
        RECT -79.725 -118.485 -79.395 -118.155 ;
    END
  END vss
  PIN addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -21.24 -184.925 -20.92 -184.605 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -28.04 -184.925 -27.72 -184.605 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -34.16 -184.925 -33.84 -184.605 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -40.28 -184.925 -39.96 -184.605 ;
    END
  END addr[3]
  PIN addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -46.4 -184.925 -46.08 -184.605 ;
    END
  END addr[4]
  PIN addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -52.52 -184.925 -52.2 -184.605 ;
    END
  END addr[5]
  PIN addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -58.64 -184.925 -58.32 -184.605 ;
    END
  END addr[6]
  PIN addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -64.76 -184.925 -64.44 -184.605 ;
    END
  END addr[7]
  PIN addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -70.88 -184.925 -70.56 -184.605 ;
    END
  END addr[8]
  PIN addr[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -77.68 -184.925 -77.36 -184.605 ;
    END
  END addr[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -9.68 -184.925 -9.36 -184.605 ;
    END
  END clk
  PIN din[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 5.6 -184.925 6 -184.525 ;
    END
  END din[0]
  PIN din[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 114.6 -184.925 115 -184.525 ;
    END
  END din[10]
  PIN din[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 125.5 -184.925 125.9 -184.525 ;
    END
  END din[11]
  PIN din[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 136.4 -184.925 136.8 -184.525 ;
    END
  END din[12]
  PIN din[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 147.3 -184.925 147.7 -184.525 ;
    END
  END din[13]
  PIN din[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 158.2 -184.925 158.6 -184.525 ;
    END
  END din[14]
  PIN din[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 169.1 -184.925 169.5 -184.525 ;
    END
  END din[15]
  PIN din[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 180 -184.925 180.4 -184.525 ;
    END
  END din[16]
  PIN din[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 190.9 -184.925 191.3 -184.525 ;
    END
  END din[17]
  PIN din[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 201.8 -184.925 202.2 -184.525 ;
    END
  END din[18]
  PIN din[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 212.7 -184.925 213.1 -184.525 ;
    END
  END din[19]
  PIN din[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 16.5 -184.925 16.9 -184.525 ;
    END
  END din[1]
  PIN din[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 223.6 -184.925 224 -184.525 ;
    END
  END din[20]
  PIN din[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 234.5 -184.925 234.9 -184.525 ;
    END
  END din[21]
  PIN din[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 245.4 -184.925 245.8 -184.525 ;
    END
  END din[22]
  PIN din[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 256.3 -184.925 256.7 -184.525 ;
    END
  END din[23]
  PIN din[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 267.2 -184.925 267.6 -184.525 ;
    END
  END din[24]
  PIN din[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 278.1 -184.925 278.5 -184.525 ;
    END
  END din[25]
  PIN din[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 289 -184.925 289.4 -184.525 ;
    END
  END din[26]
  PIN din[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 299.9 -184.925 300.3 -184.525 ;
    END
  END din[27]
  PIN din[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 310.8 -184.925 311.2 -184.525 ;
    END
  END din[28]
  PIN din[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 321.7 -184.925 322.1 -184.525 ;
    END
  END din[29]
  PIN din[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 27.4 -184.925 27.8 -184.525 ;
    END
  END din[2]
  PIN din[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 332.6 -184.925 333 -184.525 ;
    END
  END din[30]
  PIN din[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 343.5 -184.925 343.9 -184.525 ;
    END
  END din[31]
  PIN din[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 38.3 -184.925 38.7 -184.525 ;
    END
  END din[3]
  PIN din[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 49.2 -184.925 49.6 -184.525 ;
    END
  END din[4]
  PIN din[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 60.1 -184.925 60.5 -184.525 ;
    END
  END din[5]
  PIN din[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 71 -184.925 71.4 -184.525 ;
    END
  END din[6]
  PIN din[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 81.9 -184.925 82.3 -184.525 ;
    END
  END din[7]
  PIN din[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 92.8 -184.925 93.2 -184.525 ;
    END
  END din[8]
  PIN din[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 103.7 -184.925 104.1 -184.525 ;
    END
  END din[9]
  PIN dout[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 4 -184.925 4.4 -184.525 ;
    END
  END dout[0]
  PIN dout[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 113 -184.925 113.4 -184.525 ;
    END
  END dout[10]
  PIN dout[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 123.9 -184.925 124.3 -184.525 ;
    END
  END dout[11]
  PIN dout[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 134.8 -184.925 135.2 -184.525 ;
    END
  END dout[12]
  PIN dout[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 145.7 -184.925 146.1 -184.525 ;
    END
  END dout[13]
  PIN dout[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 156.6 -184.925 157 -184.525 ;
    END
  END dout[14]
  PIN dout[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 167.5 -184.925 167.9 -184.525 ;
    END
  END dout[15]
  PIN dout[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 178.4 -184.925 178.8 -184.525 ;
    END
  END dout[16]
  PIN dout[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 189.3 -184.925 189.7 -184.525 ;
    END
  END dout[17]
  PIN dout[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 200.2 -184.925 200.6 -184.525 ;
    END
  END dout[18]
  PIN dout[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 211.1 -184.925 211.5 -184.525 ;
    END
  END dout[19]
  PIN dout[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 14.9 -184.925 15.3 -184.525 ;
    END
  END dout[1]
  PIN dout[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 222 -184.925 222.4 -184.525 ;
    END
  END dout[20]
  PIN dout[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 232.9 -184.925 233.3 -184.525 ;
    END
  END dout[21]
  PIN dout[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 243.8 -184.925 244.2 -184.525 ;
    END
  END dout[22]
  PIN dout[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 254.7 -184.925 255.1 -184.525 ;
    END
  END dout[23]
  PIN dout[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 265.6 -184.925 266 -184.525 ;
    END
  END dout[24]
  PIN dout[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 276.5 -184.925 276.9 -184.525 ;
    END
  END dout[25]
  PIN dout[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 287.4 -184.925 287.8 -184.525 ;
    END
  END dout[26]
  PIN dout[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 298.3 -184.925 298.7 -184.525 ;
    END
  END dout[27]
  PIN dout[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 309.2 -184.925 309.6 -184.525 ;
    END
  END dout[28]
  PIN dout[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 320.1 -184.925 320.5 -184.525 ;
    END
  END dout[29]
  PIN dout[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 25.8 -184.925 26.2 -184.525 ;
    END
  END dout[2]
  PIN dout[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 331 -184.925 331.4 -184.525 ;
    END
  END dout[30]
  PIN dout[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 341.9 -184.925 342.3 -184.525 ;
    END
  END dout[31]
  PIN dout[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 36.7 -184.925 37.1 -184.525 ;
    END
  END dout[3]
  PIN dout[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 47.6 -184.925 48 -184.525 ;
    END
  END dout[4]
  PIN dout[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 58.5 -184.925 58.9 -184.525 ;
    END
  END dout[5]
  PIN dout[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 69.4 -184.925 69.8 -184.525 ;
    END
  END dout[6]
  PIN dout[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 80.3 -184.925 80.7 -184.525 ;
    END
  END dout[7]
  PIN dout[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 91.2 -184.925 91.6 -184.525 ;
    END
  END dout[8]
  PIN dout[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 102.1 -184.925 102.5 -184.525 ;
    END
  END dout[9]
  PIN sae_int
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -9 -184.925 -8.68 -184.605 ;
    END
  END sae_int
  PIN sae_muxed
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -8.32 -184.925 -8 -184.605 ;
    END
  END sae_muxed
  PIN we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -15.12 -184.925 -14.8 -184.605 ;
    END
  END we
  PIN wmask
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 6.4 -184.925 6.8 -184.525 ;
    END
  END wmask
  OBS
    LAYER met1 SPACING 0.14 ;
      RECT -86.345 -184.925 366.505 245.445 ;
    LAYER met2 SPACING 0.14 ;
      RECT -86.345 -184.925 366.505 245.445 ;
    LAYER met3 SPACING 0.3 ;
      RECT 0.515 -40.285 0.845 -39.955 ;
      RECT 0.52 -66.805 0.84 -39.955 ;
      RECT 0.515 -66.805 0.845 -66.475 ;
      RECT -0.165 -38.245 0.165 -37.915 ;
      RECT -0.16 -49.805 0.16 -37.915 ;
      RECT -0.165 -49.805 0.165 -49.475 ;
      RECT -0.845 -36.885 -0.515 -36.555 ;
      RECT -0.84 -50.485 -0.52 -36.555 ;
      RECT -0.845 -50.485 -0.515 -50.155 ;
      RECT -7.645 -19.205 -7.315 -18.875 ;
      RECT -7.64 -105.565 -7.32 -18.875 ;
      RECT -7.645 -105.565 -7.315 -105.235 ;
      RECT -8.325 -166.765 -7.995 -166.435 ;
      RECT -8.32 -184.115 -8 -166.435 ;
      RECT -8.325 -21.925 -7.995 -21.595 ;
      RECT -8.32 -106.245 -8 -21.595 ;
      RECT -8.325 -106.245 -7.995 -105.915 ;
      RECT -9.005 -167.445 -8.675 -167.115 ;
      RECT -9 -184.115 -8.68 -167.115 ;
      RECT -9.005 -23.285 -8.675 -22.955 ;
      RECT -9 -108.965 -8.68 -22.955 ;
      RECT -9.005 -108.965 -8.675 -108.635 ;
      RECT -9.685 -168.125 -9.355 -167.795 ;
      RECT -9.68 -184.115 -9.36 -167.795 ;
      RECT -10.365 -168.805 -10.035 -168.475 ;
      RECT -10.36 -173.565 -10.04 -168.475 ;
      RECT -10.365 -173.565 -10.035 -173.235 ;
      RECT -11.725 -18.525 -11.395 -18.195 ;
      RECT -11.72 -104.885 -11.4 -18.195 ;
      RECT -11.725 -104.885 -11.395 -104.555 ;
      RECT -12.405 -15.805 -12.075 -15.475 ;
      RECT -12.4 -26.005 -12.08 -15.475 ;
      RECT -12.405 -26.005 -12.075 -25.675 ;
      RECT -14.445 -168.125 -14.115 -167.795 ;
      RECT -14.44 -172.885 -14.12 -167.795 ;
      RECT -14.445 -172.885 -14.115 -172.555 ;
      RECT -14.445 -89.925 -14.115 -89.595 ;
      RECT -14.44 -159.285 -14.12 -89.595 ;
      RECT -14.445 -159.285 -14.115 -158.955 ;
      RECT -15.12 -184.115 -14.8 -173.24 ;
      RECT -15.125 -173.7 -14.795 -173.37 ;
      RECT -15.125 -20.565 -14.795 -20.235 ;
      RECT -15.12 -104.885 -14.8 -20.235 ;
      RECT -15.125 -104.885 -14.795 -104.555 ;
      RECT -15.805 -21.245 -15.475 -20.915 ;
      RECT -15.8 -105.565 -15.48 -20.915 ;
      RECT -15.805 -105.565 -15.475 -105.235 ;
      RECT -16.485 -43.685 -16.155 -43.355 ;
      RECT -16.48 -122.565 -16.16 -43.355 ;
      RECT -16.485 -122.565 -16.155 -122.235 ;
      RECT -16.485 -13.765 -16.155 -13.435 ;
      RECT -16.48 -26.005 -16.16 -13.435 ;
      RECT -16.485 -26.005 -16.155 -25.675 ;
      RECT -17.165 -116.445 -16.835 -116.115 ;
      RECT -17.16 -174.925 -16.84 -116.115 ;
      RECT -17.165 -174.925 -16.835 -174.595 ;
      RECT -17.165 -13.085 -16.835 -12.755 ;
      RECT -17.16 -26.005 -16.84 -12.755 ;
      RECT -17.165 -26.005 -16.835 -25.675 ;
      RECT -17.845 -34.845 -17.515 -34.515 ;
      RECT -17.84 -120.525 -17.52 -34.515 ;
      RECT -17.845 -120.525 -17.515 -120.195 ;
      RECT -17.845 -12.405 -17.515 -12.075 ;
      RECT -17.84 -26.005 -17.52 -12.075 ;
      RECT -17.845 -26.005 -17.515 -25.675 ;
      RECT -18.525 -110.13 -18.195 -109.8 ;
      RECT -18.52 -113.725 -18.2 -109.8 ;
      RECT -18.525 -113.725 -18.195 -113.395 ;
      RECT -18.525 -22.49 -18.195 -22.16 ;
      RECT -18.52 -26.005 -18.2 -22.16 ;
      RECT -18.525 -26.005 -18.195 -25.675 ;
      RECT -19.205 -115.765 -18.875 -115.435 ;
      RECT -19.2 -172.885 -18.88 -115.435 ;
      RECT -19.205 -172.885 -18.875 -172.555 ;
      RECT -19.205 -110.61 -18.875 -110.28 ;
      RECT -19.2 -114.405 -18.88 -110.28 ;
      RECT -19.205 -114.405 -18.875 -114.075 ;
      RECT -19.205 -22.97 -18.875 -22.64 ;
      RECT -19.2 -26.685 -18.88 -22.64 ;
      RECT -19.205 -26.685 -18.875 -26.355 ;
      RECT -19.885 -168.125 -19.555 -167.795 ;
      RECT -19.88 -172.885 -19.56 -167.795 ;
      RECT -19.885 -172.885 -19.555 -172.555 ;
      RECT -19.885 -111.09 -19.555 -110.76 ;
      RECT -19.88 -115.085 -19.56 -110.76 ;
      RECT -19.885 -115.085 -19.555 -114.755 ;
      RECT -19.885 -23.45 -19.555 -23.12 ;
      RECT -19.88 -27.365 -19.56 -23.12 ;
      RECT -19.885 -27.365 -19.555 -27.035 ;
      RECT -20.565 -111.57 -20.235 -111.24 ;
      RECT -20.56 -174.925 -20.24 -111.24 ;
      RECT -20.565 -174.925 -20.235 -174.595 ;
      RECT -20.565 -23.93 -20.235 -23.6 ;
      RECT -20.56 -28.045 -20.24 -23.6 ;
      RECT -20.565 -28.045 -20.235 -27.715 ;
      RECT -21.24 -184.115 -20.92 -173.24 ;
      RECT -21.245 -173.7 -20.915 -173.37 ;
      RECT -21.245 -112.05 -20.915 -111.72 ;
      RECT -21.24 -115.765 -20.92 -111.72 ;
      RECT -21.245 -115.765 -20.915 -115.435 ;
      RECT -21.245 -24.41 -20.915 -24.08 ;
      RECT -21.24 -28.725 -20.92 -24.08 ;
      RECT -21.245 -28.725 -20.915 -28.395 ;
      RECT -21.925 -112.53 -21.595 -112.2 ;
      RECT -21.92 -116.445 -21.6 -112.2 ;
      RECT -21.925 -116.445 -21.595 -116.115 ;
      RECT -21.925 -24.89 -21.595 -24.56 ;
      RECT -21.92 -29.405 -21.6 -24.56 ;
      RECT -21.925 -29.405 -21.595 -29.075 ;
      RECT -23.285 -115.085 -22.955 -114.755 ;
      RECT -23.28 -172.885 -22.96 -114.755 ;
      RECT -23.285 -172.885 -22.955 -172.555 ;
      RECT -24.645 -114.405 -24.315 -114.075 ;
      RECT -24.64 -174.925 -24.32 -114.075 ;
      RECT -24.645 -174.925 -24.315 -174.595 ;
      RECT -26.685 -168.125 -26.355 -167.795 ;
      RECT -26.68 -172.885 -26.36 -167.795 ;
      RECT -26.685 -172.885 -26.355 -172.555 ;
      RECT -27.365 -11.725 -27.035 -11.395 ;
      RECT -27.36 -30.085 -27.04 -11.395 ;
      RECT -27.365 -30.085 -27.035 -29.755 ;
      RECT -28.04 -184.115 -27.72 -173.24 ;
      RECT -28.045 -173.7 -27.715 -173.37 ;
      RECT -28.725 -64.33 -28.395 -64 ;
      RECT -28.72 -68.845 -28.4 -64 ;
      RECT -28.725 -68.845 -28.395 -68.515 ;
      RECT -29.405 -113.725 -29.075 -113.395 ;
      RECT -29.4 -172.885 -29.08 -113.395 ;
      RECT -29.405 -172.885 -29.075 -172.555 ;
      RECT -29.405 -64.81 -29.075 -64.48 ;
      RECT -29.4 -68.165 -29.08 -64.48 ;
      RECT -29.405 -68.165 -29.075 -67.835 ;
      RECT -30.085 -65.29 -29.755 -64.96 ;
      RECT -30.08 -66.805 -29.76 -64.96 ;
      RECT -30.085 -66.805 -29.755 -66.475 ;
      RECT -30.765 -88.565 -30.435 -88.235 ;
      RECT -30.76 -121.205 -30.44 -88.235 ;
      RECT -30.765 -121.205 -30.435 -120.875 ;
      RECT -30.765 -65.77 -30.435 -65.44 ;
      RECT -30.76 -67.485 -30.44 -65.44 ;
      RECT -30.765 -67.485 -30.435 -67.155 ;
      RECT -32.805 -168.125 -32.475 -167.795 ;
      RECT -32.8 -172.885 -32.48 -167.795 ;
      RECT -32.805 -172.885 -32.475 -172.555 ;
      RECT -34.16 -184.115 -33.84 -173.24 ;
      RECT -34.165 -173.7 -33.835 -173.37 ;
      RECT -35.525 -114.405 -35.195 -114.075 ;
      RECT -35.52 -174.925 -35.2 -114.075 ;
      RECT -35.525 -174.925 -35.195 -174.595 ;
      RECT -38.245 -113.725 -37.915 -113.395 ;
      RECT -38.24 -172.885 -37.92 -113.395 ;
      RECT -38.245 -172.885 -37.915 -172.555 ;
      RECT -38.925 -168.125 -38.595 -167.795 ;
      RECT -38.92 -172.885 -38.6 -167.795 ;
      RECT -38.925 -172.885 -38.595 -172.555 ;
      RECT -40.28 -184.115 -39.96 -173.24 ;
      RECT -40.285 -173.7 -39.955 -173.37 ;
      RECT -43.005 -64.33 -42.675 -64 ;
      RECT -43 -66.805 -42.68 -64 ;
      RECT -43.005 -66.805 -42.675 -66.475 ;
      RECT -43.685 -113.725 -43.355 -113.395 ;
      RECT -43.68 -174.925 -43.36 -113.395 ;
      RECT -43.685 -174.925 -43.355 -174.595 ;
      RECT -43.685 -64.81 -43.355 -64.48 ;
      RECT -43.68 -67.485 -43.36 -64.48 ;
      RECT -43.685 -67.485 -43.355 -67.155 ;
      RECT -44.365 -113.725 -44.035 -113.395 ;
      RECT -44.36 -172.885 -44.04 -113.395 ;
      RECT -44.365 -172.885 -44.035 -172.555 ;
      RECT -44.365 -65.29 -44.035 -64.96 ;
      RECT -44.36 -68.165 -44.04 -64.96 ;
      RECT -44.365 -68.165 -44.035 -67.835 ;
      RECT -45.045 -168.125 -44.715 -167.795 ;
      RECT -45.04 -172.885 -44.72 -167.795 ;
      RECT -45.045 -172.885 -44.715 -172.555 ;
      RECT -45.045 -65.77 -44.715 -65.44 ;
      RECT -45.04 -68.845 -44.72 -65.44 ;
      RECT -45.045 -68.845 -44.715 -68.515 ;
      RECT -46.4 -184.115 -46.08 -173.24 ;
      RECT -46.405 -173.7 -46.075 -173.37 ;
      RECT -46.405 -2.205 -46.075 -1.875 ;
      RECT -46.4 -30.085 -46.08 -1.875 ;
      RECT -46.405 -30.085 -46.075 -29.755 ;
      RECT -47.085 -2.205 -46.755 -1.875 ;
      RECT -47.08 -30.765 -46.76 -1.875 ;
      RECT -47.085 -30.765 -46.755 -30.435 ;
      RECT -47.765 -113.725 -47.435 -113.395 ;
      RECT -47.76 -172.885 -47.44 -113.395 ;
      RECT -47.765 -172.885 -47.435 -172.555 ;
      RECT -48.445 -114.405 -48.115 -114.075 ;
      RECT -48.44 -174.925 -48.12 -114.075 ;
      RECT -48.445 -174.925 -48.115 -174.595 ;
      RECT -51.165 -168.125 -50.835 -167.795 ;
      RECT -51.16 -172.885 -50.84 -167.795 ;
      RECT -51.165 -172.885 -50.835 -172.555 ;
      RECT -52.52 -184.115 -52.2 -173.24 ;
      RECT -52.525 -173.7 -52.195 -173.37 ;
      RECT -53.48 116.48 -52.2 117.12 ;
      RECT -52.52 -119.845 -52.2 117.12 ;
      RECT -52.525 -119.845 -52.195 -119.515 ;
      RECT -53.885 -113.725 -53.555 -113.395 ;
      RECT -53.88 -172.885 -53.56 -113.395 ;
      RECT -53.885 -172.885 -53.555 -172.555 ;
      RECT -54.565 -114.405 -54.235 -114.075 ;
      RECT -54.56 -174.925 -54.24 -114.075 ;
      RECT -54.565 -174.925 -54.235 -174.595 ;
      RECT -57.285 -168.125 -56.955 -167.795 ;
      RECT -57.28 -172.885 -56.96 -167.795 ;
      RECT -57.285 -172.885 -56.955 -172.555 ;
      RECT -58.64 -184.115 -58.32 -173.24 ;
      RECT -58.645 -173.7 -58.315 -173.37 ;
      RECT -58.645 -113.725 -58.315 -113.395 ;
      RECT -58.64 -172.885 -58.32 -113.395 ;
      RECT -58.645 -172.885 -58.315 -172.555 ;
      RECT -59.325 86.875 -58.995 87.205 ;
      RECT -59.32 -1.525 -59 87.205 ;
      RECT -59.325 -1.525 -58.995 -1.195 ;
      RECT -60.005 86.195 -59.675 86.525 ;
      RECT -60 -122.565 -59.68 86.525 ;
      RECT -60.005 -122.565 -59.675 -122.235 ;
      RECT -60.685 -114.405 -60.355 -114.075 ;
      RECT -60.68 -174.925 -60.36 -114.075 ;
      RECT -60.685 -174.925 -60.355 -174.595 ;
      RECT -62.725 -113.725 -62.395 -113.395 ;
      RECT -62.72 -174.925 -62.4 -113.395 ;
      RECT -62.725 -174.925 -62.395 -174.595 ;
      RECT -64.085 -168.125 -63.755 -167.795 ;
      RECT -64.08 -172.885 -63.76 -167.795 ;
      RECT -64.085 -172.885 -63.755 -172.555 ;
      RECT -64.76 -184.115 -64.44 -173.24 ;
      RECT -64.765 -173.7 -64.435 -173.37 ;
      RECT -64.765 -113.725 -64.435 -113.395 ;
      RECT -64.76 -172.885 -64.44 -113.395 ;
      RECT -64.765 -172.885 -64.435 -172.555 ;
      RECT -68.165 -114.405 -67.835 -114.075 ;
      RECT -68.16 -174.925 -67.84 -114.075 ;
      RECT -68.165 -174.925 -67.835 -174.595 ;
      RECT -70.88 -184.115 -70.56 -173.24 ;
      RECT -70.885 -173.7 -70.555 -173.37 ;
      RECT -71.565 -172.205 -71.235 -171.875 ;
      RECT -71.56 -172.885 -71.24 -171.875 ;
      RECT -71.565 -172.885 -71.235 -172.555 ;
      RECT -71.565 -113.045 -71.235 -112.715 ;
      RECT -71.56 -121.885 -71.24 -112.715 ;
      RECT -71.565 -121.885 -71.235 -121.555 ;
      RECT -72.925 -113.725 -72.595 -113.395 ;
      RECT -72.92 -172.885 -72.6 -113.395 ;
      RECT -72.925 -172.885 -72.595 -172.555 ;
      RECT -73.605 -168.125 -73.275 -167.795 ;
      RECT -73.6 -172.885 -73.28 -167.795 ;
      RECT -73.605 -172.205 -73.275 -171.875 ;
      RECT -73.605 -172.885 -73.275 -172.555 ;
      RECT -77.68 -184.115 -77.36 -173.24 ;
      RECT -77.685 -173.7 -77.355 -173.37 ;
      RECT 345.1 -84.215 345.5 -22.12 ;
      RECT 344.3 -83.355 344.7 -22.12 ;
      RECT 343.5 -184.035 343.9 -83.445 ;
      RECT 342.7 -67.5 343.1 -52.905 ;
      RECT 342.7 -49.08 343.1 -15.74 ;
      RECT 341.9 -184.035 342.3 -77.605 ;
      RECT 341.9 -68 342.3 -53.36 ;
      RECT 341.9 -49.51 342.3 -12.47 ;
      RECT 334.2 -84.215 334.6 -22.12 ;
      RECT 333.4 -83.355 333.8 -22.12 ;
      RECT 332.6 -184.035 333 -83.445 ;
      RECT 331.8 -67.5 332.2 -52.905 ;
      RECT 331.8 -49.08 332.2 -15.74 ;
      RECT 331 -184.035 331.4 -77.605 ;
      RECT 331 -68 331.4 -53.36 ;
      RECT 331 -49.51 331.4 -12.47 ;
      RECT 323.3 -84.215 323.7 -22.12 ;
      RECT 322.5 -83.355 322.9 -22.12 ;
      RECT 321.7 -184.035 322.1 -83.445 ;
      RECT 320.9 -67.5 321.3 -52.905 ;
      RECT 320.9 -49.08 321.3 -15.74 ;
      RECT 320.1 -184.035 320.5 -77.605 ;
      RECT 320.1 -68 320.5 -53.36 ;
      RECT 320.1 -49.51 320.5 -12.47 ;
      RECT 312.4 -84.215 312.8 -22.12 ;
      RECT 311.6 -83.355 312 -22.12 ;
      RECT 310.8 -184.035 311.2 -83.445 ;
      RECT 310 -67.5 310.4 -52.905 ;
      RECT 310 -49.08 310.4 -15.74 ;
      RECT 309.2 -184.035 309.6 -77.605 ;
      RECT 309.2 -68 309.6 -53.36 ;
      RECT 309.2 -49.51 309.6 -12.47 ;
      RECT 301.5 -84.215 301.9 -22.12 ;
      RECT 300.7 -83.355 301.1 -22.12 ;
      RECT 299.9 -184.035 300.3 -83.445 ;
      RECT 299.1 -67.5 299.5 -52.905 ;
      RECT 299.1 -49.08 299.5 -15.74 ;
      RECT 298.3 -184.035 298.7 -77.605 ;
      RECT 298.3 -68 298.7 -53.36 ;
      RECT 298.3 -49.51 298.7 -12.47 ;
      RECT 290.6 -84.215 291 -22.12 ;
      RECT 289.8 -83.355 290.2 -22.12 ;
      RECT 289 -184.035 289.4 -83.445 ;
      RECT 288.2 -67.5 288.6 -52.905 ;
      RECT 288.2 -49.08 288.6 -15.74 ;
      RECT 287.4 -184.035 287.8 -77.605 ;
      RECT 287.4 -68 287.8 -53.36 ;
      RECT 287.4 -49.51 287.8 -12.47 ;
      RECT 279.7 -84.215 280.1 -22.12 ;
      RECT 278.9 -83.355 279.3 -22.12 ;
      RECT 278.1 -184.035 278.5 -83.445 ;
      RECT 277.3 -67.5 277.7 -52.905 ;
      RECT 277.3 -49.08 277.7 -15.74 ;
      RECT 276.5 -184.035 276.9 -77.605 ;
      RECT 276.5 -68 276.9 -53.36 ;
      RECT 276.5 -49.51 276.9 -12.47 ;
      RECT 268.8 -84.215 269.2 -22.12 ;
      RECT 268 -83.355 268.4 -22.12 ;
      RECT 267.2 -184.035 267.6 -83.445 ;
      RECT 266.4 -67.5 266.8 -52.905 ;
      RECT 266.4 -49.08 266.8 -15.74 ;
      RECT 265.6 -184.035 266 -77.605 ;
      RECT 265.6 -68 266 -53.36 ;
      RECT 265.6 -49.51 266 -12.47 ;
      RECT 257.9 -84.215 258.3 -22.12 ;
      RECT 257.1 -83.355 257.5 -22.12 ;
      RECT 256.3 -184.035 256.7 -83.445 ;
      RECT 255.5 -67.5 255.9 -52.905 ;
      RECT 255.5 -49.08 255.9 -15.74 ;
      RECT 254.7 -184.035 255.1 -77.605 ;
      RECT 254.7 -68 255.1 -53.36 ;
      RECT 254.7 -49.51 255.1 -12.47 ;
      RECT 247 -84.215 247.4 -22.12 ;
      RECT 246.2 -83.355 246.6 -22.12 ;
      RECT 245.4 -184.035 245.8 -83.445 ;
      RECT 244.6 -67.5 245 -52.905 ;
      RECT 244.6 -49.08 245 -15.74 ;
      RECT 243.8 -184.035 244.2 -77.605 ;
      RECT 243.8 -68 244.2 -53.36 ;
      RECT 243.8 -49.51 244.2 -12.47 ;
      RECT 236.1 -84.215 236.5 -22.12 ;
      RECT 235.3 -83.355 235.7 -22.12 ;
      RECT 234.5 -184.035 234.9 -83.445 ;
      RECT 233.7 -67.5 234.1 -52.905 ;
      RECT 233.7 -49.08 234.1 -15.74 ;
      RECT 232.9 -184.035 233.3 -77.605 ;
      RECT 232.9 -68 233.3 -53.36 ;
      RECT 232.9 -49.51 233.3 -12.47 ;
      RECT 225.2 -84.215 225.6 -22.12 ;
      RECT 224.4 -83.355 224.8 -22.12 ;
      RECT 223.6 -184.035 224 -83.445 ;
      RECT 222.8 -67.5 223.2 -52.905 ;
      RECT 222.8 -49.08 223.2 -15.74 ;
      RECT 222 -184.035 222.4 -77.605 ;
      RECT 222 -68 222.4 -53.36 ;
      RECT 222 -49.51 222.4 -12.47 ;
      RECT 214.3 -84.215 214.7 -22.12 ;
      RECT 213.5 -83.355 213.9 -22.12 ;
      RECT 212.7 -184.035 213.1 -83.445 ;
      RECT 211.9 -67.5 212.3 -52.905 ;
      RECT 211.9 -49.08 212.3 -15.74 ;
      RECT 211.1 -184.035 211.5 -77.605 ;
      RECT 211.1 -68 211.5 -53.36 ;
      RECT 211.1 -49.51 211.5 -12.47 ;
      RECT 203.4 -84.215 203.8 -22.12 ;
      RECT 202.6 -83.355 203 -22.12 ;
      RECT 201.8 -184.035 202.2 -83.445 ;
      RECT 201 -67.5 201.4 -52.905 ;
      RECT 201 -49.08 201.4 -15.74 ;
      RECT 200.2 -184.035 200.6 -77.605 ;
      RECT 200.2 -68 200.6 -53.36 ;
      RECT 200.2 -49.51 200.6 -12.47 ;
      RECT 192.5 -84.215 192.9 -22.12 ;
      RECT 191.7 -83.355 192.1 -22.12 ;
      RECT 190.9 -184.035 191.3 -83.445 ;
      RECT 190.1 -67.5 190.5 -52.905 ;
      RECT 190.1 -49.08 190.5 -15.74 ;
      RECT 189.3 -184.035 189.7 -77.605 ;
      RECT 189.3 -68 189.7 -53.36 ;
      RECT 189.3 -49.51 189.7 -12.47 ;
      RECT 181.6 -84.215 182 -22.12 ;
      RECT 180.8 -83.355 181.2 -22.12 ;
      RECT 180 -184.035 180.4 -83.445 ;
      RECT 179.2 -67.5 179.6 -52.905 ;
      RECT 179.2 -49.08 179.6 -15.74 ;
      RECT 178.4 -184.035 178.8 -77.605 ;
      RECT 178.4 -68 178.8 -53.36 ;
      RECT 178.4 -49.51 178.8 -12.47 ;
      RECT 170.7 -84.215 171.1 -22.12 ;
      RECT 169.9 -83.355 170.3 -22.12 ;
      RECT 169.1 -184.035 169.5 -83.445 ;
      RECT 168.3 -67.5 168.7 -52.905 ;
      RECT 168.3 -49.08 168.7 -15.74 ;
      RECT 167.5 -184.035 167.9 -77.605 ;
      RECT 167.5 -68 167.9 -53.36 ;
      RECT 167.5 -49.51 167.9 -12.47 ;
      RECT 159.8 -84.215 160.2 -22.12 ;
      RECT 159 -83.355 159.4 -22.12 ;
      RECT 158.2 -184.035 158.6 -83.445 ;
      RECT 157.4 -67.5 157.8 -52.905 ;
      RECT 157.4 -49.08 157.8 -15.74 ;
      RECT 156.6 -184.035 157 -77.605 ;
      RECT 156.6 -68 157 -53.36 ;
      RECT 156.6 -49.51 157 -12.47 ;
      RECT 148.9 -84.215 149.3 -22.12 ;
      RECT 148.1 -83.355 148.5 -22.12 ;
      RECT 147.3 -184.035 147.7 -83.445 ;
      RECT 146.5 -67.5 146.9 -52.905 ;
      RECT 146.5 -49.08 146.9 -15.74 ;
      RECT 145.7 -184.035 146.1 -77.605 ;
      RECT 145.7 -68 146.1 -53.36 ;
      RECT 145.7 -49.51 146.1 -12.47 ;
      RECT 138 -84.215 138.4 -22.12 ;
      RECT 137.2 -83.355 137.6 -22.12 ;
      RECT 136.4 -184.035 136.8 -83.445 ;
      RECT 135.6 -67.5 136 -52.905 ;
      RECT 135.6 -49.08 136 -15.74 ;
      RECT 134.8 -184.035 135.2 -77.605 ;
      RECT 134.8 -68 135.2 -53.36 ;
      RECT 134.8 -49.51 135.2 -12.47 ;
      RECT 127.1 -84.215 127.5 -22.12 ;
      RECT 126.3 -83.355 126.7 -22.12 ;
      RECT 125.5 -184.035 125.9 -83.445 ;
      RECT 124.7 -67.5 125.1 -52.905 ;
      RECT 124.7 -49.08 125.1 -15.74 ;
      RECT 123.9 -184.035 124.3 -77.605 ;
      RECT 123.9 -68 124.3 -53.36 ;
      RECT 123.9 -49.51 124.3 -12.47 ;
      RECT 116.2 -84.215 116.6 -22.12 ;
      RECT 115.4 -83.355 115.8 -22.12 ;
      RECT 114.6 -184.035 115 -83.445 ;
      RECT 113.8 -67.5 114.2 -52.905 ;
      RECT 113.8 -49.08 114.2 -15.74 ;
      RECT 113 -184.035 113.4 -77.605 ;
      RECT 113 -68 113.4 -53.36 ;
      RECT 113 -49.51 113.4 -12.47 ;
      RECT 105.3 -84.215 105.7 -22.12 ;
      RECT 104.5 -83.355 104.9 -22.12 ;
      RECT 103.7 -184.035 104.1 -83.445 ;
      RECT 102.9 -67.5 103.3 -52.905 ;
      RECT 102.9 -49.08 103.3 -15.74 ;
      RECT 102.1 -184.035 102.5 -77.605 ;
      RECT 102.1 -68 102.5 -53.36 ;
      RECT 102.1 -49.51 102.5 -12.47 ;
      RECT 94.4 -84.215 94.8 -22.12 ;
      RECT 93.6 -83.355 94 -22.12 ;
      RECT 92.8 -184.035 93.2 -83.445 ;
      RECT 92 -67.5 92.4 -52.905 ;
      RECT 92 -49.08 92.4 -15.74 ;
      RECT 91.2 -184.035 91.6 -77.605 ;
      RECT 91.2 -68 91.6 -53.36 ;
      RECT 91.2 -49.51 91.6 -12.47 ;
      RECT 83.5 -84.215 83.9 -22.12 ;
      RECT 82.7 -83.355 83.1 -22.12 ;
      RECT 81.9 -184.035 82.3 -83.445 ;
      RECT 81.1 -67.5 81.5 -52.905 ;
      RECT 81.1 -49.08 81.5 -15.74 ;
      RECT 80.3 -184.035 80.7 -77.605 ;
      RECT 80.3 -68 80.7 -53.36 ;
      RECT 80.3 -49.51 80.7 -12.47 ;
      RECT 72.6 -84.215 73 -22.12 ;
      RECT 71.8 -83.355 72.2 -22.12 ;
      RECT 71 -184.035 71.4 -83.445 ;
      RECT 70.2 -67.5 70.6 -52.905 ;
      RECT 70.2 -49.08 70.6 -15.74 ;
      RECT 69.4 -184.035 69.8 -77.605 ;
      RECT 69.4 -68 69.8 -53.36 ;
      RECT 69.4 -49.51 69.8 -12.47 ;
      RECT 61.7 -84.215 62.1 -22.12 ;
      RECT 60.9 -83.355 61.3 -22.12 ;
      RECT 60.1 -184.035 60.5 -83.445 ;
      RECT 59.3 -67.5 59.7 -52.905 ;
      RECT 59.3 -49.08 59.7 -15.74 ;
      RECT 58.5 -184.035 58.9 -77.605 ;
      RECT 58.5 -68 58.9 -53.36 ;
      RECT 58.5 -49.51 58.9 -12.47 ;
      RECT 50.8 -84.215 51.2 -22.12 ;
      RECT 50 -83.355 50.4 -22.12 ;
      RECT 49.2 -184.035 49.6 -83.445 ;
      RECT 48.4 -67.5 48.8 -52.905 ;
      RECT 48.4 -49.08 48.8 -15.74 ;
      RECT 47.6 -184.035 48 -77.605 ;
      RECT 47.6 -68 48 -53.36 ;
      RECT 47.6 -49.51 48 -12.47 ;
      RECT 39.9 -84.215 40.3 -22.12 ;
      RECT 39.1 -83.355 39.5 -22.12 ;
      RECT 38.3 -184.035 38.7 -83.445 ;
      RECT 37.5 -67.5 37.9 -52.905 ;
      RECT 37.5 -49.08 37.9 -15.74 ;
      RECT 36.7 -184.035 37.1 -77.605 ;
      RECT 36.7 -68 37.1 -53.36 ;
      RECT 36.7 -49.51 37.1 -12.47 ;
      RECT 29 -84.215 29.4 -22.12 ;
      RECT 28.2 -83.355 28.6 -22.12 ;
      RECT 27.4 -184.035 27.8 -83.445 ;
      RECT 26.6 -67.5 27 -52.905 ;
      RECT 26.6 -49.08 27 -15.74 ;
      RECT 25.8 -184.035 26.2 -77.605 ;
      RECT 25.8 -68 26.2 -53.36 ;
      RECT 25.8 -49.51 26.2 -12.47 ;
      RECT 18.1 -84.215 18.5 -22.12 ;
      RECT 17.3 -83.355 17.7 -22.12 ;
      RECT 16.5 -184.035 16.9 -83.445 ;
      RECT 15.7 -67.5 16.1 -52.905 ;
      RECT 15.7 -49.08 16.1 -15.74 ;
      RECT 14.9 -184.035 15.3 -77.605 ;
      RECT 14.9 -68 15.3 -53.36 ;
      RECT 14.9 -49.51 15.3 -12.47 ;
      RECT 8 -91.06 8.4 -22.12 ;
      RECT 7.2 -84.215 7.6 -22.12 ;
      RECT 6.4 -184.035 6.8 -91.15 ;
      RECT 6.4 -83.355 6.8 -22.12 ;
      RECT 5.6 -184.035 6 -83.445 ;
      RECT 4.8 -67.5 5.2 -52.905 ;
      RECT 4.8 -49.08 5.2 -15.74 ;
      RECT 4 -184.035 4.4 -77.605 ;
      RECT 4 -68 4.4 -53.36 ;
      RECT 4 -49.51 4.4 -12.47 ;
  END
END sram22_1024x32m8w32

END LIBRARY
