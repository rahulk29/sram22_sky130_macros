* circuit.Package sramgen_sramgen_sram_4096x8m8w8_replica_v1
* Written by SpiceNetlister
* 

.SUBCKT hierarchical_decoder_nand_2 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder_inv_3 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder_nand_92 
+ gnd vdd a b c y 

xn1 
+ x1 a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ x2 b x1 gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn3 
+ y c x2 gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp3 
+ y c vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT hierarchical_decoder 
+ vdd gnd addr[8] addr[7] addr[6] addr[5] addr[4] addr[3] addr[2] addr[1] addr[0] addr_b[8] addr_b[7] addr_b[6] addr_b[5] addr_b[4] addr_b[3] addr_b[2] addr_b[1] addr_b[0] decode[511] decode[510] decode[509] decode[508] decode[507] decode[506] decode[505] decode[504] decode[503] decode[502] decode[501] decode[500] decode[499] decode[498] decode[497] decode[496] decode[495] decode[494] decode[493] decode[492] decode[491] decode[490] decode[489] decode[488] decode[487] decode[486] decode[485] decode[484] decode[483] decode[482] decode[481] decode[480] decode[479] decode[478] decode[477] decode[476] decode[475] decode[474] decode[473] decode[472] decode[471] decode[470] decode[469] decode[468] decode[467] decode[466] decode[465] decode[464] decode[463] decode[462] decode[461] decode[460] decode[459] decode[458] decode[457] decode[456] decode[455] decode[454] decode[453] decode[452] decode[451] decode[450] decode[449] decode[448] decode[447] decode[446] decode[445] decode[444] decode[443] decode[442] decode[441] decode[440] decode[439] decode[438] decode[437] decode[436] decode[435] decode[434] decode[433] decode[432] decode[431] decode[430] decode[429] decode[428] decode[427] decode[426] decode[425] decode[424] decode[423] decode[422] decode[421] decode[420] decode[419] decode[418] decode[417] decode[416] decode[415] decode[414] decode[413] decode[412] decode[411] decode[410] decode[409] decode[408] decode[407] decode[406] decode[405] decode[404] decode[403] decode[402] decode[401] decode[400] decode[399] decode[398] decode[397] decode[396] decode[395] decode[394] decode[393] decode[392] decode[391] decode[390] decode[389] decode[388] decode[387] decode[386] decode[385] decode[384] decode[383] decode[382] decode[381] decode[380] decode[379] decode[378] decode[377] decode[376] decode[375] decode[374] decode[373] decode[372] decode[371] decode[370] decode[369] decode[368] decode[367] decode[366] decode[365] decode[364] decode[363] decode[362] decode[361] decode[360] decode[359] decode[358] decode[357] decode[356] decode[355] decode[354] decode[353] decode[352] decode[351] decode[350] decode[349] decode[348] decode[347] decode[346] decode[345] decode[344] decode[343] decode[342] decode[341] decode[340] decode[339] decode[338] decode[337] decode[336] decode[335] decode[334] decode[333] decode[332] decode[331] decode[330] decode[329] decode[328] decode[327] decode[326] decode[325] decode[324] decode[323] decode[322] decode[321] decode[320] decode[319] decode[318] decode[317] decode[316] decode[315] decode[314] decode[313] decode[312] decode[311] decode[310] decode[309] decode[308] decode[307] decode[306] decode[305] decode[304] decode[303] decode[302] decode[301] decode[300] decode[299] decode[298] decode[297] decode[296] decode[295] decode[294] decode[293] decode[292] decode[291] decode[290] decode[289] decode[288] decode[287] decode[286] decode[285] decode[284] decode[283] decode[282] decode[281] decode[280] decode[279] decode[278] decode[277] decode[276] decode[275] decode[274] decode[273] decode[272] decode[271] decode[270] decode[269] decode[268] decode[267] decode[266] decode[265] decode[264] decode[263] decode[262] decode[261] decode[260] decode[259] decode[258] decode[257] decode[256] decode[255] decode[254] decode[253] decode[252] decode[251] decode[250] decode[249] decode[248] decode[247] decode[246] decode[245] decode[244] decode[243] decode[242] decode[241] decode[240] decode[239] decode[238] decode[237] decode[236] decode[235] decode[234] decode[233] decode[232] decode[231] decode[230] decode[229] decode[228] decode[227] decode[226] decode[225] decode[224] decode[223] decode[222] decode[221] decode[220] decode[219] decode[218] decode[217] decode[216] decode[215] decode[214] decode[213] decode[212] decode[211] decode[210] decode[209] decode[208] decode[207] decode[206] decode[205] decode[204] decode[203] decode[202] decode[201] decode[200] decode[199] decode[198] decode[197] decode[196] decode[195] decode[194] decode[193] decode[192] decode[191] decode[190] decode[189] decode[188] decode[187] decode[186] decode[185] decode[184] decode[183] decode[182] decode[181] decode[180] decode[179] decode[178] decode[177] decode[176] decode[175] decode[174] decode[173] decode[172] decode[171] decode[170] decode[169] decode[168] decode[167] decode[166] decode[165] decode[164] decode[163] decode[162] decode[161] decode[160] decode[159] decode[158] decode[157] decode[156] decode[155] decode[154] decode[153] decode[152] decode[151] decode[150] decode[149] decode[148] decode[147] decode[146] decode[145] decode[144] decode[143] decode[142] decode[141] decode[140] decode[139] decode[138] decode[137] decode[136] decode[135] decode[134] decode[133] decode[132] decode[131] decode[130] decode[129] decode[128] decode[127] decode[126] decode[125] decode[124] decode[123] decode[122] decode[121] decode[120] decode[119] decode[118] decode[117] decode[116] decode[115] decode[114] decode[113] decode[112] decode[111] decode[110] decode[109] decode[108] decode[107] decode[106] decode[105] decode[104] decode[103] decode[102] decode[101] decode[100] decode[99] decode[98] decode[97] decode[96] decode[95] decode[94] decode[93] decode[92] decode[91] decode[90] decode[89] decode[88] decode[87] decode[86] decode[85] decode[84] decode[83] decode[82] decode[81] decode[80] decode[79] decode[78] decode[77] decode[76] decode[75] decode[74] decode[73] decode[72] decode[71] decode[70] decode[69] decode[68] decode[67] decode[66] decode[65] decode[64] decode[63] decode[62] decode[61] decode[60] decode[59] decode[58] decode[57] decode[56] decode[55] decode[54] decode[53] decode[52] decode[51] decode[50] decode[49] decode[48] decode[47] decode[46] decode[45] decode[44] decode[43] decode[42] decode[41] decode[40] decode[39] decode[38] decode[37] decode[36] decode[35] decode[34] decode[33] decode[32] decode[31] decode[30] decode[29] decode[28] decode[27] decode[26] decode[25] decode[24] decode[23] decode[22] decode[21] decode[20] decode[19] decode[18] decode[17] decode[16] decode[15] decode[14] decode[13] decode[12] decode[11] decode[10] decode[9] decode[8] decode[7] decode[6] decode[5] decode[4] decode[3] decode[2] decode[1] decode[0] decode_b[511] decode_b[510] decode_b[509] decode_b[508] decode_b[507] decode_b[506] decode_b[505] decode_b[504] decode_b[503] decode_b[502] decode_b[501] decode_b[500] decode_b[499] decode_b[498] decode_b[497] decode_b[496] decode_b[495] decode_b[494] decode_b[493] decode_b[492] decode_b[491] decode_b[490] decode_b[489] decode_b[488] decode_b[487] decode_b[486] decode_b[485] decode_b[484] decode_b[483] decode_b[482] decode_b[481] decode_b[480] decode_b[479] decode_b[478] decode_b[477] decode_b[476] decode_b[475] decode_b[474] decode_b[473] decode_b[472] decode_b[471] decode_b[470] decode_b[469] decode_b[468] decode_b[467] decode_b[466] decode_b[465] decode_b[464] decode_b[463] decode_b[462] decode_b[461] decode_b[460] decode_b[459] decode_b[458] decode_b[457] decode_b[456] decode_b[455] decode_b[454] decode_b[453] decode_b[452] decode_b[451] decode_b[450] decode_b[449] decode_b[448] decode_b[447] decode_b[446] decode_b[445] decode_b[444] decode_b[443] decode_b[442] decode_b[441] decode_b[440] decode_b[439] decode_b[438] decode_b[437] decode_b[436] decode_b[435] decode_b[434] decode_b[433] decode_b[432] decode_b[431] decode_b[430] decode_b[429] decode_b[428] decode_b[427] decode_b[426] decode_b[425] decode_b[424] decode_b[423] decode_b[422] decode_b[421] decode_b[420] decode_b[419] decode_b[418] decode_b[417] decode_b[416] decode_b[415] decode_b[414] decode_b[413] decode_b[412] decode_b[411] decode_b[410] decode_b[409] decode_b[408] decode_b[407] decode_b[406] decode_b[405] decode_b[404] decode_b[403] decode_b[402] decode_b[401] decode_b[400] decode_b[399] decode_b[398] decode_b[397] decode_b[396] decode_b[395] decode_b[394] decode_b[393] decode_b[392] decode_b[391] decode_b[390] decode_b[389] decode_b[388] decode_b[387] decode_b[386] decode_b[385] decode_b[384] decode_b[383] decode_b[382] decode_b[381] decode_b[380] decode_b[379] decode_b[378] decode_b[377] decode_b[376] decode_b[375] decode_b[374] decode_b[373] decode_b[372] decode_b[371] decode_b[370] decode_b[369] decode_b[368] decode_b[367] decode_b[366] decode_b[365] decode_b[364] decode_b[363] decode_b[362] decode_b[361] decode_b[360] decode_b[359] decode_b[358] decode_b[357] decode_b[356] decode_b[355] decode_b[354] decode_b[353] decode_b[352] decode_b[351] decode_b[350] decode_b[349] decode_b[348] decode_b[347] decode_b[346] decode_b[345] decode_b[344] decode_b[343] decode_b[342] decode_b[341] decode_b[340] decode_b[339] decode_b[338] decode_b[337] decode_b[336] decode_b[335] decode_b[334] decode_b[333] decode_b[332] decode_b[331] decode_b[330] decode_b[329] decode_b[328] decode_b[327] decode_b[326] decode_b[325] decode_b[324] decode_b[323] decode_b[322] decode_b[321] decode_b[320] decode_b[319] decode_b[318] decode_b[317] decode_b[316] decode_b[315] decode_b[314] decode_b[313] decode_b[312] decode_b[311] decode_b[310] decode_b[309] decode_b[308] decode_b[307] decode_b[306] decode_b[305] decode_b[304] decode_b[303] decode_b[302] decode_b[301] decode_b[300] decode_b[299] decode_b[298] decode_b[297] decode_b[296] decode_b[295] decode_b[294] decode_b[293] decode_b[292] decode_b[291] decode_b[290] decode_b[289] decode_b[288] decode_b[287] decode_b[286] decode_b[285] decode_b[284] decode_b[283] decode_b[282] decode_b[281] decode_b[280] decode_b[279] decode_b[278] decode_b[277] decode_b[276] decode_b[275] decode_b[274] decode_b[273] decode_b[272] decode_b[271] decode_b[270] decode_b[269] decode_b[268] decode_b[267] decode_b[266] decode_b[265] decode_b[264] decode_b[263] decode_b[262] decode_b[261] decode_b[260] decode_b[259] decode_b[258] decode_b[257] decode_b[256] decode_b[255] decode_b[254] decode_b[253] decode_b[252] decode_b[251] decode_b[250] decode_b[249] decode_b[248] decode_b[247] decode_b[246] decode_b[245] decode_b[244] decode_b[243] decode_b[242] decode_b[241] decode_b[240] decode_b[239] decode_b[238] decode_b[237] decode_b[236] decode_b[235] decode_b[234] decode_b[233] decode_b[232] decode_b[231] decode_b[230] decode_b[229] decode_b[228] decode_b[227] decode_b[226] decode_b[225] decode_b[224] decode_b[223] decode_b[222] decode_b[221] decode_b[220] decode_b[219] decode_b[218] decode_b[217] decode_b[216] decode_b[215] decode_b[214] decode_b[213] decode_b[212] decode_b[211] decode_b[210] decode_b[209] decode_b[208] decode_b[207] decode_b[206] decode_b[205] decode_b[204] decode_b[203] decode_b[202] decode_b[201] decode_b[200] decode_b[199] decode_b[198] decode_b[197] decode_b[196] decode_b[195] decode_b[194] decode_b[193] decode_b[192] decode_b[191] decode_b[190] decode_b[189] decode_b[188] decode_b[187] decode_b[186] decode_b[185] decode_b[184] decode_b[183] decode_b[182] decode_b[181] decode_b[180] decode_b[179] decode_b[178] decode_b[177] decode_b[176] decode_b[175] decode_b[174] decode_b[173] decode_b[172] decode_b[171] decode_b[170] decode_b[169] decode_b[168] decode_b[167] decode_b[166] decode_b[165] decode_b[164] decode_b[163] decode_b[162] decode_b[161] decode_b[160] decode_b[159] decode_b[158] decode_b[157] decode_b[156] decode_b[155] decode_b[154] decode_b[153] decode_b[152] decode_b[151] decode_b[150] decode_b[149] decode_b[148] decode_b[147] decode_b[146] decode_b[145] decode_b[144] decode_b[143] decode_b[142] decode_b[141] decode_b[140] decode_b[139] decode_b[138] decode_b[137] decode_b[136] decode_b[135] decode_b[134] decode_b[133] decode_b[132] decode_b[131] decode_b[130] decode_b[129] decode_b[128] decode_b[127] decode_b[126] decode_b[125] decode_b[124] decode_b[123] decode_b[122] decode_b[121] decode_b[120] decode_b[119] decode_b[118] decode_b[117] decode_b[116] decode_b[115] decode_b[114] decode_b[113] decode_b[112] decode_b[111] decode_b[110] decode_b[109] decode_b[108] decode_b[107] decode_b[106] decode_b[105] decode_b[104] decode_b[103] decode_b[102] decode_b[101] decode_b[100] decode_b[99] decode_b[98] decode_b[97] decode_b[96] decode_b[95] decode_b[94] decode_b[93] decode_b[92] decode_b[91] decode_b[90] decode_b[89] decode_b[88] decode_b[87] decode_b[86] decode_b[85] decode_b[84] decode_b[83] decode_b[82] decode_b[81] decode_b[80] decode_b[79] decode_b[78] decode_b[77] decode_b[76] decode_b[75] decode_b[74] decode_b[73] decode_b[72] decode_b[71] decode_b[70] decode_b[69] decode_b[68] decode_b[67] decode_b[66] decode_b[65] decode_b[64] decode_b[63] decode_b[62] decode_b[61] decode_b[60] decode_b[59] decode_b[58] decode_b[57] decode_b[56] decode_b[55] decode_b[54] decode_b[53] decode_b[52] decode_b[51] decode_b[50] decode_b[49] decode_b[48] decode_b[47] decode_b[46] decode_b[45] decode_b[44] decode_b[43] decode_b[42] decode_b[41] decode_b[40] decode_b[39] decode_b[38] decode_b[37] decode_b[36] decode_b[35] decode_b[34] decode_b[33] decode_b[32] decode_b[31] decode_b[30] decode_b[29] decode_b[28] decode_b[27] decode_b[26] decode_b[25] decode_b[24] decode_b[23] decode_b[22] decode_b[21] decode_b[20] decode_b[19] decode_b[18] decode_b[17] decode_b[16] decode_b[15] decode_b[14] decode_b[13] decode_b[12] decode_b[11] decode_b[10] decode_b[9] decode_b[8] decode_b[7] decode_b[6] decode_b[5] decode_b[4] decode_b[3] decode_b[2] decode_b[1] decode_b[0] 

xnand_5 
+ gnd vdd addr_b[8] addr_b[7] net_4 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_6 
+ gnd vdd net_4 predecode_1[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_8 
+ gnd vdd addr_b[8] addr[7] net_7 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_9 
+ gnd vdd net_7 predecode_1[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_11 
+ gnd vdd addr[8] addr_b[7] net_10 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_12 
+ gnd vdd net_10 predecode_1[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_14 
+ gnd vdd addr[8] addr[7] net_13 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_15 
+ gnd vdd net_13 predecode_1[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_18 
+ gnd vdd addr_b[6] addr_b[5] net_17 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_19 
+ gnd vdd net_17 predecode_16[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_21 
+ gnd vdd addr_b[6] addr[5] net_20 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_22 
+ gnd vdd net_20 predecode_16[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_24 
+ gnd vdd addr[6] addr_b[5] net_23 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_25 
+ gnd vdd net_23 predecode_16[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_27 
+ gnd vdd addr[6] addr[5] net_26 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_28 
+ gnd vdd net_26 predecode_16[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_31 
+ gnd vdd predecode_1[0] predecode_16[0] net_30 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_32 
+ gnd vdd net_30 predecode_29[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_34 
+ gnd vdd predecode_1[0] predecode_16[1] net_33 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_35 
+ gnd vdd net_33 predecode_29[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_37 
+ gnd vdd predecode_1[0] predecode_16[2] net_36 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_38 
+ gnd vdd net_36 predecode_29[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_40 
+ gnd vdd predecode_1[0] predecode_16[3] net_39 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_41 
+ gnd vdd net_39 predecode_29[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_43 
+ gnd vdd predecode_1[1] predecode_16[0] net_42 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_44 
+ gnd vdd net_42 predecode_29[4] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_46 
+ gnd vdd predecode_1[1] predecode_16[1] net_45 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_47 
+ gnd vdd net_45 predecode_29[5] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_49 
+ gnd vdd predecode_1[1] predecode_16[2] net_48 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_50 
+ gnd vdd net_48 predecode_29[6] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_52 
+ gnd vdd predecode_1[1] predecode_16[3] net_51 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_53 
+ gnd vdd net_51 predecode_29[7] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_55 
+ gnd vdd predecode_1[2] predecode_16[0] net_54 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_56 
+ gnd vdd net_54 predecode_29[8] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_58 
+ gnd vdd predecode_1[2] predecode_16[1] net_57 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_59 
+ gnd vdd net_57 predecode_29[9] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_61 
+ gnd vdd predecode_1[2] predecode_16[2] net_60 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_62 
+ gnd vdd net_60 predecode_29[10] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_64 
+ gnd vdd predecode_1[2] predecode_16[3] net_63 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_65 
+ gnd vdd net_63 predecode_29[11] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_67 
+ gnd vdd predecode_1[3] predecode_16[0] net_66 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_68 
+ gnd vdd net_66 predecode_29[12] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_70 
+ gnd vdd predecode_1[3] predecode_16[1] net_69 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_71 
+ gnd vdd net_69 predecode_29[13] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_73 
+ gnd vdd predecode_1[3] predecode_16[2] net_72 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_74 
+ gnd vdd net_72 predecode_29[14] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_76 
+ gnd vdd predecode_1[3] predecode_16[3] net_75 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_77 
+ gnd vdd net_75 predecode_29[15] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_80 
+ gnd vdd addr_b[4] addr_b[3] net_79 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_81 
+ gnd vdd net_79 predecode_78[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_83 
+ gnd vdd addr_b[4] addr[3] net_82 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_84 
+ gnd vdd net_82 predecode_78[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_86 
+ gnd vdd addr[4] addr_b[3] net_85 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_87 
+ gnd vdd net_85 predecode_78[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_89 
+ gnd vdd addr[4] addr[3] net_88 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_90 
+ gnd vdd net_88 predecode_78[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_94 
+ gnd vdd addr_b[2] addr_b[1] addr_b[0] net_93 
+ hierarchical_decoder_nand_92 
* No parameters

xinv_95 
+ gnd vdd net_93 predecode_91[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_97 
+ gnd vdd addr_b[2] addr_b[1] addr[0] net_96 
+ hierarchical_decoder_nand_92 
* No parameters

xinv_98 
+ gnd vdd net_96 predecode_91[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_100 
+ gnd vdd addr_b[2] addr[1] addr_b[0] net_99 
+ hierarchical_decoder_nand_92 
* No parameters

xinv_101 
+ gnd vdd net_99 predecode_91[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_103 
+ gnd vdd addr_b[2] addr[1] addr[0] net_102 
+ hierarchical_decoder_nand_92 
* No parameters

xinv_104 
+ gnd vdd net_102 predecode_91[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_106 
+ gnd vdd addr[2] addr_b[1] addr_b[0] net_105 
+ hierarchical_decoder_nand_92 
* No parameters

xinv_107 
+ gnd vdd net_105 predecode_91[4] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_109 
+ gnd vdd addr[2] addr_b[1] addr[0] net_108 
+ hierarchical_decoder_nand_92 
* No parameters

xinv_110 
+ gnd vdd net_108 predecode_91[5] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_112 
+ gnd vdd addr[2] addr[1] addr_b[0] net_111 
+ hierarchical_decoder_nand_92 
* No parameters

xinv_113 
+ gnd vdd net_111 predecode_91[6] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_115 
+ gnd vdd addr[2] addr[1] addr[0] net_114 
+ hierarchical_decoder_nand_92 
* No parameters

xinv_116 
+ gnd vdd net_114 predecode_91[7] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_119 
+ gnd vdd predecode_78[0] predecode_91[0] net_118 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_120 
+ gnd vdd net_118 predecode_117[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_122 
+ gnd vdd predecode_78[0] predecode_91[1] net_121 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_123 
+ gnd vdd net_121 predecode_117[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_125 
+ gnd vdd predecode_78[0] predecode_91[2] net_124 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_126 
+ gnd vdd net_124 predecode_117[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_128 
+ gnd vdd predecode_78[0] predecode_91[3] net_127 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_129 
+ gnd vdd net_127 predecode_117[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_131 
+ gnd vdd predecode_78[0] predecode_91[4] net_130 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_132 
+ gnd vdd net_130 predecode_117[4] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_134 
+ gnd vdd predecode_78[0] predecode_91[5] net_133 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_135 
+ gnd vdd net_133 predecode_117[5] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_137 
+ gnd vdd predecode_78[0] predecode_91[6] net_136 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_138 
+ gnd vdd net_136 predecode_117[6] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_140 
+ gnd vdd predecode_78[0] predecode_91[7] net_139 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_141 
+ gnd vdd net_139 predecode_117[7] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_143 
+ gnd vdd predecode_78[1] predecode_91[0] net_142 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_144 
+ gnd vdd net_142 predecode_117[8] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_146 
+ gnd vdd predecode_78[1] predecode_91[1] net_145 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_147 
+ gnd vdd net_145 predecode_117[9] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_149 
+ gnd vdd predecode_78[1] predecode_91[2] net_148 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_150 
+ gnd vdd net_148 predecode_117[10] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_152 
+ gnd vdd predecode_78[1] predecode_91[3] net_151 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_153 
+ gnd vdd net_151 predecode_117[11] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_155 
+ gnd vdd predecode_78[1] predecode_91[4] net_154 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_156 
+ gnd vdd net_154 predecode_117[12] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_158 
+ gnd vdd predecode_78[1] predecode_91[5] net_157 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_159 
+ gnd vdd net_157 predecode_117[13] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_161 
+ gnd vdd predecode_78[1] predecode_91[6] net_160 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_162 
+ gnd vdd net_160 predecode_117[14] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_164 
+ gnd vdd predecode_78[1] predecode_91[7] net_163 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_165 
+ gnd vdd net_163 predecode_117[15] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_167 
+ gnd vdd predecode_78[2] predecode_91[0] net_166 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_168 
+ gnd vdd net_166 predecode_117[16] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_170 
+ gnd vdd predecode_78[2] predecode_91[1] net_169 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_171 
+ gnd vdd net_169 predecode_117[17] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_173 
+ gnd vdd predecode_78[2] predecode_91[2] net_172 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_174 
+ gnd vdd net_172 predecode_117[18] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_176 
+ gnd vdd predecode_78[2] predecode_91[3] net_175 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_177 
+ gnd vdd net_175 predecode_117[19] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_179 
+ gnd vdd predecode_78[2] predecode_91[4] net_178 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_180 
+ gnd vdd net_178 predecode_117[20] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_182 
+ gnd vdd predecode_78[2] predecode_91[5] net_181 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_183 
+ gnd vdd net_181 predecode_117[21] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_185 
+ gnd vdd predecode_78[2] predecode_91[6] net_184 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_186 
+ gnd vdd net_184 predecode_117[22] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_188 
+ gnd vdd predecode_78[2] predecode_91[7] net_187 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_189 
+ gnd vdd net_187 predecode_117[23] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_191 
+ gnd vdd predecode_78[3] predecode_91[0] net_190 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_192 
+ gnd vdd net_190 predecode_117[24] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_194 
+ gnd vdd predecode_78[3] predecode_91[1] net_193 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_195 
+ gnd vdd net_193 predecode_117[25] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_197 
+ gnd vdd predecode_78[3] predecode_91[2] net_196 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_198 
+ gnd vdd net_196 predecode_117[26] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_200 
+ gnd vdd predecode_78[3] predecode_91[3] net_199 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_201 
+ gnd vdd net_199 predecode_117[27] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_203 
+ gnd vdd predecode_78[3] predecode_91[4] net_202 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_204 
+ gnd vdd net_202 predecode_117[28] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_206 
+ gnd vdd predecode_78[3] predecode_91[5] net_205 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_207 
+ gnd vdd net_205 predecode_117[29] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_209 
+ gnd vdd predecode_78[3] predecode_91[6] net_208 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_210 
+ gnd vdd net_208 predecode_117[30] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_212 
+ gnd vdd predecode_78[3] predecode_91[7] net_211 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_213 
+ gnd vdd net_211 predecode_117[31] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_214 
+ gnd vdd predecode_29[0] predecode_117[0] decode_b[0] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_215 
+ gnd vdd decode_b[0] decode[0] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_216 
+ gnd vdd predecode_29[0] predecode_117[1] decode_b[1] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_217 
+ gnd vdd decode_b[1] decode[1] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_218 
+ gnd vdd predecode_29[0] predecode_117[2] decode_b[2] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_219 
+ gnd vdd decode_b[2] decode[2] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_220 
+ gnd vdd predecode_29[0] predecode_117[3] decode_b[3] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_221 
+ gnd vdd decode_b[3] decode[3] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_222 
+ gnd vdd predecode_29[0] predecode_117[4] decode_b[4] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_223 
+ gnd vdd decode_b[4] decode[4] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_224 
+ gnd vdd predecode_29[0] predecode_117[5] decode_b[5] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_225 
+ gnd vdd decode_b[5] decode[5] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_226 
+ gnd vdd predecode_29[0] predecode_117[6] decode_b[6] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_227 
+ gnd vdd decode_b[6] decode[6] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_228 
+ gnd vdd predecode_29[0] predecode_117[7] decode_b[7] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_229 
+ gnd vdd decode_b[7] decode[7] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_230 
+ gnd vdd predecode_29[0] predecode_117[8] decode_b[8] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_231 
+ gnd vdd decode_b[8] decode[8] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_232 
+ gnd vdd predecode_29[0] predecode_117[9] decode_b[9] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_233 
+ gnd vdd decode_b[9] decode[9] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_234 
+ gnd vdd predecode_29[0] predecode_117[10] decode_b[10] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_235 
+ gnd vdd decode_b[10] decode[10] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_236 
+ gnd vdd predecode_29[0] predecode_117[11] decode_b[11] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_237 
+ gnd vdd decode_b[11] decode[11] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_238 
+ gnd vdd predecode_29[0] predecode_117[12] decode_b[12] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_239 
+ gnd vdd decode_b[12] decode[12] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_240 
+ gnd vdd predecode_29[0] predecode_117[13] decode_b[13] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_241 
+ gnd vdd decode_b[13] decode[13] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_242 
+ gnd vdd predecode_29[0] predecode_117[14] decode_b[14] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_243 
+ gnd vdd decode_b[14] decode[14] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_244 
+ gnd vdd predecode_29[0] predecode_117[15] decode_b[15] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_245 
+ gnd vdd decode_b[15] decode[15] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_246 
+ gnd vdd predecode_29[0] predecode_117[16] decode_b[16] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_247 
+ gnd vdd decode_b[16] decode[16] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_248 
+ gnd vdd predecode_29[0] predecode_117[17] decode_b[17] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_249 
+ gnd vdd decode_b[17] decode[17] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_250 
+ gnd vdd predecode_29[0] predecode_117[18] decode_b[18] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_251 
+ gnd vdd decode_b[18] decode[18] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_252 
+ gnd vdd predecode_29[0] predecode_117[19] decode_b[19] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_253 
+ gnd vdd decode_b[19] decode[19] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_254 
+ gnd vdd predecode_29[0] predecode_117[20] decode_b[20] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_255 
+ gnd vdd decode_b[20] decode[20] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_256 
+ gnd vdd predecode_29[0] predecode_117[21] decode_b[21] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_257 
+ gnd vdd decode_b[21] decode[21] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_258 
+ gnd vdd predecode_29[0] predecode_117[22] decode_b[22] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_259 
+ gnd vdd decode_b[22] decode[22] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_260 
+ gnd vdd predecode_29[0] predecode_117[23] decode_b[23] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_261 
+ gnd vdd decode_b[23] decode[23] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_262 
+ gnd vdd predecode_29[0] predecode_117[24] decode_b[24] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_263 
+ gnd vdd decode_b[24] decode[24] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_264 
+ gnd vdd predecode_29[0] predecode_117[25] decode_b[25] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_265 
+ gnd vdd decode_b[25] decode[25] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_266 
+ gnd vdd predecode_29[0] predecode_117[26] decode_b[26] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_267 
+ gnd vdd decode_b[26] decode[26] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_268 
+ gnd vdd predecode_29[0] predecode_117[27] decode_b[27] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_269 
+ gnd vdd decode_b[27] decode[27] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_270 
+ gnd vdd predecode_29[0] predecode_117[28] decode_b[28] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_271 
+ gnd vdd decode_b[28] decode[28] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_272 
+ gnd vdd predecode_29[0] predecode_117[29] decode_b[29] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_273 
+ gnd vdd decode_b[29] decode[29] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_274 
+ gnd vdd predecode_29[0] predecode_117[30] decode_b[30] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_275 
+ gnd vdd decode_b[30] decode[30] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_276 
+ gnd vdd predecode_29[0] predecode_117[31] decode_b[31] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_277 
+ gnd vdd decode_b[31] decode[31] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_278 
+ gnd vdd predecode_29[1] predecode_117[0] decode_b[32] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_279 
+ gnd vdd decode_b[32] decode[32] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_280 
+ gnd vdd predecode_29[1] predecode_117[1] decode_b[33] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_281 
+ gnd vdd decode_b[33] decode[33] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_282 
+ gnd vdd predecode_29[1] predecode_117[2] decode_b[34] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_283 
+ gnd vdd decode_b[34] decode[34] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_284 
+ gnd vdd predecode_29[1] predecode_117[3] decode_b[35] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_285 
+ gnd vdd decode_b[35] decode[35] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_286 
+ gnd vdd predecode_29[1] predecode_117[4] decode_b[36] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_287 
+ gnd vdd decode_b[36] decode[36] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_288 
+ gnd vdd predecode_29[1] predecode_117[5] decode_b[37] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_289 
+ gnd vdd decode_b[37] decode[37] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_290 
+ gnd vdd predecode_29[1] predecode_117[6] decode_b[38] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_291 
+ gnd vdd decode_b[38] decode[38] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_292 
+ gnd vdd predecode_29[1] predecode_117[7] decode_b[39] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_293 
+ gnd vdd decode_b[39] decode[39] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_294 
+ gnd vdd predecode_29[1] predecode_117[8] decode_b[40] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_295 
+ gnd vdd decode_b[40] decode[40] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_296 
+ gnd vdd predecode_29[1] predecode_117[9] decode_b[41] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_297 
+ gnd vdd decode_b[41] decode[41] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_298 
+ gnd vdd predecode_29[1] predecode_117[10] decode_b[42] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_299 
+ gnd vdd decode_b[42] decode[42] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_300 
+ gnd vdd predecode_29[1] predecode_117[11] decode_b[43] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_301 
+ gnd vdd decode_b[43] decode[43] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_302 
+ gnd vdd predecode_29[1] predecode_117[12] decode_b[44] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_303 
+ gnd vdd decode_b[44] decode[44] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_304 
+ gnd vdd predecode_29[1] predecode_117[13] decode_b[45] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_305 
+ gnd vdd decode_b[45] decode[45] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_306 
+ gnd vdd predecode_29[1] predecode_117[14] decode_b[46] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_307 
+ gnd vdd decode_b[46] decode[46] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_308 
+ gnd vdd predecode_29[1] predecode_117[15] decode_b[47] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_309 
+ gnd vdd decode_b[47] decode[47] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_310 
+ gnd vdd predecode_29[1] predecode_117[16] decode_b[48] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_311 
+ gnd vdd decode_b[48] decode[48] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_312 
+ gnd vdd predecode_29[1] predecode_117[17] decode_b[49] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_313 
+ gnd vdd decode_b[49] decode[49] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_314 
+ gnd vdd predecode_29[1] predecode_117[18] decode_b[50] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_315 
+ gnd vdd decode_b[50] decode[50] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_316 
+ gnd vdd predecode_29[1] predecode_117[19] decode_b[51] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_317 
+ gnd vdd decode_b[51] decode[51] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_318 
+ gnd vdd predecode_29[1] predecode_117[20] decode_b[52] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_319 
+ gnd vdd decode_b[52] decode[52] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_320 
+ gnd vdd predecode_29[1] predecode_117[21] decode_b[53] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_321 
+ gnd vdd decode_b[53] decode[53] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_322 
+ gnd vdd predecode_29[1] predecode_117[22] decode_b[54] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_323 
+ gnd vdd decode_b[54] decode[54] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_324 
+ gnd vdd predecode_29[1] predecode_117[23] decode_b[55] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_325 
+ gnd vdd decode_b[55] decode[55] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_326 
+ gnd vdd predecode_29[1] predecode_117[24] decode_b[56] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_327 
+ gnd vdd decode_b[56] decode[56] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_328 
+ gnd vdd predecode_29[1] predecode_117[25] decode_b[57] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_329 
+ gnd vdd decode_b[57] decode[57] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_330 
+ gnd vdd predecode_29[1] predecode_117[26] decode_b[58] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_331 
+ gnd vdd decode_b[58] decode[58] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_332 
+ gnd vdd predecode_29[1] predecode_117[27] decode_b[59] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_333 
+ gnd vdd decode_b[59] decode[59] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_334 
+ gnd vdd predecode_29[1] predecode_117[28] decode_b[60] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_335 
+ gnd vdd decode_b[60] decode[60] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_336 
+ gnd vdd predecode_29[1] predecode_117[29] decode_b[61] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_337 
+ gnd vdd decode_b[61] decode[61] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_338 
+ gnd vdd predecode_29[1] predecode_117[30] decode_b[62] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_339 
+ gnd vdd decode_b[62] decode[62] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_340 
+ gnd vdd predecode_29[1] predecode_117[31] decode_b[63] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_341 
+ gnd vdd decode_b[63] decode[63] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_342 
+ gnd vdd predecode_29[2] predecode_117[0] decode_b[64] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_343 
+ gnd vdd decode_b[64] decode[64] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_344 
+ gnd vdd predecode_29[2] predecode_117[1] decode_b[65] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_345 
+ gnd vdd decode_b[65] decode[65] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_346 
+ gnd vdd predecode_29[2] predecode_117[2] decode_b[66] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_347 
+ gnd vdd decode_b[66] decode[66] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_348 
+ gnd vdd predecode_29[2] predecode_117[3] decode_b[67] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_349 
+ gnd vdd decode_b[67] decode[67] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_350 
+ gnd vdd predecode_29[2] predecode_117[4] decode_b[68] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_351 
+ gnd vdd decode_b[68] decode[68] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_352 
+ gnd vdd predecode_29[2] predecode_117[5] decode_b[69] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_353 
+ gnd vdd decode_b[69] decode[69] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_354 
+ gnd vdd predecode_29[2] predecode_117[6] decode_b[70] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_355 
+ gnd vdd decode_b[70] decode[70] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_356 
+ gnd vdd predecode_29[2] predecode_117[7] decode_b[71] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_357 
+ gnd vdd decode_b[71] decode[71] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_358 
+ gnd vdd predecode_29[2] predecode_117[8] decode_b[72] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_359 
+ gnd vdd decode_b[72] decode[72] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_360 
+ gnd vdd predecode_29[2] predecode_117[9] decode_b[73] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_361 
+ gnd vdd decode_b[73] decode[73] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_362 
+ gnd vdd predecode_29[2] predecode_117[10] decode_b[74] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_363 
+ gnd vdd decode_b[74] decode[74] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_364 
+ gnd vdd predecode_29[2] predecode_117[11] decode_b[75] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_365 
+ gnd vdd decode_b[75] decode[75] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_366 
+ gnd vdd predecode_29[2] predecode_117[12] decode_b[76] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_367 
+ gnd vdd decode_b[76] decode[76] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_368 
+ gnd vdd predecode_29[2] predecode_117[13] decode_b[77] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_369 
+ gnd vdd decode_b[77] decode[77] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_370 
+ gnd vdd predecode_29[2] predecode_117[14] decode_b[78] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_371 
+ gnd vdd decode_b[78] decode[78] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_372 
+ gnd vdd predecode_29[2] predecode_117[15] decode_b[79] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_373 
+ gnd vdd decode_b[79] decode[79] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_374 
+ gnd vdd predecode_29[2] predecode_117[16] decode_b[80] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_375 
+ gnd vdd decode_b[80] decode[80] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_376 
+ gnd vdd predecode_29[2] predecode_117[17] decode_b[81] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_377 
+ gnd vdd decode_b[81] decode[81] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_378 
+ gnd vdd predecode_29[2] predecode_117[18] decode_b[82] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_379 
+ gnd vdd decode_b[82] decode[82] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_380 
+ gnd vdd predecode_29[2] predecode_117[19] decode_b[83] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_381 
+ gnd vdd decode_b[83] decode[83] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_382 
+ gnd vdd predecode_29[2] predecode_117[20] decode_b[84] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_383 
+ gnd vdd decode_b[84] decode[84] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_384 
+ gnd vdd predecode_29[2] predecode_117[21] decode_b[85] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_385 
+ gnd vdd decode_b[85] decode[85] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_386 
+ gnd vdd predecode_29[2] predecode_117[22] decode_b[86] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_387 
+ gnd vdd decode_b[86] decode[86] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_388 
+ gnd vdd predecode_29[2] predecode_117[23] decode_b[87] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_389 
+ gnd vdd decode_b[87] decode[87] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_390 
+ gnd vdd predecode_29[2] predecode_117[24] decode_b[88] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_391 
+ gnd vdd decode_b[88] decode[88] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_392 
+ gnd vdd predecode_29[2] predecode_117[25] decode_b[89] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_393 
+ gnd vdd decode_b[89] decode[89] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_394 
+ gnd vdd predecode_29[2] predecode_117[26] decode_b[90] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_395 
+ gnd vdd decode_b[90] decode[90] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_396 
+ gnd vdd predecode_29[2] predecode_117[27] decode_b[91] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_397 
+ gnd vdd decode_b[91] decode[91] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_398 
+ gnd vdd predecode_29[2] predecode_117[28] decode_b[92] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_399 
+ gnd vdd decode_b[92] decode[92] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_400 
+ gnd vdd predecode_29[2] predecode_117[29] decode_b[93] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_401 
+ gnd vdd decode_b[93] decode[93] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_402 
+ gnd vdd predecode_29[2] predecode_117[30] decode_b[94] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_403 
+ gnd vdd decode_b[94] decode[94] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_404 
+ gnd vdd predecode_29[2] predecode_117[31] decode_b[95] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_405 
+ gnd vdd decode_b[95] decode[95] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_406 
+ gnd vdd predecode_29[3] predecode_117[0] decode_b[96] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_407 
+ gnd vdd decode_b[96] decode[96] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_408 
+ gnd vdd predecode_29[3] predecode_117[1] decode_b[97] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_409 
+ gnd vdd decode_b[97] decode[97] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_410 
+ gnd vdd predecode_29[3] predecode_117[2] decode_b[98] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_411 
+ gnd vdd decode_b[98] decode[98] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_412 
+ gnd vdd predecode_29[3] predecode_117[3] decode_b[99] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_413 
+ gnd vdd decode_b[99] decode[99] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_414 
+ gnd vdd predecode_29[3] predecode_117[4] decode_b[100] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_415 
+ gnd vdd decode_b[100] decode[100] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_416 
+ gnd vdd predecode_29[3] predecode_117[5] decode_b[101] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_417 
+ gnd vdd decode_b[101] decode[101] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_418 
+ gnd vdd predecode_29[3] predecode_117[6] decode_b[102] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_419 
+ gnd vdd decode_b[102] decode[102] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_420 
+ gnd vdd predecode_29[3] predecode_117[7] decode_b[103] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_421 
+ gnd vdd decode_b[103] decode[103] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_422 
+ gnd vdd predecode_29[3] predecode_117[8] decode_b[104] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_423 
+ gnd vdd decode_b[104] decode[104] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_424 
+ gnd vdd predecode_29[3] predecode_117[9] decode_b[105] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_425 
+ gnd vdd decode_b[105] decode[105] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_426 
+ gnd vdd predecode_29[3] predecode_117[10] decode_b[106] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_427 
+ gnd vdd decode_b[106] decode[106] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_428 
+ gnd vdd predecode_29[3] predecode_117[11] decode_b[107] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_429 
+ gnd vdd decode_b[107] decode[107] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_430 
+ gnd vdd predecode_29[3] predecode_117[12] decode_b[108] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_431 
+ gnd vdd decode_b[108] decode[108] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_432 
+ gnd vdd predecode_29[3] predecode_117[13] decode_b[109] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_433 
+ gnd vdd decode_b[109] decode[109] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_434 
+ gnd vdd predecode_29[3] predecode_117[14] decode_b[110] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_435 
+ gnd vdd decode_b[110] decode[110] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_436 
+ gnd vdd predecode_29[3] predecode_117[15] decode_b[111] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_437 
+ gnd vdd decode_b[111] decode[111] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_438 
+ gnd vdd predecode_29[3] predecode_117[16] decode_b[112] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_439 
+ gnd vdd decode_b[112] decode[112] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_440 
+ gnd vdd predecode_29[3] predecode_117[17] decode_b[113] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_441 
+ gnd vdd decode_b[113] decode[113] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_442 
+ gnd vdd predecode_29[3] predecode_117[18] decode_b[114] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_443 
+ gnd vdd decode_b[114] decode[114] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_444 
+ gnd vdd predecode_29[3] predecode_117[19] decode_b[115] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_445 
+ gnd vdd decode_b[115] decode[115] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_446 
+ gnd vdd predecode_29[3] predecode_117[20] decode_b[116] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_447 
+ gnd vdd decode_b[116] decode[116] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_448 
+ gnd vdd predecode_29[3] predecode_117[21] decode_b[117] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_449 
+ gnd vdd decode_b[117] decode[117] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_450 
+ gnd vdd predecode_29[3] predecode_117[22] decode_b[118] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_451 
+ gnd vdd decode_b[118] decode[118] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_452 
+ gnd vdd predecode_29[3] predecode_117[23] decode_b[119] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_453 
+ gnd vdd decode_b[119] decode[119] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_454 
+ gnd vdd predecode_29[3] predecode_117[24] decode_b[120] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_455 
+ gnd vdd decode_b[120] decode[120] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_456 
+ gnd vdd predecode_29[3] predecode_117[25] decode_b[121] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_457 
+ gnd vdd decode_b[121] decode[121] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_458 
+ gnd vdd predecode_29[3] predecode_117[26] decode_b[122] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_459 
+ gnd vdd decode_b[122] decode[122] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_460 
+ gnd vdd predecode_29[3] predecode_117[27] decode_b[123] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_461 
+ gnd vdd decode_b[123] decode[123] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_462 
+ gnd vdd predecode_29[3] predecode_117[28] decode_b[124] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_463 
+ gnd vdd decode_b[124] decode[124] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_464 
+ gnd vdd predecode_29[3] predecode_117[29] decode_b[125] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_465 
+ gnd vdd decode_b[125] decode[125] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_466 
+ gnd vdd predecode_29[3] predecode_117[30] decode_b[126] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_467 
+ gnd vdd decode_b[126] decode[126] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_468 
+ gnd vdd predecode_29[3] predecode_117[31] decode_b[127] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_469 
+ gnd vdd decode_b[127] decode[127] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_470 
+ gnd vdd predecode_29[4] predecode_117[0] decode_b[128] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_471 
+ gnd vdd decode_b[128] decode[128] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_472 
+ gnd vdd predecode_29[4] predecode_117[1] decode_b[129] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_473 
+ gnd vdd decode_b[129] decode[129] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_474 
+ gnd vdd predecode_29[4] predecode_117[2] decode_b[130] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_475 
+ gnd vdd decode_b[130] decode[130] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_476 
+ gnd vdd predecode_29[4] predecode_117[3] decode_b[131] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_477 
+ gnd vdd decode_b[131] decode[131] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_478 
+ gnd vdd predecode_29[4] predecode_117[4] decode_b[132] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_479 
+ gnd vdd decode_b[132] decode[132] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_480 
+ gnd vdd predecode_29[4] predecode_117[5] decode_b[133] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_481 
+ gnd vdd decode_b[133] decode[133] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_482 
+ gnd vdd predecode_29[4] predecode_117[6] decode_b[134] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_483 
+ gnd vdd decode_b[134] decode[134] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_484 
+ gnd vdd predecode_29[4] predecode_117[7] decode_b[135] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_485 
+ gnd vdd decode_b[135] decode[135] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_486 
+ gnd vdd predecode_29[4] predecode_117[8] decode_b[136] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_487 
+ gnd vdd decode_b[136] decode[136] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_488 
+ gnd vdd predecode_29[4] predecode_117[9] decode_b[137] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_489 
+ gnd vdd decode_b[137] decode[137] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_490 
+ gnd vdd predecode_29[4] predecode_117[10] decode_b[138] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_491 
+ gnd vdd decode_b[138] decode[138] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_492 
+ gnd vdd predecode_29[4] predecode_117[11] decode_b[139] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_493 
+ gnd vdd decode_b[139] decode[139] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_494 
+ gnd vdd predecode_29[4] predecode_117[12] decode_b[140] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_495 
+ gnd vdd decode_b[140] decode[140] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_496 
+ gnd vdd predecode_29[4] predecode_117[13] decode_b[141] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_497 
+ gnd vdd decode_b[141] decode[141] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_498 
+ gnd vdd predecode_29[4] predecode_117[14] decode_b[142] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_499 
+ gnd vdd decode_b[142] decode[142] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_500 
+ gnd vdd predecode_29[4] predecode_117[15] decode_b[143] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_501 
+ gnd vdd decode_b[143] decode[143] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_502 
+ gnd vdd predecode_29[4] predecode_117[16] decode_b[144] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_503 
+ gnd vdd decode_b[144] decode[144] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_504 
+ gnd vdd predecode_29[4] predecode_117[17] decode_b[145] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_505 
+ gnd vdd decode_b[145] decode[145] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_506 
+ gnd vdd predecode_29[4] predecode_117[18] decode_b[146] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_507 
+ gnd vdd decode_b[146] decode[146] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_508 
+ gnd vdd predecode_29[4] predecode_117[19] decode_b[147] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_509 
+ gnd vdd decode_b[147] decode[147] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_510 
+ gnd vdd predecode_29[4] predecode_117[20] decode_b[148] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_511 
+ gnd vdd decode_b[148] decode[148] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_512 
+ gnd vdd predecode_29[4] predecode_117[21] decode_b[149] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_513 
+ gnd vdd decode_b[149] decode[149] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_514 
+ gnd vdd predecode_29[4] predecode_117[22] decode_b[150] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_515 
+ gnd vdd decode_b[150] decode[150] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_516 
+ gnd vdd predecode_29[4] predecode_117[23] decode_b[151] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_517 
+ gnd vdd decode_b[151] decode[151] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_518 
+ gnd vdd predecode_29[4] predecode_117[24] decode_b[152] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_519 
+ gnd vdd decode_b[152] decode[152] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_520 
+ gnd vdd predecode_29[4] predecode_117[25] decode_b[153] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_521 
+ gnd vdd decode_b[153] decode[153] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_522 
+ gnd vdd predecode_29[4] predecode_117[26] decode_b[154] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_523 
+ gnd vdd decode_b[154] decode[154] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_524 
+ gnd vdd predecode_29[4] predecode_117[27] decode_b[155] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_525 
+ gnd vdd decode_b[155] decode[155] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_526 
+ gnd vdd predecode_29[4] predecode_117[28] decode_b[156] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_527 
+ gnd vdd decode_b[156] decode[156] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_528 
+ gnd vdd predecode_29[4] predecode_117[29] decode_b[157] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_529 
+ gnd vdd decode_b[157] decode[157] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_530 
+ gnd vdd predecode_29[4] predecode_117[30] decode_b[158] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_531 
+ gnd vdd decode_b[158] decode[158] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_532 
+ gnd vdd predecode_29[4] predecode_117[31] decode_b[159] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_533 
+ gnd vdd decode_b[159] decode[159] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_534 
+ gnd vdd predecode_29[5] predecode_117[0] decode_b[160] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_535 
+ gnd vdd decode_b[160] decode[160] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_536 
+ gnd vdd predecode_29[5] predecode_117[1] decode_b[161] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_537 
+ gnd vdd decode_b[161] decode[161] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_538 
+ gnd vdd predecode_29[5] predecode_117[2] decode_b[162] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_539 
+ gnd vdd decode_b[162] decode[162] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_540 
+ gnd vdd predecode_29[5] predecode_117[3] decode_b[163] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_541 
+ gnd vdd decode_b[163] decode[163] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_542 
+ gnd vdd predecode_29[5] predecode_117[4] decode_b[164] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_543 
+ gnd vdd decode_b[164] decode[164] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_544 
+ gnd vdd predecode_29[5] predecode_117[5] decode_b[165] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_545 
+ gnd vdd decode_b[165] decode[165] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_546 
+ gnd vdd predecode_29[5] predecode_117[6] decode_b[166] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_547 
+ gnd vdd decode_b[166] decode[166] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_548 
+ gnd vdd predecode_29[5] predecode_117[7] decode_b[167] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_549 
+ gnd vdd decode_b[167] decode[167] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_550 
+ gnd vdd predecode_29[5] predecode_117[8] decode_b[168] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_551 
+ gnd vdd decode_b[168] decode[168] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_552 
+ gnd vdd predecode_29[5] predecode_117[9] decode_b[169] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_553 
+ gnd vdd decode_b[169] decode[169] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_554 
+ gnd vdd predecode_29[5] predecode_117[10] decode_b[170] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_555 
+ gnd vdd decode_b[170] decode[170] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_556 
+ gnd vdd predecode_29[5] predecode_117[11] decode_b[171] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_557 
+ gnd vdd decode_b[171] decode[171] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_558 
+ gnd vdd predecode_29[5] predecode_117[12] decode_b[172] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_559 
+ gnd vdd decode_b[172] decode[172] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_560 
+ gnd vdd predecode_29[5] predecode_117[13] decode_b[173] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_561 
+ gnd vdd decode_b[173] decode[173] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_562 
+ gnd vdd predecode_29[5] predecode_117[14] decode_b[174] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_563 
+ gnd vdd decode_b[174] decode[174] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_564 
+ gnd vdd predecode_29[5] predecode_117[15] decode_b[175] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_565 
+ gnd vdd decode_b[175] decode[175] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_566 
+ gnd vdd predecode_29[5] predecode_117[16] decode_b[176] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_567 
+ gnd vdd decode_b[176] decode[176] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_568 
+ gnd vdd predecode_29[5] predecode_117[17] decode_b[177] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_569 
+ gnd vdd decode_b[177] decode[177] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_570 
+ gnd vdd predecode_29[5] predecode_117[18] decode_b[178] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_571 
+ gnd vdd decode_b[178] decode[178] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_572 
+ gnd vdd predecode_29[5] predecode_117[19] decode_b[179] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_573 
+ gnd vdd decode_b[179] decode[179] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_574 
+ gnd vdd predecode_29[5] predecode_117[20] decode_b[180] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_575 
+ gnd vdd decode_b[180] decode[180] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_576 
+ gnd vdd predecode_29[5] predecode_117[21] decode_b[181] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_577 
+ gnd vdd decode_b[181] decode[181] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_578 
+ gnd vdd predecode_29[5] predecode_117[22] decode_b[182] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_579 
+ gnd vdd decode_b[182] decode[182] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_580 
+ gnd vdd predecode_29[5] predecode_117[23] decode_b[183] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_581 
+ gnd vdd decode_b[183] decode[183] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_582 
+ gnd vdd predecode_29[5] predecode_117[24] decode_b[184] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_583 
+ gnd vdd decode_b[184] decode[184] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_584 
+ gnd vdd predecode_29[5] predecode_117[25] decode_b[185] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_585 
+ gnd vdd decode_b[185] decode[185] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_586 
+ gnd vdd predecode_29[5] predecode_117[26] decode_b[186] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_587 
+ gnd vdd decode_b[186] decode[186] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_588 
+ gnd vdd predecode_29[5] predecode_117[27] decode_b[187] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_589 
+ gnd vdd decode_b[187] decode[187] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_590 
+ gnd vdd predecode_29[5] predecode_117[28] decode_b[188] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_591 
+ gnd vdd decode_b[188] decode[188] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_592 
+ gnd vdd predecode_29[5] predecode_117[29] decode_b[189] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_593 
+ gnd vdd decode_b[189] decode[189] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_594 
+ gnd vdd predecode_29[5] predecode_117[30] decode_b[190] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_595 
+ gnd vdd decode_b[190] decode[190] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_596 
+ gnd vdd predecode_29[5] predecode_117[31] decode_b[191] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_597 
+ gnd vdd decode_b[191] decode[191] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_598 
+ gnd vdd predecode_29[6] predecode_117[0] decode_b[192] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_599 
+ gnd vdd decode_b[192] decode[192] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_600 
+ gnd vdd predecode_29[6] predecode_117[1] decode_b[193] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_601 
+ gnd vdd decode_b[193] decode[193] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_602 
+ gnd vdd predecode_29[6] predecode_117[2] decode_b[194] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_603 
+ gnd vdd decode_b[194] decode[194] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_604 
+ gnd vdd predecode_29[6] predecode_117[3] decode_b[195] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_605 
+ gnd vdd decode_b[195] decode[195] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_606 
+ gnd vdd predecode_29[6] predecode_117[4] decode_b[196] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_607 
+ gnd vdd decode_b[196] decode[196] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_608 
+ gnd vdd predecode_29[6] predecode_117[5] decode_b[197] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_609 
+ gnd vdd decode_b[197] decode[197] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_610 
+ gnd vdd predecode_29[6] predecode_117[6] decode_b[198] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_611 
+ gnd vdd decode_b[198] decode[198] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_612 
+ gnd vdd predecode_29[6] predecode_117[7] decode_b[199] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_613 
+ gnd vdd decode_b[199] decode[199] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_614 
+ gnd vdd predecode_29[6] predecode_117[8] decode_b[200] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_615 
+ gnd vdd decode_b[200] decode[200] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_616 
+ gnd vdd predecode_29[6] predecode_117[9] decode_b[201] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_617 
+ gnd vdd decode_b[201] decode[201] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_618 
+ gnd vdd predecode_29[6] predecode_117[10] decode_b[202] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_619 
+ gnd vdd decode_b[202] decode[202] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_620 
+ gnd vdd predecode_29[6] predecode_117[11] decode_b[203] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_621 
+ gnd vdd decode_b[203] decode[203] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_622 
+ gnd vdd predecode_29[6] predecode_117[12] decode_b[204] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_623 
+ gnd vdd decode_b[204] decode[204] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_624 
+ gnd vdd predecode_29[6] predecode_117[13] decode_b[205] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_625 
+ gnd vdd decode_b[205] decode[205] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_626 
+ gnd vdd predecode_29[6] predecode_117[14] decode_b[206] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_627 
+ gnd vdd decode_b[206] decode[206] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_628 
+ gnd vdd predecode_29[6] predecode_117[15] decode_b[207] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_629 
+ gnd vdd decode_b[207] decode[207] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_630 
+ gnd vdd predecode_29[6] predecode_117[16] decode_b[208] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_631 
+ gnd vdd decode_b[208] decode[208] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_632 
+ gnd vdd predecode_29[6] predecode_117[17] decode_b[209] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_633 
+ gnd vdd decode_b[209] decode[209] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_634 
+ gnd vdd predecode_29[6] predecode_117[18] decode_b[210] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_635 
+ gnd vdd decode_b[210] decode[210] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_636 
+ gnd vdd predecode_29[6] predecode_117[19] decode_b[211] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_637 
+ gnd vdd decode_b[211] decode[211] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_638 
+ gnd vdd predecode_29[6] predecode_117[20] decode_b[212] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_639 
+ gnd vdd decode_b[212] decode[212] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_640 
+ gnd vdd predecode_29[6] predecode_117[21] decode_b[213] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_641 
+ gnd vdd decode_b[213] decode[213] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_642 
+ gnd vdd predecode_29[6] predecode_117[22] decode_b[214] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_643 
+ gnd vdd decode_b[214] decode[214] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_644 
+ gnd vdd predecode_29[6] predecode_117[23] decode_b[215] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_645 
+ gnd vdd decode_b[215] decode[215] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_646 
+ gnd vdd predecode_29[6] predecode_117[24] decode_b[216] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_647 
+ gnd vdd decode_b[216] decode[216] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_648 
+ gnd vdd predecode_29[6] predecode_117[25] decode_b[217] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_649 
+ gnd vdd decode_b[217] decode[217] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_650 
+ gnd vdd predecode_29[6] predecode_117[26] decode_b[218] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_651 
+ gnd vdd decode_b[218] decode[218] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_652 
+ gnd vdd predecode_29[6] predecode_117[27] decode_b[219] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_653 
+ gnd vdd decode_b[219] decode[219] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_654 
+ gnd vdd predecode_29[6] predecode_117[28] decode_b[220] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_655 
+ gnd vdd decode_b[220] decode[220] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_656 
+ gnd vdd predecode_29[6] predecode_117[29] decode_b[221] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_657 
+ gnd vdd decode_b[221] decode[221] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_658 
+ gnd vdd predecode_29[6] predecode_117[30] decode_b[222] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_659 
+ gnd vdd decode_b[222] decode[222] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_660 
+ gnd vdd predecode_29[6] predecode_117[31] decode_b[223] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_661 
+ gnd vdd decode_b[223] decode[223] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_662 
+ gnd vdd predecode_29[7] predecode_117[0] decode_b[224] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_663 
+ gnd vdd decode_b[224] decode[224] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_664 
+ gnd vdd predecode_29[7] predecode_117[1] decode_b[225] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_665 
+ gnd vdd decode_b[225] decode[225] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_666 
+ gnd vdd predecode_29[7] predecode_117[2] decode_b[226] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_667 
+ gnd vdd decode_b[226] decode[226] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_668 
+ gnd vdd predecode_29[7] predecode_117[3] decode_b[227] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_669 
+ gnd vdd decode_b[227] decode[227] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_670 
+ gnd vdd predecode_29[7] predecode_117[4] decode_b[228] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_671 
+ gnd vdd decode_b[228] decode[228] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_672 
+ gnd vdd predecode_29[7] predecode_117[5] decode_b[229] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_673 
+ gnd vdd decode_b[229] decode[229] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_674 
+ gnd vdd predecode_29[7] predecode_117[6] decode_b[230] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_675 
+ gnd vdd decode_b[230] decode[230] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_676 
+ gnd vdd predecode_29[7] predecode_117[7] decode_b[231] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_677 
+ gnd vdd decode_b[231] decode[231] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_678 
+ gnd vdd predecode_29[7] predecode_117[8] decode_b[232] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_679 
+ gnd vdd decode_b[232] decode[232] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_680 
+ gnd vdd predecode_29[7] predecode_117[9] decode_b[233] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_681 
+ gnd vdd decode_b[233] decode[233] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_682 
+ gnd vdd predecode_29[7] predecode_117[10] decode_b[234] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_683 
+ gnd vdd decode_b[234] decode[234] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_684 
+ gnd vdd predecode_29[7] predecode_117[11] decode_b[235] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_685 
+ gnd vdd decode_b[235] decode[235] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_686 
+ gnd vdd predecode_29[7] predecode_117[12] decode_b[236] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_687 
+ gnd vdd decode_b[236] decode[236] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_688 
+ gnd vdd predecode_29[7] predecode_117[13] decode_b[237] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_689 
+ gnd vdd decode_b[237] decode[237] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_690 
+ gnd vdd predecode_29[7] predecode_117[14] decode_b[238] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_691 
+ gnd vdd decode_b[238] decode[238] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_692 
+ gnd vdd predecode_29[7] predecode_117[15] decode_b[239] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_693 
+ gnd vdd decode_b[239] decode[239] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_694 
+ gnd vdd predecode_29[7] predecode_117[16] decode_b[240] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_695 
+ gnd vdd decode_b[240] decode[240] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_696 
+ gnd vdd predecode_29[7] predecode_117[17] decode_b[241] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_697 
+ gnd vdd decode_b[241] decode[241] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_698 
+ gnd vdd predecode_29[7] predecode_117[18] decode_b[242] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_699 
+ gnd vdd decode_b[242] decode[242] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_700 
+ gnd vdd predecode_29[7] predecode_117[19] decode_b[243] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_701 
+ gnd vdd decode_b[243] decode[243] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_702 
+ gnd vdd predecode_29[7] predecode_117[20] decode_b[244] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_703 
+ gnd vdd decode_b[244] decode[244] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_704 
+ gnd vdd predecode_29[7] predecode_117[21] decode_b[245] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_705 
+ gnd vdd decode_b[245] decode[245] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_706 
+ gnd vdd predecode_29[7] predecode_117[22] decode_b[246] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_707 
+ gnd vdd decode_b[246] decode[246] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_708 
+ gnd vdd predecode_29[7] predecode_117[23] decode_b[247] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_709 
+ gnd vdd decode_b[247] decode[247] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_710 
+ gnd vdd predecode_29[7] predecode_117[24] decode_b[248] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_711 
+ gnd vdd decode_b[248] decode[248] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_712 
+ gnd vdd predecode_29[7] predecode_117[25] decode_b[249] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_713 
+ gnd vdd decode_b[249] decode[249] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_714 
+ gnd vdd predecode_29[7] predecode_117[26] decode_b[250] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_715 
+ gnd vdd decode_b[250] decode[250] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_716 
+ gnd vdd predecode_29[7] predecode_117[27] decode_b[251] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_717 
+ gnd vdd decode_b[251] decode[251] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_718 
+ gnd vdd predecode_29[7] predecode_117[28] decode_b[252] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_719 
+ gnd vdd decode_b[252] decode[252] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_720 
+ gnd vdd predecode_29[7] predecode_117[29] decode_b[253] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_721 
+ gnd vdd decode_b[253] decode[253] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_722 
+ gnd vdd predecode_29[7] predecode_117[30] decode_b[254] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_723 
+ gnd vdd decode_b[254] decode[254] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_724 
+ gnd vdd predecode_29[7] predecode_117[31] decode_b[255] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_725 
+ gnd vdd decode_b[255] decode[255] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_726 
+ gnd vdd predecode_29[8] predecode_117[0] decode_b[256] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_727 
+ gnd vdd decode_b[256] decode[256] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_728 
+ gnd vdd predecode_29[8] predecode_117[1] decode_b[257] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_729 
+ gnd vdd decode_b[257] decode[257] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_730 
+ gnd vdd predecode_29[8] predecode_117[2] decode_b[258] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_731 
+ gnd vdd decode_b[258] decode[258] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_732 
+ gnd vdd predecode_29[8] predecode_117[3] decode_b[259] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_733 
+ gnd vdd decode_b[259] decode[259] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_734 
+ gnd vdd predecode_29[8] predecode_117[4] decode_b[260] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_735 
+ gnd vdd decode_b[260] decode[260] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_736 
+ gnd vdd predecode_29[8] predecode_117[5] decode_b[261] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_737 
+ gnd vdd decode_b[261] decode[261] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_738 
+ gnd vdd predecode_29[8] predecode_117[6] decode_b[262] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_739 
+ gnd vdd decode_b[262] decode[262] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_740 
+ gnd vdd predecode_29[8] predecode_117[7] decode_b[263] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_741 
+ gnd vdd decode_b[263] decode[263] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_742 
+ gnd vdd predecode_29[8] predecode_117[8] decode_b[264] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_743 
+ gnd vdd decode_b[264] decode[264] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_744 
+ gnd vdd predecode_29[8] predecode_117[9] decode_b[265] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_745 
+ gnd vdd decode_b[265] decode[265] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_746 
+ gnd vdd predecode_29[8] predecode_117[10] decode_b[266] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_747 
+ gnd vdd decode_b[266] decode[266] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_748 
+ gnd vdd predecode_29[8] predecode_117[11] decode_b[267] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_749 
+ gnd vdd decode_b[267] decode[267] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_750 
+ gnd vdd predecode_29[8] predecode_117[12] decode_b[268] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_751 
+ gnd vdd decode_b[268] decode[268] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_752 
+ gnd vdd predecode_29[8] predecode_117[13] decode_b[269] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_753 
+ gnd vdd decode_b[269] decode[269] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_754 
+ gnd vdd predecode_29[8] predecode_117[14] decode_b[270] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_755 
+ gnd vdd decode_b[270] decode[270] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_756 
+ gnd vdd predecode_29[8] predecode_117[15] decode_b[271] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_757 
+ gnd vdd decode_b[271] decode[271] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_758 
+ gnd vdd predecode_29[8] predecode_117[16] decode_b[272] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_759 
+ gnd vdd decode_b[272] decode[272] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_760 
+ gnd vdd predecode_29[8] predecode_117[17] decode_b[273] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_761 
+ gnd vdd decode_b[273] decode[273] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_762 
+ gnd vdd predecode_29[8] predecode_117[18] decode_b[274] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_763 
+ gnd vdd decode_b[274] decode[274] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_764 
+ gnd vdd predecode_29[8] predecode_117[19] decode_b[275] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_765 
+ gnd vdd decode_b[275] decode[275] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_766 
+ gnd vdd predecode_29[8] predecode_117[20] decode_b[276] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_767 
+ gnd vdd decode_b[276] decode[276] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_768 
+ gnd vdd predecode_29[8] predecode_117[21] decode_b[277] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_769 
+ gnd vdd decode_b[277] decode[277] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_770 
+ gnd vdd predecode_29[8] predecode_117[22] decode_b[278] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_771 
+ gnd vdd decode_b[278] decode[278] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_772 
+ gnd vdd predecode_29[8] predecode_117[23] decode_b[279] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_773 
+ gnd vdd decode_b[279] decode[279] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_774 
+ gnd vdd predecode_29[8] predecode_117[24] decode_b[280] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_775 
+ gnd vdd decode_b[280] decode[280] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_776 
+ gnd vdd predecode_29[8] predecode_117[25] decode_b[281] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_777 
+ gnd vdd decode_b[281] decode[281] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_778 
+ gnd vdd predecode_29[8] predecode_117[26] decode_b[282] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_779 
+ gnd vdd decode_b[282] decode[282] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_780 
+ gnd vdd predecode_29[8] predecode_117[27] decode_b[283] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_781 
+ gnd vdd decode_b[283] decode[283] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_782 
+ gnd vdd predecode_29[8] predecode_117[28] decode_b[284] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_783 
+ gnd vdd decode_b[284] decode[284] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_784 
+ gnd vdd predecode_29[8] predecode_117[29] decode_b[285] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_785 
+ gnd vdd decode_b[285] decode[285] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_786 
+ gnd vdd predecode_29[8] predecode_117[30] decode_b[286] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_787 
+ gnd vdd decode_b[286] decode[286] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_788 
+ gnd vdd predecode_29[8] predecode_117[31] decode_b[287] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_789 
+ gnd vdd decode_b[287] decode[287] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_790 
+ gnd vdd predecode_29[9] predecode_117[0] decode_b[288] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_791 
+ gnd vdd decode_b[288] decode[288] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_792 
+ gnd vdd predecode_29[9] predecode_117[1] decode_b[289] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_793 
+ gnd vdd decode_b[289] decode[289] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_794 
+ gnd vdd predecode_29[9] predecode_117[2] decode_b[290] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_795 
+ gnd vdd decode_b[290] decode[290] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_796 
+ gnd vdd predecode_29[9] predecode_117[3] decode_b[291] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_797 
+ gnd vdd decode_b[291] decode[291] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_798 
+ gnd vdd predecode_29[9] predecode_117[4] decode_b[292] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_799 
+ gnd vdd decode_b[292] decode[292] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_800 
+ gnd vdd predecode_29[9] predecode_117[5] decode_b[293] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_801 
+ gnd vdd decode_b[293] decode[293] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_802 
+ gnd vdd predecode_29[9] predecode_117[6] decode_b[294] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_803 
+ gnd vdd decode_b[294] decode[294] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_804 
+ gnd vdd predecode_29[9] predecode_117[7] decode_b[295] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_805 
+ gnd vdd decode_b[295] decode[295] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_806 
+ gnd vdd predecode_29[9] predecode_117[8] decode_b[296] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_807 
+ gnd vdd decode_b[296] decode[296] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_808 
+ gnd vdd predecode_29[9] predecode_117[9] decode_b[297] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_809 
+ gnd vdd decode_b[297] decode[297] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_810 
+ gnd vdd predecode_29[9] predecode_117[10] decode_b[298] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_811 
+ gnd vdd decode_b[298] decode[298] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_812 
+ gnd vdd predecode_29[9] predecode_117[11] decode_b[299] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_813 
+ gnd vdd decode_b[299] decode[299] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_814 
+ gnd vdd predecode_29[9] predecode_117[12] decode_b[300] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_815 
+ gnd vdd decode_b[300] decode[300] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_816 
+ gnd vdd predecode_29[9] predecode_117[13] decode_b[301] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_817 
+ gnd vdd decode_b[301] decode[301] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_818 
+ gnd vdd predecode_29[9] predecode_117[14] decode_b[302] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_819 
+ gnd vdd decode_b[302] decode[302] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_820 
+ gnd vdd predecode_29[9] predecode_117[15] decode_b[303] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_821 
+ gnd vdd decode_b[303] decode[303] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_822 
+ gnd vdd predecode_29[9] predecode_117[16] decode_b[304] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_823 
+ gnd vdd decode_b[304] decode[304] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_824 
+ gnd vdd predecode_29[9] predecode_117[17] decode_b[305] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_825 
+ gnd vdd decode_b[305] decode[305] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_826 
+ gnd vdd predecode_29[9] predecode_117[18] decode_b[306] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_827 
+ gnd vdd decode_b[306] decode[306] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_828 
+ gnd vdd predecode_29[9] predecode_117[19] decode_b[307] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_829 
+ gnd vdd decode_b[307] decode[307] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_830 
+ gnd vdd predecode_29[9] predecode_117[20] decode_b[308] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_831 
+ gnd vdd decode_b[308] decode[308] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_832 
+ gnd vdd predecode_29[9] predecode_117[21] decode_b[309] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_833 
+ gnd vdd decode_b[309] decode[309] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_834 
+ gnd vdd predecode_29[9] predecode_117[22] decode_b[310] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_835 
+ gnd vdd decode_b[310] decode[310] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_836 
+ gnd vdd predecode_29[9] predecode_117[23] decode_b[311] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_837 
+ gnd vdd decode_b[311] decode[311] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_838 
+ gnd vdd predecode_29[9] predecode_117[24] decode_b[312] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_839 
+ gnd vdd decode_b[312] decode[312] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_840 
+ gnd vdd predecode_29[9] predecode_117[25] decode_b[313] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_841 
+ gnd vdd decode_b[313] decode[313] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_842 
+ gnd vdd predecode_29[9] predecode_117[26] decode_b[314] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_843 
+ gnd vdd decode_b[314] decode[314] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_844 
+ gnd vdd predecode_29[9] predecode_117[27] decode_b[315] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_845 
+ gnd vdd decode_b[315] decode[315] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_846 
+ gnd vdd predecode_29[9] predecode_117[28] decode_b[316] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_847 
+ gnd vdd decode_b[316] decode[316] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_848 
+ gnd vdd predecode_29[9] predecode_117[29] decode_b[317] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_849 
+ gnd vdd decode_b[317] decode[317] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_850 
+ gnd vdd predecode_29[9] predecode_117[30] decode_b[318] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_851 
+ gnd vdd decode_b[318] decode[318] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_852 
+ gnd vdd predecode_29[9] predecode_117[31] decode_b[319] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_853 
+ gnd vdd decode_b[319] decode[319] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_854 
+ gnd vdd predecode_29[10] predecode_117[0] decode_b[320] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_855 
+ gnd vdd decode_b[320] decode[320] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_856 
+ gnd vdd predecode_29[10] predecode_117[1] decode_b[321] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_857 
+ gnd vdd decode_b[321] decode[321] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_858 
+ gnd vdd predecode_29[10] predecode_117[2] decode_b[322] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_859 
+ gnd vdd decode_b[322] decode[322] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_860 
+ gnd vdd predecode_29[10] predecode_117[3] decode_b[323] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_861 
+ gnd vdd decode_b[323] decode[323] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_862 
+ gnd vdd predecode_29[10] predecode_117[4] decode_b[324] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_863 
+ gnd vdd decode_b[324] decode[324] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_864 
+ gnd vdd predecode_29[10] predecode_117[5] decode_b[325] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_865 
+ gnd vdd decode_b[325] decode[325] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_866 
+ gnd vdd predecode_29[10] predecode_117[6] decode_b[326] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_867 
+ gnd vdd decode_b[326] decode[326] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_868 
+ gnd vdd predecode_29[10] predecode_117[7] decode_b[327] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_869 
+ gnd vdd decode_b[327] decode[327] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_870 
+ gnd vdd predecode_29[10] predecode_117[8] decode_b[328] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_871 
+ gnd vdd decode_b[328] decode[328] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_872 
+ gnd vdd predecode_29[10] predecode_117[9] decode_b[329] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_873 
+ gnd vdd decode_b[329] decode[329] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_874 
+ gnd vdd predecode_29[10] predecode_117[10] decode_b[330] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_875 
+ gnd vdd decode_b[330] decode[330] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_876 
+ gnd vdd predecode_29[10] predecode_117[11] decode_b[331] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_877 
+ gnd vdd decode_b[331] decode[331] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_878 
+ gnd vdd predecode_29[10] predecode_117[12] decode_b[332] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_879 
+ gnd vdd decode_b[332] decode[332] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_880 
+ gnd vdd predecode_29[10] predecode_117[13] decode_b[333] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_881 
+ gnd vdd decode_b[333] decode[333] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_882 
+ gnd vdd predecode_29[10] predecode_117[14] decode_b[334] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_883 
+ gnd vdd decode_b[334] decode[334] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_884 
+ gnd vdd predecode_29[10] predecode_117[15] decode_b[335] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_885 
+ gnd vdd decode_b[335] decode[335] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_886 
+ gnd vdd predecode_29[10] predecode_117[16] decode_b[336] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_887 
+ gnd vdd decode_b[336] decode[336] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_888 
+ gnd vdd predecode_29[10] predecode_117[17] decode_b[337] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_889 
+ gnd vdd decode_b[337] decode[337] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_890 
+ gnd vdd predecode_29[10] predecode_117[18] decode_b[338] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_891 
+ gnd vdd decode_b[338] decode[338] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_892 
+ gnd vdd predecode_29[10] predecode_117[19] decode_b[339] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_893 
+ gnd vdd decode_b[339] decode[339] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_894 
+ gnd vdd predecode_29[10] predecode_117[20] decode_b[340] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_895 
+ gnd vdd decode_b[340] decode[340] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_896 
+ gnd vdd predecode_29[10] predecode_117[21] decode_b[341] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_897 
+ gnd vdd decode_b[341] decode[341] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_898 
+ gnd vdd predecode_29[10] predecode_117[22] decode_b[342] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_899 
+ gnd vdd decode_b[342] decode[342] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_900 
+ gnd vdd predecode_29[10] predecode_117[23] decode_b[343] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_901 
+ gnd vdd decode_b[343] decode[343] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_902 
+ gnd vdd predecode_29[10] predecode_117[24] decode_b[344] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_903 
+ gnd vdd decode_b[344] decode[344] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_904 
+ gnd vdd predecode_29[10] predecode_117[25] decode_b[345] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_905 
+ gnd vdd decode_b[345] decode[345] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_906 
+ gnd vdd predecode_29[10] predecode_117[26] decode_b[346] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_907 
+ gnd vdd decode_b[346] decode[346] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_908 
+ gnd vdd predecode_29[10] predecode_117[27] decode_b[347] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_909 
+ gnd vdd decode_b[347] decode[347] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_910 
+ gnd vdd predecode_29[10] predecode_117[28] decode_b[348] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_911 
+ gnd vdd decode_b[348] decode[348] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_912 
+ gnd vdd predecode_29[10] predecode_117[29] decode_b[349] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_913 
+ gnd vdd decode_b[349] decode[349] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_914 
+ gnd vdd predecode_29[10] predecode_117[30] decode_b[350] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_915 
+ gnd vdd decode_b[350] decode[350] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_916 
+ gnd vdd predecode_29[10] predecode_117[31] decode_b[351] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_917 
+ gnd vdd decode_b[351] decode[351] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_918 
+ gnd vdd predecode_29[11] predecode_117[0] decode_b[352] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_919 
+ gnd vdd decode_b[352] decode[352] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_920 
+ gnd vdd predecode_29[11] predecode_117[1] decode_b[353] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_921 
+ gnd vdd decode_b[353] decode[353] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_922 
+ gnd vdd predecode_29[11] predecode_117[2] decode_b[354] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_923 
+ gnd vdd decode_b[354] decode[354] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_924 
+ gnd vdd predecode_29[11] predecode_117[3] decode_b[355] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_925 
+ gnd vdd decode_b[355] decode[355] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_926 
+ gnd vdd predecode_29[11] predecode_117[4] decode_b[356] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_927 
+ gnd vdd decode_b[356] decode[356] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_928 
+ gnd vdd predecode_29[11] predecode_117[5] decode_b[357] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_929 
+ gnd vdd decode_b[357] decode[357] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_930 
+ gnd vdd predecode_29[11] predecode_117[6] decode_b[358] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_931 
+ gnd vdd decode_b[358] decode[358] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_932 
+ gnd vdd predecode_29[11] predecode_117[7] decode_b[359] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_933 
+ gnd vdd decode_b[359] decode[359] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_934 
+ gnd vdd predecode_29[11] predecode_117[8] decode_b[360] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_935 
+ gnd vdd decode_b[360] decode[360] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_936 
+ gnd vdd predecode_29[11] predecode_117[9] decode_b[361] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_937 
+ gnd vdd decode_b[361] decode[361] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_938 
+ gnd vdd predecode_29[11] predecode_117[10] decode_b[362] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_939 
+ gnd vdd decode_b[362] decode[362] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_940 
+ gnd vdd predecode_29[11] predecode_117[11] decode_b[363] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_941 
+ gnd vdd decode_b[363] decode[363] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_942 
+ gnd vdd predecode_29[11] predecode_117[12] decode_b[364] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_943 
+ gnd vdd decode_b[364] decode[364] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_944 
+ gnd vdd predecode_29[11] predecode_117[13] decode_b[365] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_945 
+ gnd vdd decode_b[365] decode[365] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_946 
+ gnd vdd predecode_29[11] predecode_117[14] decode_b[366] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_947 
+ gnd vdd decode_b[366] decode[366] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_948 
+ gnd vdd predecode_29[11] predecode_117[15] decode_b[367] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_949 
+ gnd vdd decode_b[367] decode[367] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_950 
+ gnd vdd predecode_29[11] predecode_117[16] decode_b[368] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_951 
+ gnd vdd decode_b[368] decode[368] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_952 
+ gnd vdd predecode_29[11] predecode_117[17] decode_b[369] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_953 
+ gnd vdd decode_b[369] decode[369] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_954 
+ gnd vdd predecode_29[11] predecode_117[18] decode_b[370] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_955 
+ gnd vdd decode_b[370] decode[370] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_956 
+ gnd vdd predecode_29[11] predecode_117[19] decode_b[371] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_957 
+ gnd vdd decode_b[371] decode[371] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_958 
+ gnd vdd predecode_29[11] predecode_117[20] decode_b[372] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_959 
+ gnd vdd decode_b[372] decode[372] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_960 
+ gnd vdd predecode_29[11] predecode_117[21] decode_b[373] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_961 
+ gnd vdd decode_b[373] decode[373] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_962 
+ gnd vdd predecode_29[11] predecode_117[22] decode_b[374] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_963 
+ gnd vdd decode_b[374] decode[374] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_964 
+ gnd vdd predecode_29[11] predecode_117[23] decode_b[375] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_965 
+ gnd vdd decode_b[375] decode[375] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_966 
+ gnd vdd predecode_29[11] predecode_117[24] decode_b[376] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_967 
+ gnd vdd decode_b[376] decode[376] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_968 
+ gnd vdd predecode_29[11] predecode_117[25] decode_b[377] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_969 
+ gnd vdd decode_b[377] decode[377] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_970 
+ gnd vdd predecode_29[11] predecode_117[26] decode_b[378] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_971 
+ gnd vdd decode_b[378] decode[378] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_972 
+ gnd vdd predecode_29[11] predecode_117[27] decode_b[379] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_973 
+ gnd vdd decode_b[379] decode[379] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_974 
+ gnd vdd predecode_29[11] predecode_117[28] decode_b[380] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_975 
+ gnd vdd decode_b[380] decode[380] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_976 
+ gnd vdd predecode_29[11] predecode_117[29] decode_b[381] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_977 
+ gnd vdd decode_b[381] decode[381] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_978 
+ gnd vdd predecode_29[11] predecode_117[30] decode_b[382] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_979 
+ gnd vdd decode_b[382] decode[382] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_980 
+ gnd vdd predecode_29[11] predecode_117[31] decode_b[383] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_981 
+ gnd vdd decode_b[383] decode[383] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_982 
+ gnd vdd predecode_29[12] predecode_117[0] decode_b[384] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_983 
+ gnd vdd decode_b[384] decode[384] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_984 
+ gnd vdd predecode_29[12] predecode_117[1] decode_b[385] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_985 
+ gnd vdd decode_b[385] decode[385] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_986 
+ gnd vdd predecode_29[12] predecode_117[2] decode_b[386] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_987 
+ gnd vdd decode_b[386] decode[386] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_988 
+ gnd vdd predecode_29[12] predecode_117[3] decode_b[387] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_989 
+ gnd vdd decode_b[387] decode[387] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_990 
+ gnd vdd predecode_29[12] predecode_117[4] decode_b[388] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_991 
+ gnd vdd decode_b[388] decode[388] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_992 
+ gnd vdd predecode_29[12] predecode_117[5] decode_b[389] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_993 
+ gnd vdd decode_b[389] decode[389] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_994 
+ gnd vdd predecode_29[12] predecode_117[6] decode_b[390] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_995 
+ gnd vdd decode_b[390] decode[390] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_996 
+ gnd vdd predecode_29[12] predecode_117[7] decode_b[391] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_997 
+ gnd vdd decode_b[391] decode[391] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_998 
+ gnd vdd predecode_29[12] predecode_117[8] decode_b[392] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_999 
+ gnd vdd decode_b[392] decode[392] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1000 
+ gnd vdd predecode_29[12] predecode_117[9] decode_b[393] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1001 
+ gnd vdd decode_b[393] decode[393] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1002 
+ gnd vdd predecode_29[12] predecode_117[10] decode_b[394] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1003 
+ gnd vdd decode_b[394] decode[394] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1004 
+ gnd vdd predecode_29[12] predecode_117[11] decode_b[395] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1005 
+ gnd vdd decode_b[395] decode[395] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1006 
+ gnd vdd predecode_29[12] predecode_117[12] decode_b[396] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1007 
+ gnd vdd decode_b[396] decode[396] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1008 
+ gnd vdd predecode_29[12] predecode_117[13] decode_b[397] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1009 
+ gnd vdd decode_b[397] decode[397] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1010 
+ gnd vdd predecode_29[12] predecode_117[14] decode_b[398] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1011 
+ gnd vdd decode_b[398] decode[398] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1012 
+ gnd vdd predecode_29[12] predecode_117[15] decode_b[399] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1013 
+ gnd vdd decode_b[399] decode[399] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1014 
+ gnd vdd predecode_29[12] predecode_117[16] decode_b[400] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1015 
+ gnd vdd decode_b[400] decode[400] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1016 
+ gnd vdd predecode_29[12] predecode_117[17] decode_b[401] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1017 
+ gnd vdd decode_b[401] decode[401] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1018 
+ gnd vdd predecode_29[12] predecode_117[18] decode_b[402] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1019 
+ gnd vdd decode_b[402] decode[402] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1020 
+ gnd vdd predecode_29[12] predecode_117[19] decode_b[403] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1021 
+ gnd vdd decode_b[403] decode[403] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1022 
+ gnd vdd predecode_29[12] predecode_117[20] decode_b[404] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1023 
+ gnd vdd decode_b[404] decode[404] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1024 
+ gnd vdd predecode_29[12] predecode_117[21] decode_b[405] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1025 
+ gnd vdd decode_b[405] decode[405] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1026 
+ gnd vdd predecode_29[12] predecode_117[22] decode_b[406] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1027 
+ gnd vdd decode_b[406] decode[406] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1028 
+ gnd vdd predecode_29[12] predecode_117[23] decode_b[407] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1029 
+ gnd vdd decode_b[407] decode[407] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1030 
+ gnd vdd predecode_29[12] predecode_117[24] decode_b[408] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1031 
+ gnd vdd decode_b[408] decode[408] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1032 
+ gnd vdd predecode_29[12] predecode_117[25] decode_b[409] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1033 
+ gnd vdd decode_b[409] decode[409] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1034 
+ gnd vdd predecode_29[12] predecode_117[26] decode_b[410] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1035 
+ gnd vdd decode_b[410] decode[410] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1036 
+ gnd vdd predecode_29[12] predecode_117[27] decode_b[411] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1037 
+ gnd vdd decode_b[411] decode[411] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1038 
+ gnd vdd predecode_29[12] predecode_117[28] decode_b[412] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1039 
+ gnd vdd decode_b[412] decode[412] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1040 
+ gnd vdd predecode_29[12] predecode_117[29] decode_b[413] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1041 
+ gnd vdd decode_b[413] decode[413] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1042 
+ gnd vdd predecode_29[12] predecode_117[30] decode_b[414] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1043 
+ gnd vdd decode_b[414] decode[414] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1044 
+ gnd vdd predecode_29[12] predecode_117[31] decode_b[415] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1045 
+ gnd vdd decode_b[415] decode[415] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1046 
+ gnd vdd predecode_29[13] predecode_117[0] decode_b[416] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1047 
+ gnd vdd decode_b[416] decode[416] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1048 
+ gnd vdd predecode_29[13] predecode_117[1] decode_b[417] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1049 
+ gnd vdd decode_b[417] decode[417] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1050 
+ gnd vdd predecode_29[13] predecode_117[2] decode_b[418] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1051 
+ gnd vdd decode_b[418] decode[418] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1052 
+ gnd vdd predecode_29[13] predecode_117[3] decode_b[419] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1053 
+ gnd vdd decode_b[419] decode[419] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1054 
+ gnd vdd predecode_29[13] predecode_117[4] decode_b[420] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1055 
+ gnd vdd decode_b[420] decode[420] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1056 
+ gnd vdd predecode_29[13] predecode_117[5] decode_b[421] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1057 
+ gnd vdd decode_b[421] decode[421] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1058 
+ gnd vdd predecode_29[13] predecode_117[6] decode_b[422] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1059 
+ gnd vdd decode_b[422] decode[422] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1060 
+ gnd vdd predecode_29[13] predecode_117[7] decode_b[423] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1061 
+ gnd vdd decode_b[423] decode[423] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1062 
+ gnd vdd predecode_29[13] predecode_117[8] decode_b[424] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1063 
+ gnd vdd decode_b[424] decode[424] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1064 
+ gnd vdd predecode_29[13] predecode_117[9] decode_b[425] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1065 
+ gnd vdd decode_b[425] decode[425] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1066 
+ gnd vdd predecode_29[13] predecode_117[10] decode_b[426] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1067 
+ gnd vdd decode_b[426] decode[426] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1068 
+ gnd vdd predecode_29[13] predecode_117[11] decode_b[427] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1069 
+ gnd vdd decode_b[427] decode[427] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1070 
+ gnd vdd predecode_29[13] predecode_117[12] decode_b[428] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1071 
+ gnd vdd decode_b[428] decode[428] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1072 
+ gnd vdd predecode_29[13] predecode_117[13] decode_b[429] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1073 
+ gnd vdd decode_b[429] decode[429] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1074 
+ gnd vdd predecode_29[13] predecode_117[14] decode_b[430] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1075 
+ gnd vdd decode_b[430] decode[430] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1076 
+ gnd vdd predecode_29[13] predecode_117[15] decode_b[431] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1077 
+ gnd vdd decode_b[431] decode[431] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1078 
+ gnd vdd predecode_29[13] predecode_117[16] decode_b[432] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1079 
+ gnd vdd decode_b[432] decode[432] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1080 
+ gnd vdd predecode_29[13] predecode_117[17] decode_b[433] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1081 
+ gnd vdd decode_b[433] decode[433] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1082 
+ gnd vdd predecode_29[13] predecode_117[18] decode_b[434] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1083 
+ gnd vdd decode_b[434] decode[434] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1084 
+ gnd vdd predecode_29[13] predecode_117[19] decode_b[435] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1085 
+ gnd vdd decode_b[435] decode[435] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1086 
+ gnd vdd predecode_29[13] predecode_117[20] decode_b[436] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1087 
+ gnd vdd decode_b[436] decode[436] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1088 
+ gnd vdd predecode_29[13] predecode_117[21] decode_b[437] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1089 
+ gnd vdd decode_b[437] decode[437] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1090 
+ gnd vdd predecode_29[13] predecode_117[22] decode_b[438] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1091 
+ gnd vdd decode_b[438] decode[438] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1092 
+ gnd vdd predecode_29[13] predecode_117[23] decode_b[439] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1093 
+ gnd vdd decode_b[439] decode[439] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1094 
+ gnd vdd predecode_29[13] predecode_117[24] decode_b[440] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1095 
+ gnd vdd decode_b[440] decode[440] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1096 
+ gnd vdd predecode_29[13] predecode_117[25] decode_b[441] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1097 
+ gnd vdd decode_b[441] decode[441] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1098 
+ gnd vdd predecode_29[13] predecode_117[26] decode_b[442] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1099 
+ gnd vdd decode_b[442] decode[442] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1100 
+ gnd vdd predecode_29[13] predecode_117[27] decode_b[443] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1101 
+ gnd vdd decode_b[443] decode[443] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1102 
+ gnd vdd predecode_29[13] predecode_117[28] decode_b[444] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1103 
+ gnd vdd decode_b[444] decode[444] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1104 
+ gnd vdd predecode_29[13] predecode_117[29] decode_b[445] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1105 
+ gnd vdd decode_b[445] decode[445] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1106 
+ gnd vdd predecode_29[13] predecode_117[30] decode_b[446] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1107 
+ gnd vdd decode_b[446] decode[446] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1108 
+ gnd vdd predecode_29[13] predecode_117[31] decode_b[447] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1109 
+ gnd vdd decode_b[447] decode[447] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1110 
+ gnd vdd predecode_29[14] predecode_117[0] decode_b[448] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1111 
+ gnd vdd decode_b[448] decode[448] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1112 
+ gnd vdd predecode_29[14] predecode_117[1] decode_b[449] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1113 
+ gnd vdd decode_b[449] decode[449] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1114 
+ gnd vdd predecode_29[14] predecode_117[2] decode_b[450] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1115 
+ gnd vdd decode_b[450] decode[450] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1116 
+ gnd vdd predecode_29[14] predecode_117[3] decode_b[451] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1117 
+ gnd vdd decode_b[451] decode[451] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1118 
+ gnd vdd predecode_29[14] predecode_117[4] decode_b[452] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1119 
+ gnd vdd decode_b[452] decode[452] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1120 
+ gnd vdd predecode_29[14] predecode_117[5] decode_b[453] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1121 
+ gnd vdd decode_b[453] decode[453] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1122 
+ gnd vdd predecode_29[14] predecode_117[6] decode_b[454] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1123 
+ gnd vdd decode_b[454] decode[454] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1124 
+ gnd vdd predecode_29[14] predecode_117[7] decode_b[455] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1125 
+ gnd vdd decode_b[455] decode[455] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1126 
+ gnd vdd predecode_29[14] predecode_117[8] decode_b[456] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1127 
+ gnd vdd decode_b[456] decode[456] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1128 
+ gnd vdd predecode_29[14] predecode_117[9] decode_b[457] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1129 
+ gnd vdd decode_b[457] decode[457] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1130 
+ gnd vdd predecode_29[14] predecode_117[10] decode_b[458] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1131 
+ gnd vdd decode_b[458] decode[458] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1132 
+ gnd vdd predecode_29[14] predecode_117[11] decode_b[459] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1133 
+ gnd vdd decode_b[459] decode[459] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1134 
+ gnd vdd predecode_29[14] predecode_117[12] decode_b[460] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1135 
+ gnd vdd decode_b[460] decode[460] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1136 
+ gnd vdd predecode_29[14] predecode_117[13] decode_b[461] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1137 
+ gnd vdd decode_b[461] decode[461] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1138 
+ gnd vdd predecode_29[14] predecode_117[14] decode_b[462] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1139 
+ gnd vdd decode_b[462] decode[462] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1140 
+ gnd vdd predecode_29[14] predecode_117[15] decode_b[463] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1141 
+ gnd vdd decode_b[463] decode[463] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1142 
+ gnd vdd predecode_29[14] predecode_117[16] decode_b[464] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1143 
+ gnd vdd decode_b[464] decode[464] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1144 
+ gnd vdd predecode_29[14] predecode_117[17] decode_b[465] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1145 
+ gnd vdd decode_b[465] decode[465] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1146 
+ gnd vdd predecode_29[14] predecode_117[18] decode_b[466] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1147 
+ gnd vdd decode_b[466] decode[466] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1148 
+ gnd vdd predecode_29[14] predecode_117[19] decode_b[467] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1149 
+ gnd vdd decode_b[467] decode[467] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1150 
+ gnd vdd predecode_29[14] predecode_117[20] decode_b[468] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1151 
+ gnd vdd decode_b[468] decode[468] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1152 
+ gnd vdd predecode_29[14] predecode_117[21] decode_b[469] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1153 
+ gnd vdd decode_b[469] decode[469] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1154 
+ gnd vdd predecode_29[14] predecode_117[22] decode_b[470] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1155 
+ gnd vdd decode_b[470] decode[470] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1156 
+ gnd vdd predecode_29[14] predecode_117[23] decode_b[471] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1157 
+ gnd vdd decode_b[471] decode[471] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1158 
+ gnd vdd predecode_29[14] predecode_117[24] decode_b[472] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1159 
+ gnd vdd decode_b[472] decode[472] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1160 
+ gnd vdd predecode_29[14] predecode_117[25] decode_b[473] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1161 
+ gnd vdd decode_b[473] decode[473] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1162 
+ gnd vdd predecode_29[14] predecode_117[26] decode_b[474] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1163 
+ gnd vdd decode_b[474] decode[474] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1164 
+ gnd vdd predecode_29[14] predecode_117[27] decode_b[475] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1165 
+ gnd vdd decode_b[475] decode[475] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1166 
+ gnd vdd predecode_29[14] predecode_117[28] decode_b[476] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1167 
+ gnd vdd decode_b[476] decode[476] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1168 
+ gnd vdd predecode_29[14] predecode_117[29] decode_b[477] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1169 
+ gnd vdd decode_b[477] decode[477] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1170 
+ gnd vdd predecode_29[14] predecode_117[30] decode_b[478] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1171 
+ gnd vdd decode_b[478] decode[478] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1172 
+ gnd vdd predecode_29[14] predecode_117[31] decode_b[479] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1173 
+ gnd vdd decode_b[479] decode[479] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1174 
+ gnd vdd predecode_29[15] predecode_117[0] decode_b[480] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1175 
+ gnd vdd decode_b[480] decode[480] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1176 
+ gnd vdd predecode_29[15] predecode_117[1] decode_b[481] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1177 
+ gnd vdd decode_b[481] decode[481] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1178 
+ gnd vdd predecode_29[15] predecode_117[2] decode_b[482] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1179 
+ gnd vdd decode_b[482] decode[482] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1180 
+ gnd vdd predecode_29[15] predecode_117[3] decode_b[483] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1181 
+ gnd vdd decode_b[483] decode[483] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1182 
+ gnd vdd predecode_29[15] predecode_117[4] decode_b[484] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1183 
+ gnd vdd decode_b[484] decode[484] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1184 
+ gnd vdd predecode_29[15] predecode_117[5] decode_b[485] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1185 
+ gnd vdd decode_b[485] decode[485] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1186 
+ gnd vdd predecode_29[15] predecode_117[6] decode_b[486] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1187 
+ gnd vdd decode_b[486] decode[486] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1188 
+ gnd vdd predecode_29[15] predecode_117[7] decode_b[487] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1189 
+ gnd vdd decode_b[487] decode[487] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1190 
+ gnd vdd predecode_29[15] predecode_117[8] decode_b[488] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1191 
+ gnd vdd decode_b[488] decode[488] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1192 
+ gnd vdd predecode_29[15] predecode_117[9] decode_b[489] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1193 
+ gnd vdd decode_b[489] decode[489] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1194 
+ gnd vdd predecode_29[15] predecode_117[10] decode_b[490] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1195 
+ gnd vdd decode_b[490] decode[490] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1196 
+ gnd vdd predecode_29[15] predecode_117[11] decode_b[491] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1197 
+ gnd vdd decode_b[491] decode[491] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1198 
+ gnd vdd predecode_29[15] predecode_117[12] decode_b[492] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1199 
+ gnd vdd decode_b[492] decode[492] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1200 
+ gnd vdd predecode_29[15] predecode_117[13] decode_b[493] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1201 
+ gnd vdd decode_b[493] decode[493] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1202 
+ gnd vdd predecode_29[15] predecode_117[14] decode_b[494] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1203 
+ gnd vdd decode_b[494] decode[494] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1204 
+ gnd vdd predecode_29[15] predecode_117[15] decode_b[495] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1205 
+ gnd vdd decode_b[495] decode[495] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1206 
+ gnd vdd predecode_29[15] predecode_117[16] decode_b[496] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1207 
+ gnd vdd decode_b[496] decode[496] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1208 
+ gnd vdd predecode_29[15] predecode_117[17] decode_b[497] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1209 
+ gnd vdd decode_b[497] decode[497] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1210 
+ gnd vdd predecode_29[15] predecode_117[18] decode_b[498] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1211 
+ gnd vdd decode_b[498] decode[498] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1212 
+ gnd vdd predecode_29[15] predecode_117[19] decode_b[499] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1213 
+ gnd vdd decode_b[499] decode[499] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1214 
+ gnd vdd predecode_29[15] predecode_117[20] decode_b[500] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1215 
+ gnd vdd decode_b[500] decode[500] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1216 
+ gnd vdd predecode_29[15] predecode_117[21] decode_b[501] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1217 
+ gnd vdd decode_b[501] decode[501] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1218 
+ gnd vdd predecode_29[15] predecode_117[22] decode_b[502] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1219 
+ gnd vdd decode_b[502] decode[502] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1220 
+ gnd vdd predecode_29[15] predecode_117[23] decode_b[503] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1221 
+ gnd vdd decode_b[503] decode[503] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1222 
+ gnd vdd predecode_29[15] predecode_117[24] decode_b[504] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1223 
+ gnd vdd decode_b[504] decode[504] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1224 
+ gnd vdd predecode_29[15] predecode_117[25] decode_b[505] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1225 
+ gnd vdd decode_b[505] decode[505] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1226 
+ gnd vdd predecode_29[15] predecode_117[26] decode_b[506] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1227 
+ gnd vdd decode_b[506] decode[506] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1228 
+ gnd vdd predecode_29[15] predecode_117[27] decode_b[507] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1229 
+ gnd vdd decode_b[507] decode[507] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1230 
+ gnd vdd predecode_29[15] predecode_117[28] decode_b[508] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1231 
+ gnd vdd decode_b[508] decode[508] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1232 
+ gnd vdd predecode_29[15] predecode_117[29] decode_b[509] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1233 
+ gnd vdd decode_b[509] decode[509] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1234 
+ gnd vdd predecode_29[15] predecode_117[30] decode_b[510] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1235 
+ gnd vdd decode_b[510] decode[510] 
+ hierarchical_decoder_inv_3 
* No parameters

xnand_1236 
+ gnd vdd predecode_29[15] predecode_117[31] decode_b[511] 
+ hierarchical_decoder_nand_2 
* No parameters

xinv_1237 
+ gnd vdd decode_b[511] decode[511] 
+ hierarchical_decoder_inv_3 
* No parameters

.ENDS

.SUBCKT column_decoder_nand_1 
+ gnd vdd a b c y 

xn1 
+ x1 a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ x2 b x1 gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn3 
+ y c x2 gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp3 
+ y c vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT column_decoder_inv_2 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT column_decoder 
+ vdd gnd addr[2] addr[1] addr[0] addr_b[2] addr_b[1] addr_b[0] decode[7] decode[6] decode[5] decode[4] decode[3] decode[2] decode[1] decode[0] decode_b[7] decode_b[6] decode_b[5] decode_b[4] decode_b[3] decode_b[2] decode_b[1] decode_b[0] 

xnand_3 
+ gnd vdd addr_b[2] addr_b[1] addr_b[0] decode_b[0] 
+ column_decoder_nand_1 
* No parameters

xinv_4 
+ gnd vdd decode_b[0] decode[0] 
+ column_decoder_inv_2 
* No parameters

xnand_5 
+ gnd vdd addr_b[2] addr_b[1] addr[0] decode_b[1] 
+ column_decoder_nand_1 
* No parameters

xinv_6 
+ gnd vdd decode_b[1] decode[1] 
+ column_decoder_inv_2 
* No parameters

xnand_7 
+ gnd vdd addr_b[2] addr[1] addr_b[0] decode_b[2] 
+ column_decoder_nand_1 
* No parameters

xinv_8 
+ gnd vdd decode_b[2] decode[2] 
+ column_decoder_inv_2 
* No parameters

xnand_9 
+ gnd vdd addr_b[2] addr[1] addr[0] decode_b[3] 
+ column_decoder_nand_1 
* No parameters

xinv_10 
+ gnd vdd decode_b[3] decode[3] 
+ column_decoder_inv_2 
* No parameters

xnand_11 
+ gnd vdd addr[2] addr_b[1] addr_b[0] decode_b[4] 
+ column_decoder_nand_1 
* No parameters

xinv_12 
+ gnd vdd decode_b[4] decode[4] 
+ column_decoder_inv_2 
* No parameters

xnand_13 
+ gnd vdd addr[2] addr_b[1] addr[0] decode_b[5] 
+ column_decoder_nand_1 
* No parameters

xinv_14 
+ gnd vdd decode_b[5] decode[5] 
+ column_decoder_inv_2 
* No parameters

xnand_15 
+ gnd vdd addr[2] addr[1] addr_b[0] decode_b[6] 
+ column_decoder_nand_1 
* No parameters

xinv_16 
+ gnd vdd decode_b[6] decode[6] 
+ column_decoder_inv_2 
* No parameters

xnand_17 
+ gnd vdd addr[2] addr[1] addr[0] decode_b[7] 
+ column_decoder_nand_1 
* No parameters

xinv_18 
+ gnd vdd decode_b[7] decode[7] 
+ column_decoder_inv_2 
* No parameters

.ENDS

.SUBCKT wordline_driver_and2_nand 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.2' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT wordline_driver_and2_inv 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='1.6' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.4' l='0.15' 

.ENDS

.SUBCKT wordline_driver_and2 
+ a b y vdd vss 

xnand 
+ vss vdd a b tmp 
+ wordline_driver_and2_nand 
* No parameters

xinv 
+ vss vdd tmp y 
+ wordline_driver_and2_inv 
* No parameters

.ENDS

.SUBCKT wordline_driver 
+ vdd vss din wl_en wl 

xand2 
+ din wl_en wl vdd vss 
+ wordline_driver_and2 
* No parameters

.ENDS

.SUBCKT wordline_driver_array 
+ vdd vss din[511] din[510] din[509] din[508] din[507] din[506] din[505] din[504] din[503] din[502] din[501] din[500] din[499] din[498] din[497] din[496] din[495] din[494] din[493] din[492] din[491] din[490] din[489] din[488] din[487] din[486] din[485] din[484] din[483] din[482] din[481] din[480] din[479] din[478] din[477] din[476] din[475] din[474] din[473] din[472] din[471] din[470] din[469] din[468] din[467] din[466] din[465] din[464] din[463] din[462] din[461] din[460] din[459] din[458] din[457] din[456] din[455] din[454] din[453] din[452] din[451] din[450] din[449] din[448] din[447] din[446] din[445] din[444] din[443] din[442] din[441] din[440] din[439] din[438] din[437] din[436] din[435] din[434] din[433] din[432] din[431] din[430] din[429] din[428] din[427] din[426] din[425] din[424] din[423] din[422] din[421] din[420] din[419] din[418] din[417] din[416] din[415] din[414] din[413] din[412] din[411] din[410] din[409] din[408] din[407] din[406] din[405] din[404] din[403] din[402] din[401] din[400] din[399] din[398] din[397] din[396] din[395] din[394] din[393] din[392] din[391] din[390] din[389] din[388] din[387] din[386] din[385] din[384] din[383] din[382] din[381] din[380] din[379] din[378] din[377] din[376] din[375] din[374] din[373] din[372] din[371] din[370] din[369] din[368] din[367] din[366] din[365] din[364] din[363] din[362] din[361] din[360] din[359] din[358] din[357] din[356] din[355] din[354] din[353] din[352] din[351] din[350] din[349] din[348] din[347] din[346] din[345] din[344] din[343] din[342] din[341] din[340] din[339] din[338] din[337] din[336] din[335] din[334] din[333] din[332] din[331] din[330] din[329] din[328] din[327] din[326] din[325] din[324] din[323] din[322] din[321] din[320] din[319] din[318] din[317] din[316] din[315] din[314] din[313] din[312] din[311] din[310] din[309] din[308] din[307] din[306] din[305] din[304] din[303] din[302] din[301] din[300] din[299] din[298] din[297] din[296] din[295] din[294] din[293] din[292] din[291] din[290] din[289] din[288] din[287] din[286] din[285] din[284] din[283] din[282] din[281] din[280] din[279] din[278] din[277] din[276] din[275] din[274] din[273] din[272] din[271] din[270] din[269] din[268] din[267] din[266] din[265] din[264] din[263] din[262] din[261] din[260] din[259] din[258] din[257] din[256] din[255] din[254] din[253] din[252] din[251] din[250] din[249] din[248] din[247] din[246] din[245] din[244] din[243] din[242] din[241] din[240] din[239] din[238] din[237] din[236] din[235] din[234] din[233] din[232] din[231] din[230] din[229] din[228] din[227] din[226] din[225] din[224] din[223] din[222] din[221] din[220] din[219] din[218] din[217] din[216] din[215] din[214] din[213] din[212] din[211] din[210] din[209] din[208] din[207] din[206] din[205] din[204] din[203] din[202] din[201] din[200] din[199] din[198] din[197] din[196] din[195] din[194] din[193] din[192] din[191] din[190] din[189] din[188] din[187] din[186] din[185] din[184] din[183] din[182] din[181] din[180] din[179] din[178] din[177] din[176] din[175] din[174] din[173] din[172] din[171] din[170] din[169] din[168] din[167] din[166] din[165] din[164] din[163] din[162] din[161] din[160] din[159] din[158] din[157] din[156] din[155] din[154] din[153] din[152] din[151] din[150] din[149] din[148] din[147] din[146] din[145] din[144] din[143] din[142] din[141] din[140] din[139] din[138] din[137] din[136] din[135] din[134] din[133] din[132] din[131] din[130] din[129] din[128] din[127] din[126] din[125] din[124] din[123] din[122] din[121] din[120] din[119] din[118] din[117] din[116] din[115] din[114] din[113] din[112] din[111] din[110] din[109] din[108] din[107] din[106] din[105] din[104] din[103] din[102] din[101] din[100] din[99] din[98] din[97] din[96] din[95] din[94] din[93] din[92] din[91] din[90] din[89] din[88] din[87] din[86] din[85] din[84] din[83] din[82] din[81] din[80] din[79] din[78] din[77] din[76] din[75] din[74] din[73] din[72] din[71] din[70] din[69] din[68] din[67] din[66] din[65] din[64] din[63] din[62] din[61] din[60] din[59] din[58] din[57] din[56] din[55] din[54] din[53] din[52] din[51] din[50] din[49] din[48] din[47] din[46] din[45] din[44] din[43] din[42] din[41] din[40] din[39] din[38] din[37] din[36] din[35] din[34] din[33] din[32] din[31] din[30] din[29] din[28] din[27] din[26] din[25] din[24] din[23] din[22] din[21] din[20] din[19] din[18] din[17] din[16] din[15] din[14] din[13] din[12] din[11] din[10] din[9] din[8] din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] wl_en wl[511] wl[510] wl[509] wl[508] wl[507] wl[506] wl[505] wl[504] wl[503] wl[502] wl[501] wl[500] wl[499] wl[498] wl[497] wl[496] wl[495] wl[494] wl[493] wl[492] wl[491] wl[490] wl[489] wl[488] wl[487] wl[486] wl[485] wl[484] wl[483] wl[482] wl[481] wl[480] wl[479] wl[478] wl[477] wl[476] wl[475] wl[474] wl[473] wl[472] wl[471] wl[470] wl[469] wl[468] wl[467] wl[466] wl[465] wl[464] wl[463] wl[462] wl[461] wl[460] wl[459] wl[458] wl[457] wl[456] wl[455] wl[454] wl[453] wl[452] wl[451] wl[450] wl[449] wl[448] wl[447] wl[446] wl[445] wl[444] wl[443] wl[442] wl[441] wl[440] wl[439] wl[438] wl[437] wl[436] wl[435] wl[434] wl[433] wl[432] wl[431] wl[430] wl[429] wl[428] wl[427] wl[426] wl[425] wl[424] wl[423] wl[422] wl[421] wl[420] wl[419] wl[418] wl[417] wl[416] wl[415] wl[414] wl[413] wl[412] wl[411] wl[410] wl[409] wl[408] wl[407] wl[406] wl[405] wl[404] wl[403] wl[402] wl[401] wl[400] wl[399] wl[398] wl[397] wl[396] wl[395] wl[394] wl[393] wl[392] wl[391] wl[390] wl[389] wl[388] wl[387] wl[386] wl[385] wl[384] wl[383] wl[382] wl[381] wl[380] wl[379] wl[378] wl[377] wl[376] wl[375] wl[374] wl[373] wl[372] wl[371] wl[370] wl[369] wl[368] wl[367] wl[366] wl[365] wl[364] wl[363] wl[362] wl[361] wl[360] wl[359] wl[358] wl[357] wl[356] wl[355] wl[354] wl[353] wl[352] wl[351] wl[350] wl[349] wl[348] wl[347] wl[346] wl[345] wl[344] wl[343] wl[342] wl[341] wl[340] wl[339] wl[338] wl[337] wl[336] wl[335] wl[334] wl[333] wl[332] wl[331] wl[330] wl[329] wl[328] wl[327] wl[326] wl[325] wl[324] wl[323] wl[322] wl[321] wl[320] wl[319] wl[318] wl[317] wl[316] wl[315] wl[314] wl[313] wl[312] wl[311] wl[310] wl[309] wl[308] wl[307] wl[306] wl[305] wl[304] wl[303] wl[302] wl[301] wl[300] wl[299] wl[298] wl[297] wl[296] wl[295] wl[294] wl[293] wl[292] wl[291] wl[290] wl[289] wl[288] wl[287] wl[286] wl[285] wl[284] wl[283] wl[282] wl[281] wl[280] wl[279] wl[278] wl[277] wl[276] wl[275] wl[274] wl[273] wl[272] wl[271] wl[270] wl[269] wl[268] wl[267] wl[266] wl[265] wl[264] wl[263] wl[262] wl[261] wl[260] wl[259] wl[258] wl[257] wl[256] wl[255] wl[254] wl[253] wl[252] wl[251] wl[250] wl[249] wl[248] wl[247] wl[246] wl[245] wl[244] wl[243] wl[242] wl[241] wl[240] wl[239] wl[238] wl[237] wl[236] wl[235] wl[234] wl[233] wl[232] wl[231] wl[230] wl[229] wl[228] wl[227] wl[226] wl[225] wl[224] wl[223] wl[222] wl[221] wl[220] wl[219] wl[218] wl[217] wl[216] wl[215] wl[214] wl[213] wl[212] wl[211] wl[210] wl[209] wl[208] wl[207] wl[206] wl[205] wl[204] wl[203] wl[202] wl[201] wl[200] wl[199] wl[198] wl[197] wl[196] wl[195] wl[194] wl[193] wl[192] wl[191] wl[190] wl[189] wl[188] wl[187] wl[186] wl[185] wl[184] wl[183] wl[182] wl[181] wl[180] wl[179] wl[178] wl[177] wl[176] wl[175] wl[174] wl[173] wl[172] wl[171] wl[170] wl[169] wl[168] wl[167] wl[166] wl[165] wl[164] wl[163] wl[162] wl[161] wl[160] wl[159] wl[158] wl[157] wl[156] wl[155] wl[154] wl[153] wl[152] wl[151] wl[150] wl[149] wl[148] wl[147] wl[146] wl[145] wl[144] wl[143] wl[142] wl[141] wl[140] wl[139] wl[138] wl[137] wl[136] wl[135] wl[134] wl[133] wl[132] wl[131] wl[130] wl[129] wl[128] wl[127] wl[126] wl[125] wl[124] wl[123] wl[122] wl[121] wl[120] wl[119] wl[118] wl[117] wl[116] wl[115] wl[114] wl[113] wl[112] wl[111] wl[110] wl[109] wl[108] wl[107] wl[106] wl[105] wl[104] wl[103] wl[102] wl[101] wl[100] wl[99] wl[98] wl[97] wl[96] wl[95] wl[94] wl[93] wl[92] wl[91] wl[90] wl[89] wl[88] wl[87] wl[86] wl[85] wl[84] wl[83] wl[82] wl[81] wl[80] wl[79] wl[78] wl[77] wl[76] wl[75] wl[74] wl[73] wl[72] wl[71] wl[70] wl[69] wl[68] wl[67] wl[66] wl[65] wl[64] wl[63] wl[62] wl[61] wl[60] wl[59] wl[58] wl[57] wl[56] wl[55] wl[54] wl[53] wl[52] wl[51] wl[50] wl[49] wl[48] wl[47] wl[46] wl[45] wl[44] wl[43] wl[42] wl[41] wl[40] wl[39] wl[38] wl[37] wl[36] wl[35] wl[34] wl[33] wl[32] wl[31] wl[30] wl[29] wl[28] wl[27] wl[26] wl[25] wl[24] wl[23] wl[22] wl[21] wl[20] wl[19] wl[18] wl[17] wl[16] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] 

xwl_driver_0 
+ vdd vss din[0] wl_en wl[0] 
+ wordline_driver 
* No parameters

xwl_driver_1 
+ vdd vss din[1] wl_en wl[1] 
+ wordline_driver 
* No parameters

xwl_driver_2 
+ vdd vss din[2] wl_en wl[2] 
+ wordline_driver 
* No parameters

xwl_driver_3 
+ vdd vss din[3] wl_en wl[3] 
+ wordline_driver 
* No parameters

xwl_driver_4 
+ vdd vss din[4] wl_en wl[4] 
+ wordline_driver 
* No parameters

xwl_driver_5 
+ vdd vss din[5] wl_en wl[5] 
+ wordline_driver 
* No parameters

xwl_driver_6 
+ vdd vss din[6] wl_en wl[6] 
+ wordline_driver 
* No parameters

xwl_driver_7 
+ vdd vss din[7] wl_en wl[7] 
+ wordline_driver 
* No parameters

xwl_driver_8 
+ vdd vss din[8] wl_en wl[8] 
+ wordline_driver 
* No parameters

xwl_driver_9 
+ vdd vss din[9] wl_en wl[9] 
+ wordline_driver 
* No parameters

xwl_driver_10 
+ vdd vss din[10] wl_en wl[10] 
+ wordline_driver 
* No parameters

xwl_driver_11 
+ vdd vss din[11] wl_en wl[11] 
+ wordline_driver 
* No parameters

xwl_driver_12 
+ vdd vss din[12] wl_en wl[12] 
+ wordline_driver 
* No parameters

xwl_driver_13 
+ vdd vss din[13] wl_en wl[13] 
+ wordline_driver 
* No parameters

xwl_driver_14 
+ vdd vss din[14] wl_en wl[14] 
+ wordline_driver 
* No parameters

xwl_driver_15 
+ vdd vss din[15] wl_en wl[15] 
+ wordline_driver 
* No parameters

xwl_driver_16 
+ vdd vss din[16] wl_en wl[16] 
+ wordline_driver 
* No parameters

xwl_driver_17 
+ vdd vss din[17] wl_en wl[17] 
+ wordline_driver 
* No parameters

xwl_driver_18 
+ vdd vss din[18] wl_en wl[18] 
+ wordline_driver 
* No parameters

xwl_driver_19 
+ vdd vss din[19] wl_en wl[19] 
+ wordline_driver 
* No parameters

xwl_driver_20 
+ vdd vss din[20] wl_en wl[20] 
+ wordline_driver 
* No parameters

xwl_driver_21 
+ vdd vss din[21] wl_en wl[21] 
+ wordline_driver 
* No parameters

xwl_driver_22 
+ vdd vss din[22] wl_en wl[22] 
+ wordline_driver 
* No parameters

xwl_driver_23 
+ vdd vss din[23] wl_en wl[23] 
+ wordline_driver 
* No parameters

xwl_driver_24 
+ vdd vss din[24] wl_en wl[24] 
+ wordline_driver 
* No parameters

xwl_driver_25 
+ vdd vss din[25] wl_en wl[25] 
+ wordline_driver 
* No parameters

xwl_driver_26 
+ vdd vss din[26] wl_en wl[26] 
+ wordline_driver 
* No parameters

xwl_driver_27 
+ vdd vss din[27] wl_en wl[27] 
+ wordline_driver 
* No parameters

xwl_driver_28 
+ vdd vss din[28] wl_en wl[28] 
+ wordline_driver 
* No parameters

xwl_driver_29 
+ vdd vss din[29] wl_en wl[29] 
+ wordline_driver 
* No parameters

xwl_driver_30 
+ vdd vss din[30] wl_en wl[30] 
+ wordline_driver 
* No parameters

xwl_driver_31 
+ vdd vss din[31] wl_en wl[31] 
+ wordline_driver 
* No parameters

xwl_driver_32 
+ vdd vss din[32] wl_en wl[32] 
+ wordline_driver 
* No parameters

xwl_driver_33 
+ vdd vss din[33] wl_en wl[33] 
+ wordline_driver 
* No parameters

xwl_driver_34 
+ vdd vss din[34] wl_en wl[34] 
+ wordline_driver 
* No parameters

xwl_driver_35 
+ vdd vss din[35] wl_en wl[35] 
+ wordline_driver 
* No parameters

xwl_driver_36 
+ vdd vss din[36] wl_en wl[36] 
+ wordline_driver 
* No parameters

xwl_driver_37 
+ vdd vss din[37] wl_en wl[37] 
+ wordline_driver 
* No parameters

xwl_driver_38 
+ vdd vss din[38] wl_en wl[38] 
+ wordline_driver 
* No parameters

xwl_driver_39 
+ vdd vss din[39] wl_en wl[39] 
+ wordline_driver 
* No parameters

xwl_driver_40 
+ vdd vss din[40] wl_en wl[40] 
+ wordline_driver 
* No parameters

xwl_driver_41 
+ vdd vss din[41] wl_en wl[41] 
+ wordline_driver 
* No parameters

xwl_driver_42 
+ vdd vss din[42] wl_en wl[42] 
+ wordline_driver 
* No parameters

xwl_driver_43 
+ vdd vss din[43] wl_en wl[43] 
+ wordline_driver 
* No parameters

xwl_driver_44 
+ vdd vss din[44] wl_en wl[44] 
+ wordline_driver 
* No parameters

xwl_driver_45 
+ vdd vss din[45] wl_en wl[45] 
+ wordline_driver 
* No parameters

xwl_driver_46 
+ vdd vss din[46] wl_en wl[46] 
+ wordline_driver 
* No parameters

xwl_driver_47 
+ vdd vss din[47] wl_en wl[47] 
+ wordline_driver 
* No parameters

xwl_driver_48 
+ vdd vss din[48] wl_en wl[48] 
+ wordline_driver 
* No parameters

xwl_driver_49 
+ vdd vss din[49] wl_en wl[49] 
+ wordline_driver 
* No parameters

xwl_driver_50 
+ vdd vss din[50] wl_en wl[50] 
+ wordline_driver 
* No parameters

xwl_driver_51 
+ vdd vss din[51] wl_en wl[51] 
+ wordline_driver 
* No parameters

xwl_driver_52 
+ vdd vss din[52] wl_en wl[52] 
+ wordline_driver 
* No parameters

xwl_driver_53 
+ vdd vss din[53] wl_en wl[53] 
+ wordline_driver 
* No parameters

xwl_driver_54 
+ vdd vss din[54] wl_en wl[54] 
+ wordline_driver 
* No parameters

xwl_driver_55 
+ vdd vss din[55] wl_en wl[55] 
+ wordline_driver 
* No parameters

xwl_driver_56 
+ vdd vss din[56] wl_en wl[56] 
+ wordline_driver 
* No parameters

xwl_driver_57 
+ vdd vss din[57] wl_en wl[57] 
+ wordline_driver 
* No parameters

xwl_driver_58 
+ vdd vss din[58] wl_en wl[58] 
+ wordline_driver 
* No parameters

xwl_driver_59 
+ vdd vss din[59] wl_en wl[59] 
+ wordline_driver 
* No parameters

xwl_driver_60 
+ vdd vss din[60] wl_en wl[60] 
+ wordline_driver 
* No parameters

xwl_driver_61 
+ vdd vss din[61] wl_en wl[61] 
+ wordline_driver 
* No parameters

xwl_driver_62 
+ vdd vss din[62] wl_en wl[62] 
+ wordline_driver 
* No parameters

xwl_driver_63 
+ vdd vss din[63] wl_en wl[63] 
+ wordline_driver 
* No parameters

xwl_driver_64 
+ vdd vss din[64] wl_en wl[64] 
+ wordline_driver 
* No parameters

xwl_driver_65 
+ vdd vss din[65] wl_en wl[65] 
+ wordline_driver 
* No parameters

xwl_driver_66 
+ vdd vss din[66] wl_en wl[66] 
+ wordline_driver 
* No parameters

xwl_driver_67 
+ vdd vss din[67] wl_en wl[67] 
+ wordline_driver 
* No parameters

xwl_driver_68 
+ vdd vss din[68] wl_en wl[68] 
+ wordline_driver 
* No parameters

xwl_driver_69 
+ vdd vss din[69] wl_en wl[69] 
+ wordline_driver 
* No parameters

xwl_driver_70 
+ vdd vss din[70] wl_en wl[70] 
+ wordline_driver 
* No parameters

xwl_driver_71 
+ vdd vss din[71] wl_en wl[71] 
+ wordline_driver 
* No parameters

xwl_driver_72 
+ vdd vss din[72] wl_en wl[72] 
+ wordline_driver 
* No parameters

xwl_driver_73 
+ vdd vss din[73] wl_en wl[73] 
+ wordline_driver 
* No parameters

xwl_driver_74 
+ vdd vss din[74] wl_en wl[74] 
+ wordline_driver 
* No parameters

xwl_driver_75 
+ vdd vss din[75] wl_en wl[75] 
+ wordline_driver 
* No parameters

xwl_driver_76 
+ vdd vss din[76] wl_en wl[76] 
+ wordline_driver 
* No parameters

xwl_driver_77 
+ vdd vss din[77] wl_en wl[77] 
+ wordline_driver 
* No parameters

xwl_driver_78 
+ vdd vss din[78] wl_en wl[78] 
+ wordline_driver 
* No parameters

xwl_driver_79 
+ vdd vss din[79] wl_en wl[79] 
+ wordline_driver 
* No parameters

xwl_driver_80 
+ vdd vss din[80] wl_en wl[80] 
+ wordline_driver 
* No parameters

xwl_driver_81 
+ vdd vss din[81] wl_en wl[81] 
+ wordline_driver 
* No parameters

xwl_driver_82 
+ vdd vss din[82] wl_en wl[82] 
+ wordline_driver 
* No parameters

xwl_driver_83 
+ vdd vss din[83] wl_en wl[83] 
+ wordline_driver 
* No parameters

xwl_driver_84 
+ vdd vss din[84] wl_en wl[84] 
+ wordline_driver 
* No parameters

xwl_driver_85 
+ vdd vss din[85] wl_en wl[85] 
+ wordline_driver 
* No parameters

xwl_driver_86 
+ vdd vss din[86] wl_en wl[86] 
+ wordline_driver 
* No parameters

xwl_driver_87 
+ vdd vss din[87] wl_en wl[87] 
+ wordline_driver 
* No parameters

xwl_driver_88 
+ vdd vss din[88] wl_en wl[88] 
+ wordline_driver 
* No parameters

xwl_driver_89 
+ vdd vss din[89] wl_en wl[89] 
+ wordline_driver 
* No parameters

xwl_driver_90 
+ vdd vss din[90] wl_en wl[90] 
+ wordline_driver 
* No parameters

xwl_driver_91 
+ vdd vss din[91] wl_en wl[91] 
+ wordline_driver 
* No parameters

xwl_driver_92 
+ vdd vss din[92] wl_en wl[92] 
+ wordline_driver 
* No parameters

xwl_driver_93 
+ vdd vss din[93] wl_en wl[93] 
+ wordline_driver 
* No parameters

xwl_driver_94 
+ vdd vss din[94] wl_en wl[94] 
+ wordline_driver 
* No parameters

xwl_driver_95 
+ vdd vss din[95] wl_en wl[95] 
+ wordline_driver 
* No parameters

xwl_driver_96 
+ vdd vss din[96] wl_en wl[96] 
+ wordline_driver 
* No parameters

xwl_driver_97 
+ vdd vss din[97] wl_en wl[97] 
+ wordline_driver 
* No parameters

xwl_driver_98 
+ vdd vss din[98] wl_en wl[98] 
+ wordline_driver 
* No parameters

xwl_driver_99 
+ vdd vss din[99] wl_en wl[99] 
+ wordline_driver 
* No parameters

xwl_driver_100 
+ vdd vss din[100] wl_en wl[100] 
+ wordline_driver 
* No parameters

xwl_driver_101 
+ vdd vss din[101] wl_en wl[101] 
+ wordline_driver 
* No parameters

xwl_driver_102 
+ vdd vss din[102] wl_en wl[102] 
+ wordline_driver 
* No parameters

xwl_driver_103 
+ vdd vss din[103] wl_en wl[103] 
+ wordline_driver 
* No parameters

xwl_driver_104 
+ vdd vss din[104] wl_en wl[104] 
+ wordline_driver 
* No parameters

xwl_driver_105 
+ vdd vss din[105] wl_en wl[105] 
+ wordline_driver 
* No parameters

xwl_driver_106 
+ vdd vss din[106] wl_en wl[106] 
+ wordline_driver 
* No parameters

xwl_driver_107 
+ vdd vss din[107] wl_en wl[107] 
+ wordline_driver 
* No parameters

xwl_driver_108 
+ vdd vss din[108] wl_en wl[108] 
+ wordline_driver 
* No parameters

xwl_driver_109 
+ vdd vss din[109] wl_en wl[109] 
+ wordline_driver 
* No parameters

xwl_driver_110 
+ vdd vss din[110] wl_en wl[110] 
+ wordline_driver 
* No parameters

xwl_driver_111 
+ vdd vss din[111] wl_en wl[111] 
+ wordline_driver 
* No parameters

xwl_driver_112 
+ vdd vss din[112] wl_en wl[112] 
+ wordline_driver 
* No parameters

xwl_driver_113 
+ vdd vss din[113] wl_en wl[113] 
+ wordline_driver 
* No parameters

xwl_driver_114 
+ vdd vss din[114] wl_en wl[114] 
+ wordline_driver 
* No parameters

xwl_driver_115 
+ vdd vss din[115] wl_en wl[115] 
+ wordline_driver 
* No parameters

xwl_driver_116 
+ vdd vss din[116] wl_en wl[116] 
+ wordline_driver 
* No parameters

xwl_driver_117 
+ vdd vss din[117] wl_en wl[117] 
+ wordline_driver 
* No parameters

xwl_driver_118 
+ vdd vss din[118] wl_en wl[118] 
+ wordline_driver 
* No parameters

xwl_driver_119 
+ vdd vss din[119] wl_en wl[119] 
+ wordline_driver 
* No parameters

xwl_driver_120 
+ vdd vss din[120] wl_en wl[120] 
+ wordline_driver 
* No parameters

xwl_driver_121 
+ vdd vss din[121] wl_en wl[121] 
+ wordline_driver 
* No parameters

xwl_driver_122 
+ vdd vss din[122] wl_en wl[122] 
+ wordline_driver 
* No parameters

xwl_driver_123 
+ vdd vss din[123] wl_en wl[123] 
+ wordline_driver 
* No parameters

xwl_driver_124 
+ vdd vss din[124] wl_en wl[124] 
+ wordline_driver 
* No parameters

xwl_driver_125 
+ vdd vss din[125] wl_en wl[125] 
+ wordline_driver 
* No parameters

xwl_driver_126 
+ vdd vss din[126] wl_en wl[126] 
+ wordline_driver 
* No parameters

xwl_driver_127 
+ vdd vss din[127] wl_en wl[127] 
+ wordline_driver 
* No parameters

xwl_driver_128 
+ vdd vss din[128] wl_en wl[128] 
+ wordline_driver 
* No parameters

xwl_driver_129 
+ vdd vss din[129] wl_en wl[129] 
+ wordline_driver 
* No parameters

xwl_driver_130 
+ vdd vss din[130] wl_en wl[130] 
+ wordline_driver 
* No parameters

xwl_driver_131 
+ vdd vss din[131] wl_en wl[131] 
+ wordline_driver 
* No parameters

xwl_driver_132 
+ vdd vss din[132] wl_en wl[132] 
+ wordline_driver 
* No parameters

xwl_driver_133 
+ vdd vss din[133] wl_en wl[133] 
+ wordline_driver 
* No parameters

xwl_driver_134 
+ vdd vss din[134] wl_en wl[134] 
+ wordline_driver 
* No parameters

xwl_driver_135 
+ vdd vss din[135] wl_en wl[135] 
+ wordline_driver 
* No parameters

xwl_driver_136 
+ vdd vss din[136] wl_en wl[136] 
+ wordline_driver 
* No parameters

xwl_driver_137 
+ vdd vss din[137] wl_en wl[137] 
+ wordline_driver 
* No parameters

xwl_driver_138 
+ vdd vss din[138] wl_en wl[138] 
+ wordline_driver 
* No parameters

xwl_driver_139 
+ vdd vss din[139] wl_en wl[139] 
+ wordline_driver 
* No parameters

xwl_driver_140 
+ vdd vss din[140] wl_en wl[140] 
+ wordline_driver 
* No parameters

xwl_driver_141 
+ vdd vss din[141] wl_en wl[141] 
+ wordline_driver 
* No parameters

xwl_driver_142 
+ vdd vss din[142] wl_en wl[142] 
+ wordline_driver 
* No parameters

xwl_driver_143 
+ vdd vss din[143] wl_en wl[143] 
+ wordline_driver 
* No parameters

xwl_driver_144 
+ vdd vss din[144] wl_en wl[144] 
+ wordline_driver 
* No parameters

xwl_driver_145 
+ vdd vss din[145] wl_en wl[145] 
+ wordline_driver 
* No parameters

xwl_driver_146 
+ vdd vss din[146] wl_en wl[146] 
+ wordline_driver 
* No parameters

xwl_driver_147 
+ vdd vss din[147] wl_en wl[147] 
+ wordline_driver 
* No parameters

xwl_driver_148 
+ vdd vss din[148] wl_en wl[148] 
+ wordline_driver 
* No parameters

xwl_driver_149 
+ vdd vss din[149] wl_en wl[149] 
+ wordline_driver 
* No parameters

xwl_driver_150 
+ vdd vss din[150] wl_en wl[150] 
+ wordline_driver 
* No parameters

xwl_driver_151 
+ vdd vss din[151] wl_en wl[151] 
+ wordline_driver 
* No parameters

xwl_driver_152 
+ vdd vss din[152] wl_en wl[152] 
+ wordline_driver 
* No parameters

xwl_driver_153 
+ vdd vss din[153] wl_en wl[153] 
+ wordline_driver 
* No parameters

xwl_driver_154 
+ vdd vss din[154] wl_en wl[154] 
+ wordline_driver 
* No parameters

xwl_driver_155 
+ vdd vss din[155] wl_en wl[155] 
+ wordline_driver 
* No parameters

xwl_driver_156 
+ vdd vss din[156] wl_en wl[156] 
+ wordline_driver 
* No parameters

xwl_driver_157 
+ vdd vss din[157] wl_en wl[157] 
+ wordline_driver 
* No parameters

xwl_driver_158 
+ vdd vss din[158] wl_en wl[158] 
+ wordline_driver 
* No parameters

xwl_driver_159 
+ vdd vss din[159] wl_en wl[159] 
+ wordline_driver 
* No parameters

xwl_driver_160 
+ vdd vss din[160] wl_en wl[160] 
+ wordline_driver 
* No parameters

xwl_driver_161 
+ vdd vss din[161] wl_en wl[161] 
+ wordline_driver 
* No parameters

xwl_driver_162 
+ vdd vss din[162] wl_en wl[162] 
+ wordline_driver 
* No parameters

xwl_driver_163 
+ vdd vss din[163] wl_en wl[163] 
+ wordline_driver 
* No parameters

xwl_driver_164 
+ vdd vss din[164] wl_en wl[164] 
+ wordline_driver 
* No parameters

xwl_driver_165 
+ vdd vss din[165] wl_en wl[165] 
+ wordline_driver 
* No parameters

xwl_driver_166 
+ vdd vss din[166] wl_en wl[166] 
+ wordline_driver 
* No parameters

xwl_driver_167 
+ vdd vss din[167] wl_en wl[167] 
+ wordline_driver 
* No parameters

xwl_driver_168 
+ vdd vss din[168] wl_en wl[168] 
+ wordline_driver 
* No parameters

xwl_driver_169 
+ vdd vss din[169] wl_en wl[169] 
+ wordline_driver 
* No parameters

xwl_driver_170 
+ vdd vss din[170] wl_en wl[170] 
+ wordline_driver 
* No parameters

xwl_driver_171 
+ vdd vss din[171] wl_en wl[171] 
+ wordline_driver 
* No parameters

xwl_driver_172 
+ vdd vss din[172] wl_en wl[172] 
+ wordline_driver 
* No parameters

xwl_driver_173 
+ vdd vss din[173] wl_en wl[173] 
+ wordline_driver 
* No parameters

xwl_driver_174 
+ vdd vss din[174] wl_en wl[174] 
+ wordline_driver 
* No parameters

xwl_driver_175 
+ vdd vss din[175] wl_en wl[175] 
+ wordline_driver 
* No parameters

xwl_driver_176 
+ vdd vss din[176] wl_en wl[176] 
+ wordline_driver 
* No parameters

xwl_driver_177 
+ vdd vss din[177] wl_en wl[177] 
+ wordline_driver 
* No parameters

xwl_driver_178 
+ vdd vss din[178] wl_en wl[178] 
+ wordline_driver 
* No parameters

xwl_driver_179 
+ vdd vss din[179] wl_en wl[179] 
+ wordline_driver 
* No parameters

xwl_driver_180 
+ vdd vss din[180] wl_en wl[180] 
+ wordline_driver 
* No parameters

xwl_driver_181 
+ vdd vss din[181] wl_en wl[181] 
+ wordline_driver 
* No parameters

xwl_driver_182 
+ vdd vss din[182] wl_en wl[182] 
+ wordline_driver 
* No parameters

xwl_driver_183 
+ vdd vss din[183] wl_en wl[183] 
+ wordline_driver 
* No parameters

xwl_driver_184 
+ vdd vss din[184] wl_en wl[184] 
+ wordline_driver 
* No parameters

xwl_driver_185 
+ vdd vss din[185] wl_en wl[185] 
+ wordline_driver 
* No parameters

xwl_driver_186 
+ vdd vss din[186] wl_en wl[186] 
+ wordline_driver 
* No parameters

xwl_driver_187 
+ vdd vss din[187] wl_en wl[187] 
+ wordline_driver 
* No parameters

xwl_driver_188 
+ vdd vss din[188] wl_en wl[188] 
+ wordline_driver 
* No parameters

xwl_driver_189 
+ vdd vss din[189] wl_en wl[189] 
+ wordline_driver 
* No parameters

xwl_driver_190 
+ vdd vss din[190] wl_en wl[190] 
+ wordline_driver 
* No parameters

xwl_driver_191 
+ vdd vss din[191] wl_en wl[191] 
+ wordline_driver 
* No parameters

xwl_driver_192 
+ vdd vss din[192] wl_en wl[192] 
+ wordline_driver 
* No parameters

xwl_driver_193 
+ vdd vss din[193] wl_en wl[193] 
+ wordline_driver 
* No parameters

xwl_driver_194 
+ vdd vss din[194] wl_en wl[194] 
+ wordline_driver 
* No parameters

xwl_driver_195 
+ vdd vss din[195] wl_en wl[195] 
+ wordline_driver 
* No parameters

xwl_driver_196 
+ vdd vss din[196] wl_en wl[196] 
+ wordline_driver 
* No parameters

xwl_driver_197 
+ vdd vss din[197] wl_en wl[197] 
+ wordline_driver 
* No parameters

xwl_driver_198 
+ vdd vss din[198] wl_en wl[198] 
+ wordline_driver 
* No parameters

xwl_driver_199 
+ vdd vss din[199] wl_en wl[199] 
+ wordline_driver 
* No parameters

xwl_driver_200 
+ vdd vss din[200] wl_en wl[200] 
+ wordline_driver 
* No parameters

xwl_driver_201 
+ vdd vss din[201] wl_en wl[201] 
+ wordline_driver 
* No parameters

xwl_driver_202 
+ vdd vss din[202] wl_en wl[202] 
+ wordline_driver 
* No parameters

xwl_driver_203 
+ vdd vss din[203] wl_en wl[203] 
+ wordline_driver 
* No parameters

xwl_driver_204 
+ vdd vss din[204] wl_en wl[204] 
+ wordline_driver 
* No parameters

xwl_driver_205 
+ vdd vss din[205] wl_en wl[205] 
+ wordline_driver 
* No parameters

xwl_driver_206 
+ vdd vss din[206] wl_en wl[206] 
+ wordline_driver 
* No parameters

xwl_driver_207 
+ vdd vss din[207] wl_en wl[207] 
+ wordline_driver 
* No parameters

xwl_driver_208 
+ vdd vss din[208] wl_en wl[208] 
+ wordline_driver 
* No parameters

xwl_driver_209 
+ vdd vss din[209] wl_en wl[209] 
+ wordline_driver 
* No parameters

xwl_driver_210 
+ vdd vss din[210] wl_en wl[210] 
+ wordline_driver 
* No parameters

xwl_driver_211 
+ vdd vss din[211] wl_en wl[211] 
+ wordline_driver 
* No parameters

xwl_driver_212 
+ vdd vss din[212] wl_en wl[212] 
+ wordline_driver 
* No parameters

xwl_driver_213 
+ vdd vss din[213] wl_en wl[213] 
+ wordline_driver 
* No parameters

xwl_driver_214 
+ vdd vss din[214] wl_en wl[214] 
+ wordline_driver 
* No parameters

xwl_driver_215 
+ vdd vss din[215] wl_en wl[215] 
+ wordline_driver 
* No parameters

xwl_driver_216 
+ vdd vss din[216] wl_en wl[216] 
+ wordline_driver 
* No parameters

xwl_driver_217 
+ vdd vss din[217] wl_en wl[217] 
+ wordline_driver 
* No parameters

xwl_driver_218 
+ vdd vss din[218] wl_en wl[218] 
+ wordline_driver 
* No parameters

xwl_driver_219 
+ vdd vss din[219] wl_en wl[219] 
+ wordline_driver 
* No parameters

xwl_driver_220 
+ vdd vss din[220] wl_en wl[220] 
+ wordline_driver 
* No parameters

xwl_driver_221 
+ vdd vss din[221] wl_en wl[221] 
+ wordline_driver 
* No parameters

xwl_driver_222 
+ vdd vss din[222] wl_en wl[222] 
+ wordline_driver 
* No parameters

xwl_driver_223 
+ vdd vss din[223] wl_en wl[223] 
+ wordline_driver 
* No parameters

xwl_driver_224 
+ vdd vss din[224] wl_en wl[224] 
+ wordline_driver 
* No parameters

xwl_driver_225 
+ vdd vss din[225] wl_en wl[225] 
+ wordline_driver 
* No parameters

xwl_driver_226 
+ vdd vss din[226] wl_en wl[226] 
+ wordline_driver 
* No parameters

xwl_driver_227 
+ vdd vss din[227] wl_en wl[227] 
+ wordline_driver 
* No parameters

xwl_driver_228 
+ vdd vss din[228] wl_en wl[228] 
+ wordline_driver 
* No parameters

xwl_driver_229 
+ vdd vss din[229] wl_en wl[229] 
+ wordline_driver 
* No parameters

xwl_driver_230 
+ vdd vss din[230] wl_en wl[230] 
+ wordline_driver 
* No parameters

xwl_driver_231 
+ vdd vss din[231] wl_en wl[231] 
+ wordline_driver 
* No parameters

xwl_driver_232 
+ vdd vss din[232] wl_en wl[232] 
+ wordline_driver 
* No parameters

xwl_driver_233 
+ vdd vss din[233] wl_en wl[233] 
+ wordline_driver 
* No parameters

xwl_driver_234 
+ vdd vss din[234] wl_en wl[234] 
+ wordline_driver 
* No parameters

xwl_driver_235 
+ vdd vss din[235] wl_en wl[235] 
+ wordline_driver 
* No parameters

xwl_driver_236 
+ vdd vss din[236] wl_en wl[236] 
+ wordline_driver 
* No parameters

xwl_driver_237 
+ vdd vss din[237] wl_en wl[237] 
+ wordline_driver 
* No parameters

xwl_driver_238 
+ vdd vss din[238] wl_en wl[238] 
+ wordline_driver 
* No parameters

xwl_driver_239 
+ vdd vss din[239] wl_en wl[239] 
+ wordline_driver 
* No parameters

xwl_driver_240 
+ vdd vss din[240] wl_en wl[240] 
+ wordline_driver 
* No parameters

xwl_driver_241 
+ vdd vss din[241] wl_en wl[241] 
+ wordline_driver 
* No parameters

xwl_driver_242 
+ vdd vss din[242] wl_en wl[242] 
+ wordline_driver 
* No parameters

xwl_driver_243 
+ vdd vss din[243] wl_en wl[243] 
+ wordline_driver 
* No parameters

xwl_driver_244 
+ vdd vss din[244] wl_en wl[244] 
+ wordline_driver 
* No parameters

xwl_driver_245 
+ vdd vss din[245] wl_en wl[245] 
+ wordline_driver 
* No parameters

xwl_driver_246 
+ vdd vss din[246] wl_en wl[246] 
+ wordline_driver 
* No parameters

xwl_driver_247 
+ vdd vss din[247] wl_en wl[247] 
+ wordline_driver 
* No parameters

xwl_driver_248 
+ vdd vss din[248] wl_en wl[248] 
+ wordline_driver 
* No parameters

xwl_driver_249 
+ vdd vss din[249] wl_en wl[249] 
+ wordline_driver 
* No parameters

xwl_driver_250 
+ vdd vss din[250] wl_en wl[250] 
+ wordline_driver 
* No parameters

xwl_driver_251 
+ vdd vss din[251] wl_en wl[251] 
+ wordline_driver 
* No parameters

xwl_driver_252 
+ vdd vss din[252] wl_en wl[252] 
+ wordline_driver 
* No parameters

xwl_driver_253 
+ vdd vss din[253] wl_en wl[253] 
+ wordline_driver 
* No parameters

xwl_driver_254 
+ vdd vss din[254] wl_en wl[254] 
+ wordline_driver 
* No parameters

xwl_driver_255 
+ vdd vss din[255] wl_en wl[255] 
+ wordline_driver 
* No parameters

xwl_driver_256 
+ vdd vss din[256] wl_en wl[256] 
+ wordline_driver 
* No parameters

xwl_driver_257 
+ vdd vss din[257] wl_en wl[257] 
+ wordline_driver 
* No parameters

xwl_driver_258 
+ vdd vss din[258] wl_en wl[258] 
+ wordline_driver 
* No parameters

xwl_driver_259 
+ vdd vss din[259] wl_en wl[259] 
+ wordline_driver 
* No parameters

xwl_driver_260 
+ vdd vss din[260] wl_en wl[260] 
+ wordline_driver 
* No parameters

xwl_driver_261 
+ vdd vss din[261] wl_en wl[261] 
+ wordline_driver 
* No parameters

xwl_driver_262 
+ vdd vss din[262] wl_en wl[262] 
+ wordline_driver 
* No parameters

xwl_driver_263 
+ vdd vss din[263] wl_en wl[263] 
+ wordline_driver 
* No parameters

xwl_driver_264 
+ vdd vss din[264] wl_en wl[264] 
+ wordline_driver 
* No parameters

xwl_driver_265 
+ vdd vss din[265] wl_en wl[265] 
+ wordline_driver 
* No parameters

xwl_driver_266 
+ vdd vss din[266] wl_en wl[266] 
+ wordline_driver 
* No parameters

xwl_driver_267 
+ vdd vss din[267] wl_en wl[267] 
+ wordline_driver 
* No parameters

xwl_driver_268 
+ vdd vss din[268] wl_en wl[268] 
+ wordline_driver 
* No parameters

xwl_driver_269 
+ vdd vss din[269] wl_en wl[269] 
+ wordline_driver 
* No parameters

xwl_driver_270 
+ vdd vss din[270] wl_en wl[270] 
+ wordline_driver 
* No parameters

xwl_driver_271 
+ vdd vss din[271] wl_en wl[271] 
+ wordline_driver 
* No parameters

xwl_driver_272 
+ vdd vss din[272] wl_en wl[272] 
+ wordline_driver 
* No parameters

xwl_driver_273 
+ vdd vss din[273] wl_en wl[273] 
+ wordline_driver 
* No parameters

xwl_driver_274 
+ vdd vss din[274] wl_en wl[274] 
+ wordline_driver 
* No parameters

xwl_driver_275 
+ vdd vss din[275] wl_en wl[275] 
+ wordline_driver 
* No parameters

xwl_driver_276 
+ vdd vss din[276] wl_en wl[276] 
+ wordline_driver 
* No parameters

xwl_driver_277 
+ vdd vss din[277] wl_en wl[277] 
+ wordline_driver 
* No parameters

xwl_driver_278 
+ vdd vss din[278] wl_en wl[278] 
+ wordline_driver 
* No parameters

xwl_driver_279 
+ vdd vss din[279] wl_en wl[279] 
+ wordline_driver 
* No parameters

xwl_driver_280 
+ vdd vss din[280] wl_en wl[280] 
+ wordline_driver 
* No parameters

xwl_driver_281 
+ vdd vss din[281] wl_en wl[281] 
+ wordline_driver 
* No parameters

xwl_driver_282 
+ vdd vss din[282] wl_en wl[282] 
+ wordline_driver 
* No parameters

xwl_driver_283 
+ vdd vss din[283] wl_en wl[283] 
+ wordline_driver 
* No parameters

xwl_driver_284 
+ vdd vss din[284] wl_en wl[284] 
+ wordline_driver 
* No parameters

xwl_driver_285 
+ vdd vss din[285] wl_en wl[285] 
+ wordline_driver 
* No parameters

xwl_driver_286 
+ vdd vss din[286] wl_en wl[286] 
+ wordline_driver 
* No parameters

xwl_driver_287 
+ vdd vss din[287] wl_en wl[287] 
+ wordline_driver 
* No parameters

xwl_driver_288 
+ vdd vss din[288] wl_en wl[288] 
+ wordline_driver 
* No parameters

xwl_driver_289 
+ vdd vss din[289] wl_en wl[289] 
+ wordline_driver 
* No parameters

xwl_driver_290 
+ vdd vss din[290] wl_en wl[290] 
+ wordline_driver 
* No parameters

xwl_driver_291 
+ vdd vss din[291] wl_en wl[291] 
+ wordline_driver 
* No parameters

xwl_driver_292 
+ vdd vss din[292] wl_en wl[292] 
+ wordline_driver 
* No parameters

xwl_driver_293 
+ vdd vss din[293] wl_en wl[293] 
+ wordline_driver 
* No parameters

xwl_driver_294 
+ vdd vss din[294] wl_en wl[294] 
+ wordline_driver 
* No parameters

xwl_driver_295 
+ vdd vss din[295] wl_en wl[295] 
+ wordline_driver 
* No parameters

xwl_driver_296 
+ vdd vss din[296] wl_en wl[296] 
+ wordline_driver 
* No parameters

xwl_driver_297 
+ vdd vss din[297] wl_en wl[297] 
+ wordline_driver 
* No parameters

xwl_driver_298 
+ vdd vss din[298] wl_en wl[298] 
+ wordline_driver 
* No parameters

xwl_driver_299 
+ vdd vss din[299] wl_en wl[299] 
+ wordline_driver 
* No parameters

xwl_driver_300 
+ vdd vss din[300] wl_en wl[300] 
+ wordline_driver 
* No parameters

xwl_driver_301 
+ vdd vss din[301] wl_en wl[301] 
+ wordline_driver 
* No parameters

xwl_driver_302 
+ vdd vss din[302] wl_en wl[302] 
+ wordline_driver 
* No parameters

xwl_driver_303 
+ vdd vss din[303] wl_en wl[303] 
+ wordline_driver 
* No parameters

xwl_driver_304 
+ vdd vss din[304] wl_en wl[304] 
+ wordline_driver 
* No parameters

xwl_driver_305 
+ vdd vss din[305] wl_en wl[305] 
+ wordline_driver 
* No parameters

xwl_driver_306 
+ vdd vss din[306] wl_en wl[306] 
+ wordline_driver 
* No parameters

xwl_driver_307 
+ vdd vss din[307] wl_en wl[307] 
+ wordline_driver 
* No parameters

xwl_driver_308 
+ vdd vss din[308] wl_en wl[308] 
+ wordline_driver 
* No parameters

xwl_driver_309 
+ vdd vss din[309] wl_en wl[309] 
+ wordline_driver 
* No parameters

xwl_driver_310 
+ vdd vss din[310] wl_en wl[310] 
+ wordline_driver 
* No parameters

xwl_driver_311 
+ vdd vss din[311] wl_en wl[311] 
+ wordline_driver 
* No parameters

xwl_driver_312 
+ vdd vss din[312] wl_en wl[312] 
+ wordline_driver 
* No parameters

xwl_driver_313 
+ vdd vss din[313] wl_en wl[313] 
+ wordline_driver 
* No parameters

xwl_driver_314 
+ vdd vss din[314] wl_en wl[314] 
+ wordline_driver 
* No parameters

xwl_driver_315 
+ vdd vss din[315] wl_en wl[315] 
+ wordline_driver 
* No parameters

xwl_driver_316 
+ vdd vss din[316] wl_en wl[316] 
+ wordline_driver 
* No parameters

xwl_driver_317 
+ vdd vss din[317] wl_en wl[317] 
+ wordline_driver 
* No parameters

xwl_driver_318 
+ vdd vss din[318] wl_en wl[318] 
+ wordline_driver 
* No parameters

xwl_driver_319 
+ vdd vss din[319] wl_en wl[319] 
+ wordline_driver 
* No parameters

xwl_driver_320 
+ vdd vss din[320] wl_en wl[320] 
+ wordline_driver 
* No parameters

xwl_driver_321 
+ vdd vss din[321] wl_en wl[321] 
+ wordline_driver 
* No parameters

xwl_driver_322 
+ vdd vss din[322] wl_en wl[322] 
+ wordline_driver 
* No parameters

xwl_driver_323 
+ vdd vss din[323] wl_en wl[323] 
+ wordline_driver 
* No parameters

xwl_driver_324 
+ vdd vss din[324] wl_en wl[324] 
+ wordline_driver 
* No parameters

xwl_driver_325 
+ vdd vss din[325] wl_en wl[325] 
+ wordline_driver 
* No parameters

xwl_driver_326 
+ vdd vss din[326] wl_en wl[326] 
+ wordline_driver 
* No parameters

xwl_driver_327 
+ vdd vss din[327] wl_en wl[327] 
+ wordline_driver 
* No parameters

xwl_driver_328 
+ vdd vss din[328] wl_en wl[328] 
+ wordline_driver 
* No parameters

xwl_driver_329 
+ vdd vss din[329] wl_en wl[329] 
+ wordline_driver 
* No parameters

xwl_driver_330 
+ vdd vss din[330] wl_en wl[330] 
+ wordline_driver 
* No parameters

xwl_driver_331 
+ vdd vss din[331] wl_en wl[331] 
+ wordline_driver 
* No parameters

xwl_driver_332 
+ vdd vss din[332] wl_en wl[332] 
+ wordline_driver 
* No parameters

xwl_driver_333 
+ vdd vss din[333] wl_en wl[333] 
+ wordline_driver 
* No parameters

xwl_driver_334 
+ vdd vss din[334] wl_en wl[334] 
+ wordline_driver 
* No parameters

xwl_driver_335 
+ vdd vss din[335] wl_en wl[335] 
+ wordline_driver 
* No parameters

xwl_driver_336 
+ vdd vss din[336] wl_en wl[336] 
+ wordline_driver 
* No parameters

xwl_driver_337 
+ vdd vss din[337] wl_en wl[337] 
+ wordline_driver 
* No parameters

xwl_driver_338 
+ vdd vss din[338] wl_en wl[338] 
+ wordline_driver 
* No parameters

xwl_driver_339 
+ vdd vss din[339] wl_en wl[339] 
+ wordline_driver 
* No parameters

xwl_driver_340 
+ vdd vss din[340] wl_en wl[340] 
+ wordline_driver 
* No parameters

xwl_driver_341 
+ vdd vss din[341] wl_en wl[341] 
+ wordline_driver 
* No parameters

xwl_driver_342 
+ vdd vss din[342] wl_en wl[342] 
+ wordline_driver 
* No parameters

xwl_driver_343 
+ vdd vss din[343] wl_en wl[343] 
+ wordline_driver 
* No parameters

xwl_driver_344 
+ vdd vss din[344] wl_en wl[344] 
+ wordline_driver 
* No parameters

xwl_driver_345 
+ vdd vss din[345] wl_en wl[345] 
+ wordline_driver 
* No parameters

xwl_driver_346 
+ vdd vss din[346] wl_en wl[346] 
+ wordline_driver 
* No parameters

xwl_driver_347 
+ vdd vss din[347] wl_en wl[347] 
+ wordline_driver 
* No parameters

xwl_driver_348 
+ vdd vss din[348] wl_en wl[348] 
+ wordline_driver 
* No parameters

xwl_driver_349 
+ vdd vss din[349] wl_en wl[349] 
+ wordline_driver 
* No parameters

xwl_driver_350 
+ vdd vss din[350] wl_en wl[350] 
+ wordline_driver 
* No parameters

xwl_driver_351 
+ vdd vss din[351] wl_en wl[351] 
+ wordline_driver 
* No parameters

xwl_driver_352 
+ vdd vss din[352] wl_en wl[352] 
+ wordline_driver 
* No parameters

xwl_driver_353 
+ vdd vss din[353] wl_en wl[353] 
+ wordline_driver 
* No parameters

xwl_driver_354 
+ vdd vss din[354] wl_en wl[354] 
+ wordline_driver 
* No parameters

xwl_driver_355 
+ vdd vss din[355] wl_en wl[355] 
+ wordline_driver 
* No parameters

xwl_driver_356 
+ vdd vss din[356] wl_en wl[356] 
+ wordline_driver 
* No parameters

xwl_driver_357 
+ vdd vss din[357] wl_en wl[357] 
+ wordline_driver 
* No parameters

xwl_driver_358 
+ vdd vss din[358] wl_en wl[358] 
+ wordline_driver 
* No parameters

xwl_driver_359 
+ vdd vss din[359] wl_en wl[359] 
+ wordline_driver 
* No parameters

xwl_driver_360 
+ vdd vss din[360] wl_en wl[360] 
+ wordline_driver 
* No parameters

xwl_driver_361 
+ vdd vss din[361] wl_en wl[361] 
+ wordline_driver 
* No parameters

xwl_driver_362 
+ vdd vss din[362] wl_en wl[362] 
+ wordline_driver 
* No parameters

xwl_driver_363 
+ vdd vss din[363] wl_en wl[363] 
+ wordline_driver 
* No parameters

xwl_driver_364 
+ vdd vss din[364] wl_en wl[364] 
+ wordline_driver 
* No parameters

xwl_driver_365 
+ vdd vss din[365] wl_en wl[365] 
+ wordline_driver 
* No parameters

xwl_driver_366 
+ vdd vss din[366] wl_en wl[366] 
+ wordline_driver 
* No parameters

xwl_driver_367 
+ vdd vss din[367] wl_en wl[367] 
+ wordline_driver 
* No parameters

xwl_driver_368 
+ vdd vss din[368] wl_en wl[368] 
+ wordline_driver 
* No parameters

xwl_driver_369 
+ vdd vss din[369] wl_en wl[369] 
+ wordline_driver 
* No parameters

xwl_driver_370 
+ vdd vss din[370] wl_en wl[370] 
+ wordline_driver 
* No parameters

xwl_driver_371 
+ vdd vss din[371] wl_en wl[371] 
+ wordline_driver 
* No parameters

xwl_driver_372 
+ vdd vss din[372] wl_en wl[372] 
+ wordline_driver 
* No parameters

xwl_driver_373 
+ vdd vss din[373] wl_en wl[373] 
+ wordline_driver 
* No parameters

xwl_driver_374 
+ vdd vss din[374] wl_en wl[374] 
+ wordline_driver 
* No parameters

xwl_driver_375 
+ vdd vss din[375] wl_en wl[375] 
+ wordline_driver 
* No parameters

xwl_driver_376 
+ vdd vss din[376] wl_en wl[376] 
+ wordline_driver 
* No parameters

xwl_driver_377 
+ vdd vss din[377] wl_en wl[377] 
+ wordline_driver 
* No parameters

xwl_driver_378 
+ vdd vss din[378] wl_en wl[378] 
+ wordline_driver 
* No parameters

xwl_driver_379 
+ vdd vss din[379] wl_en wl[379] 
+ wordline_driver 
* No parameters

xwl_driver_380 
+ vdd vss din[380] wl_en wl[380] 
+ wordline_driver 
* No parameters

xwl_driver_381 
+ vdd vss din[381] wl_en wl[381] 
+ wordline_driver 
* No parameters

xwl_driver_382 
+ vdd vss din[382] wl_en wl[382] 
+ wordline_driver 
* No parameters

xwl_driver_383 
+ vdd vss din[383] wl_en wl[383] 
+ wordline_driver 
* No parameters

xwl_driver_384 
+ vdd vss din[384] wl_en wl[384] 
+ wordline_driver 
* No parameters

xwl_driver_385 
+ vdd vss din[385] wl_en wl[385] 
+ wordline_driver 
* No parameters

xwl_driver_386 
+ vdd vss din[386] wl_en wl[386] 
+ wordline_driver 
* No parameters

xwl_driver_387 
+ vdd vss din[387] wl_en wl[387] 
+ wordline_driver 
* No parameters

xwl_driver_388 
+ vdd vss din[388] wl_en wl[388] 
+ wordline_driver 
* No parameters

xwl_driver_389 
+ vdd vss din[389] wl_en wl[389] 
+ wordline_driver 
* No parameters

xwl_driver_390 
+ vdd vss din[390] wl_en wl[390] 
+ wordline_driver 
* No parameters

xwl_driver_391 
+ vdd vss din[391] wl_en wl[391] 
+ wordline_driver 
* No parameters

xwl_driver_392 
+ vdd vss din[392] wl_en wl[392] 
+ wordline_driver 
* No parameters

xwl_driver_393 
+ vdd vss din[393] wl_en wl[393] 
+ wordline_driver 
* No parameters

xwl_driver_394 
+ vdd vss din[394] wl_en wl[394] 
+ wordline_driver 
* No parameters

xwl_driver_395 
+ vdd vss din[395] wl_en wl[395] 
+ wordline_driver 
* No parameters

xwl_driver_396 
+ vdd vss din[396] wl_en wl[396] 
+ wordline_driver 
* No parameters

xwl_driver_397 
+ vdd vss din[397] wl_en wl[397] 
+ wordline_driver 
* No parameters

xwl_driver_398 
+ vdd vss din[398] wl_en wl[398] 
+ wordline_driver 
* No parameters

xwl_driver_399 
+ vdd vss din[399] wl_en wl[399] 
+ wordline_driver 
* No parameters

xwl_driver_400 
+ vdd vss din[400] wl_en wl[400] 
+ wordline_driver 
* No parameters

xwl_driver_401 
+ vdd vss din[401] wl_en wl[401] 
+ wordline_driver 
* No parameters

xwl_driver_402 
+ vdd vss din[402] wl_en wl[402] 
+ wordline_driver 
* No parameters

xwl_driver_403 
+ vdd vss din[403] wl_en wl[403] 
+ wordline_driver 
* No parameters

xwl_driver_404 
+ vdd vss din[404] wl_en wl[404] 
+ wordline_driver 
* No parameters

xwl_driver_405 
+ vdd vss din[405] wl_en wl[405] 
+ wordline_driver 
* No parameters

xwl_driver_406 
+ vdd vss din[406] wl_en wl[406] 
+ wordline_driver 
* No parameters

xwl_driver_407 
+ vdd vss din[407] wl_en wl[407] 
+ wordline_driver 
* No parameters

xwl_driver_408 
+ vdd vss din[408] wl_en wl[408] 
+ wordline_driver 
* No parameters

xwl_driver_409 
+ vdd vss din[409] wl_en wl[409] 
+ wordline_driver 
* No parameters

xwl_driver_410 
+ vdd vss din[410] wl_en wl[410] 
+ wordline_driver 
* No parameters

xwl_driver_411 
+ vdd vss din[411] wl_en wl[411] 
+ wordline_driver 
* No parameters

xwl_driver_412 
+ vdd vss din[412] wl_en wl[412] 
+ wordline_driver 
* No parameters

xwl_driver_413 
+ vdd vss din[413] wl_en wl[413] 
+ wordline_driver 
* No parameters

xwl_driver_414 
+ vdd vss din[414] wl_en wl[414] 
+ wordline_driver 
* No parameters

xwl_driver_415 
+ vdd vss din[415] wl_en wl[415] 
+ wordline_driver 
* No parameters

xwl_driver_416 
+ vdd vss din[416] wl_en wl[416] 
+ wordline_driver 
* No parameters

xwl_driver_417 
+ vdd vss din[417] wl_en wl[417] 
+ wordline_driver 
* No parameters

xwl_driver_418 
+ vdd vss din[418] wl_en wl[418] 
+ wordline_driver 
* No parameters

xwl_driver_419 
+ vdd vss din[419] wl_en wl[419] 
+ wordline_driver 
* No parameters

xwl_driver_420 
+ vdd vss din[420] wl_en wl[420] 
+ wordline_driver 
* No parameters

xwl_driver_421 
+ vdd vss din[421] wl_en wl[421] 
+ wordline_driver 
* No parameters

xwl_driver_422 
+ vdd vss din[422] wl_en wl[422] 
+ wordline_driver 
* No parameters

xwl_driver_423 
+ vdd vss din[423] wl_en wl[423] 
+ wordline_driver 
* No parameters

xwl_driver_424 
+ vdd vss din[424] wl_en wl[424] 
+ wordline_driver 
* No parameters

xwl_driver_425 
+ vdd vss din[425] wl_en wl[425] 
+ wordline_driver 
* No parameters

xwl_driver_426 
+ vdd vss din[426] wl_en wl[426] 
+ wordline_driver 
* No parameters

xwl_driver_427 
+ vdd vss din[427] wl_en wl[427] 
+ wordline_driver 
* No parameters

xwl_driver_428 
+ vdd vss din[428] wl_en wl[428] 
+ wordline_driver 
* No parameters

xwl_driver_429 
+ vdd vss din[429] wl_en wl[429] 
+ wordline_driver 
* No parameters

xwl_driver_430 
+ vdd vss din[430] wl_en wl[430] 
+ wordline_driver 
* No parameters

xwl_driver_431 
+ vdd vss din[431] wl_en wl[431] 
+ wordline_driver 
* No parameters

xwl_driver_432 
+ vdd vss din[432] wl_en wl[432] 
+ wordline_driver 
* No parameters

xwl_driver_433 
+ vdd vss din[433] wl_en wl[433] 
+ wordline_driver 
* No parameters

xwl_driver_434 
+ vdd vss din[434] wl_en wl[434] 
+ wordline_driver 
* No parameters

xwl_driver_435 
+ vdd vss din[435] wl_en wl[435] 
+ wordline_driver 
* No parameters

xwl_driver_436 
+ vdd vss din[436] wl_en wl[436] 
+ wordline_driver 
* No parameters

xwl_driver_437 
+ vdd vss din[437] wl_en wl[437] 
+ wordline_driver 
* No parameters

xwl_driver_438 
+ vdd vss din[438] wl_en wl[438] 
+ wordline_driver 
* No parameters

xwl_driver_439 
+ vdd vss din[439] wl_en wl[439] 
+ wordline_driver 
* No parameters

xwl_driver_440 
+ vdd vss din[440] wl_en wl[440] 
+ wordline_driver 
* No parameters

xwl_driver_441 
+ vdd vss din[441] wl_en wl[441] 
+ wordline_driver 
* No parameters

xwl_driver_442 
+ vdd vss din[442] wl_en wl[442] 
+ wordline_driver 
* No parameters

xwl_driver_443 
+ vdd vss din[443] wl_en wl[443] 
+ wordline_driver 
* No parameters

xwl_driver_444 
+ vdd vss din[444] wl_en wl[444] 
+ wordline_driver 
* No parameters

xwl_driver_445 
+ vdd vss din[445] wl_en wl[445] 
+ wordline_driver 
* No parameters

xwl_driver_446 
+ vdd vss din[446] wl_en wl[446] 
+ wordline_driver 
* No parameters

xwl_driver_447 
+ vdd vss din[447] wl_en wl[447] 
+ wordline_driver 
* No parameters

xwl_driver_448 
+ vdd vss din[448] wl_en wl[448] 
+ wordline_driver 
* No parameters

xwl_driver_449 
+ vdd vss din[449] wl_en wl[449] 
+ wordline_driver 
* No parameters

xwl_driver_450 
+ vdd vss din[450] wl_en wl[450] 
+ wordline_driver 
* No parameters

xwl_driver_451 
+ vdd vss din[451] wl_en wl[451] 
+ wordline_driver 
* No parameters

xwl_driver_452 
+ vdd vss din[452] wl_en wl[452] 
+ wordline_driver 
* No parameters

xwl_driver_453 
+ vdd vss din[453] wl_en wl[453] 
+ wordline_driver 
* No parameters

xwl_driver_454 
+ vdd vss din[454] wl_en wl[454] 
+ wordline_driver 
* No parameters

xwl_driver_455 
+ vdd vss din[455] wl_en wl[455] 
+ wordline_driver 
* No parameters

xwl_driver_456 
+ vdd vss din[456] wl_en wl[456] 
+ wordline_driver 
* No parameters

xwl_driver_457 
+ vdd vss din[457] wl_en wl[457] 
+ wordline_driver 
* No parameters

xwl_driver_458 
+ vdd vss din[458] wl_en wl[458] 
+ wordline_driver 
* No parameters

xwl_driver_459 
+ vdd vss din[459] wl_en wl[459] 
+ wordline_driver 
* No parameters

xwl_driver_460 
+ vdd vss din[460] wl_en wl[460] 
+ wordline_driver 
* No parameters

xwl_driver_461 
+ vdd vss din[461] wl_en wl[461] 
+ wordline_driver 
* No parameters

xwl_driver_462 
+ vdd vss din[462] wl_en wl[462] 
+ wordline_driver 
* No parameters

xwl_driver_463 
+ vdd vss din[463] wl_en wl[463] 
+ wordline_driver 
* No parameters

xwl_driver_464 
+ vdd vss din[464] wl_en wl[464] 
+ wordline_driver 
* No parameters

xwl_driver_465 
+ vdd vss din[465] wl_en wl[465] 
+ wordline_driver 
* No parameters

xwl_driver_466 
+ vdd vss din[466] wl_en wl[466] 
+ wordline_driver 
* No parameters

xwl_driver_467 
+ vdd vss din[467] wl_en wl[467] 
+ wordline_driver 
* No parameters

xwl_driver_468 
+ vdd vss din[468] wl_en wl[468] 
+ wordline_driver 
* No parameters

xwl_driver_469 
+ vdd vss din[469] wl_en wl[469] 
+ wordline_driver 
* No parameters

xwl_driver_470 
+ vdd vss din[470] wl_en wl[470] 
+ wordline_driver 
* No parameters

xwl_driver_471 
+ vdd vss din[471] wl_en wl[471] 
+ wordline_driver 
* No parameters

xwl_driver_472 
+ vdd vss din[472] wl_en wl[472] 
+ wordline_driver 
* No parameters

xwl_driver_473 
+ vdd vss din[473] wl_en wl[473] 
+ wordline_driver 
* No parameters

xwl_driver_474 
+ vdd vss din[474] wl_en wl[474] 
+ wordline_driver 
* No parameters

xwl_driver_475 
+ vdd vss din[475] wl_en wl[475] 
+ wordline_driver 
* No parameters

xwl_driver_476 
+ vdd vss din[476] wl_en wl[476] 
+ wordline_driver 
* No parameters

xwl_driver_477 
+ vdd vss din[477] wl_en wl[477] 
+ wordline_driver 
* No parameters

xwl_driver_478 
+ vdd vss din[478] wl_en wl[478] 
+ wordline_driver 
* No parameters

xwl_driver_479 
+ vdd vss din[479] wl_en wl[479] 
+ wordline_driver 
* No parameters

xwl_driver_480 
+ vdd vss din[480] wl_en wl[480] 
+ wordline_driver 
* No parameters

xwl_driver_481 
+ vdd vss din[481] wl_en wl[481] 
+ wordline_driver 
* No parameters

xwl_driver_482 
+ vdd vss din[482] wl_en wl[482] 
+ wordline_driver 
* No parameters

xwl_driver_483 
+ vdd vss din[483] wl_en wl[483] 
+ wordline_driver 
* No parameters

xwl_driver_484 
+ vdd vss din[484] wl_en wl[484] 
+ wordline_driver 
* No parameters

xwl_driver_485 
+ vdd vss din[485] wl_en wl[485] 
+ wordline_driver 
* No parameters

xwl_driver_486 
+ vdd vss din[486] wl_en wl[486] 
+ wordline_driver 
* No parameters

xwl_driver_487 
+ vdd vss din[487] wl_en wl[487] 
+ wordline_driver 
* No parameters

xwl_driver_488 
+ vdd vss din[488] wl_en wl[488] 
+ wordline_driver 
* No parameters

xwl_driver_489 
+ vdd vss din[489] wl_en wl[489] 
+ wordline_driver 
* No parameters

xwl_driver_490 
+ vdd vss din[490] wl_en wl[490] 
+ wordline_driver 
* No parameters

xwl_driver_491 
+ vdd vss din[491] wl_en wl[491] 
+ wordline_driver 
* No parameters

xwl_driver_492 
+ vdd vss din[492] wl_en wl[492] 
+ wordline_driver 
* No parameters

xwl_driver_493 
+ vdd vss din[493] wl_en wl[493] 
+ wordline_driver 
* No parameters

xwl_driver_494 
+ vdd vss din[494] wl_en wl[494] 
+ wordline_driver 
* No parameters

xwl_driver_495 
+ vdd vss din[495] wl_en wl[495] 
+ wordline_driver 
* No parameters

xwl_driver_496 
+ vdd vss din[496] wl_en wl[496] 
+ wordline_driver 
* No parameters

xwl_driver_497 
+ vdd vss din[497] wl_en wl[497] 
+ wordline_driver 
* No parameters

xwl_driver_498 
+ vdd vss din[498] wl_en wl[498] 
+ wordline_driver 
* No parameters

xwl_driver_499 
+ vdd vss din[499] wl_en wl[499] 
+ wordline_driver 
* No parameters

xwl_driver_500 
+ vdd vss din[500] wl_en wl[500] 
+ wordline_driver 
* No parameters

xwl_driver_501 
+ vdd vss din[501] wl_en wl[501] 
+ wordline_driver 
* No parameters

xwl_driver_502 
+ vdd vss din[502] wl_en wl[502] 
+ wordline_driver 
* No parameters

xwl_driver_503 
+ vdd vss din[503] wl_en wl[503] 
+ wordline_driver 
* No parameters

xwl_driver_504 
+ vdd vss din[504] wl_en wl[504] 
+ wordline_driver 
* No parameters

xwl_driver_505 
+ vdd vss din[505] wl_en wl[505] 
+ wordline_driver 
* No parameters

xwl_driver_506 
+ vdd vss din[506] wl_en wl[506] 
+ wordline_driver 
* No parameters

xwl_driver_507 
+ vdd vss din[507] wl_en wl[507] 
+ wordline_driver 
* No parameters

xwl_driver_508 
+ vdd vss din[508] wl_en wl[508] 
+ wordline_driver 
* No parameters

xwl_driver_509 
+ vdd vss din[509] wl_en wl[509] 
+ wordline_driver 
* No parameters

xwl_driver_510 
+ vdd vss din[510] wl_en wl[510] 
+ wordline_driver 
* No parameters

xwl_driver_511 
+ vdd vss din[511] wl_en wl[511] 
+ wordline_driver 
* No parameters

.ENDS

.SUBCKT bitcell_array 
+ vdd vss bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] wl[511] wl[510] wl[509] wl[508] wl[507] wl[506] wl[505] wl[504] wl[503] wl[502] wl[501] wl[500] wl[499] wl[498] wl[497] wl[496] wl[495] wl[494] wl[493] wl[492] wl[491] wl[490] wl[489] wl[488] wl[487] wl[486] wl[485] wl[484] wl[483] wl[482] wl[481] wl[480] wl[479] wl[478] wl[477] wl[476] wl[475] wl[474] wl[473] wl[472] wl[471] wl[470] wl[469] wl[468] wl[467] wl[466] wl[465] wl[464] wl[463] wl[462] wl[461] wl[460] wl[459] wl[458] wl[457] wl[456] wl[455] wl[454] wl[453] wl[452] wl[451] wl[450] wl[449] wl[448] wl[447] wl[446] wl[445] wl[444] wl[443] wl[442] wl[441] wl[440] wl[439] wl[438] wl[437] wl[436] wl[435] wl[434] wl[433] wl[432] wl[431] wl[430] wl[429] wl[428] wl[427] wl[426] wl[425] wl[424] wl[423] wl[422] wl[421] wl[420] wl[419] wl[418] wl[417] wl[416] wl[415] wl[414] wl[413] wl[412] wl[411] wl[410] wl[409] wl[408] wl[407] wl[406] wl[405] wl[404] wl[403] wl[402] wl[401] wl[400] wl[399] wl[398] wl[397] wl[396] wl[395] wl[394] wl[393] wl[392] wl[391] wl[390] wl[389] wl[388] wl[387] wl[386] wl[385] wl[384] wl[383] wl[382] wl[381] wl[380] wl[379] wl[378] wl[377] wl[376] wl[375] wl[374] wl[373] wl[372] wl[371] wl[370] wl[369] wl[368] wl[367] wl[366] wl[365] wl[364] wl[363] wl[362] wl[361] wl[360] wl[359] wl[358] wl[357] wl[356] wl[355] wl[354] wl[353] wl[352] wl[351] wl[350] wl[349] wl[348] wl[347] wl[346] wl[345] wl[344] wl[343] wl[342] wl[341] wl[340] wl[339] wl[338] wl[337] wl[336] wl[335] wl[334] wl[333] wl[332] wl[331] wl[330] wl[329] wl[328] wl[327] wl[326] wl[325] wl[324] wl[323] wl[322] wl[321] wl[320] wl[319] wl[318] wl[317] wl[316] wl[315] wl[314] wl[313] wl[312] wl[311] wl[310] wl[309] wl[308] wl[307] wl[306] wl[305] wl[304] wl[303] wl[302] wl[301] wl[300] wl[299] wl[298] wl[297] wl[296] wl[295] wl[294] wl[293] wl[292] wl[291] wl[290] wl[289] wl[288] wl[287] wl[286] wl[285] wl[284] wl[283] wl[282] wl[281] wl[280] wl[279] wl[278] wl[277] wl[276] wl[275] wl[274] wl[273] wl[272] wl[271] wl[270] wl[269] wl[268] wl[267] wl[266] wl[265] wl[264] wl[263] wl[262] wl[261] wl[260] wl[259] wl[258] wl[257] wl[256] wl[255] wl[254] wl[253] wl[252] wl[251] wl[250] wl[249] wl[248] wl[247] wl[246] wl[245] wl[244] wl[243] wl[242] wl[241] wl[240] wl[239] wl[238] wl[237] wl[236] wl[235] wl[234] wl[233] wl[232] wl[231] wl[230] wl[229] wl[228] wl[227] wl[226] wl[225] wl[224] wl[223] wl[222] wl[221] wl[220] wl[219] wl[218] wl[217] wl[216] wl[215] wl[214] wl[213] wl[212] wl[211] wl[210] wl[209] wl[208] wl[207] wl[206] wl[205] wl[204] wl[203] wl[202] wl[201] wl[200] wl[199] wl[198] wl[197] wl[196] wl[195] wl[194] wl[193] wl[192] wl[191] wl[190] wl[189] wl[188] wl[187] wl[186] wl[185] wl[184] wl[183] wl[182] wl[181] wl[180] wl[179] wl[178] wl[177] wl[176] wl[175] wl[174] wl[173] wl[172] wl[171] wl[170] wl[169] wl[168] wl[167] wl[166] wl[165] wl[164] wl[163] wl[162] wl[161] wl[160] wl[159] wl[158] wl[157] wl[156] wl[155] wl[154] wl[153] wl[152] wl[151] wl[150] wl[149] wl[148] wl[147] wl[146] wl[145] wl[144] wl[143] wl[142] wl[141] wl[140] wl[139] wl[138] wl[137] wl[136] wl[135] wl[134] wl[133] wl[132] wl[131] wl[130] wl[129] wl[128] wl[127] wl[126] wl[125] wl[124] wl[123] wl[122] wl[121] wl[120] wl[119] wl[118] wl[117] wl[116] wl[115] wl[114] wl[113] wl[112] wl[111] wl[110] wl[109] wl[108] wl[107] wl[106] wl[105] wl[104] wl[103] wl[102] wl[101] wl[100] wl[99] wl[98] wl[97] wl[96] wl[95] wl[94] wl[93] wl[92] wl[91] wl[90] wl[89] wl[88] wl[87] wl[86] wl[85] wl[84] wl[83] wl[82] wl[81] wl[80] wl[79] wl[78] wl[77] wl[76] wl[75] wl[74] wl[73] wl[72] wl[71] wl[70] wl[69] wl[68] wl[67] wl[66] wl[65] wl[64] wl[63] wl[62] wl[61] wl[60] wl[59] wl[58] wl[57] wl[56] wl[55] wl[54] wl[53] wl[52] wl[51] wl[50] wl[49] wl[48] wl[47] wl[46] wl[45] wl[44] wl[43] wl[42] wl[41] wl[40] wl[39] wl[38] wl[37] wl[36] wl[35] wl[34] wl[33] wl[32] wl[31] wl[30] wl[29] wl[28] wl[27] wl[26] wl[25] wl[24] wl[23] wl[22] wl[21] wl[20] wl[19] wl[18] wl[17] wl[16] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] vnb vpb rbl rbr 

xbitcell_0_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_66 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_0_67 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_66 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_1_67 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_0 
+ vdd vdd vss vdd vpb vnb wl[0] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_2_1 
+ rbl rbr vss vdd vpb vnb wl[0] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_2_2 
+ bl[0] br[0] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_3 
+ bl[1] br[1] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_4 
+ bl[2] br[2] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_5 
+ bl[3] br[3] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_6 
+ bl[4] br[4] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_7 
+ bl[5] br[5] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_8 
+ bl[6] br[6] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_9 
+ bl[7] br[7] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_10 
+ bl[8] br[8] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_11 
+ bl[9] br[9] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_12 
+ bl[10] br[10] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_13 
+ bl[11] br[11] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_14 
+ bl[12] br[12] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_15 
+ bl[13] br[13] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_16 
+ bl[14] br[14] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_17 
+ bl[15] br[15] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_18 
+ bl[16] br[16] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_19 
+ bl[17] br[17] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_20 
+ bl[18] br[18] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_21 
+ bl[19] br[19] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_22 
+ bl[20] br[20] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_23 
+ bl[21] br[21] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_24 
+ bl[22] br[22] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_25 
+ bl[23] br[23] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_26 
+ bl[24] br[24] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_27 
+ bl[25] br[25] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_28 
+ bl[26] br[26] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_29 
+ bl[27] br[27] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_30 
+ bl[28] br[28] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_31 
+ bl[29] br[29] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_32 
+ bl[30] br[30] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_33 
+ bl[31] br[31] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_34 
+ bl[32] br[32] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_35 
+ bl[33] br[33] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_36 
+ bl[34] br[34] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_37 
+ bl[35] br[35] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_38 
+ bl[36] br[36] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_39 
+ bl[37] br[37] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_40 
+ bl[38] br[38] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_41 
+ bl[39] br[39] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_42 
+ bl[40] br[40] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_43 
+ bl[41] br[41] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_44 
+ bl[42] br[42] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_45 
+ bl[43] br[43] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_46 
+ bl[44] br[44] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_47 
+ bl[45] br[45] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_48 
+ bl[46] br[46] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_49 
+ bl[47] br[47] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_50 
+ bl[48] br[48] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_51 
+ bl[49] br[49] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_52 
+ bl[50] br[50] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_53 
+ bl[51] br[51] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_54 
+ bl[52] br[52] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_55 
+ bl[53] br[53] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_56 
+ bl[54] br[54] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_57 
+ bl[55] br[55] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_58 
+ bl[56] br[56] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_59 
+ bl[57] br[57] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_60 
+ bl[58] br[58] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_61 
+ bl[59] br[59] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_62 
+ bl[60] br[60] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_63 
+ bl[61] br[61] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_64 
+ bl[62] br[62] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_65 
+ bl[63] br[63] vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_66 
+ vdd vdd vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_2_67 
+ vdd vdd vdd vss wl[0] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_0 
+ vdd vdd vss vdd vpb vnb wl[1] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_3_1 
+ rbl rbr vss vdd vpb vnb wl[1] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_3_2 
+ bl[0] br[0] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_3 
+ bl[1] br[1] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_4 
+ bl[2] br[2] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_5 
+ bl[3] br[3] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_6 
+ bl[4] br[4] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_7 
+ bl[5] br[5] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_8 
+ bl[6] br[6] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_9 
+ bl[7] br[7] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_10 
+ bl[8] br[8] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_11 
+ bl[9] br[9] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_12 
+ bl[10] br[10] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_13 
+ bl[11] br[11] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_14 
+ bl[12] br[12] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_15 
+ bl[13] br[13] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_16 
+ bl[14] br[14] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_17 
+ bl[15] br[15] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_18 
+ bl[16] br[16] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_19 
+ bl[17] br[17] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_20 
+ bl[18] br[18] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_21 
+ bl[19] br[19] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_22 
+ bl[20] br[20] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_23 
+ bl[21] br[21] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_24 
+ bl[22] br[22] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_25 
+ bl[23] br[23] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_26 
+ bl[24] br[24] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_27 
+ bl[25] br[25] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_28 
+ bl[26] br[26] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_29 
+ bl[27] br[27] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_30 
+ bl[28] br[28] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_31 
+ bl[29] br[29] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_32 
+ bl[30] br[30] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_33 
+ bl[31] br[31] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_34 
+ bl[32] br[32] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_35 
+ bl[33] br[33] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_36 
+ bl[34] br[34] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_37 
+ bl[35] br[35] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_38 
+ bl[36] br[36] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_39 
+ bl[37] br[37] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_40 
+ bl[38] br[38] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_41 
+ bl[39] br[39] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_42 
+ bl[40] br[40] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_43 
+ bl[41] br[41] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_44 
+ bl[42] br[42] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_45 
+ bl[43] br[43] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_46 
+ bl[44] br[44] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_47 
+ bl[45] br[45] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_48 
+ bl[46] br[46] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_49 
+ bl[47] br[47] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_50 
+ bl[48] br[48] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_51 
+ bl[49] br[49] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_52 
+ bl[50] br[50] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_53 
+ bl[51] br[51] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_54 
+ bl[52] br[52] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_55 
+ bl[53] br[53] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_56 
+ bl[54] br[54] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_57 
+ bl[55] br[55] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_58 
+ bl[56] br[56] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_59 
+ bl[57] br[57] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_60 
+ bl[58] br[58] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_61 
+ bl[59] br[59] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_62 
+ bl[60] br[60] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_63 
+ bl[61] br[61] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_64 
+ bl[62] br[62] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_65 
+ bl[63] br[63] vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_66 
+ vdd vdd vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_3_67 
+ vdd vdd vdd vss wl[1] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_0 
+ vdd vdd vss vdd vpb vnb wl[2] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_4_1 
+ rbl rbr vss vdd vpb vnb wl[2] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_4_2 
+ bl[0] br[0] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_3 
+ bl[1] br[1] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_4 
+ bl[2] br[2] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_5 
+ bl[3] br[3] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_6 
+ bl[4] br[4] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_7 
+ bl[5] br[5] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_8 
+ bl[6] br[6] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_9 
+ bl[7] br[7] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_10 
+ bl[8] br[8] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_11 
+ bl[9] br[9] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_12 
+ bl[10] br[10] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_13 
+ bl[11] br[11] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_14 
+ bl[12] br[12] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_15 
+ bl[13] br[13] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_16 
+ bl[14] br[14] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_17 
+ bl[15] br[15] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_18 
+ bl[16] br[16] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_19 
+ bl[17] br[17] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_20 
+ bl[18] br[18] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_21 
+ bl[19] br[19] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_22 
+ bl[20] br[20] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_23 
+ bl[21] br[21] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_24 
+ bl[22] br[22] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_25 
+ bl[23] br[23] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_26 
+ bl[24] br[24] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_27 
+ bl[25] br[25] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_28 
+ bl[26] br[26] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_29 
+ bl[27] br[27] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_30 
+ bl[28] br[28] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_31 
+ bl[29] br[29] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_32 
+ bl[30] br[30] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_33 
+ bl[31] br[31] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_34 
+ bl[32] br[32] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_35 
+ bl[33] br[33] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_36 
+ bl[34] br[34] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_37 
+ bl[35] br[35] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_38 
+ bl[36] br[36] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_39 
+ bl[37] br[37] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_40 
+ bl[38] br[38] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_41 
+ bl[39] br[39] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_42 
+ bl[40] br[40] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_43 
+ bl[41] br[41] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_44 
+ bl[42] br[42] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_45 
+ bl[43] br[43] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_46 
+ bl[44] br[44] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_47 
+ bl[45] br[45] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_48 
+ bl[46] br[46] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_49 
+ bl[47] br[47] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_50 
+ bl[48] br[48] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_51 
+ bl[49] br[49] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_52 
+ bl[50] br[50] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_53 
+ bl[51] br[51] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_54 
+ bl[52] br[52] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_55 
+ bl[53] br[53] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_56 
+ bl[54] br[54] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_57 
+ bl[55] br[55] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_58 
+ bl[56] br[56] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_59 
+ bl[57] br[57] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_60 
+ bl[58] br[58] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_61 
+ bl[59] br[59] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_62 
+ bl[60] br[60] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_63 
+ bl[61] br[61] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_64 
+ bl[62] br[62] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_65 
+ bl[63] br[63] vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_66 
+ vdd vdd vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_4_67 
+ vdd vdd vdd vss wl[2] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_0 
+ vdd vdd vss vdd vpb vnb wl[3] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_5_1 
+ rbl rbr vss vdd vpb vnb wl[3] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_5_2 
+ bl[0] br[0] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_3 
+ bl[1] br[1] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_4 
+ bl[2] br[2] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_5 
+ bl[3] br[3] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_6 
+ bl[4] br[4] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_7 
+ bl[5] br[5] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_8 
+ bl[6] br[6] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_9 
+ bl[7] br[7] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_10 
+ bl[8] br[8] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_11 
+ bl[9] br[9] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_12 
+ bl[10] br[10] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_13 
+ bl[11] br[11] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_14 
+ bl[12] br[12] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_15 
+ bl[13] br[13] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_16 
+ bl[14] br[14] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_17 
+ bl[15] br[15] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_18 
+ bl[16] br[16] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_19 
+ bl[17] br[17] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_20 
+ bl[18] br[18] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_21 
+ bl[19] br[19] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_22 
+ bl[20] br[20] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_23 
+ bl[21] br[21] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_24 
+ bl[22] br[22] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_25 
+ bl[23] br[23] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_26 
+ bl[24] br[24] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_27 
+ bl[25] br[25] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_28 
+ bl[26] br[26] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_29 
+ bl[27] br[27] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_30 
+ bl[28] br[28] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_31 
+ bl[29] br[29] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_32 
+ bl[30] br[30] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_33 
+ bl[31] br[31] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_34 
+ bl[32] br[32] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_35 
+ bl[33] br[33] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_36 
+ bl[34] br[34] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_37 
+ bl[35] br[35] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_38 
+ bl[36] br[36] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_39 
+ bl[37] br[37] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_40 
+ bl[38] br[38] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_41 
+ bl[39] br[39] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_42 
+ bl[40] br[40] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_43 
+ bl[41] br[41] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_44 
+ bl[42] br[42] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_45 
+ bl[43] br[43] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_46 
+ bl[44] br[44] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_47 
+ bl[45] br[45] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_48 
+ bl[46] br[46] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_49 
+ bl[47] br[47] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_50 
+ bl[48] br[48] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_51 
+ bl[49] br[49] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_52 
+ bl[50] br[50] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_53 
+ bl[51] br[51] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_54 
+ bl[52] br[52] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_55 
+ bl[53] br[53] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_56 
+ bl[54] br[54] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_57 
+ bl[55] br[55] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_58 
+ bl[56] br[56] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_59 
+ bl[57] br[57] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_60 
+ bl[58] br[58] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_61 
+ bl[59] br[59] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_62 
+ bl[60] br[60] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_63 
+ bl[61] br[61] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_64 
+ bl[62] br[62] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_65 
+ bl[63] br[63] vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_66 
+ vdd vdd vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_5_67 
+ vdd vdd vdd vss wl[3] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_0 
+ vdd vdd vss vdd vpb vnb wl[4] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_6_1 
+ rbl rbr vss vdd vpb vnb wl[4] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_6_2 
+ bl[0] br[0] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_3 
+ bl[1] br[1] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_4 
+ bl[2] br[2] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_5 
+ bl[3] br[3] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_6 
+ bl[4] br[4] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_7 
+ bl[5] br[5] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_8 
+ bl[6] br[6] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_9 
+ bl[7] br[7] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_10 
+ bl[8] br[8] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_11 
+ bl[9] br[9] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_12 
+ bl[10] br[10] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_13 
+ bl[11] br[11] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_14 
+ bl[12] br[12] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_15 
+ bl[13] br[13] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_16 
+ bl[14] br[14] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_17 
+ bl[15] br[15] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_18 
+ bl[16] br[16] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_19 
+ bl[17] br[17] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_20 
+ bl[18] br[18] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_21 
+ bl[19] br[19] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_22 
+ bl[20] br[20] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_23 
+ bl[21] br[21] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_24 
+ bl[22] br[22] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_25 
+ bl[23] br[23] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_26 
+ bl[24] br[24] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_27 
+ bl[25] br[25] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_28 
+ bl[26] br[26] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_29 
+ bl[27] br[27] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_30 
+ bl[28] br[28] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_31 
+ bl[29] br[29] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_32 
+ bl[30] br[30] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_33 
+ bl[31] br[31] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_34 
+ bl[32] br[32] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_35 
+ bl[33] br[33] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_36 
+ bl[34] br[34] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_37 
+ bl[35] br[35] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_38 
+ bl[36] br[36] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_39 
+ bl[37] br[37] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_40 
+ bl[38] br[38] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_41 
+ bl[39] br[39] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_42 
+ bl[40] br[40] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_43 
+ bl[41] br[41] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_44 
+ bl[42] br[42] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_45 
+ bl[43] br[43] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_46 
+ bl[44] br[44] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_47 
+ bl[45] br[45] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_48 
+ bl[46] br[46] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_49 
+ bl[47] br[47] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_50 
+ bl[48] br[48] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_51 
+ bl[49] br[49] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_52 
+ bl[50] br[50] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_53 
+ bl[51] br[51] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_54 
+ bl[52] br[52] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_55 
+ bl[53] br[53] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_56 
+ bl[54] br[54] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_57 
+ bl[55] br[55] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_58 
+ bl[56] br[56] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_59 
+ bl[57] br[57] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_60 
+ bl[58] br[58] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_61 
+ bl[59] br[59] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_62 
+ bl[60] br[60] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_63 
+ bl[61] br[61] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_64 
+ bl[62] br[62] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_65 
+ bl[63] br[63] vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_66 
+ vdd vdd vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_6_67 
+ vdd vdd vdd vss wl[4] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_0 
+ vdd vdd vss vdd vpb vnb wl[5] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_7_1 
+ rbl rbr vss vdd vpb vnb wl[5] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_7_2 
+ bl[0] br[0] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_3 
+ bl[1] br[1] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_4 
+ bl[2] br[2] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_5 
+ bl[3] br[3] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_6 
+ bl[4] br[4] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_7 
+ bl[5] br[5] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_8 
+ bl[6] br[6] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_9 
+ bl[7] br[7] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_10 
+ bl[8] br[8] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_11 
+ bl[9] br[9] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_12 
+ bl[10] br[10] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_13 
+ bl[11] br[11] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_14 
+ bl[12] br[12] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_15 
+ bl[13] br[13] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_16 
+ bl[14] br[14] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_17 
+ bl[15] br[15] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_18 
+ bl[16] br[16] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_19 
+ bl[17] br[17] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_20 
+ bl[18] br[18] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_21 
+ bl[19] br[19] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_22 
+ bl[20] br[20] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_23 
+ bl[21] br[21] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_24 
+ bl[22] br[22] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_25 
+ bl[23] br[23] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_26 
+ bl[24] br[24] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_27 
+ bl[25] br[25] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_28 
+ bl[26] br[26] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_29 
+ bl[27] br[27] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_30 
+ bl[28] br[28] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_31 
+ bl[29] br[29] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_32 
+ bl[30] br[30] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_33 
+ bl[31] br[31] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_34 
+ bl[32] br[32] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_35 
+ bl[33] br[33] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_36 
+ bl[34] br[34] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_37 
+ bl[35] br[35] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_38 
+ bl[36] br[36] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_39 
+ bl[37] br[37] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_40 
+ bl[38] br[38] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_41 
+ bl[39] br[39] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_42 
+ bl[40] br[40] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_43 
+ bl[41] br[41] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_44 
+ bl[42] br[42] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_45 
+ bl[43] br[43] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_46 
+ bl[44] br[44] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_47 
+ bl[45] br[45] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_48 
+ bl[46] br[46] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_49 
+ bl[47] br[47] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_50 
+ bl[48] br[48] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_51 
+ bl[49] br[49] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_52 
+ bl[50] br[50] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_53 
+ bl[51] br[51] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_54 
+ bl[52] br[52] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_55 
+ bl[53] br[53] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_56 
+ bl[54] br[54] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_57 
+ bl[55] br[55] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_58 
+ bl[56] br[56] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_59 
+ bl[57] br[57] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_60 
+ bl[58] br[58] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_61 
+ bl[59] br[59] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_62 
+ bl[60] br[60] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_63 
+ bl[61] br[61] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_64 
+ bl[62] br[62] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_65 
+ bl[63] br[63] vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_66 
+ vdd vdd vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_7_67 
+ vdd vdd vdd vss wl[5] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_0 
+ vdd vdd vss vdd vpb vnb wl[6] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_8_1 
+ rbl rbr vss vdd vpb vnb wl[6] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_8_2 
+ bl[0] br[0] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_3 
+ bl[1] br[1] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_4 
+ bl[2] br[2] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_5 
+ bl[3] br[3] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_6 
+ bl[4] br[4] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_7 
+ bl[5] br[5] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_8 
+ bl[6] br[6] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_9 
+ bl[7] br[7] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_10 
+ bl[8] br[8] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_11 
+ bl[9] br[9] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_12 
+ bl[10] br[10] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_13 
+ bl[11] br[11] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_14 
+ bl[12] br[12] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_15 
+ bl[13] br[13] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_16 
+ bl[14] br[14] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_17 
+ bl[15] br[15] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_18 
+ bl[16] br[16] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_19 
+ bl[17] br[17] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_20 
+ bl[18] br[18] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_21 
+ bl[19] br[19] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_22 
+ bl[20] br[20] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_23 
+ bl[21] br[21] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_24 
+ bl[22] br[22] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_25 
+ bl[23] br[23] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_26 
+ bl[24] br[24] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_27 
+ bl[25] br[25] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_28 
+ bl[26] br[26] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_29 
+ bl[27] br[27] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_30 
+ bl[28] br[28] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_31 
+ bl[29] br[29] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_32 
+ bl[30] br[30] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_33 
+ bl[31] br[31] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_34 
+ bl[32] br[32] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_35 
+ bl[33] br[33] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_36 
+ bl[34] br[34] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_37 
+ bl[35] br[35] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_38 
+ bl[36] br[36] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_39 
+ bl[37] br[37] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_40 
+ bl[38] br[38] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_41 
+ bl[39] br[39] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_42 
+ bl[40] br[40] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_43 
+ bl[41] br[41] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_44 
+ bl[42] br[42] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_45 
+ bl[43] br[43] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_46 
+ bl[44] br[44] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_47 
+ bl[45] br[45] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_48 
+ bl[46] br[46] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_49 
+ bl[47] br[47] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_50 
+ bl[48] br[48] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_51 
+ bl[49] br[49] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_52 
+ bl[50] br[50] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_53 
+ bl[51] br[51] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_54 
+ bl[52] br[52] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_55 
+ bl[53] br[53] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_56 
+ bl[54] br[54] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_57 
+ bl[55] br[55] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_58 
+ bl[56] br[56] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_59 
+ bl[57] br[57] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_60 
+ bl[58] br[58] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_61 
+ bl[59] br[59] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_62 
+ bl[60] br[60] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_63 
+ bl[61] br[61] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_64 
+ bl[62] br[62] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_65 
+ bl[63] br[63] vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_66 
+ vdd vdd vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_8_67 
+ vdd vdd vdd vss wl[6] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_0 
+ vdd vdd vss vdd vpb vnb wl[7] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_9_1 
+ rbl rbr vss vdd vpb vnb wl[7] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_9_2 
+ bl[0] br[0] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_3 
+ bl[1] br[1] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_4 
+ bl[2] br[2] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_5 
+ bl[3] br[3] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_6 
+ bl[4] br[4] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_7 
+ bl[5] br[5] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_8 
+ bl[6] br[6] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_9 
+ bl[7] br[7] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_10 
+ bl[8] br[8] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_11 
+ bl[9] br[9] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_12 
+ bl[10] br[10] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_13 
+ bl[11] br[11] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_14 
+ bl[12] br[12] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_15 
+ bl[13] br[13] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_16 
+ bl[14] br[14] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_17 
+ bl[15] br[15] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_18 
+ bl[16] br[16] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_19 
+ bl[17] br[17] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_20 
+ bl[18] br[18] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_21 
+ bl[19] br[19] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_22 
+ bl[20] br[20] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_23 
+ bl[21] br[21] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_24 
+ bl[22] br[22] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_25 
+ bl[23] br[23] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_26 
+ bl[24] br[24] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_27 
+ bl[25] br[25] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_28 
+ bl[26] br[26] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_29 
+ bl[27] br[27] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_30 
+ bl[28] br[28] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_31 
+ bl[29] br[29] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_32 
+ bl[30] br[30] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_33 
+ bl[31] br[31] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_34 
+ bl[32] br[32] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_35 
+ bl[33] br[33] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_36 
+ bl[34] br[34] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_37 
+ bl[35] br[35] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_38 
+ bl[36] br[36] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_39 
+ bl[37] br[37] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_40 
+ bl[38] br[38] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_41 
+ bl[39] br[39] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_42 
+ bl[40] br[40] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_43 
+ bl[41] br[41] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_44 
+ bl[42] br[42] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_45 
+ bl[43] br[43] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_46 
+ bl[44] br[44] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_47 
+ bl[45] br[45] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_48 
+ bl[46] br[46] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_49 
+ bl[47] br[47] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_50 
+ bl[48] br[48] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_51 
+ bl[49] br[49] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_52 
+ bl[50] br[50] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_53 
+ bl[51] br[51] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_54 
+ bl[52] br[52] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_55 
+ bl[53] br[53] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_56 
+ bl[54] br[54] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_57 
+ bl[55] br[55] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_58 
+ bl[56] br[56] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_59 
+ bl[57] br[57] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_60 
+ bl[58] br[58] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_61 
+ bl[59] br[59] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_62 
+ bl[60] br[60] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_63 
+ bl[61] br[61] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_64 
+ bl[62] br[62] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_65 
+ bl[63] br[63] vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_66 
+ vdd vdd vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_9_67 
+ vdd vdd vdd vss wl[7] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_0 
+ vdd vdd vss vdd vpb vnb wl[8] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_10_1 
+ rbl rbr vss vdd vpb vnb wl[8] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_10_2 
+ bl[0] br[0] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_3 
+ bl[1] br[1] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_4 
+ bl[2] br[2] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_5 
+ bl[3] br[3] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_6 
+ bl[4] br[4] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_7 
+ bl[5] br[5] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_8 
+ bl[6] br[6] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_9 
+ bl[7] br[7] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_10 
+ bl[8] br[8] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_11 
+ bl[9] br[9] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_12 
+ bl[10] br[10] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_13 
+ bl[11] br[11] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_14 
+ bl[12] br[12] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_15 
+ bl[13] br[13] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_16 
+ bl[14] br[14] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_17 
+ bl[15] br[15] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_18 
+ bl[16] br[16] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_19 
+ bl[17] br[17] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_20 
+ bl[18] br[18] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_21 
+ bl[19] br[19] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_22 
+ bl[20] br[20] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_23 
+ bl[21] br[21] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_24 
+ bl[22] br[22] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_25 
+ bl[23] br[23] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_26 
+ bl[24] br[24] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_27 
+ bl[25] br[25] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_28 
+ bl[26] br[26] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_29 
+ bl[27] br[27] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_30 
+ bl[28] br[28] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_31 
+ bl[29] br[29] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_32 
+ bl[30] br[30] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_33 
+ bl[31] br[31] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_34 
+ bl[32] br[32] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_35 
+ bl[33] br[33] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_36 
+ bl[34] br[34] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_37 
+ bl[35] br[35] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_38 
+ bl[36] br[36] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_39 
+ bl[37] br[37] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_40 
+ bl[38] br[38] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_41 
+ bl[39] br[39] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_42 
+ bl[40] br[40] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_43 
+ bl[41] br[41] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_44 
+ bl[42] br[42] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_45 
+ bl[43] br[43] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_46 
+ bl[44] br[44] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_47 
+ bl[45] br[45] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_48 
+ bl[46] br[46] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_49 
+ bl[47] br[47] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_50 
+ bl[48] br[48] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_51 
+ bl[49] br[49] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_52 
+ bl[50] br[50] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_53 
+ bl[51] br[51] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_54 
+ bl[52] br[52] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_55 
+ bl[53] br[53] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_56 
+ bl[54] br[54] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_57 
+ bl[55] br[55] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_58 
+ bl[56] br[56] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_59 
+ bl[57] br[57] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_60 
+ bl[58] br[58] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_61 
+ bl[59] br[59] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_62 
+ bl[60] br[60] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_63 
+ bl[61] br[61] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_64 
+ bl[62] br[62] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_65 
+ bl[63] br[63] vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_66 
+ vdd vdd vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_10_67 
+ vdd vdd vdd vss wl[8] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_0 
+ vdd vdd vss vdd vpb vnb wl[9] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_11_1 
+ rbl rbr vss vdd vpb vnb wl[9] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_11_2 
+ bl[0] br[0] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_3 
+ bl[1] br[1] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_4 
+ bl[2] br[2] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_5 
+ bl[3] br[3] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_6 
+ bl[4] br[4] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_7 
+ bl[5] br[5] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_8 
+ bl[6] br[6] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_9 
+ bl[7] br[7] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_10 
+ bl[8] br[8] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_11 
+ bl[9] br[9] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_12 
+ bl[10] br[10] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_13 
+ bl[11] br[11] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_14 
+ bl[12] br[12] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_15 
+ bl[13] br[13] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_16 
+ bl[14] br[14] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_17 
+ bl[15] br[15] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_18 
+ bl[16] br[16] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_19 
+ bl[17] br[17] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_20 
+ bl[18] br[18] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_21 
+ bl[19] br[19] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_22 
+ bl[20] br[20] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_23 
+ bl[21] br[21] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_24 
+ bl[22] br[22] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_25 
+ bl[23] br[23] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_26 
+ bl[24] br[24] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_27 
+ bl[25] br[25] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_28 
+ bl[26] br[26] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_29 
+ bl[27] br[27] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_30 
+ bl[28] br[28] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_31 
+ bl[29] br[29] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_32 
+ bl[30] br[30] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_33 
+ bl[31] br[31] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_34 
+ bl[32] br[32] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_35 
+ bl[33] br[33] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_36 
+ bl[34] br[34] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_37 
+ bl[35] br[35] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_38 
+ bl[36] br[36] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_39 
+ bl[37] br[37] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_40 
+ bl[38] br[38] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_41 
+ bl[39] br[39] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_42 
+ bl[40] br[40] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_43 
+ bl[41] br[41] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_44 
+ bl[42] br[42] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_45 
+ bl[43] br[43] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_46 
+ bl[44] br[44] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_47 
+ bl[45] br[45] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_48 
+ bl[46] br[46] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_49 
+ bl[47] br[47] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_50 
+ bl[48] br[48] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_51 
+ bl[49] br[49] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_52 
+ bl[50] br[50] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_53 
+ bl[51] br[51] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_54 
+ bl[52] br[52] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_55 
+ bl[53] br[53] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_56 
+ bl[54] br[54] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_57 
+ bl[55] br[55] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_58 
+ bl[56] br[56] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_59 
+ bl[57] br[57] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_60 
+ bl[58] br[58] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_61 
+ bl[59] br[59] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_62 
+ bl[60] br[60] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_63 
+ bl[61] br[61] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_64 
+ bl[62] br[62] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_65 
+ bl[63] br[63] vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_66 
+ vdd vdd vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_11_67 
+ vdd vdd vdd vss wl[9] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_0 
+ vdd vdd vss vdd vpb vnb wl[10] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_12_1 
+ rbl rbr vss vdd vpb vnb wl[10] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_12_2 
+ bl[0] br[0] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_3 
+ bl[1] br[1] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_4 
+ bl[2] br[2] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_5 
+ bl[3] br[3] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_6 
+ bl[4] br[4] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_7 
+ bl[5] br[5] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_8 
+ bl[6] br[6] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_9 
+ bl[7] br[7] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_10 
+ bl[8] br[8] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_11 
+ bl[9] br[9] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_12 
+ bl[10] br[10] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_13 
+ bl[11] br[11] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_14 
+ bl[12] br[12] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_15 
+ bl[13] br[13] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_16 
+ bl[14] br[14] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_17 
+ bl[15] br[15] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_18 
+ bl[16] br[16] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_19 
+ bl[17] br[17] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_20 
+ bl[18] br[18] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_21 
+ bl[19] br[19] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_22 
+ bl[20] br[20] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_23 
+ bl[21] br[21] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_24 
+ bl[22] br[22] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_25 
+ bl[23] br[23] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_26 
+ bl[24] br[24] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_27 
+ bl[25] br[25] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_28 
+ bl[26] br[26] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_29 
+ bl[27] br[27] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_30 
+ bl[28] br[28] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_31 
+ bl[29] br[29] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_32 
+ bl[30] br[30] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_33 
+ bl[31] br[31] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_34 
+ bl[32] br[32] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_35 
+ bl[33] br[33] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_36 
+ bl[34] br[34] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_37 
+ bl[35] br[35] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_38 
+ bl[36] br[36] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_39 
+ bl[37] br[37] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_40 
+ bl[38] br[38] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_41 
+ bl[39] br[39] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_42 
+ bl[40] br[40] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_43 
+ bl[41] br[41] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_44 
+ bl[42] br[42] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_45 
+ bl[43] br[43] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_46 
+ bl[44] br[44] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_47 
+ bl[45] br[45] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_48 
+ bl[46] br[46] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_49 
+ bl[47] br[47] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_50 
+ bl[48] br[48] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_51 
+ bl[49] br[49] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_52 
+ bl[50] br[50] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_53 
+ bl[51] br[51] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_54 
+ bl[52] br[52] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_55 
+ bl[53] br[53] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_56 
+ bl[54] br[54] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_57 
+ bl[55] br[55] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_58 
+ bl[56] br[56] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_59 
+ bl[57] br[57] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_60 
+ bl[58] br[58] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_61 
+ bl[59] br[59] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_62 
+ bl[60] br[60] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_63 
+ bl[61] br[61] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_64 
+ bl[62] br[62] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_65 
+ bl[63] br[63] vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_66 
+ vdd vdd vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_12_67 
+ vdd vdd vdd vss wl[10] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_0 
+ vdd vdd vss vdd vpb vnb wl[11] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_13_1 
+ rbl rbr vss vdd vpb vnb wl[11] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_13_2 
+ bl[0] br[0] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_3 
+ bl[1] br[1] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_4 
+ bl[2] br[2] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_5 
+ bl[3] br[3] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_6 
+ bl[4] br[4] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_7 
+ bl[5] br[5] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_8 
+ bl[6] br[6] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_9 
+ bl[7] br[7] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_10 
+ bl[8] br[8] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_11 
+ bl[9] br[9] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_12 
+ bl[10] br[10] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_13 
+ bl[11] br[11] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_14 
+ bl[12] br[12] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_15 
+ bl[13] br[13] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_16 
+ bl[14] br[14] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_17 
+ bl[15] br[15] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_18 
+ bl[16] br[16] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_19 
+ bl[17] br[17] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_20 
+ bl[18] br[18] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_21 
+ bl[19] br[19] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_22 
+ bl[20] br[20] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_23 
+ bl[21] br[21] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_24 
+ bl[22] br[22] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_25 
+ bl[23] br[23] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_26 
+ bl[24] br[24] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_27 
+ bl[25] br[25] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_28 
+ bl[26] br[26] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_29 
+ bl[27] br[27] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_30 
+ bl[28] br[28] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_31 
+ bl[29] br[29] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_32 
+ bl[30] br[30] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_33 
+ bl[31] br[31] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_34 
+ bl[32] br[32] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_35 
+ bl[33] br[33] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_36 
+ bl[34] br[34] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_37 
+ bl[35] br[35] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_38 
+ bl[36] br[36] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_39 
+ bl[37] br[37] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_40 
+ bl[38] br[38] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_41 
+ bl[39] br[39] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_42 
+ bl[40] br[40] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_43 
+ bl[41] br[41] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_44 
+ bl[42] br[42] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_45 
+ bl[43] br[43] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_46 
+ bl[44] br[44] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_47 
+ bl[45] br[45] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_48 
+ bl[46] br[46] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_49 
+ bl[47] br[47] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_50 
+ bl[48] br[48] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_51 
+ bl[49] br[49] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_52 
+ bl[50] br[50] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_53 
+ bl[51] br[51] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_54 
+ bl[52] br[52] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_55 
+ bl[53] br[53] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_56 
+ bl[54] br[54] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_57 
+ bl[55] br[55] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_58 
+ bl[56] br[56] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_59 
+ bl[57] br[57] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_60 
+ bl[58] br[58] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_61 
+ bl[59] br[59] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_62 
+ bl[60] br[60] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_63 
+ bl[61] br[61] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_64 
+ bl[62] br[62] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_65 
+ bl[63] br[63] vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_66 
+ vdd vdd vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_13_67 
+ vdd vdd vdd vss wl[11] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_0 
+ vdd vdd vss vdd vpb vnb wl[12] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_14_1 
+ rbl rbr vss vdd vpb vnb wl[12] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_14_2 
+ bl[0] br[0] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_3 
+ bl[1] br[1] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_4 
+ bl[2] br[2] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_5 
+ bl[3] br[3] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_6 
+ bl[4] br[4] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_7 
+ bl[5] br[5] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_8 
+ bl[6] br[6] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_9 
+ bl[7] br[7] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_10 
+ bl[8] br[8] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_11 
+ bl[9] br[9] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_12 
+ bl[10] br[10] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_13 
+ bl[11] br[11] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_14 
+ bl[12] br[12] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_15 
+ bl[13] br[13] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_16 
+ bl[14] br[14] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_17 
+ bl[15] br[15] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_18 
+ bl[16] br[16] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_19 
+ bl[17] br[17] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_20 
+ bl[18] br[18] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_21 
+ bl[19] br[19] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_22 
+ bl[20] br[20] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_23 
+ bl[21] br[21] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_24 
+ bl[22] br[22] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_25 
+ bl[23] br[23] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_26 
+ bl[24] br[24] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_27 
+ bl[25] br[25] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_28 
+ bl[26] br[26] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_29 
+ bl[27] br[27] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_30 
+ bl[28] br[28] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_31 
+ bl[29] br[29] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_32 
+ bl[30] br[30] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_33 
+ bl[31] br[31] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_34 
+ bl[32] br[32] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_35 
+ bl[33] br[33] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_36 
+ bl[34] br[34] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_37 
+ bl[35] br[35] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_38 
+ bl[36] br[36] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_39 
+ bl[37] br[37] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_40 
+ bl[38] br[38] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_41 
+ bl[39] br[39] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_42 
+ bl[40] br[40] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_43 
+ bl[41] br[41] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_44 
+ bl[42] br[42] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_45 
+ bl[43] br[43] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_46 
+ bl[44] br[44] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_47 
+ bl[45] br[45] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_48 
+ bl[46] br[46] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_49 
+ bl[47] br[47] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_50 
+ bl[48] br[48] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_51 
+ bl[49] br[49] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_52 
+ bl[50] br[50] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_53 
+ bl[51] br[51] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_54 
+ bl[52] br[52] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_55 
+ bl[53] br[53] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_56 
+ bl[54] br[54] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_57 
+ bl[55] br[55] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_58 
+ bl[56] br[56] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_59 
+ bl[57] br[57] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_60 
+ bl[58] br[58] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_61 
+ bl[59] br[59] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_62 
+ bl[60] br[60] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_63 
+ bl[61] br[61] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_64 
+ bl[62] br[62] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_65 
+ bl[63] br[63] vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_66 
+ vdd vdd vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_14_67 
+ vdd vdd vdd vss wl[12] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_0 
+ vdd vdd vss vdd vpb vnb wl[13] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_15_1 
+ rbl rbr vss vdd vpb vnb wl[13] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_15_2 
+ bl[0] br[0] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_3 
+ bl[1] br[1] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_4 
+ bl[2] br[2] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_5 
+ bl[3] br[3] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_6 
+ bl[4] br[4] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_7 
+ bl[5] br[5] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_8 
+ bl[6] br[6] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_9 
+ bl[7] br[7] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_10 
+ bl[8] br[8] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_11 
+ bl[9] br[9] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_12 
+ bl[10] br[10] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_13 
+ bl[11] br[11] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_14 
+ bl[12] br[12] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_15 
+ bl[13] br[13] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_16 
+ bl[14] br[14] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_17 
+ bl[15] br[15] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_18 
+ bl[16] br[16] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_19 
+ bl[17] br[17] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_20 
+ bl[18] br[18] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_21 
+ bl[19] br[19] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_22 
+ bl[20] br[20] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_23 
+ bl[21] br[21] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_24 
+ bl[22] br[22] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_25 
+ bl[23] br[23] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_26 
+ bl[24] br[24] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_27 
+ bl[25] br[25] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_28 
+ bl[26] br[26] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_29 
+ bl[27] br[27] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_30 
+ bl[28] br[28] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_31 
+ bl[29] br[29] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_32 
+ bl[30] br[30] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_33 
+ bl[31] br[31] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_34 
+ bl[32] br[32] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_35 
+ bl[33] br[33] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_36 
+ bl[34] br[34] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_37 
+ bl[35] br[35] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_38 
+ bl[36] br[36] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_39 
+ bl[37] br[37] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_40 
+ bl[38] br[38] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_41 
+ bl[39] br[39] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_42 
+ bl[40] br[40] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_43 
+ bl[41] br[41] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_44 
+ bl[42] br[42] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_45 
+ bl[43] br[43] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_46 
+ bl[44] br[44] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_47 
+ bl[45] br[45] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_48 
+ bl[46] br[46] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_49 
+ bl[47] br[47] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_50 
+ bl[48] br[48] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_51 
+ bl[49] br[49] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_52 
+ bl[50] br[50] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_53 
+ bl[51] br[51] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_54 
+ bl[52] br[52] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_55 
+ bl[53] br[53] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_56 
+ bl[54] br[54] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_57 
+ bl[55] br[55] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_58 
+ bl[56] br[56] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_59 
+ bl[57] br[57] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_60 
+ bl[58] br[58] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_61 
+ bl[59] br[59] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_62 
+ bl[60] br[60] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_63 
+ bl[61] br[61] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_64 
+ bl[62] br[62] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_65 
+ bl[63] br[63] vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_66 
+ vdd vdd vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_15_67 
+ vdd vdd vdd vss wl[13] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_0 
+ vdd vdd vss vdd vpb vnb wl[14] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_16_1 
+ rbl rbr vss vdd vpb vnb wl[14] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_16_2 
+ bl[0] br[0] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_3 
+ bl[1] br[1] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_4 
+ bl[2] br[2] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_5 
+ bl[3] br[3] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_6 
+ bl[4] br[4] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_7 
+ bl[5] br[5] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_8 
+ bl[6] br[6] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_9 
+ bl[7] br[7] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_10 
+ bl[8] br[8] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_11 
+ bl[9] br[9] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_12 
+ bl[10] br[10] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_13 
+ bl[11] br[11] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_14 
+ bl[12] br[12] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_15 
+ bl[13] br[13] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_16 
+ bl[14] br[14] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_17 
+ bl[15] br[15] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_18 
+ bl[16] br[16] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_19 
+ bl[17] br[17] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_20 
+ bl[18] br[18] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_21 
+ bl[19] br[19] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_22 
+ bl[20] br[20] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_23 
+ bl[21] br[21] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_24 
+ bl[22] br[22] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_25 
+ bl[23] br[23] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_26 
+ bl[24] br[24] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_27 
+ bl[25] br[25] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_28 
+ bl[26] br[26] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_29 
+ bl[27] br[27] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_30 
+ bl[28] br[28] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_31 
+ bl[29] br[29] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_32 
+ bl[30] br[30] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_33 
+ bl[31] br[31] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_34 
+ bl[32] br[32] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_35 
+ bl[33] br[33] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_36 
+ bl[34] br[34] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_37 
+ bl[35] br[35] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_38 
+ bl[36] br[36] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_39 
+ bl[37] br[37] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_40 
+ bl[38] br[38] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_41 
+ bl[39] br[39] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_42 
+ bl[40] br[40] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_43 
+ bl[41] br[41] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_44 
+ bl[42] br[42] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_45 
+ bl[43] br[43] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_46 
+ bl[44] br[44] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_47 
+ bl[45] br[45] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_48 
+ bl[46] br[46] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_49 
+ bl[47] br[47] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_50 
+ bl[48] br[48] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_51 
+ bl[49] br[49] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_52 
+ bl[50] br[50] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_53 
+ bl[51] br[51] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_54 
+ bl[52] br[52] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_55 
+ bl[53] br[53] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_56 
+ bl[54] br[54] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_57 
+ bl[55] br[55] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_58 
+ bl[56] br[56] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_59 
+ bl[57] br[57] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_60 
+ bl[58] br[58] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_61 
+ bl[59] br[59] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_62 
+ bl[60] br[60] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_63 
+ bl[61] br[61] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_64 
+ bl[62] br[62] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_65 
+ bl[63] br[63] vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_66 
+ vdd vdd vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_16_67 
+ vdd vdd vdd vss wl[14] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_0 
+ vdd vdd vss vdd vpb vnb wl[15] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_17_1 
+ rbl rbr vss vdd vpb vnb wl[15] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_17_2 
+ bl[0] br[0] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_3 
+ bl[1] br[1] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_4 
+ bl[2] br[2] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_5 
+ bl[3] br[3] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_6 
+ bl[4] br[4] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_7 
+ bl[5] br[5] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_8 
+ bl[6] br[6] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_9 
+ bl[7] br[7] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_10 
+ bl[8] br[8] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_11 
+ bl[9] br[9] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_12 
+ bl[10] br[10] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_13 
+ bl[11] br[11] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_14 
+ bl[12] br[12] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_15 
+ bl[13] br[13] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_16 
+ bl[14] br[14] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_17 
+ bl[15] br[15] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_18 
+ bl[16] br[16] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_19 
+ bl[17] br[17] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_20 
+ bl[18] br[18] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_21 
+ bl[19] br[19] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_22 
+ bl[20] br[20] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_23 
+ bl[21] br[21] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_24 
+ bl[22] br[22] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_25 
+ bl[23] br[23] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_26 
+ bl[24] br[24] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_27 
+ bl[25] br[25] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_28 
+ bl[26] br[26] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_29 
+ bl[27] br[27] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_30 
+ bl[28] br[28] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_31 
+ bl[29] br[29] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_32 
+ bl[30] br[30] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_33 
+ bl[31] br[31] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_34 
+ bl[32] br[32] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_35 
+ bl[33] br[33] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_36 
+ bl[34] br[34] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_37 
+ bl[35] br[35] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_38 
+ bl[36] br[36] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_39 
+ bl[37] br[37] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_40 
+ bl[38] br[38] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_41 
+ bl[39] br[39] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_42 
+ bl[40] br[40] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_43 
+ bl[41] br[41] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_44 
+ bl[42] br[42] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_45 
+ bl[43] br[43] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_46 
+ bl[44] br[44] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_47 
+ bl[45] br[45] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_48 
+ bl[46] br[46] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_49 
+ bl[47] br[47] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_50 
+ bl[48] br[48] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_51 
+ bl[49] br[49] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_52 
+ bl[50] br[50] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_53 
+ bl[51] br[51] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_54 
+ bl[52] br[52] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_55 
+ bl[53] br[53] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_56 
+ bl[54] br[54] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_57 
+ bl[55] br[55] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_58 
+ bl[56] br[56] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_59 
+ bl[57] br[57] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_60 
+ bl[58] br[58] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_61 
+ bl[59] br[59] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_62 
+ bl[60] br[60] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_63 
+ bl[61] br[61] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_64 
+ bl[62] br[62] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_65 
+ bl[63] br[63] vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_66 
+ vdd vdd vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_17_67 
+ vdd vdd vdd vss wl[15] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_0 
+ vdd vdd vss vdd vpb vnb wl[16] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_18_1 
+ rbl rbr vss vdd vpb vnb wl[16] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_18_2 
+ bl[0] br[0] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_3 
+ bl[1] br[1] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_4 
+ bl[2] br[2] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_5 
+ bl[3] br[3] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_6 
+ bl[4] br[4] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_7 
+ bl[5] br[5] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_8 
+ bl[6] br[6] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_9 
+ bl[7] br[7] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_10 
+ bl[8] br[8] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_11 
+ bl[9] br[9] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_12 
+ bl[10] br[10] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_13 
+ bl[11] br[11] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_14 
+ bl[12] br[12] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_15 
+ bl[13] br[13] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_16 
+ bl[14] br[14] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_17 
+ bl[15] br[15] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_18 
+ bl[16] br[16] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_19 
+ bl[17] br[17] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_20 
+ bl[18] br[18] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_21 
+ bl[19] br[19] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_22 
+ bl[20] br[20] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_23 
+ bl[21] br[21] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_24 
+ bl[22] br[22] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_25 
+ bl[23] br[23] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_26 
+ bl[24] br[24] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_27 
+ bl[25] br[25] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_28 
+ bl[26] br[26] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_29 
+ bl[27] br[27] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_30 
+ bl[28] br[28] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_31 
+ bl[29] br[29] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_32 
+ bl[30] br[30] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_33 
+ bl[31] br[31] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_34 
+ bl[32] br[32] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_35 
+ bl[33] br[33] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_36 
+ bl[34] br[34] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_37 
+ bl[35] br[35] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_38 
+ bl[36] br[36] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_39 
+ bl[37] br[37] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_40 
+ bl[38] br[38] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_41 
+ bl[39] br[39] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_42 
+ bl[40] br[40] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_43 
+ bl[41] br[41] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_44 
+ bl[42] br[42] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_45 
+ bl[43] br[43] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_46 
+ bl[44] br[44] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_47 
+ bl[45] br[45] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_48 
+ bl[46] br[46] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_49 
+ bl[47] br[47] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_50 
+ bl[48] br[48] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_51 
+ bl[49] br[49] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_52 
+ bl[50] br[50] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_53 
+ bl[51] br[51] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_54 
+ bl[52] br[52] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_55 
+ bl[53] br[53] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_56 
+ bl[54] br[54] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_57 
+ bl[55] br[55] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_58 
+ bl[56] br[56] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_59 
+ bl[57] br[57] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_60 
+ bl[58] br[58] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_61 
+ bl[59] br[59] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_62 
+ bl[60] br[60] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_63 
+ bl[61] br[61] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_64 
+ bl[62] br[62] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_65 
+ bl[63] br[63] vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_66 
+ vdd vdd vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_18_67 
+ vdd vdd vdd vss wl[16] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_0 
+ vdd vdd vss vdd vpb vnb wl[17] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_19_1 
+ rbl rbr vss vdd vpb vnb wl[17] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_19_2 
+ bl[0] br[0] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_3 
+ bl[1] br[1] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_4 
+ bl[2] br[2] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_5 
+ bl[3] br[3] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_6 
+ bl[4] br[4] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_7 
+ bl[5] br[5] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_8 
+ bl[6] br[6] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_9 
+ bl[7] br[7] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_10 
+ bl[8] br[8] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_11 
+ bl[9] br[9] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_12 
+ bl[10] br[10] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_13 
+ bl[11] br[11] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_14 
+ bl[12] br[12] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_15 
+ bl[13] br[13] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_16 
+ bl[14] br[14] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_17 
+ bl[15] br[15] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_18 
+ bl[16] br[16] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_19 
+ bl[17] br[17] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_20 
+ bl[18] br[18] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_21 
+ bl[19] br[19] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_22 
+ bl[20] br[20] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_23 
+ bl[21] br[21] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_24 
+ bl[22] br[22] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_25 
+ bl[23] br[23] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_26 
+ bl[24] br[24] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_27 
+ bl[25] br[25] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_28 
+ bl[26] br[26] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_29 
+ bl[27] br[27] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_30 
+ bl[28] br[28] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_31 
+ bl[29] br[29] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_32 
+ bl[30] br[30] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_33 
+ bl[31] br[31] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_34 
+ bl[32] br[32] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_35 
+ bl[33] br[33] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_36 
+ bl[34] br[34] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_37 
+ bl[35] br[35] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_38 
+ bl[36] br[36] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_39 
+ bl[37] br[37] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_40 
+ bl[38] br[38] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_41 
+ bl[39] br[39] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_42 
+ bl[40] br[40] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_43 
+ bl[41] br[41] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_44 
+ bl[42] br[42] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_45 
+ bl[43] br[43] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_46 
+ bl[44] br[44] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_47 
+ bl[45] br[45] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_48 
+ bl[46] br[46] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_49 
+ bl[47] br[47] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_50 
+ bl[48] br[48] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_51 
+ bl[49] br[49] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_52 
+ bl[50] br[50] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_53 
+ bl[51] br[51] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_54 
+ bl[52] br[52] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_55 
+ bl[53] br[53] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_56 
+ bl[54] br[54] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_57 
+ bl[55] br[55] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_58 
+ bl[56] br[56] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_59 
+ bl[57] br[57] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_60 
+ bl[58] br[58] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_61 
+ bl[59] br[59] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_62 
+ bl[60] br[60] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_63 
+ bl[61] br[61] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_64 
+ bl[62] br[62] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_65 
+ bl[63] br[63] vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_66 
+ vdd vdd vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_19_67 
+ vdd vdd vdd vss wl[17] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_0 
+ vdd vdd vss vdd vpb vnb wl[18] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_20_1 
+ rbl rbr vss vdd vpb vnb wl[18] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_20_2 
+ bl[0] br[0] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_3 
+ bl[1] br[1] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_4 
+ bl[2] br[2] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_5 
+ bl[3] br[3] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_6 
+ bl[4] br[4] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_7 
+ bl[5] br[5] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_8 
+ bl[6] br[6] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_9 
+ bl[7] br[7] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_10 
+ bl[8] br[8] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_11 
+ bl[9] br[9] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_12 
+ bl[10] br[10] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_13 
+ bl[11] br[11] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_14 
+ bl[12] br[12] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_15 
+ bl[13] br[13] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_16 
+ bl[14] br[14] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_17 
+ bl[15] br[15] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_18 
+ bl[16] br[16] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_19 
+ bl[17] br[17] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_20 
+ bl[18] br[18] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_21 
+ bl[19] br[19] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_22 
+ bl[20] br[20] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_23 
+ bl[21] br[21] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_24 
+ bl[22] br[22] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_25 
+ bl[23] br[23] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_26 
+ bl[24] br[24] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_27 
+ bl[25] br[25] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_28 
+ bl[26] br[26] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_29 
+ bl[27] br[27] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_30 
+ bl[28] br[28] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_31 
+ bl[29] br[29] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_32 
+ bl[30] br[30] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_33 
+ bl[31] br[31] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_34 
+ bl[32] br[32] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_35 
+ bl[33] br[33] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_36 
+ bl[34] br[34] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_37 
+ bl[35] br[35] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_38 
+ bl[36] br[36] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_39 
+ bl[37] br[37] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_40 
+ bl[38] br[38] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_41 
+ bl[39] br[39] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_42 
+ bl[40] br[40] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_43 
+ bl[41] br[41] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_44 
+ bl[42] br[42] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_45 
+ bl[43] br[43] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_46 
+ bl[44] br[44] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_47 
+ bl[45] br[45] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_48 
+ bl[46] br[46] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_49 
+ bl[47] br[47] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_50 
+ bl[48] br[48] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_51 
+ bl[49] br[49] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_52 
+ bl[50] br[50] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_53 
+ bl[51] br[51] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_54 
+ bl[52] br[52] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_55 
+ bl[53] br[53] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_56 
+ bl[54] br[54] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_57 
+ bl[55] br[55] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_58 
+ bl[56] br[56] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_59 
+ bl[57] br[57] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_60 
+ bl[58] br[58] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_61 
+ bl[59] br[59] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_62 
+ bl[60] br[60] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_63 
+ bl[61] br[61] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_64 
+ bl[62] br[62] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_65 
+ bl[63] br[63] vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_66 
+ vdd vdd vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_20_67 
+ vdd vdd vdd vss wl[18] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_0 
+ vdd vdd vss vdd vpb vnb wl[19] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_21_1 
+ rbl rbr vss vdd vpb vnb wl[19] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_21_2 
+ bl[0] br[0] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_3 
+ bl[1] br[1] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_4 
+ bl[2] br[2] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_5 
+ bl[3] br[3] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_6 
+ bl[4] br[4] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_7 
+ bl[5] br[5] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_8 
+ bl[6] br[6] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_9 
+ bl[7] br[7] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_10 
+ bl[8] br[8] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_11 
+ bl[9] br[9] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_12 
+ bl[10] br[10] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_13 
+ bl[11] br[11] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_14 
+ bl[12] br[12] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_15 
+ bl[13] br[13] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_16 
+ bl[14] br[14] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_17 
+ bl[15] br[15] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_18 
+ bl[16] br[16] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_19 
+ bl[17] br[17] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_20 
+ bl[18] br[18] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_21 
+ bl[19] br[19] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_22 
+ bl[20] br[20] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_23 
+ bl[21] br[21] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_24 
+ bl[22] br[22] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_25 
+ bl[23] br[23] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_26 
+ bl[24] br[24] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_27 
+ bl[25] br[25] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_28 
+ bl[26] br[26] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_29 
+ bl[27] br[27] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_30 
+ bl[28] br[28] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_31 
+ bl[29] br[29] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_32 
+ bl[30] br[30] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_33 
+ bl[31] br[31] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_34 
+ bl[32] br[32] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_35 
+ bl[33] br[33] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_36 
+ bl[34] br[34] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_37 
+ bl[35] br[35] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_38 
+ bl[36] br[36] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_39 
+ bl[37] br[37] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_40 
+ bl[38] br[38] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_41 
+ bl[39] br[39] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_42 
+ bl[40] br[40] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_43 
+ bl[41] br[41] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_44 
+ bl[42] br[42] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_45 
+ bl[43] br[43] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_46 
+ bl[44] br[44] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_47 
+ bl[45] br[45] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_48 
+ bl[46] br[46] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_49 
+ bl[47] br[47] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_50 
+ bl[48] br[48] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_51 
+ bl[49] br[49] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_52 
+ bl[50] br[50] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_53 
+ bl[51] br[51] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_54 
+ bl[52] br[52] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_55 
+ bl[53] br[53] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_56 
+ bl[54] br[54] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_57 
+ bl[55] br[55] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_58 
+ bl[56] br[56] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_59 
+ bl[57] br[57] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_60 
+ bl[58] br[58] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_61 
+ bl[59] br[59] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_62 
+ bl[60] br[60] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_63 
+ bl[61] br[61] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_64 
+ bl[62] br[62] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_65 
+ bl[63] br[63] vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_66 
+ vdd vdd vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_21_67 
+ vdd vdd vdd vss wl[19] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_0 
+ vdd vdd vss vdd vpb vnb wl[20] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_22_1 
+ rbl rbr vss vdd vpb vnb wl[20] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_22_2 
+ bl[0] br[0] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_3 
+ bl[1] br[1] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_4 
+ bl[2] br[2] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_5 
+ bl[3] br[3] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_6 
+ bl[4] br[4] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_7 
+ bl[5] br[5] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_8 
+ bl[6] br[6] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_9 
+ bl[7] br[7] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_10 
+ bl[8] br[8] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_11 
+ bl[9] br[9] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_12 
+ bl[10] br[10] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_13 
+ bl[11] br[11] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_14 
+ bl[12] br[12] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_15 
+ bl[13] br[13] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_16 
+ bl[14] br[14] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_17 
+ bl[15] br[15] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_18 
+ bl[16] br[16] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_19 
+ bl[17] br[17] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_20 
+ bl[18] br[18] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_21 
+ bl[19] br[19] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_22 
+ bl[20] br[20] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_23 
+ bl[21] br[21] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_24 
+ bl[22] br[22] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_25 
+ bl[23] br[23] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_26 
+ bl[24] br[24] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_27 
+ bl[25] br[25] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_28 
+ bl[26] br[26] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_29 
+ bl[27] br[27] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_30 
+ bl[28] br[28] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_31 
+ bl[29] br[29] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_32 
+ bl[30] br[30] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_33 
+ bl[31] br[31] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_34 
+ bl[32] br[32] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_35 
+ bl[33] br[33] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_36 
+ bl[34] br[34] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_37 
+ bl[35] br[35] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_38 
+ bl[36] br[36] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_39 
+ bl[37] br[37] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_40 
+ bl[38] br[38] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_41 
+ bl[39] br[39] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_42 
+ bl[40] br[40] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_43 
+ bl[41] br[41] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_44 
+ bl[42] br[42] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_45 
+ bl[43] br[43] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_46 
+ bl[44] br[44] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_47 
+ bl[45] br[45] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_48 
+ bl[46] br[46] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_49 
+ bl[47] br[47] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_50 
+ bl[48] br[48] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_51 
+ bl[49] br[49] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_52 
+ bl[50] br[50] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_53 
+ bl[51] br[51] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_54 
+ bl[52] br[52] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_55 
+ bl[53] br[53] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_56 
+ bl[54] br[54] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_57 
+ bl[55] br[55] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_58 
+ bl[56] br[56] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_59 
+ bl[57] br[57] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_60 
+ bl[58] br[58] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_61 
+ bl[59] br[59] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_62 
+ bl[60] br[60] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_63 
+ bl[61] br[61] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_64 
+ bl[62] br[62] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_65 
+ bl[63] br[63] vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_66 
+ vdd vdd vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_22_67 
+ vdd vdd vdd vss wl[20] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_0 
+ vdd vdd vss vdd vpb vnb wl[21] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_23_1 
+ rbl rbr vss vdd vpb vnb wl[21] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_23_2 
+ bl[0] br[0] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_3 
+ bl[1] br[1] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_4 
+ bl[2] br[2] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_5 
+ bl[3] br[3] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_6 
+ bl[4] br[4] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_7 
+ bl[5] br[5] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_8 
+ bl[6] br[6] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_9 
+ bl[7] br[7] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_10 
+ bl[8] br[8] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_11 
+ bl[9] br[9] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_12 
+ bl[10] br[10] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_13 
+ bl[11] br[11] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_14 
+ bl[12] br[12] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_15 
+ bl[13] br[13] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_16 
+ bl[14] br[14] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_17 
+ bl[15] br[15] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_18 
+ bl[16] br[16] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_19 
+ bl[17] br[17] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_20 
+ bl[18] br[18] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_21 
+ bl[19] br[19] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_22 
+ bl[20] br[20] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_23 
+ bl[21] br[21] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_24 
+ bl[22] br[22] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_25 
+ bl[23] br[23] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_26 
+ bl[24] br[24] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_27 
+ bl[25] br[25] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_28 
+ bl[26] br[26] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_29 
+ bl[27] br[27] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_30 
+ bl[28] br[28] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_31 
+ bl[29] br[29] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_32 
+ bl[30] br[30] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_33 
+ bl[31] br[31] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_34 
+ bl[32] br[32] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_35 
+ bl[33] br[33] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_36 
+ bl[34] br[34] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_37 
+ bl[35] br[35] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_38 
+ bl[36] br[36] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_39 
+ bl[37] br[37] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_40 
+ bl[38] br[38] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_41 
+ bl[39] br[39] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_42 
+ bl[40] br[40] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_43 
+ bl[41] br[41] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_44 
+ bl[42] br[42] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_45 
+ bl[43] br[43] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_46 
+ bl[44] br[44] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_47 
+ bl[45] br[45] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_48 
+ bl[46] br[46] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_49 
+ bl[47] br[47] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_50 
+ bl[48] br[48] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_51 
+ bl[49] br[49] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_52 
+ bl[50] br[50] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_53 
+ bl[51] br[51] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_54 
+ bl[52] br[52] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_55 
+ bl[53] br[53] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_56 
+ bl[54] br[54] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_57 
+ bl[55] br[55] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_58 
+ bl[56] br[56] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_59 
+ bl[57] br[57] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_60 
+ bl[58] br[58] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_61 
+ bl[59] br[59] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_62 
+ bl[60] br[60] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_63 
+ bl[61] br[61] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_64 
+ bl[62] br[62] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_65 
+ bl[63] br[63] vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_66 
+ vdd vdd vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_23_67 
+ vdd vdd vdd vss wl[21] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_0 
+ vdd vdd vss vdd vpb vnb wl[22] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_24_1 
+ rbl rbr vss vdd vpb vnb wl[22] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_24_2 
+ bl[0] br[0] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_3 
+ bl[1] br[1] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_4 
+ bl[2] br[2] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_5 
+ bl[3] br[3] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_6 
+ bl[4] br[4] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_7 
+ bl[5] br[5] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_8 
+ bl[6] br[6] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_9 
+ bl[7] br[7] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_10 
+ bl[8] br[8] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_11 
+ bl[9] br[9] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_12 
+ bl[10] br[10] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_13 
+ bl[11] br[11] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_14 
+ bl[12] br[12] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_15 
+ bl[13] br[13] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_16 
+ bl[14] br[14] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_17 
+ bl[15] br[15] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_18 
+ bl[16] br[16] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_19 
+ bl[17] br[17] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_20 
+ bl[18] br[18] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_21 
+ bl[19] br[19] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_22 
+ bl[20] br[20] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_23 
+ bl[21] br[21] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_24 
+ bl[22] br[22] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_25 
+ bl[23] br[23] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_26 
+ bl[24] br[24] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_27 
+ bl[25] br[25] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_28 
+ bl[26] br[26] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_29 
+ bl[27] br[27] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_30 
+ bl[28] br[28] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_31 
+ bl[29] br[29] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_32 
+ bl[30] br[30] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_33 
+ bl[31] br[31] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_34 
+ bl[32] br[32] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_35 
+ bl[33] br[33] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_36 
+ bl[34] br[34] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_37 
+ bl[35] br[35] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_38 
+ bl[36] br[36] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_39 
+ bl[37] br[37] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_40 
+ bl[38] br[38] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_41 
+ bl[39] br[39] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_42 
+ bl[40] br[40] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_43 
+ bl[41] br[41] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_44 
+ bl[42] br[42] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_45 
+ bl[43] br[43] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_46 
+ bl[44] br[44] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_47 
+ bl[45] br[45] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_48 
+ bl[46] br[46] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_49 
+ bl[47] br[47] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_50 
+ bl[48] br[48] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_51 
+ bl[49] br[49] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_52 
+ bl[50] br[50] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_53 
+ bl[51] br[51] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_54 
+ bl[52] br[52] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_55 
+ bl[53] br[53] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_56 
+ bl[54] br[54] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_57 
+ bl[55] br[55] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_58 
+ bl[56] br[56] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_59 
+ bl[57] br[57] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_60 
+ bl[58] br[58] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_61 
+ bl[59] br[59] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_62 
+ bl[60] br[60] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_63 
+ bl[61] br[61] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_64 
+ bl[62] br[62] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_65 
+ bl[63] br[63] vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_66 
+ vdd vdd vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_24_67 
+ vdd vdd vdd vss wl[22] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_0 
+ vdd vdd vss vdd vpb vnb wl[23] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_25_1 
+ rbl rbr vss vdd vpb vnb wl[23] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_25_2 
+ bl[0] br[0] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_3 
+ bl[1] br[1] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_4 
+ bl[2] br[2] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_5 
+ bl[3] br[3] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_6 
+ bl[4] br[4] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_7 
+ bl[5] br[5] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_8 
+ bl[6] br[6] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_9 
+ bl[7] br[7] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_10 
+ bl[8] br[8] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_11 
+ bl[9] br[9] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_12 
+ bl[10] br[10] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_13 
+ bl[11] br[11] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_14 
+ bl[12] br[12] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_15 
+ bl[13] br[13] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_16 
+ bl[14] br[14] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_17 
+ bl[15] br[15] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_18 
+ bl[16] br[16] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_19 
+ bl[17] br[17] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_20 
+ bl[18] br[18] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_21 
+ bl[19] br[19] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_22 
+ bl[20] br[20] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_23 
+ bl[21] br[21] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_24 
+ bl[22] br[22] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_25 
+ bl[23] br[23] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_26 
+ bl[24] br[24] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_27 
+ bl[25] br[25] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_28 
+ bl[26] br[26] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_29 
+ bl[27] br[27] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_30 
+ bl[28] br[28] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_31 
+ bl[29] br[29] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_32 
+ bl[30] br[30] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_33 
+ bl[31] br[31] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_34 
+ bl[32] br[32] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_35 
+ bl[33] br[33] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_36 
+ bl[34] br[34] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_37 
+ bl[35] br[35] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_38 
+ bl[36] br[36] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_39 
+ bl[37] br[37] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_40 
+ bl[38] br[38] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_41 
+ bl[39] br[39] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_42 
+ bl[40] br[40] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_43 
+ bl[41] br[41] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_44 
+ bl[42] br[42] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_45 
+ bl[43] br[43] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_46 
+ bl[44] br[44] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_47 
+ bl[45] br[45] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_48 
+ bl[46] br[46] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_49 
+ bl[47] br[47] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_50 
+ bl[48] br[48] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_51 
+ bl[49] br[49] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_52 
+ bl[50] br[50] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_53 
+ bl[51] br[51] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_54 
+ bl[52] br[52] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_55 
+ bl[53] br[53] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_56 
+ bl[54] br[54] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_57 
+ bl[55] br[55] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_58 
+ bl[56] br[56] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_59 
+ bl[57] br[57] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_60 
+ bl[58] br[58] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_61 
+ bl[59] br[59] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_62 
+ bl[60] br[60] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_63 
+ bl[61] br[61] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_64 
+ bl[62] br[62] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_65 
+ bl[63] br[63] vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_66 
+ vdd vdd vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_25_67 
+ vdd vdd vdd vss wl[23] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_0 
+ vdd vdd vss vdd vpb vnb wl[24] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_26_1 
+ rbl rbr vss vdd vpb vnb wl[24] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_26_2 
+ bl[0] br[0] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_3 
+ bl[1] br[1] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_4 
+ bl[2] br[2] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_5 
+ bl[3] br[3] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_6 
+ bl[4] br[4] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_7 
+ bl[5] br[5] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_8 
+ bl[6] br[6] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_9 
+ bl[7] br[7] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_10 
+ bl[8] br[8] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_11 
+ bl[9] br[9] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_12 
+ bl[10] br[10] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_13 
+ bl[11] br[11] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_14 
+ bl[12] br[12] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_15 
+ bl[13] br[13] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_16 
+ bl[14] br[14] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_17 
+ bl[15] br[15] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_18 
+ bl[16] br[16] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_19 
+ bl[17] br[17] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_20 
+ bl[18] br[18] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_21 
+ bl[19] br[19] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_22 
+ bl[20] br[20] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_23 
+ bl[21] br[21] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_24 
+ bl[22] br[22] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_25 
+ bl[23] br[23] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_26 
+ bl[24] br[24] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_27 
+ bl[25] br[25] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_28 
+ bl[26] br[26] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_29 
+ bl[27] br[27] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_30 
+ bl[28] br[28] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_31 
+ bl[29] br[29] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_32 
+ bl[30] br[30] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_33 
+ bl[31] br[31] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_34 
+ bl[32] br[32] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_35 
+ bl[33] br[33] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_36 
+ bl[34] br[34] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_37 
+ bl[35] br[35] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_38 
+ bl[36] br[36] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_39 
+ bl[37] br[37] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_40 
+ bl[38] br[38] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_41 
+ bl[39] br[39] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_42 
+ bl[40] br[40] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_43 
+ bl[41] br[41] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_44 
+ bl[42] br[42] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_45 
+ bl[43] br[43] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_46 
+ bl[44] br[44] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_47 
+ bl[45] br[45] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_48 
+ bl[46] br[46] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_49 
+ bl[47] br[47] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_50 
+ bl[48] br[48] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_51 
+ bl[49] br[49] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_52 
+ bl[50] br[50] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_53 
+ bl[51] br[51] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_54 
+ bl[52] br[52] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_55 
+ bl[53] br[53] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_56 
+ bl[54] br[54] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_57 
+ bl[55] br[55] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_58 
+ bl[56] br[56] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_59 
+ bl[57] br[57] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_60 
+ bl[58] br[58] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_61 
+ bl[59] br[59] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_62 
+ bl[60] br[60] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_63 
+ bl[61] br[61] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_64 
+ bl[62] br[62] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_65 
+ bl[63] br[63] vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_66 
+ vdd vdd vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_26_67 
+ vdd vdd vdd vss wl[24] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_0 
+ vdd vdd vss vdd vpb vnb wl[25] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_27_1 
+ rbl rbr vss vdd vpb vnb wl[25] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_27_2 
+ bl[0] br[0] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_3 
+ bl[1] br[1] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_4 
+ bl[2] br[2] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_5 
+ bl[3] br[3] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_6 
+ bl[4] br[4] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_7 
+ bl[5] br[5] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_8 
+ bl[6] br[6] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_9 
+ bl[7] br[7] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_10 
+ bl[8] br[8] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_11 
+ bl[9] br[9] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_12 
+ bl[10] br[10] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_13 
+ bl[11] br[11] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_14 
+ bl[12] br[12] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_15 
+ bl[13] br[13] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_16 
+ bl[14] br[14] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_17 
+ bl[15] br[15] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_18 
+ bl[16] br[16] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_19 
+ bl[17] br[17] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_20 
+ bl[18] br[18] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_21 
+ bl[19] br[19] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_22 
+ bl[20] br[20] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_23 
+ bl[21] br[21] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_24 
+ bl[22] br[22] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_25 
+ bl[23] br[23] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_26 
+ bl[24] br[24] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_27 
+ bl[25] br[25] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_28 
+ bl[26] br[26] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_29 
+ bl[27] br[27] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_30 
+ bl[28] br[28] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_31 
+ bl[29] br[29] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_32 
+ bl[30] br[30] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_33 
+ bl[31] br[31] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_34 
+ bl[32] br[32] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_35 
+ bl[33] br[33] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_36 
+ bl[34] br[34] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_37 
+ bl[35] br[35] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_38 
+ bl[36] br[36] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_39 
+ bl[37] br[37] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_40 
+ bl[38] br[38] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_41 
+ bl[39] br[39] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_42 
+ bl[40] br[40] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_43 
+ bl[41] br[41] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_44 
+ bl[42] br[42] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_45 
+ bl[43] br[43] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_46 
+ bl[44] br[44] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_47 
+ bl[45] br[45] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_48 
+ bl[46] br[46] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_49 
+ bl[47] br[47] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_50 
+ bl[48] br[48] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_51 
+ bl[49] br[49] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_52 
+ bl[50] br[50] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_53 
+ bl[51] br[51] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_54 
+ bl[52] br[52] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_55 
+ bl[53] br[53] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_56 
+ bl[54] br[54] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_57 
+ bl[55] br[55] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_58 
+ bl[56] br[56] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_59 
+ bl[57] br[57] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_60 
+ bl[58] br[58] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_61 
+ bl[59] br[59] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_62 
+ bl[60] br[60] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_63 
+ bl[61] br[61] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_64 
+ bl[62] br[62] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_65 
+ bl[63] br[63] vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_66 
+ vdd vdd vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_27_67 
+ vdd vdd vdd vss wl[25] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_0 
+ vdd vdd vss vdd vpb vnb wl[26] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_28_1 
+ rbl rbr vss vdd vpb vnb wl[26] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_28_2 
+ bl[0] br[0] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_3 
+ bl[1] br[1] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_4 
+ bl[2] br[2] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_5 
+ bl[3] br[3] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_6 
+ bl[4] br[4] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_7 
+ bl[5] br[5] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_8 
+ bl[6] br[6] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_9 
+ bl[7] br[7] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_10 
+ bl[8] br[8] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_11 
+ bl[9] br[9] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_12 
+ bl[10] br[10] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_13 
+ bl[11] br[11] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_14 
+ bl[12] br[12] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_15 
+ bl[13] br[13] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_16 
+ bl[14] br[14] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_17 
+ bl[15] br[15] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_18 
+ bl[16] br[16] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_19 
+ bl[17] br[17] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_20 
+ bl[18] br[18] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_21 
+ bl[19] br[19] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_22 
+ bl[20] br[20] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_23 
+ bl[21] br[21] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_24 
+ bl[22] br[22] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_25 
+ bl[23] br[23] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_26 
+ bl[24] br[24] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_27 
+ bl[25] br[25] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_28 
+ bl[26] br[26] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_29 
+ bl[27] br[27] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_30 
+ bl[28] br[28] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_31 
+ bl[29] br[29] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_32 
+ bl[30] br[30] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_33 
+ bl[31] br[31] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_34 
+ bl[32] br[32] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_35 
+ bl[33] br[33] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_36 
+ bl[34] br[34] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_37 
+ bl[35] br[35] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_38 
+ bl[36] br[36] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_39 
+ bl[37] br[37] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_40 
+ bl[38] br[38] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_41 
+ bl[39] br[39] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_42 
+ bl[40] br[40] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_43 
+ bl[41] br[41] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_44 
+ bl[42] br[42] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_45 
+ bl[43] br[43] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_46 
+ bl[44] br[44] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_47 
+ bl[45] br[45] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_48 
+ bl[46] br[46] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_49 
+ bl[47] br[47] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_50 
+ bl[48] br[48] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_51 
+ bl[49] br[49] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_52 
+ bl[50] br[50] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_53 
+ bl[51] br[51] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_54 
+ bl[52] br[52] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_55 
+ bl[53] br[53] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_56 
+ bl[54] br[54] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_57 
+ bl[55] br[55] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_58 
+ bl[56] br[56] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_59 
+ bl[57] br[57] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_60 
+ bl[58] br[58] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_61 
+ bl[59] br[59] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_62 
+ bl[60] br[60] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_63 
+ bl[61] br[61] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_64 
+ bl[62] br[62] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_65 
+ bl[63] br[63] vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_66 
+ vdd vdd vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_28_67 
+ vdd vdd vdd vss wl[26] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_0 
+ vdd vdd vss vdd vpb vnb wl[27] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_29_1 
+ rbl rbr vss vdd vpb vnb wl[27] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_29_2 
+ bl[0] br[0] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_3 
+ bl[1] br[1] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_4 
+ bl[2] br[2] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_5 
+ bl[3] br[3] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_6 
+ bl[4] br[4] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_7 
+ bl[5] br[5] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_8 
+ bl[6] br[6] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_9 
+ bl[7] br[7] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_10 
+ bl[8] br[8] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_11 
+ bl[9] br[9] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_12 
+ bl[10] br[10] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_13 
+ bl[11] br[11] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_14 
+ bl[12] br[12] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_15 
+ bl[13] br[13] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_16 
+ bl[14] br[14] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_17 
+ bl[15] br[15] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_18 
+ bl[16] br[16] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_19 
+ bl[17] br[17] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_20 
+ bl[18] br[18] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_21 
+ bl[19] br[19] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_22 
+ bl[20] br[20] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_23 
+ bl[21] br[21] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_24 
+ bl[22] br[22] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_25 
+ bl[23] br[23] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_26 
+ bl[24] br[24] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_27 
+ bl[25] br[25] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_28 
+ bl[26] br[26] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_29 
+ bl[27] br[27] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_30 
+ bl[28] br[28] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_31 
+ bl[29] br[29] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_32 
+ bl[30] br[30] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_33 
+ bl[31] br[31] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_34 
+ bl[32] br[32] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_35 
+ bl[33] br[33] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_36 
+ bl[34] br[34] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_37 
+ bl[35] br[35] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_38 
+ bl[36] br[36] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_39 
+ bl[37] br[37] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_40 
+ bl[38] br[38] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_41 
+ bl[39] br[39] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_42 
+ bl[40] br[40] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_43 
+ bl[41] br[41] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_44 
+ bl[42] br[42] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_45 
+ bl[43] br[43] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_46 
+ bl[44] br[44] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_47 
+ bl[45] br[45] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_48 
+ bl[46] br[46] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_49 
+ bl[47] br[47] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_50 
+ bl[48] br[48] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_51 
+ bl[49] br[49] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_52 
+ bl[50] br[50] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_53 
+ bl[51] br[51] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_54 
+ bl[52] br[52] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_55 
+ bl[53] br[53] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_56 
+ bl[54] br[54] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_57 
+ bl[55] br[55] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_58 
+ bl[56] br[56] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_59 
+ bl[57] br[57] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_60 
+ bl[58] br[58] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_61 
+ bl[59] br[59] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_62 
+ bl[60] br[60] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_63 
+ bl[61] br[61] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_64 
+ bl[62] br[62] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_65 
+ bl[63] br[63] vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_66 
+ vdd vdd vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_29_67 
+ vdd vdd vdd vss wl[27] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_0 
+ vdd vdd vss vdd vpb vnb wl[28] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_30_1 
+ rbl rbr vss vdd vpb vnb wl[28] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_30_2 
+ bl[0] br[0] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_3 
+ bl[1] br[1] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_4 
+ bl[2] br[2] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_5 
+ bl[3] br[3] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_6 
+ bl[4] br[4] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_7 
+ bl[5] br[5] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_8 
+ bl[6] br[6] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_9 
+ bl[7] br[7] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_10 
+ bl[8] br[8] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_11 
+ bl[9] br[9] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_12 
+ bl[10] br[10] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_13 
+ bl[11] br[11] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_14 
+ bl[12] br[12] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_15 
+ bl[13] br[13] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_16 
+ bl[14] br[14] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_17 
+ bl[15] br[15] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_18 
+ bl[16] br[16] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_19 
+ bl[17] br[17] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_20 
+ bl[18] br[18] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_21 
+ bl[19] br[19] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_22 
+ bl[20] br[20] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_23 
+ bl[21] br[21] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_24 
+ bl[22] br[22] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_25 
+ bl[23] br[23] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_26 
+ bl[24] br[24] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_27 
+ bl[25] br[25] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_28 
+ bl[26] br[26] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_29 
+ bl[27] br[27] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_30 
+ bl[28] br[28] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_31 
+ bl[29] br[29] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_32 
+ bl[30] br[30] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_33 
+ bl[31] br[31] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_34 
+ bl[32] br[32] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_35 
+ bl[33] br[33] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_36 
+ bl[34] br[34] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_37 
+ bl[35] br[35] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_38 
+ bl[36] br[36] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_39 
+ bl[37] br[37] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_40 
+ bl[38] br[38] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_41 
+ bl[39] br[39] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_42 
+ bl[40] br[40] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_43 
+ bl[41] br[41] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_44 
+ bl[42] br[42] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_45 
+ bl[43] br[43] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_46 
+ bl[44] br[44] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_47 
+ bl[45] br[45] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_48 
+ bl[46] br[46] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_49 
+ bl[47] br[47] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_50 
+ bl[48] br[48] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_51 
+ bl[49] br[49] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_52 
+ bl[50] br[50] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_53 
+ bl[51] br[51] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_54 
+ bl[52] br[52] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_55 
+ bl[53] br[53] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_56 
+ bl[54] br[54] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_57 
+ bl[55] br[55] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_58 
+ bl[56] br[56] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_59 
+ bl[57] br[57] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_60 
+ bl[58] br[58] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_61 
+ bl[59] br[59] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_62 
+ bl[60] br[60] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_63 
+ bl[61] br[61] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_64 
+ bl[62] br[62] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_65 
+ bl[63] br[63] vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_66 
+ vdd vdd vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_30_67 
+ vdd vdd vdd vss wl[28] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_0 
+ vdd vdd vss vdd vpb vnb wl[29] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_31_1 
+ rbl rbr vss vdd vpb vnb wl[29] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_31_2 
+ bl[0] br[0] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_3 
+ bl[1] br[1] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_4 
+ bl[2] br[2] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_5 
+ bl[3] br[3] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_6 
+ bl[4] br[4] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_7 
+ bl[5] br[5] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_8 
+ bl[6] br[6] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_9 
+ bl[7] br[7] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_10 
+ bl[8] br[8] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_11 
+ bl[9] br[9] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_12 
+ bl[10] br[10] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_13 
+ bl[11] br[11] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_14 
+ bl[12] br[12] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_15 
+ bl[13] br[13] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_16 
+ bl[14] br[14] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_17 
+ bl[15] br[15] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_18 
+ bl[16] br[16] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_19 
+ bl[17] br[17] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_20 
+ bl[18] br[18] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_21 
+ bl[19] br[19] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_22 
+ bl[20] br[20] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_23 
+ bl[21] br[21] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_24 
+ bl[22] br[22] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_25 
+ bl[23] br[23] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_26 
+ bl[24] br[24] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_27 
+ bl[25] br[25] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_28 
+ bl[26] br[26] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_29 
+ bl[27] br[27] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_30 
+ bl[28] br[28] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_31 
+ bl[29] br[29] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_32 
+ bl[30] br[30] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_33 
+ bl[31] br[31] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_34 
+ bl[32] br[32] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_35 
+ bl[33] br[33] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_36 
+ bl[34] br[34] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_37 
+ bl[35] br[35] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_38 
+ bl[36] br[36] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_39 
+ bl[37] br[37] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_40 
+ bl[38] br[38] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_41 
+ bl[39] br[39] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_42 
+ bl[40] br[40] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_43 
+ bl[41] br[41] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_44 
+ bl[42] br[42] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_45 
+ bl[43] br[43] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_46 
+ bl[44] br[44] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_47 
+ bl[45] br[45] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_48 
+ bl[46] br[46] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_49 
+ bl[47] br[47] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_50 
+ bl[48] br[48] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_51 
+ bl[49] br[49] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_52 
+ bl[50] br[50] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_53 
+ bl[51] br[51] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_54 
+ bl[52] br[52] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_55 
+ bl[53] br[53] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_56 
+ bl[54] br[54] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_57 
+ bl[55] br[55] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_58 
+ bl[56] br[56] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_59 
+ bl[57] br[57] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_60 
+ bl[58] br[58] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_61 
+ bl[59] br[59] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_62 
+ bl[60] br[60] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_63 
+ bl[61] br[61] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_64 
+ bl[62] br[62] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_65 
+ bl[63] br[63] vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_66 
+ vdd vdd vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_31_67 
+ vdd vdd vdd vss wl[29] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_0 
+ vdd vdd vss vdd vpb vnb wl[30] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_32_1 
+ rbl rbr vss vdd vpb vnb wl[30] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_32_2 
+ bl[0] br[0] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_3 
+ bl[1] br[1] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_4 
+ bl[2] br[2] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_5 
+ bl[3] br[3] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_6 
+ bl[4] br[4] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_7 
+ bl[5] br[5] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_8 
+ bl[6] br[6] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_9 
+ bl[7] br[7] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_10 
+ bl[8] br[8] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_11 
+ bl[9] br[9] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_12 
+ bl[10] br[10] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_13 
+ bl[11] br[11] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_14 
+ bl[12] br[12] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_15 
+ bl[13] br[13] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_16 
+ bl[14] br[14] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_17 
+ bl[15] br[15] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_18 
+ bl[16] br[16] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_19 
+ bl[17] br[17] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_20 
+ bl[18] br[18] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_21 
+ bl[19] br[19] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_22 
+ bl[20] br[20] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_23 
+ bl[21] br[21] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_24 
+ bl[22] br[22] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_25 
+ bl[23] br[23] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_26 
+ bl[24] br[24] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_27 
+ bl[25] br[25] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_28 
+ bl[26] br[26] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_29 
+ bl[27] br[27] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_30 
+ bl[28] br[28] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_31 
+ bl[29] br[29] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_32 
+ bl[30] br[30] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_33 
+ bl[31] br[31] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_34 
+ bl[32] br[32] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_35 
+ bl[33] br[33] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_36 
+ bl[34] br[34] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_37 
+ bl[35] br[35] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_38 
+ bl[36] br[36] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_39 
+ bl[37] br[37] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_40 
+ bl[38] br[38] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_41 
+ bl[39] br[39] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_42 
+ bl[40] br[40] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_43 
+ bl[41] br[41] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_44 
+ bl[42] br[42] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_45 
+ bl[43] br[43] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_46 
+ bl[44] br[44] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_47 
+ bl[45] br[45] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_48 
+ bl[46] br[46] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_49 
+ bl[47] br[47] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_50 
+ bl[48] br[48] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_51 
+ bl[49] br[49] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_52 
+ bl[50] br[50] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_53 
+ bl[51] br[51] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_54 
+ bl[52] br[52] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_55 
+ bl[53] br[53] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_56 
+ bl[54] br[54] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_57 
+ bl[55] br[55] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_58 
+ bl[56] br[56] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_59 
+ bl[57] br[57] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_60 
+ bl[58] br[58] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_61 
+ bl[59] br[59] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_62 
+ bl[60] br[60] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_63 
+ bl[61] br[61] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_64 
+ bl[62] br[62] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_65 
+ bl[63] br[63] vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_66 
+ vdd vdd vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_32_67 
+ vdd vdd vdd vss wl[30] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_0 
+ vdd vdd vss vdd vpb vnb wl[31] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_33_1 
+ rbl rbr vss vdd vpb vnb wl[31] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_33_2 
+ bl[0] br[0] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_3 
+ bl[1] br[1] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_4 
+ bl[2] br[2] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_5 
+ bl[3] br[3] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_6 
+ bl[4] br[4] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_7 
+ bl[5] br[5] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_8 
+ bl[6] br[6] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_9 
+ bl[7] br[7] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_10 
+ bl[8] br[8] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_11 
+ bl[9] br[9] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_12 
+ bl[10] br[10] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_13 
+ bl[11] br[11] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_14 
+ bl[12] br[12] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_15 
+ bl[13] br[13] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_16 
+ bl[14] br[14] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_17 
+ bl[15] br[15] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_18 
+ bl[16] br[16] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_19 
+ bl[17] br[17] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_20 
+ bl[18] br[18] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_21 
+ bl[19] br[19] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_22 
+ bl[20] br[20] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_23 
+ bl[21] br[21] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_24 
+ bl[22] br[22] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_25 
+ bl[23] br[23] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_26 
+ bl[24] br[24] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_27 
+ bl[25] br[25] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_28 
+ bl[26] br[26] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_29 
+ bl[27] br[27] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_30 
+ bl[28] br[28] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_31 
+ bl[29] br[29] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_32 
+ bl[30] br[30] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_33 
+ bl[31] br[31] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_34 
+ bl[32] br[32] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_35 
+ bl[33] br[33] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_36 
+ bl[34] br[34] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_37 
+ bl[35] br[35] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_38 
+ bl[36] br[36] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_39 
+ bl[37] br[37] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_40 
+ bl[38] br[38] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_41 
+ bl[39] br[39] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_42 
+ bl[40] br[40] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_43 
+ bl[41] br[41] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_44 
+ bl[42] br[42] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_45 
+ bl[43] br[43] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_46 
+ bl[44] br[44] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_47 
+ bl[45] br[45] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_48 
+ bl[46] br[46] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_49 
+ bl[47] br[47] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_50 
+ bl[48] br[48] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_51 
+ bl[49] br[49] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_52 
+ bl[50] br[50] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_53 
+ bl[51] br[51] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_54 
+ bl[52] br[52] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_55 
+ bl[53] br[53] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_56 
+ bl[54] br[54] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_57 
+ bl[55] br[55] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_58 
+ bl[56] br[56] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_59 
+ bl[57] br[57] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_60 
+ bl[58] br[58] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_61 
+ bl[59] br[59] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_62 
+ bl[60] br[60] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_63 
+ bl[61] br[61] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_64 
+ bl[62] br[62] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_65 
+ bl[63] br[63] vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_66 
+ vdd vdd vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_33_67 
+ vdd vdd vdd vss wl[31] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_0 
+ vdd vdd vss vdd vpb vnb wl[32] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_34_1 
+ rbl rbr vss vdd vpb vnb wl[32] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_34_2 
+ bl[0] br[0] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_3 
+ bl[1] br[1] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_4 
+ bl[2] br[2] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_5 
+ bl[3] br[3] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_6 
+ bl[4] br[4] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_7 
+ bl[5] br[5] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_8 
+ bl[6] br[6] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_9 
+ bl[7] br[7] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_10 
+ bl[8] br[8] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_11 
+ bl[9] br[9] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_12 
+ bl[10] br[10] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_13 
+ bl[11] br[11] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_14 
+ bl[12] br[12] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_15 
+ bl[13] br[13] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_16 
+ bl[14] br[14] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_17 
+ bl[15] br[15] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_18 
+ bl[16] br[16] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_19 
+ bl[17] br[17] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_20 
+ bl[18] br[18] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_21 
+ bl[19] br[19] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_22 
+ bl[20] br[20] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_23 
+ bl[21] br[21] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_24 
+ bl[22] br[22] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_25 
+ bl[23] br[23] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_26 
+ bl[24] br[24] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_27 
+ bl[25] br[25] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_28 
+ bl[26] br[26] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_29 
+ bl[27] br[27] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_30 
+ bl[28] br[28] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_31 
+ bl[29] br[29] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_32 
+ bl[30] br[30] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_33 
+ bl[31] br[31] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_34 
+ bl[32] br[32] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_35 
+ bl[33] br[33] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_36 
+ bl[34] br[34] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_37 
+ bl[35] br[35] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_38 
+ bl[36] br[36] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_39 
+ bl[37] br[37] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_40 
+ bl[38] br[38] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_41 
+ bl[39] br[39] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_42 
+ bl[40] br[40] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_43 
+ bl[41] br[41] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_44 
+ bl[42] br[42] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_45 
+ bl[43] br[43] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_46 
+ bl[44] br[44] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_47 
+ bl[45] br[45] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_48 
+ bl[46] br[46] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_49 
+ bl[47] br[47] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_50 
+ bl[48] br[48] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_51 
+ bl[49] br[49] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_52 
+ bl[50] br[50] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_53 
+ bl[51] br[51] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_54 
+ bl[52] br[52] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_55 
+ bl[53] br[53] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_56 
+ bl[54] br[54] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_57 
+ bl[55] br[55] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_58 
+ bl[56] br[56] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_59 
+ bl[57] br[57] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_60 
+ bl[58] br[58] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_61 
+ bl[59] br[59] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_62 
+ bl[60] br[60] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_63 
+ bl[61] br[61] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_64 
+ bl[62] br[62] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_65 
+ bl[63] br[63] vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_66 
+ vdd vdd vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_34_67 
+ vdd vdd vdd vss wl[32] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_0 
+ vdd vdd vss vdd vpb vnb wl[33] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_35_1 
+ rbl rbr vss vdd vpb vnb wl[33] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_35_2 
+ bl[0] br[0] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_3 
+ bl[1] br[1] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_4 
+ bl[2] br[2] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_5 
+ bl[3] br[3] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_6 
+ bl[4] br[4] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_7 
+ bl[5] br[5] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_8 
+ bl[6] br[6] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_9 
+ bl[7] br[7] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_10 
+ bl[8] br[8] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_11 
+ bl[9] br[9] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_12 
+ bl[10] br[10] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_13 
+ bl[11] br[11] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_14 
+ bl[12] br[12] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_15 
+ bl[13] br[13] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_16 
+ bl[14] br[14] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_17 
+ bl[15] br[15] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_18 
+ bl[16] br[16] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_19 
+ bl[17] br[17] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_20 
+ bl[18] br[18] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_21 
+ bl[19] br[19] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_22 
+ bl[20] br[20] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_23 
+ bl[21] br[21] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_24 
+ bl[22] br[22] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_25 
+ bl[23] br[23] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_26 
+ bl[24] br[24] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_27 
+ bl[25] br[25] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_28 
+ bl[26] br[26] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_29 
+ bl[27] br[27] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_30 
+ bl[28] br[28] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_31 
+ bl[29] br[29] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_32 
+ bl[30] br[30] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_33 
+ bl[31] br[31] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_34 
+ bl[32] br[32] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_35 
+ bl[33] br[33] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_36 
+ bl[34] br[34] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_37 
+ bl[35] br[35] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_38 
+ bl[36] br[36] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_39 
+ bl[37] br[37] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_40 
+ bl[38] br[38] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_41 
+ bl[39] br[39] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_42 
+ bl[40] br[40] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_43 
+ bl[41] br[41] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_44 
+ bl[42] br[42] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_45 
+ bl[43] br[43] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_46 
+ bl[44] br[44] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_47 
+ bl[45] br[45] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_48 
+ bl[46] br[46] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_49 
+ bl[47] br[47] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_50 
+ bl[48] br[48] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_51 
+ bl[49] br[49] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_52 
+ bl[50] br[50] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_53 
+ bl[51] br[51] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_54 
+ bl[52] br[52] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_55 
+ bl[53] br[53] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_56 
+ bl[54] br[54] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_57 
+ bl[55] br[55] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_58 
+ bl[56] br[56] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_59 
+ bl[57] br[57] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_60 
+ bl[58] br[58] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_61 
+ bl[59] br[59] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_62 
+ bl[60] br[60] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_63 
+ bl[61] br[61] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_64 
+ bl[62] br[62] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_65 
+ bl[63] br[63] vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_66 
+ vdd vdd vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_35_67 
+ vdd vdd vdd vss wl[33] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_0 
+ vdd vdd vss vdd vpb vnb wl[34] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_36_1 
+ rbl rbr vss vdd vpb vnb wl[34] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_36_2 
+ bl[0] br[0] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_3 
+ bl[1] br[1] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_4 
+ bl[2] br[2] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_5 
+ bl[3] br[3] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_6 
+ bl[4] br[4] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_7 
+ bl[5] br[5] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_8 
+ bl[6] br[6] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_9 
+ bl[7] br[7] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_10 
+ bl[8] br[8] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_11 
+ bl[9] br[9] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_12 
+ bl[10] br[10] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_13 
+ bl[11] br[11] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_14 
+ bl[12] br[12] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_15 
+ bl[13] br[13] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_16 
+ bl[14] br[14] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_17 
+ bl[15] br[15] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_18 
+ bl[16] br[16] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_19 
+ bl[17] br[17] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_20 
+ bl[18] br[18] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_21 
+ bl[19] br[19] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_22 
+ bl[20] br[20] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_23 
+ bl[21] br[21] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_24 
+ bl[22] br[22] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_25 
+ bl[23] br[23] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_26 
+ bl[24] br[24] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_27 
+ bl[25] br[25] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_28 
+ bl[26] br[26] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_29 
+ bl[27] br[27] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_30 
+ bl[28] br[28] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_31 
+ bl[29] br[29] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_32 
+ bl[30] br[30] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_33 
+ bl[31] br[31] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_34 
+ bl[32] br[32] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_35 
+ bl[33] br[33] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_36 
+ bl[34] br[34] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_37 
+ bl[35] br[35] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_38 
+ bl[36] br[36] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_39 
+ bl[37] br[37] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_40 
+ bl[38] br[38] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_41 
+ bl[39] br[39] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_42 
+ bl[40] br[40] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_43 
+ bl[41] br[41] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_44 
+ bl[42] br[42] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_45 
+ bl[43] br[43] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_46 
+ bl[44] br[44] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_47 
+ bl[45] br[45] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_48 
+ bl[46] br[46] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_49 
+ bl[47] br[47] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_50 
+ bl[48] br[48] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_51 
+ bl[49] br[49] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_52 
+ bl[50] br[50] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_53 
+ bl[51] br[51] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_54 
+ bl[52] br[52] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_55 
+ bl[53] br[53] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_56 
+ bl[54] br[54] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_57 
+ bl[55] br[55] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_58 
+ bl[56] br[56] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_59 
+ bl[57] br[57] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_60 
+ bl[58] br[58] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_61 
+ bl[59] br[59] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_62 
+ bl[60] br[60] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_63 
+ bl[61] br[61] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_64 
+ bl[62] br[62] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_65 
+ bl[63] br[63] vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_66 
+ vdd vdd vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_36_67 
+ vdd vdd vdd vss wl[34] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_0 
+ vdd vdd vss vdd vpb vnb wl[35] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_37_1 
+ rbl rbr vss vdd vpb vnb wl[35] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_37_2 
+ bl[0] br[0] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_3 
+ bl[1] br[1] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_4 
+ bl[2] br[2] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_5 
+ bl[3] br[3] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_6 
+ bl[4] br[4] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_7 
+ bl[5] br[5] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_8 
+ bl[6] br[6] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_9 
+ bl[7] br[7] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_10 
+ bl[8] br[8] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_11 
+ bl[9] br[9] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_12 
+ bl[10] br[10] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_13 
+ bl[11] br[11] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_14 
+ bl[12] br[12] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_15 
+ bl[13] br[13] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_16 
+ bl[14] br[14] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_17 
+ bl[15] br[15] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_18 
+ bl[16] br[16] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_19 
+ bl[17] br[17] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_20 
+ bl[18] br[18] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_21 
+ bl[19] br[19] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_22 
+ bl[20] br[20] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_23 
+ bl[21] br[21] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_24 
+ bl[22] br[22] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_25 
+ bl[23] br[23] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_26 
+ bl[24] br[24] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_27 
+ bl[25] br[25] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_28 
+ bl[26] br[26] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_29 
+ bl[27] br[27] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_30 
+ bl[28] br[28] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_31 
+ bl[29] br[29] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_32 
+ bl[30] br[30] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_33 
+ bl[31] br[31] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_34 
+ bl[32] br[32] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_35 
+ bl[33] br[33] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_36 
+ bl[34] br[34] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_37 
+ bl[35] br[35] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_38 
+ bl[36] br[36] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_39 
+ bl[37] br[37] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_40 
+ bl[38] br[38] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_41 
+ bl[39] br[39] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_42 
+ bl[40] br[40] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_43 
+ bl[41] br[41] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_44 
+ bl[42] br[42] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_45 
+ bl[43] br[43] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_46 
+ bl[44] br[44] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_47 
+ bl[45] br[45] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_48 
+ bl[46] br[46] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_49 
+ bl[47] br[47] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_50 
+ bl[48] br[48] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_51 
+ bl[49] br[49] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_52 
+ bl[50] br[50] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_53 
+ bl[51] br[51] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_54 
+ bl[52] br[52] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_55 
+ bl[53] br[53] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_56 
+ bl[54] br[54] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_57 
+ bl[55] br[55] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_58 
+ bl[56] br[56] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_59 
+ bl[57] br[57] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_60 
+ bl[58] br[58] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_61 
+ bl[59] br[59] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_62 
+ bl[60] br[60] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_63 
+ bl[61] br[61] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_64 
+ bl[62] br[62] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_65 
+ bl[63] br[63] vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_66 
+ vdd vdd vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_37_67 
+ vdd vdd vdd vss wl[35] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_0 
+ vdd vdd vss vdd vpb vnb wl[36] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_38_1 
+ rbl rbr vss vdd vpb vnb wl[36] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_38_2 
+ bl[0] br[0] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_3 
+ bl[1] br[1] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_4 
+ bl[2] br[2] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_5 
+ bl[3] br[3] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_6 
+ bl[4] br[4] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_7 
+ bl[5] br[5] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_8 
+ bl[6] br[6] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_9 
+ bl[7] br[7] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_10 
+ bl[8] br[8] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_11 
+ bl[9] br[9] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_12 
+ bl[10] br[10] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_13 
+ bl[11] br[11] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_14 
+ bl[12] br[12] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_15 
+ bl[13] br[13] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_16 
+ bl[14] br[14] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_17 
+ bl[15] br[15] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_18 
+ bl[16] br[16] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_19 
+ bl[17] br[17] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_20 
+ bl[18] br[18] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_21 
+ bl[19] br[19] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_22 
+ bl[20] br[20] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_23 
+ bl[21] br[21] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_24 
+ bl[22] br[22] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_25 
+ bl[23] br[23] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_26 
+ bl[24] br[24] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_27 
+ bl[25] br[25] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_28 
+ bl[26] br[26] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_29 
+ bl[27] br[27] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_30 
+ bl[28] br[28] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_31 
+ bl[29] br[29] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_32 
+ bl[30] br[30] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_33 
+ bl[31] br[31] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_34 
+ bl[32] br[32] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_35 
+ bl[33] br[33] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_36 
+ bl[34] br[34] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_37 
+ bl[35] br[35] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_38 
+ bl[36] br[36] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_39 
+ bl[37] br[37] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_40 
+ bl[38] br[38] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_41 
+ bl[39] br[39] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_42 
+ bl[40] br[40] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_43 
+ bl[41] br[41] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_44 
+ bl[42] br[42] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_45 
+ bl[43] br[43] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_46 
+ bl[44] br[44] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_47 
+ bl[45] br[45] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_48 
+ bl[46] br[46] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_49 
+ bl[47] br[47] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_50 
+ bl[48] br[48] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_51 
+ bl[49] br[49] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_52 
+ bl[50] br[50] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_53 
+ bl[51] br[51] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_54 
+ bl[52] br[52] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_55 
+ bl[53] br[53] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_56 
+ bl[54] br[54] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_57 
+ bl[55] br[55] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_58 
+ bl[56] br[56] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_59 
+ bl[57] br[57] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_60 
+ bl[58] br[58] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_61 
+ bl[59] br[59] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_62 
+ bl[60] br[60] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_63 
+ bl[61] br[61] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_64 
+ bl[62] br[62] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_65 
+ bl[63] br[63] vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_66 
+ vdd vdd vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_38_67 
+ vdd vdd vdd vss wl[36] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_0 
+ vdd vdd vss vdd vpb vnb wl[37] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_39_1 
+ rbl rbr vss vdd vpb vnb wl[37] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_39_2 
+ bl[0] br[0] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_3 
+ bl[1] br[1] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_4 
+ bl[2] br[2] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_5 
+ bl[3] br[3] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_6 
+ bl[4] br[4] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_7 
+ bl[5] br[5] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_8 
+ bl[6] br[6] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_9 
+ bl[7] br[7] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_10 
+ bl[8] br[8] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_11 
+ bl[9] br[9] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_12 
+ bl[10] br[10] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_13 
+ bl[11] br[11] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_14 
+ bl[12] br[12] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_15 
+ bl[13] br[13] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_16 
+ bl[14] br[14] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_17 
+ bl[15] br[15] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_18 
+ bl[16] br[16] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_19 
+ bl[17] br[17] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_20 
+ bl[18] br[18] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_21 
+ bl[19] br[19] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_22 
+ bl[20] br[20] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_23 
+ bl[21] br[21] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_24 
+ bl[22] br[22] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_25 
+ bl[23] br[23] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_26 
+ bl[24] br[24] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_27 
+ bl[25] br[25] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_28 
+ bl[26] br[26] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_29 
+ bl[27] br[27] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_30 
+ bl[28] br[28] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_31 
+ bl[29] br[29] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_32 
+ bl[30] br[30] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_33 
+ bl[31] br[31] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_34 
+ bl[32] br[32] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_35 
+ bl[33] br[33] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_36 
+ bl[34] br[34] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_37 
+ bl[35] br[35] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_38 
+ bl[36] br[36] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_39 
+ bl[37] br[37] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_40 
+ bl[38] br[38] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_41 
+ bl[39] br[39] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_42 
+ bl[40] br[40] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_43 
+ bl[41] br[41] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_44 
+ bl[42] br[42] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_45 
+ bl[43] br[43] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_46 
+ bl[44] br[44] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_47 
+ bl[45] br[45] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_48 
+ bl[46] br[46] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_49 
+ bl[47] br[47] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_50 
+ bl[48] br[48] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_51 
+ bl[49] br[49] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_52 
+ bl[50] br[50] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_53 
+ bl[51] br[51] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_54 
+ bl[52] br[52] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_55 
+ bl[53] br[53] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_56 
+ bl[54] br[54] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_57 
+ bl[55] br[55] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_58 
+ bl[56] br[56] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_59 
+ bl[57] br[57] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_60 
+ bl[58] br[58] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_61 
+ bl[59] br[59] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_62 
+ bl[60] br[60] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_63 
+ bl[61] br[61] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_64 
+ bl[62] br[62] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_65 
+ bl[63] br[63] vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_66 
+ vdd vdd vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_39_67 
+ vdd vdd vdd vss wl[37] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_0 
+ vdd vdd vss vdd vpb vnb wl[38] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_40_1 
+ rbl rbr vss vdd vpb vnb wl[38] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_40_2 
+ bl[0] br[0] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_3 
+ bl[1] br[1] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_4 
+ bl[2] br[2] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_5 
+ bl[3] br[3] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_6 
+ bl[4] br[4] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_7 
+ bl[5] br[5] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_8 
+ bl[6] br[6] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_9 
+ bl[7] br[7] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_10 
+ bl[8] br[8] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_11 
+ bl[9] br[9] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_12 
+ bl[10] br[10] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_13 
+ bl[11] br[11] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_14 
+ bl[12] br[12] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_15 
+ bl[13] br[13] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_16 
+ bl[14] br[14] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_17 
+ bl[15] br[15] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_18 
+ bl[16] br[16] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_19 
+ bl[17] br[17] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_20 
+ bl[18] br[18] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_21 
+ bl[19] br[19] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_22 
+ bl[20] br[20] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_23 
+ bl[21] br[21] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_24 
+ bl[22] br[22] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_25 
+ bl[23] br[23] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_26 
+ bl[24] br[24] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_27 
+ bl[25] br[25] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_28 
+ bl[26] br[26] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_29 
+ bl[27] br[27] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_30 
+ bl[28] br[28] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_31 
+ bl[29] br[29] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_32 
+ bl[30] br[30] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_33 
+ bl[31] br[31] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_34 
+ bl[32] br[32] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_35 
+ bl[33] br[33] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_36 
+ bl[34] br[34] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_37 
+ bl[35] br[35] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_38 
+ bl[36] br[36] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_39 
+ bl[37] br[37] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_40 
+ bl[38] br[38] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_41 
+ bl[39] br[39] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_42 
+ bl[40] br[40] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_43 
+ bl[41] br[41] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_44 
+ bl[42] br[42] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_45 
+ bl[43] br[43] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_46 
+ bl[44] br[44] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_47 
+ bl[45] br[45] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_48 
+ bl[46] br[46] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_49 
+ bl[47] br[47] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_50 
+ bl[48] br[48] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_51 
+ bl[49] br[49] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_52 
+ bl[50] br[50] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_53 
+ bl[51] br[51] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_54 
+ bl[52] br[52] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_55 
+ bl[53] br[53] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_56 
+ bl[54] br[54] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_57 
+ bl[55] br[55] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_58 
+ bl[56] br[56] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_59 
+ bl[57] br[57] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_60 
+ bl[58] br[58] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_61 
+ bl[59] br[59] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_62 
+ bl[60] br[60] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_63 
+ bl[61] br[61] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_64 
+ bl[62] br[62] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_65 
+ bl[63] br[63] vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_66 
+ vdd vdd vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_40_67 
+ vdd vdd vdd vss wl[38] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_0 
+ vdd vdd vss vdd vpb vnb wl[39] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_41_1 
+ rbl rbr vss vdd vpb vnb wl[39] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_41_2 
+ bl[0] br[0] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_3 
+ bl[1] br[1] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_4 
+ bl[2] br[2] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_5 
+ bl[3] br[3] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_6 
+ bl[4] br[4] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_7 
+ bl[5] br[5] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_8 
+ bl[6] br[6] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_9 
+ bl[7] br[7] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_10 
+ bl[8] br[8] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_11 
+ bl[9] br[9] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_12 
+ bl[10] br[10] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_13 
+ bl[11] br[11] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_14 
+ bl[12] br[12] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_15 
+ bl[13] br[13] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_16 
+ bl[14] br[14] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_17 
+ bl[15] br[15] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_18 
+ bl[16] br[16] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_19 
+ bl[17] br[17] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_20 
+ bl[18] br[18] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_21 
+ bl[19] br[19] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_22 
+ bl[20] br[20] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_23 
+ bl[21] br[21] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_24 
+ bl[22] br[22] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_25 
+ bl[23] br[23] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_26 
+ bl[24] br[24] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_27 
+ bl[25] br[25] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_28 
+ bl[26] br[26] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_29 
+ bl[27] br[27] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_30 
+ bl[28] br[28] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_31 
+ bl[29] br[29] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_32 
+ bl[30] br[30] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_33 
+ bl[31] br[31] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_34 
+ bl[32] br[32] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_35 
+ bl[33] br[33] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_36 
+ bl[34] br[34] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_37 
+ bl[35] br[35] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_38 
+ bl[36] br[36] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_39 
+ bl[37] br[37] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_40 
+ bl[38] br[38] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_41 
+ bl[39] br[39] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_42 
+ bl[40] br[40] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_43 
+ bl[41] br[41] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_44 
+ bl[42] br[42] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_45 
+ bl[43] br[43] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_46 
+ bl[44] br[44] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_47 
+ bl[45] br[45] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_48 
+ bl[46] br[46] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_49 
+ bl[47] br[47] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_50 
+ bl[48] br[48] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_51 
+ bl[49] br[49] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_52 
+ bl[50] br[50] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_53 
+ bl[51] br[51] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_54 
+ bl[52] br[52] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_55 
+ bl[53] br[53] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_56 
+ bl[54] br[54] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_57 
+ bl[55] br[55] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_58 
+ bl[56] br[56] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_59 
+ bl[57] br[57] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_60 
+ bl[58] br[58] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_61 
+ bl[59] br[59] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_62 
+ bl[60] br[60] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_63 
+ bl[61] br[61] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_64 
+ bl[62] br[62] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_65 
+ bl[63] br[63] vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_66 
+ vdd vdd vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_41_67 
+ vdd vdd vdd vss wl[39] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_0 
+ vdd vdd vss vdd vpb vnb wl[40] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_42_1 
+ rbl rbr vss vdd vpb vnb wl[40] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_42_2 
+ bl[0] br[0] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_3 
+ bl[1] br[1] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_4 
+ bl[2] br[2] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_5 
+ bl[3] br[3] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_6 
+ bl[4] br[4] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_7 
+ bl[5] br[5] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_8 
+ bl[6] br[6] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_9 
+ bl[7] br[7] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_10 
+ bl[8] br[8] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_11 
+ bl[9] br[9] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_12 
+ bl[10] br[10] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_13 
+ bl[11] br[11] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_14 
+ bl[12] br[12] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_15 
+ bl[13] br[13] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_16 
+ bl[14] br[14] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_17 
+ bl[15] br[15] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_18 
+ bl[16] br[16] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_19 
+ bl[17] br[17] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_20 
+ bl[18] br[18] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_21 
+ bl[19] br[19] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_22 
+ bl[20] br[20] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_23 
+ bl[21] br[21] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_24 
+ bl[22] br[22] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_25 
+ bl[23] br[23] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_26 
+ bl[24] br[24] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_27 
+ bl[25] br[25] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_28 
+ bl[26] br[26] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_29 
+ bl[27] br[27] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_30 
+ bl[28] br[28] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_31 
+ bl[29] br[29] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_32 
+ bl[30] br[30] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_33 
+ bl[31] br[31] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_34 
+ bl[32] br[32] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_35 
+ bl[33] br[33] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_36 
+ bl[34] br[34] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_37 
+ bl[35] br[35] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_38 
+ bl[36] br[36] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_39 
+ bl[37] br[37] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_40 
+ bl[38] br[38] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_41 
+ bl[39] br[39] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_42 
+ bl[40] br[40] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_43 
+ bl[41] br[41] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_44 
+ bl[42] br[42] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_45 
+ bl[43] br[43] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_46 
+ bl[44] br[44] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_47 
+ bl[45] br[45] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_48 
+ bl[46] br[46] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_49 
+ bl[47] br[47] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_50 
+ bl[48] br[48] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_51 
+ bl[49] br[49] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_52 
+ bl[50] br[50] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_53 
+ bl[51] br[51] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_54 
+ bl[52] br[52] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_55 
+ bl[53] br[53] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_56 
+ bl[54] br[54] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_57 
+ bl[55] br[55] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_58 
+ bl[56] br[56] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_59 
+ bl[57] br[57] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_60 
+ bl[58] br[58] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_61 
+ bl[59] br[59] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_62 
+ bl[60] br[60] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_63 
+ bl[61] br[61] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_64 
+ bl[62] br[62] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_65 
+ bl[63] br[63] vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_66 
+ vdd vdd vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_42_67 
+ vdd vdd vdd vss wl[40] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_0 
+ vdd vdd vss vdd vpb vnb wl[41] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_43_1 
+ rbl rbr vss vdd vpb vnb wl[41] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_43_2 
+ bl[0] br[0] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_3 
+ bl[1] br[1] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_4 
+ bl[2] br[2] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_5 
+ bl[3] br[3] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_6 
+ bl[4] br[4] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_7 
+ bl[5] br[5] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_8 
+ bl[6] br[6] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_9 
+ bl[7] br[7] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_10 
+ bl[8] br[8] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_11 
+ bl[9] br[9] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_12 
+ bl[10] br[10] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_13 
+ bl[11] br[11] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_14 
+ bl[12] br[12] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_15 
+ bl[13] br[13] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_16 
+ bl[14] br[14] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_17 
+ bl[15] br[15] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_18 
+ bl[16] br[16] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_19 
+ bl[17] br[17] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_20 
+ bl[18] br[18] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_21 
+ bl[19] br[19] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_22 
+ bl[20] br[20] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_23 
+ bl[21] br[21] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_24 
+ bl[22] br[22] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_25 
+ bl[23] br[23] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_26 
+ bl[24] br[24] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_27 
+ bl[25] br[25] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_28 
+ bl[26] br[26] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_29 
+ bl[27] br[27] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_30 
+ bl[28] br[28] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_31 
+ bl[29] br[29] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_32 
+ bl[30] br[30] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_33 
+ bl[31] br[31] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_34 
+ bl[32] br[32] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_35 
+ bl[33] br[33] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_36 
+ bl[34] br[34] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_37 
+ bl[35] br[35] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_38 
+ bl[36] br[36] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_39 
+ bl[37] br[37] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_40 
+ bl[38] br[38] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_41 
+ bl[39] br[39] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_42 
+ bl[40] br[40] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_43 
+ bl[41] br[41] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_44 
+ bl[42] br[42] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_45 
+ bl[43] br[43] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_46 
+ bl[44] br[44] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_47 
+ bl[45] br[45] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_48 
+ bl[46] br[46] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_49 
+ bl[47] br[47] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_50 
+ bl[48] br[48] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_51 
+ bl[49] br[49] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_52 
+ bl[50] br[50] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_53 
+ bl[51] br[51] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_54 
+ bl[52] br[52] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_55 
+ bl[53] br[53] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_56 
+ bl[54] br[54] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_57 
+ bl[55] br[55] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_58 
+ bl[56] br[56] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_59 
+ bl[57] br[57] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_60 
+ bl[58] br[58] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_61 
+ bl[59] br[59] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_62 
+ bl[60] br[60] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_63 
+ bl[61] br[61] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_64 
+ bl[62] br[62] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_65 
+ bl[63] br[63] vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_66 
+ vdd vdd vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_43_67 
+ vdd vdd vdd vss wl[41] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_0 
+ vdd vdd vss vdd vpb vnb wl[42] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_44_1 
+ rbl rbr vss vdd vpb vnb wl[42] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_44_2 
+ bl[0] br[0] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_3 
+ bl[1] br[1] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_4 
+ bl[2] br[2] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_5 
+ bl[3] br[3] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_6 
+ bl[4] br[4] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_7 
+ bl[5] br[5] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_8 
+ bl[6] br[6] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_9 
+ bl[7] br[7] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_10 
+ bl[8] br[8] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_11 
+ bl[9] br[9] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_12 
+ bl[10] br[10] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_13 
+ bl[11] br[11] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_14 
+ bl[12] br[12] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_15 
+ bl[13] br[13] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_16 
+ bl[14] br[14] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_17 
+ bl[15] br[15] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_18 
+ bl[16] br[16] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_19 
+ bl[17] br[17] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_20 
+ bl[18] br[18] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_21 
+ bl[19] br[19] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_22 
+ bl[20] br[20] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_23 
+ bl[21] br[21] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_24 
+ bl[22] br[22] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_25 
+ bl[23] br[23] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_26 
+ bl[24] br[24] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_27 
+ bl[25] br[25] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_28 
+ bl[26] br[26] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_29 
+ bl[27] br[27] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_30 
+ bl[28] br[28] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_31 
+ bl[29] br[29] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_32 
+ bl[30] br[30] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_33 
+ bl[31] br[31] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_34 
+ bl[32] br[32] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_35 
+ bl[33] br[33] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_36 
+ bl[34] br[34] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_37 
+ bl[35] br[35] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_38 
+ bl[36] br[36] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_39 
+ bl[37] br[37] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_40 
+ bl[38] br[38] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_41 
+ bl[39] br[39] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_42 
+ bl[40] br[40] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_43 
+ bl[41] br[41] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_44 
+ bl[42] br[42] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_45 
+ bl[43] br[43] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_46 
+ bl[44] br[44] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_47 
+ bl[45] br[45] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_48 
+ bl[46] br[46] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_49 
+ bl[47] br[47] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_50 
+ bl[48] br[48] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_51 
+ bl[49] br[49] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_52 
+ bl[50] br[50] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_53 
+ bl[51] br[51] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_54 
+ bl[52] br[52] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_55 
+ bl[53] br[53] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_56 
+ bl[54] br[54] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_57 
+ bl[55] br[55] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_58 
+ bl[56] br[56] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_59 
+ bl[57] br[57] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_60 
+ bl[58] br[58] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_61 
+ bl[59] br[59] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_62 
+ bl[60] br[60] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_63 
+ bl[61] br[61] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_64 
+ bl[62] br[62] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_65 
+ bl[63] br[63] vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_66 
+ vdd vdd vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_44_67 
+ vdd vdd vdd vss wl[42] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_0 
+ vdd vdd vss vdd vpb vnb wl[43] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_45_1 
+ rbl rbr vss vdd vpb vnb wl[43] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_45_2 
+ bl[0] br[0] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_3 
+ bl[1] br[1] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_4 
+ bl[2] br[2] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_5 
+ bl[3] br[3] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_6 
+ bl[4] br[4] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_7 
+ bl[5] br[5] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_8 
+ bl[6] br[6] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_9 
+ bl[7] br[7] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_10 
+ bl[8] br[8] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_11 
+ bl[9] br[9] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_12 
+ bl[10] br[10] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_13 
+ bl[11] br[11] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_14 
+ bl[12] br[12] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_15 
+ bl[13] br[13] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_16 
+ bl[14] br[14] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_17 
+ bl[15] br[15] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_18 
+ bl[16] br[16] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_19 
+ bl[17] br[17] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_20 
+ bl[18] br[18] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_21 
+ bl[19] br[19] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_22 
+ bl[20] br[20] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_23 
+ bl[21] br[21] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_24 
+ bl[22] br[22] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_25 
+ bl[23] br[23] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_26 
+ bl[24] br[24] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_27 
+ bl[25] br[25] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_28 
+ bl[26] br[26] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_29 
+ bl[27] br[27] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_30 
+ bl[28] br[28] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_31 
+ bl[29] br[29] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_32 
+ bl[30] br[30] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_33 
+ bl[31] br[31] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_34 
+ bl[32] br[32] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_35 
+ bl[33] br[33] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_36 
+ bl[34] br[34] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_37 
+ bl[35] br[35] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_38 
+ bl[36] br[36] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_39 
+ bl[37] br[37] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_40 
+ bl[38] br[38] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_41 
+ bl[39] br[39] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_42 
+ bl[40] br[40] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_43 
+ bl[41] br[41] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_44 
+ bl[42] br[42] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_45 
+ bl[43] br[43] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_46 
+ bl[44] br[44] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_47 
+ bl[45] br[45] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_48 
+ bl[46] br[46] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_49 
+ bl[47] br[47] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_50 
+ bl[48] br[48] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_51 
+ bl[49] br[49] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_52 
+ bl[50] br[50] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_53 
+ bl[51] br[51] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_54 
+ bl[52] br[52] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_55 
+ bl[53] br[53] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_56 
+ bl[54] br[54] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_57 
+ bl[55] br[55] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_58 
+ bl[56] br[56] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_59 
+ bl[57] br[57] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_60 
+ bl[58] br[58] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_61 
+ bl[59] br[59] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_62 
+ bl[60] br[60] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_63 
+ bl[61] br[61] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_64 
+ bl[62] br[62] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_65 
+ bl[63] br[63] vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_66 
+ vdd vdd vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_45_67 
+ vdd vdd vdd vss wl[43] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_0 
+ vdd vdd vss vdd vpb vnb wl[44] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_46_1 
+ rbl rbr vss vdd vpb vnb wl[44] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_46_2 
+ bl[0] br[0] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_3 
+ bl[1] br[1] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_4 
+ bl[2] br[2] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_5 
+ bl[3] br[3] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_6 
+ bl[4] br[4] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_7 
+ bl[5] br[5] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_8 
+ bl[6] br[6] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_9 
+ bl[7] br[7] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_10 
+ bl[8] br[8] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_11 
+ bl[9] br[9] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_12 
+ bl[10] br[10] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_13 
+ bl[11] br[11] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_14 
+ bl[12] br[12] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_15 
+ bl[13] br[13] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_16 
+ bl[14] br[14] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_17 
+ bl[15] br[15] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_18 
+ bl[16] br[16] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_19 
+ bl[17] br[17] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_20 
+ bl[18] br[18] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_21 
+ bl[19] br[19] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_22 
+ bl[20] br[20] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_23 
+ bl[21] br[21] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_24 
+ bl[22] br[22] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_25 
+ bl[23] br[23] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_26 
+ bl[24] br[24] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_27 
+ bl[25] br[25] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_28 
+ bl[26] br[26] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_29 
+ bl[27] br[27] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_30 
+ bl[28] br[28] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_31 
+ bl[29] br[29] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_32 
+ bl[30] br[30] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_33 
+ bl[31] br[31] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_34 
+ bl[32] br[32] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_35 
+ bl[33] br[33] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_36 
+ bl[34] br[34] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_37 
+ bl[35] br[35] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_38 
+ bl[36] br[36] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_39 
+ bl[37] br[37] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_40 
+ bl[38] br[38] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_41 
+ bl[39] br[39] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_42 
+ bl[40] br[40] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_43 
+ bl[41] br[41] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_44 
+ bl[42] br[42] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_45 
+ bl[43] br[43] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_46 
+ bl[44] br[44] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_47 
+ bl[45] br[45] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_48 
+ bl[46] br[46] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_49 
+ bl[47] br[47] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_50 
+ bl[48] br[48] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_51 
+ bl[49] br[49] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_52 
+ bl[50] br[50] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_53 
+ bl[51] br[51] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_54 
+ bl[52] br[52] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_55 
+ bl[53] br[53] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_56 
+ bl[54] br[54] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_57 
+ bl[55] br[55] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_58 
+ bl[56] br[56] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_59 
+ bl[57] br[57] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_60 
+ bl[58] br[58] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_61 
+ bl[59] br[59] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_62 
+ bl[60] br[60] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_63 
+ bl[61] br[61] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_64 
+ bl[62] br[62] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_65 
+ bl[63] br[63] vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_66 
+ vdd vdd vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_46_67 
+ vdd vdd vdd vss wl[44] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_0 
+ vdd vdd vss vdd vpb vnb wl[45] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_47_1 
+ rbl rbr vss vdd vpb vnb wl[45] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_47_2 
+ bl[0] br[0] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_3 
+ bl[1] br[1] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_4 
+ bl[2] br[2] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_5 
+ bl[3] br[3] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_6 
+ bl[4] br[4] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_7 
+ bl[5] br[5] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_8 
+ bl[6] br[6] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_9 
+ bl[7] br[7] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_10 
+ bl[8] br[8] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_11 
+ bl[9] br[9] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_12 
+ bl[10] br[10] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_13 
+ bl[11] br[11] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_14 
+ bl[12] br[12] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_15 
+ bl[13] br[13] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_16 
+ bl[14] br[14] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_17 
+ bl[15] br[15] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_18 
+ bl[16] br[16] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_19 
+ bl[17] br[17] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_20 
+ bl[18] br[18] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_21 
+ bl[19] br[19] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_22 
+ bl[20] br[20] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_23 
+ bl[21] br[21] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_24 
+ bl[22] br[22] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_25 
+ bl[23] br[23] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_26 
+ bl[24] br[24] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_27 
+ bl[25] br[25] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_28 
+ bl[26] br[26] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_29 
+ bl[27] br[27] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_30 
+ bl[28] br[28] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_31 
+ bl[29] br[29] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_32 
+ bl[30] br[30] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_33 
+ bl[31] br[31] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_34 
+ bl[32] br[32] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_35 
+ bl[33] br[33] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_36 
+ bl[34] br[34] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_37 
+ bl[35] br[35] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_38 
+ bl[36] br[36] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_39 
+ bl[37] br[37] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_40 
+ bl[38] br[38] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_41 
+ bl[39] br[39] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_42 
+ bl[40] br[40] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_43 
+ bl[41] br[41] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_44 
+ bl[42] br[42] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_45 
+ bl[43] br[43] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_46 
+ bl[44] br[44] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_47 
+ bl[45] br[45] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_48 
+ bl[46] br[46] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_49 
+ bl[47] br[47] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_50 
+ bl[48] br[48] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_51 
+ bl[49] br[49] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_52 
+ bl[50] br[50] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_53 
+ bl[51] br[51] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_54 
+ bl[52] br[52] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_55 
+ bl[53] br[53] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_56 
+ bl[54] br[54] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_57 
+ bl[55] br[55] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_58 
+ bl[56] br[56] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_59 
+ bl[57] br[57] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_60 
+ bl[58] br[58] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_61 
+ bl[59] br[59] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_62 
+ bl[60] br[60] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_63 
+ bl[61] br[61] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_64 
+ bl[62] br[62] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_65 
+ bl[63] br[63] vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_66 
+ vdd vdd vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_47_67 
+ vdd vdd vdd vss wl[45] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_0 
+ vdd vdd vss vdd vpb vnb wl[46] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_48_1 
+ rbl rbr vss vdd vpb vnb wl[46] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_48_2 
+ bl[0] br[0] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_3 
+ bl[1] br[1] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_4 
+ bl[2] br[2] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_5 
+ bl[3] br[3] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_6 
+ bl[4] br[4] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_7 
+ bl[5] br[5] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_8 
+ bl[6] br[6] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_9 
+ bl[7] br[7] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_10 
+ bl[8] br[8] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_11 
+ bl[9] br[9] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_12 
+ bl[10] br[10] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_13 
+ bl[11] br[11] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_14 
+ bl[12] br[12] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_15 
+ bl[13] br[13] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_16 
+ bl[14] br[14] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_17 
+ bl[15] br[15] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_18 
+ bl[16] br[16] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_19 
+ bl[17] br[17] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_20 
+ bl[18] br[18] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_21 
+ bl[19] br[19] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_22 
+ bl[20] br[20] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_23 
+ bl[21] br[21] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_24 
+ bl[22] br[22] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_25 
+ bl[23] br[23] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_26 
+ bl[24] br[24] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_27 
+ bl[25] br[25] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_28 
+ bl[26] br[26] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_29 
+ bl[27] br[27] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_30 
+ bl[28] br[28] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_31 
+ bl[29] br[29] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_32 
+ bl[30] br[30] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_33 
+ bl[31] br[31] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_34 
+ bl[32] br[32] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_35 
+ bl[33] br[33] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_36 
+ bl[34] br[34] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_37 
+ bl[35] br[35] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_38 
+ bl[36] br[36] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_39 
+ bl[37] br[37] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_40 
+ bl[38] br[38] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_41 
+ bl[39] br[39] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_42 
+ bl[40] br[40] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_43 
+ bl[41] br[41] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_44 
+ bl[42] br[42] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_45 
+ bl[43] br[43] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_46 
+ bl[44] br[44] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_47 
+ bl[45] br[45] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_48 
+ bl[46] br[46] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_49 
+ bl[47] br[47] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_50 
+ bl[48] br[48] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_51 
+ bl[49] br[49] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_52 
+ bl[50] br[50] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_53 
+ bl[51] br[51] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_54 
+ bl[52] br[52] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_55 
+ bl[53] br[53] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_56 
+ bl[54] br[54] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_57 
+ bl[55] br[55] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_58 
+ bl[56] br[56] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_59 
+ bl[57] br[57] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_60 
+ bl[58] br[58] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_61 
+ bl[59] br[59] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_62 
+ bl[60] br[60] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_63 
+ bl[61] br[61] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_64 
+ bl[62] br[62] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_65 
+ bl[63] br[63] vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_66 
+ vdd vdd vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_48_67 
+ vdd vdd vdd vss wl[46] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_0 
+ vdd vdd vss vdd vpb vnb wl[47] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_49_1 
+ rbl rbr vss vdd vpb vnb wl[47] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_49_2 
+ bl[0] br[0] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_3 
+ bl[1] br[1] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_4 
+ bl[2] br[2] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_5 
+ bl[3] br[3] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_6 
+ bl[4] br[4] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_7 
+ bl[5] br[5] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_8 
+ bl[6] br[6] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_9 
+ bl[7] br[7] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_10 
+ bl[8] br[8] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_11 
+ bl[9] br[9] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_12 
+ bl[10] br[10] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_13 
+ bl[11] br[11] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_14 
+ bl[12] br[12] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_15 
+ bl[13] br[13] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_16 
+ bl[14] br[14] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_17 
+ bl[15] br[15] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_18 
+ bl[16] br[16] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_19 
+ bl[17] br[17] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_20 
+ bl[18] br[18] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_21 
+ bl[19] br[19] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_22 
+ bl[20] br[20] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_23 
+ bl[21] br[21] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_24 
+ bl[22] br[22] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_25 
+ bl[23] br[23] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_26 
+ bl[24] br[24] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_27 
+ bl[25] br[25] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_28 
+ bl[26] br[26] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_29 
+ bl[27] br[27] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_30 
+ bl[28] br[28] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_31 
+ bl[29] br[29] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_32 
+ bl[30] br[30] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_33 
+ bl[31] br[31] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_34 
+ bl[32] br[32] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_35 
+ bl[33] br[33] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_36 
+ bl[34] br[34] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_37 
+ bl[35] br[35] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_38 
+ bl[36] br[36] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_39 
+ bl[37] br[37] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_40 
+ bl[38] br[38] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_41 
+ bl[39] br[39] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_42 
+ bl[40] br[40] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_43 
+ bl[41] br[41] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_44 
+ bl[42] br[42] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_45 
+ bl[43] br[43] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_46 
+ bl[44] br[44] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_47 
+ bl[45] br[45] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_48 
+ bl[46] br[46] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_49 
+ bl[47] br[47] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_50 
+ bl[48] br[48] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_51 
+ bl[49] br[49] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_52 
+ bl[50] br[50] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_53 
+ bl[51] br[51] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_54 
+ bl[52] br[52] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_55 
+ bl[53] br[53] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_56 
+ bl[54] br[54] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_57 
+ bl[55] br[55] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_58 
+ bl[56] br[56] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_59 
+ bl[57] br[57] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_60 
+ bl[58] br[58] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_61 
+ bl[59] br[59] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_62 
+ bl[60] br[60] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_63 
+ bl[61] br[61] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_64 
+ bl[62] br[62] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_65 
+ bl[63] br[63] vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_66 
+ vdd vdd vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_49_67 
+ vdd vdd vdd vss wl[47] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_0 
+ vdd vdd vss vdd vpb vnb wl[48] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_50_1 
+ rbl rbr vss vdd vpb vnb wl[48] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_50_2 
+ bl[0] br[0] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_3 
+ bl[1] br[1] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_4 
+ bl[2] br[2] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_5 
+ bl[3] br[3] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_6 
+ bl[4] br[4] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_7 
+ bl[5] br[5] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_8 
+ bl[6] br[6] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_9 
+ bl[7] br[7] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_10 
+ bl[8] br[8] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_11 
+ bl[9] br[9] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_12 
+ bl[10] br[10] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_13 
+ bl[11] br[11] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_14 
+ bl[12] br[12] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_15 
+ bl[13] br[13] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_16 
+ bl[14] br[14] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_17 
+ bl[15] br[15] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_18 
+ bl[16] br[16] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_19 
+ bl[17] br[17] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_20 
+ bl[18] br[18] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_21 
+ bl[19] br[19] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_22 
+ bl[20] br[20] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_23 
+ bl[21] br[21] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_24 
+ bl[22] br[22] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_25 
+ bl[23] br[23] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_26 
+ bl[24] br[24] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_27 
+ bl[25] br[25] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_28 
+ bl[26] br[26] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_29 
+ bl[27] br[27] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_30 
+ bl[28] br[28] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_31 
+ bl[29] br[29] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_32 
+ bl[30] br[30] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_33 
+ bl[31] br[31] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_34 
+ bl[32] br[32] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_35 
+ bl[33] br[33] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_36 
+ bl[34] br[34] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_37 
+ bl[35] br[35] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_38 
+ bl[36] br[36] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_39 
+ bl[37] br[37] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_40 
+ bl[38] br[38] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_41 
+ bl[39] br[39] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_42 
+ bl[40] br[40] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_43 
+ bl[41] br[41] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_44 
+ bl[42] br[42] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_45 
+ bl[43] br[43] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_46 
+ bl[44] br[44] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_47 
+ bl[45] br[45] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_48 
+ bl[46] br[46] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_49 
+ bl[47] br[47] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_50 
+ bl[48] br[48] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_51 
+ bl[49] br[49] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_52 
+ bl[50] br[50] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_53 
+ bl[51] br[51] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_54 
+ bl[52] br[52] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_55 
+ bl[53] br[53] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_56 
+ bl[54] br[54] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_57 
+ bl[55] br[55] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_58 
+ bl[56] br[56] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_59 
+ bl[57] br[57] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_60 
+ bl[58] br[58] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_61 
+ bl[59] br[59] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_62 
+ bl[60] br[60] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_63 
+ bl[61] br[61] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_64 
+ bl[62] br[62] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_65 
+ bl[63] br[63] vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_66 
+ vdd vdd vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_50_67 
+ vdd vdd vdd vss wl[48] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_0 
+ vdd vdd vss vdd vpb vnb wl[49] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_51_1 
+ rbl rbr vss vdd vpb vnb wl[49] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_51_2 
+ bl[0] br[0] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_3 
+ bl[1] br[1] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_4 
+ bl[2] br[2] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_5 
+ bl[3] br[3] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_6 
+ bl[4] br[4] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_7 
+ bl[5] br[5] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_8 
+ bl[6] br[6] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_9 
+ bl[7] br[7] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_10 
+ bl[8] br[8] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_11 
+ bl[9] br[9] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_12 
+ bl[10] br[10] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_13 
+ bl[11] br[11] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_14 
+ bl[12] br[12] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_15 
+ bl[13] br[13] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_16 
+ bl[14] br[14] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_17 
+ bl[15] br[15] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_18 
+ bl[16] br[16] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_19 
+ bl[17] br[17] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_20 
+ bl[18] br[18] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_21 
+ bl[19] br[19] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_22 
+ bl[20] br[20] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_23 
+ bl[21] br[21] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_24 
+ bl[22] br[22] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_25 
+ bl[23] br[23] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_26 
+ bl[24] br[24] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_27 
+ bl[25] br[25] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_28 
+ bl[26] br[26] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_29 
+ bl[27] br[27] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_30 
+ bl[28] br[28] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_31 
+ bl[29] br[29] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_32 
+ bl[30] br[30] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_33 
+ bl[31] br[31] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_34 
+ bl[32] br[32] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_35 
+ bl[33] br[33] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_36 
+ bl[34] br[34] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_37 
+ bl[35] br[35] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_38 
+ bl[36] br[36] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_39 
+ bl[37] br[37] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_40 
+ bl[38] br[38] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_41 
+ bl[39] br[39] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_42 
+ bl[40] br[40] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_43 
+ bl[41] br[41] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_44 
+ bl[42] br[42] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_45 
+ bl[43] br[43] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_46 
+ bl[44] br[44] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_47 
+ bl[45] br[45] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_48 
+ bl[46] br[46] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_49 
+ bl[47] br[47] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_50 
+ bl[48] br[48] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_51 
+ bl[49] br[49] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_52 
+ bl[50] br[50] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_53 
+ bl[51] br[51] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_54 
+ bl[52] br[52] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_55 
+ bl[53] br[53] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_56 
+ bl[54] br[54] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_57 
+ bl[55] br[55] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_58 
+ bl[56] br[56] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_59 
+ bl[57] br[57] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_60 
+ bl[58] br[58] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_61 
+ bl[59] br[59] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_62 
+ bl[60] br[60] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_63 
+ bl[61] br[61] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_64 
+ bl[62] br[62] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_65 
+ bl[63] br[63] vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_66 
+ vdd vdd vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_51_67 
+ vdd vdd vdd vss wl[49] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_0 
+ vdd vdd vss vdd vpb vnb wl[50] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_52_1 
+ rbl rbr vss vdd vpb vnb wl[50] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_52_2 
+ bl[0] br[0] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_3 
+ bl[1] br[1] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_4 
+ bl[2] br[2] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_5 
+ bl[3] br[3] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_6 
+ bl[4] br[4] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_7 
+ bl[5] br[5] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_8 
+ bl[6] br[6] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_9 
+ bl[7] br[7] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_10 
+ bl[8] br[8] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_11 
+ bl[9] br[9] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_12 
+ bl[10] br[10] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_13 
+ bl[11] br[11] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_14 
+ bl[12] br[12] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_15 
+ bl[13] br[13] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_16 
+ bl[14] br[14] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_17 
+ bl[15] br[15] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_18 
+ bl[16] br[16] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_19 
+ bl[17] br[17] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_20 
+ bl[18] br[18] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_21 
+ bl[19] br[19] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_22 
+ bl[20] br[20] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_23 
+ bl[21] br[21] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_24 
+ bl[22] br[22] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_25 
+ bl[23] br[23] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_26 
+ bl[24] br[24] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_27 
+ bl[25] br[25] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_28 
+ bl[26] br[26] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_29 
+ bl[27] br[27] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_30 
+ bl[28] br[28] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_31 
+ bl[29] br[29] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_32 
+ bl[30] br[30] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_33 
+ bl[31] br[31] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_34 
+ bl[32] br[32] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_35 
+ bl[33] br[33] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_36 
+ bl[34] br[34] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_37 
+ bl[35] br[35] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_38 
+ bl[36] br[36] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_39 
+ bl[37] br[37] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_40 
+ bl[38] br[38] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_41 
+ bl[39] br[39] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_42 
+ bl[40] br[40] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_43 
+ bl[41] br[41] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_44 
+ bl[42] br[42] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_45 
+ bl[43] br[43] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_46 
+ bl[44] br[44] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_47 
+ bl[45] br[45] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_48 
+ bl[46] br[46] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_49 
+ bl[47] br[47] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_50 
+ bl[48] br[48] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_51 
+ bl[49] br[49] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_52 
+ bl[50] br[50] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_53 
+ bl[51] br[51] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_54 
+ bl[52] br[52] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_55 
+ bl[53] br[53] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_56 
+ bl[54] br[54] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_57 
+ bl[55] br[55] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_58 
+ bl[56] br[56] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_59 
+ bl[57] br[57] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_60 
+ bl[58] br[58] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_61 
+ bl[59] br[59] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_62 
+ bl[60] br[60] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_63 
+ bl[61] br[61] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_64 
+ bl[62] br[62] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_65 
+ bl[63] br[63] vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_66 
+ vdd vdd vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_52_67 
+ vdd vdd vdd vss wl[50] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_0 
+ vdd vdd vss vdd vpb vnb wl[51] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_53_1 
+ rbl rbr vss vdd vpb vnb wl[51] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_53_2 
+ bl[0] br[0] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_3 
+ bl[1] br[1] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_4 
+ bl[2] br[2] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_5 
+ bl[3] br[3] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_6 
+ bl[4] br[4] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_7 
+ bl[5] br[5] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_8 
+ bl[6] br[6] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_9 
+ bl[7] br[7] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_10 
+ bl[8] br[8] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_11 
+ bl[9] br[9] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_12 
+ bl[10] br[10] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_13 
+ bl[11] br[11] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_14 
+ bl[12] br[12] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_15 
+ bl[13] br[13] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_16 
+ bl[14] br[14] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_17 
+ bl[15] br[15] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_18 
+ bl[16] br[16] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_19 
+ bl[17] br[17] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_20 
+ bl[18] br[18] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_21 
+ bl[19] br[19] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_22 
+ bl[20] br[20] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_23 
+ bl[21] br[21] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_24 
+ bl[22] br[22] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_25 
+ bl[23] br[23] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_26 
+ bl[24] br[24] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_27 
+ bl[25] br[25] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_28 
+ bl[26] br[26] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_29 
+ bl[27] br[27] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_30 
+ bl[28] br[28] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_31 
+ bl[29] br[29] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_32 
+ bl[30] br[30] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_33 
+ bl[31] br[31] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_34 
+ bl[32] br[32] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_35 
+ bl[33] br[33] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_36 
+ bl[34] br[34] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_37 
+ bl[35] br[35] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_38 
+ bl[36] br[36] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_39 
+ bl[37] br[37] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_40 
+ bl[38] br[38] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_41 
+ bl[39] br[39] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_42 
+ bl[40] br[40] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_43 
+ bl[41] br[41] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_44 
+ bl[42] br[42] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_45 
+ bl[43] br[43] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_46 
+ bl[44] br[44] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_47 
+ bl[45] br[45] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_48 
+ bl[46] br[46] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_49 
+ bl[47] br[47] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_50 
+ bl[48] br[48] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_51 
+ bl[49] br[49] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_52 
+ bl[50] br[50] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_53 
+ bl[51] br[51] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_54 
+ bl[52] br[52] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_55 
+ bl[53] br[53] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_56 
+ bl[54] br[54] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_57 
+ bl[55] br[55] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_58 
+ bl[56] br[56] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_59 
+ bl[57] br[57] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_60 
+ bl[58] br[58] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_61 
+ bl[59] br[59] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_62 
+ bl[60] br[60] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_63 
+ bl[61] br[61] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_64 
+ bl[62] br[62] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_65 
+ bl[63] br[63] vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_66 
+ vdd vdd vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_53_67 
+ vdd vdd vdd vss wl[51] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_0 
+ vdd vdd vss vdd vpb vnb wl[52] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_54_1 
+ rbl rbr vss vdd vpb vnb wl[52] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_54_2 
+ bl[0] br[0] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_3 
+ bl[1] br[1] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_4 
+ bl[2] br[2] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_5 
+ bl[3] br[3] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_6 
+ bl[4] br[4] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_7 
+ bl[5] br[5] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_8 
+ bl[6] br[6] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_9 
+ bl[7] br[7] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_10 
+ bl[8] br[8] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_11 
+ bl[9] br[9] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_12 
+ bl[10] br[10] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_13 
+ bl[11] br[11] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_14 
+ bl[12] br[12] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_15 
+ bl[13] br[13] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_16 
+ bl[14] br[14] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_17 
+ bl[15] br[15] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_18 
+ bl[16] br[16] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_19 
+ bl[17] br[17] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_20 
+ bl[18] br[18] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_21 
+ bl[19] br[19] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_22 
+ bl[20] br[20] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_23 
+ bl[21] br[21] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_24 
+ bl[22] br[22] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_25 
+ bl[23] br[23] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_26 
+ bl[24] br[24] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_27 
+ bl[25] br[25] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_28 
+ bl[26] br[26] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_29 
+ bl[27] br[27] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_30 
+ bl[28] br[28] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_31 
+ bl[29] br[29] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_32 
+ bl[30] br[30] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_33 
+ bl[31] br[31] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_34 
+ bl[32] br[32] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_35 
+ bl[33] br[33] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_36 
+ bl[34] br[34] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_37 
+ bl[35] br[35] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_38 
+ bl[36] br[36] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_39 
+ bl[37] br[37] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_40 
+ bl[38] br[38] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_41 
+ bl[39] br[39] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_42 
+ bl[40] br[40] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_43 
+ bl[41] br[41] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_44 
+ bl[42] br[42] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_45 
+ bl[43] br[43] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_46 
+ bl[44] br[44] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_47 
+ bl[45] br[45] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_48 
+ bl[46] br[46] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_49 
+ bl[47] br[47] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_50 
+ bl[48] br[48] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_51 
+ bl[49] br[49] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_52 
+ bl[50] br[50] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_53 
+ bl[51] br[51] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_54 
+ bl[52] br[52] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_55 
+ bl[53] br[53] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_56 
+ bl[54] br[54] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_57 
+ bl[55] br[55] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_58 
+ bl[56] br[56] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_59 
+ bl[57] br[57] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_60 
+ bl[58] br[58] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_61 
+ bl[59] br[59] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_62 
+ bl[60] br[60] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_63 
+ bl[61] br[61] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_64 
+ bl[62] br[62] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_65 
+ bl[63] br[63] vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_66 
+ vdd vdd vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_54_67 
+ vdd vdd vdd vss wl[52] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_0 
+ vdd vdd vss vdd vpb vnb wl[53] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_55_1 
+ rbl rbr vss vdd vpb vnb wl[53] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_55_2 
+ bl[0] br[0] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_3 
+ bl[1] br[1] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_4 
+ bl[2] br[2] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_5 
+ bl[3] br[3] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_6 
+ bl[4] br[4] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_7 
+ bl[5] br[5] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_8 
+ bl[6] br[6] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_9 
+ bl[7] br[7] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_10 
+ bl[8] br[8] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_11 
+ bl[9] br[9] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_12 
+ bl[10] br[10] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_13 
+ bl[11] br[11] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_14 
+ bl[12] br[12] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_15 
+ bl[13] br[13] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_16 
+ bl[14] br[14] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_17 
+ bl[15] br[15] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_18 
+ bl[16] br[16] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_19 
+ bl[17] br[17] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_20 
+ bl[18] br[18] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_21 
+ bl[19] br[19] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_22 
+ bl[20] br[20] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_23 
+ bl[21] br[21] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_24 
+ bl[22] br[22] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_25 
+ bl[23] br[23] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_26 
+ bl[24] br[24] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_27 
+ bl[25] br[25] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_28 
+ bl[26] br[26] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_29 
+ bl[27] br[27] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_30 
+ bl[28] br[28] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_31 
+ bl[29] br[29] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_32 
+ bl[30] br[30] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_33 
+ bl[31] br[31] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_34 
+ bl[32] br[32] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_35 
+ bl[33] br[33] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_36 
+ bl[34] br[34] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_37 
+ bl[35] br[35] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_38 
+ bl[36] br[36] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_39 
+ bl[37] br[37] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_40 
+ bl[38] br[38] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_41 
+ bl[39] br[39] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_42 
+ bl[40] br[40] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_43 
+ bl[41] br[41] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_44 
+ bl[42] br[42] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_45 
+ bl[43] br[43] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_46 
+ bl[44] br[44] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_47 
+ bl[45] br[45] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_48 
+ bl[46] br[46] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_49 
+ bl[47] br[47] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_50 
+ bl[48] br[48] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_51 
+ bl[49] br[49] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_52 
+ bl[50] br[50] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_53 
+ bl[51] br[51] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_54 
+ bl[52] br[52] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_55 
+ bl[53] br[53] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_56 
+ bl[54] br[54] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_57 
+ bl[55] br[55] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_58 
+ bl[56] br[56] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_59 
+ bl[57] br[57] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_60 
+ bl[58] br[58] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_61 
+ bl[59] br[59] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_62 
+ bl[60] br[60] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_63 
+ bl[61] br[61] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_64 
+ bl[62] br[62] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_65 
+ bl[63] br[63] vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_66 
+ vdd vdd vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_55_67 
+ vdd vdd vdd vss wl[53] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_0 
+ vdd vdd vss vdd vpb vnb wl[54] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_56_1 
+ rbl rbr vss vdd vpb vnb wl[54] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_56_2 
+ bl[0] br[0] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_3 
+ bl[1] br[1] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_4 
+ bl[2] br[2] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_5 
+ bl[3] br[3] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_6 
+ bl[4] br[4] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_7 
+ bl[5] br[5] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_8 
+ bl[6] br[6] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_9 
+ bl[7] br[7] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_10 
+ bl[8] br[8] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_11 
+ bl[9] br[9] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_12 
+ bl[10] br[10] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_13 
+ bl[11] br[11] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_14 
+ bl[12] br[12] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_15 
+ bl[13] br[13] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_16 
+ bl[14] br[14] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_17 
+ bl[15] br[15] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_18 
+ bl[16] br[16] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_19 
+ bl[17] br[17] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_20 
+ bl[18] br[18] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_21 
+ bl[19] br[19] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_22 
+ bl[20] br[20] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_23 
+ bl[21] br[21] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_24 
+ bl[22] br[22] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_25 
+ bl[23] br[23] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_26 
+ bl[24] br[24] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_27 
+ bl[25] br[25] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_28 
+ bl[26] br[26] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_29 
+ bl[27] br[27] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_30 
+ bl[28] br[28] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_31 
+ bl[29] br[29] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_32 
+ bl[30] br[30] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_33 
+ bl[31] br[31] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_34 
+ bl[32] br[32] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_35 
+ bl[33] br[33] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_36 
+ bl[34] br[34] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_37 
+ bl[35] br[35] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_38 
+ bl[36] br[36] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_39 
+ bl[37] br[37] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_40 
+ bl[38] br[38] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_41 
+ bl[39] br[39] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_42 
+ bl[40] br[40] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_43 
+ bl[41] br[41] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_44 
+ bl[42] br[42] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_45 
+ bl[43] br[43] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_46 
+ bl[44] br[44] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_47 
+ bl[45] br[45] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_48 
+ bl[46] br[46] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_49 
+ bl[47] br[47] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_50 
+ bl[48] br[48] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_51 
+ bl[49] br[49] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_52 
+ bl[50] br[50] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_53 
+ bl[51] br[51] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_54 
+ bl[52] br[52] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_55 
+ bl[53] br[53] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_56 
+ bl[54] br[54] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_57 
+ bl[55] br[55] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_58 
+ bl[56] br[56] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_59 
+ bl[57] br[57] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_60 
+ bl[58] br[58] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_61 
+ bl[59] br[59] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_62 
+ bl[60] br[60] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_63 
+ bl[61] br[61] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_64 
+ bl[62] br[62] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_65 
+ bl[63] br[63] vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_66 
+ vdd vdd vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_56_67 
+ vdd vdd vdd vss wl[54] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_0 
+ vdd vdd vss vdd vpb vnb wl[55] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_57_1 
+ rbl rbr vss vdd vpb vnb wl[55] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_57_2 
+ bl[0] br[0] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_3 
+ bl[1] br[1] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_4 
+ bl[2] br[2] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_5 
+ bl[3] br[3] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_6 
+ bl[4] br[4] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_7 
+ bl[5] br[5] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_8 
+ bl[6] br[6] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_9 
+ bl[7] br[7] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_10 
+ bl[8] br[8] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_11 
+ bl[9] br[9] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_12 
+ bl[10] br[10] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_13 
+ bl[11] br[11] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_14 
+ bl[12] br[12] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_15 
+ bl[13] br[13] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_16 
+ bl[14] br[14] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_17 
+ bl[15] br[15] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_18 
+ bl[16] br[16] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_19 
+ bl[17] br[17] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_20 
+ bl[18] br[18] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_21 
+ bl[19] br[19] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_22 
+ bl[20] br[20] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_23 
+ bl[21] br[21] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_24 
+ bl[22] br[22] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_25 
+ bl[23] br[23] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_26 
+ bl[24] br[24] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_27 
+ bl[25] br[25] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_28 
+ bl[26] br[26] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_29 
+ bl[27] br[27] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_30 
+ bl[28] br[28] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_31 
+ bl[29] br[29] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_32 
+ bl[30] br[30] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_33 
+ bl[31] br[31] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_34 
+ bl[32] br[32] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_35 
+ bl[33] br[33] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_36 
+ bl[34] br[34] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_37 
+ bl[35] br[35] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_38 
+ bl[36] br[36] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_39 
+ bl[37] br[37] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_40 
+ bl[38] br[38] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_41 
+ bl[39] br[39] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_42 
+ bl[40] br[40] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_43 
+ bl[41] br[41] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_44 
+ bl[42] br[42] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_45 
+ bl[43] br[43] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_46 
+ bl[44] br[44] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_47 
+ bl[45] br[45] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_48 
+ bl[46] br[46] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_49 
+ bl[47] br[47] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_50 
+ bl[48] br[48] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_51 
+ bl[49] br[49] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_52 
+ bl[50] br[50] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_53 
+ bl[51] br[51] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_54 
+ bl[52] br[52] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_55 
+ bl[53] br[53] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_56 
+ bl[54] br[54] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_57 
+ bl[55] br[55] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_58 
+ bl[56] br[56] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_59 
+ bl[57] br[57] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_60 
+ bl[58] br[58] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_61 
+ bl[59] br[59] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_62 
+ bl[60] br[60] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_63 
+ bl[61] br[61] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_64 
+ bl[62] br[62] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_65 
+ bl[63] br[63] vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_66 
+ vdd vdd vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_57_67 
+ vdd vdd vdd vss wl[55] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_0 
+ vdd vdd vss vdd vpb vnb wl[56] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_58_1 
+ rbl rbr vss vdd vpb vnb wl[56] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_58_2 
+ bl[0] br[0] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_3 
+ bl[1] br[1] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_4 
+ bl[2] br[2] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_5 
+ bl[3] br[3] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_6 
+ bl[4] br[4] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_7 
+ bl[5] br[5] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_8 
+ bl[6] br[6] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_9 
+ bl[7] br[7] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_10 
+ bl[8] br[8] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_11 
+ bl[9] br[9] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_12 
+ bl[10] br[10] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_13 
+ bl[11] br[11] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_14 
+ bl[12] br[12] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_15 
+ bl[13] br[13] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_16 
+ bl[14] br[14] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_17 
+ bl[15] br[15] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_18 
+ bl[16] br[16] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_19 
+ bl[17] br[17] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_20 
+ bl[18] br[18] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_21 
+ bl[19] br[19] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_22 
+ bl[20] br[20] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_23 
+ bl[21] br[21] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_24 
+ bl[22] br[22] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_25 
+ bl[23] br[23] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_26 
+ bl[24] br[24] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_27 
+ bl[25] br[25] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_28 
+ bl[26] br[26] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_29 
+ bl[27] br[27] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_30 
+ bl[28] br[28] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_31 
+ bl[29] br[29] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_32 
+ bl[30] br[30] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_33 
+ bl[31] br[31] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_34 
+ bl[32] br[32] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_35 
+ bl[33] br[33] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_36 
+ bl[34] br[34] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_37 
+ bl[35] br[35] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_38 
+ bl[36] br[36] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_39 
+ bl[37] br[37] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_40 
+ bl[38] br[38] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_41 
+ bl[39] br[39] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_42 
+ bl[40] br[40] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_43 
+ bl[41] br[41] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_44 
+ bl[42] br[42] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_45 
+ bl[43] br[43] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_46 
+ bl[44] br[44] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_47 
+ bl[45] br[45] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_48 
+ bl[46] br[46] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_49 
+ bl[47] br[47] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_50 
+ bl[48] br[48] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_51 
+ bl[49] br[49] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_52 
+ bl[50] br[50] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_53 
+ bl[51] br[51] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_54 
+ bl[52] br[52] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_55 
+ bl[53] br[53] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_56 
+ bl[54] br[54] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_57 
+ bl[55] br[55] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_58 
+ bl[56] br[56] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_59 
+ bl[57] br[57] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_60 
+ bl[58] br[58] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_61 
+ bl[59] br[59] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_62 
+ bl[60] br[60] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_63 
+ bl[61] br[61] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_64 
+ bl[62] br[62] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_65 
+ bl[63] br[63] vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_66 
+ vdd vdd vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_58_67 
+ vdd vdd vdd vss wl[56] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_0 
+ vdd vdd vss vdd vpb vnb wl[57] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_59_1 
+ rbl rbr vss vdd vpb vnb wl[57] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_59_2 
+ bl[0] br[0] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_3 
+ bl[1] br[1] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_4 
+ bl[2] br[2] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_5 
+ bl[3] br[3] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_6 
+ bl[4] br[4] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_7 
+ bl[5] br[5] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_8 
+ bl[6] br[6] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_9 
+ bl[7] br[7] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_10 
+ bl[8] br[8] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_11 
+ bl[9] br[9] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_12 
+ bl[10] br[10] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_13 
+ bl[11] br[11] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_14 
+ bl[12] br[12] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_15 
+ bl[13] br[13] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_16 
+ bl[14] br[14] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_17 
+ bl[15] br[15] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_18 
+ bl[16] br[16] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_19 
+ bl[17] br[17] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_20 
+ bl[18] br[18] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_21 
+ bl[19] br[19] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_22 
+ bl[20] br[20] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_23 
+ bl[21] br[21] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_24 
+ bl[22] br[22] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_25 
+ bl[23] br[23] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_26 
+ bl[24] br[24] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_27 
+ bl[25] br[25] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_28 
+ bl[26] br[26] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_29 
+ bl[27] br[27] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_30 
+ bl[28] br[28] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_31 
+ bl[29] br[29] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_32 
+ bl[30] br[30] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_33 
+ bl[31] br[31] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_34 
+ bl[32] br[32] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_35 
+ bl[33] br[33] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_36 
+ bl[34] br[34] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_37 
+ bl[35] br[35] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_38 
+ bl[36] br[36] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_39 
+ bl[37] br[37] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_40 
+ bl[38] br[38] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_41 
+ bl[39] br[39] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_42 
+ bl[40] br[40] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_43 
+ bl[41] br[41] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_44 
+ bl[42] br[42] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_45 
+ bl[43] br[43] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_46 
+ bl[44] br[44] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_47 
+ bl[45] br[45] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_48 
+ bl[46] br[46] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_49 
+ bl[47] br[47] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_50 
+ bl[48] br[48] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_51 
+ bl[49] br[49] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_52 
+ bl[50] br[50] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_53 
+ bl[51] br[51] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_54 
+ bl[52] br[52] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_55 
+ bl[53] br[53] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_56 
+ bl[54] br[54] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_57 
+ bl[55] br[55] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_58 
+ bl[56] br[56] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_59 
+ bl[57] br[57] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_60 
+ bl[58] br[58] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_61 
+ bl[59] br[59] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_62 
+ bl[60] br[60] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_63 
+ bl[61] br[61] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_64 
+ bl[62] br[62] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_65 
+ bl[63] br[63] vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_66 
+ vdd vdd vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_59_67 
+ vdd vdd vdd vss wl[57] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_0 
+ vdd vdd vss vdd vpb vnb wl[58] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_60_1 
+ rbl rbr vss vdd vpb vnb wl[58] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_60_2 
+ bl[0] br[0] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_3 
+ bl[1] br[1] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_4 
+ bl[2] br[2] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_5 
+ bl[3] br[3] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_6 
+ bl[4] br[4] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_7 
+ bl[5] br[5] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_8 
+ bl[6] br[6] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_9 
+ bl[7] br[7] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_10 
+ bl[8] br[8] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_11 
+ bl[9] br[9] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_12 
+ bl[10] br[10] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_13 
+ bl[11] br[11] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_14 
+ bl[12] br[12] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_15 
+ bl[13] br[13] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_16 
+ bl[14] br[14] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_17 
+ bl[15] br[15] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_18 
+ bl[16] br[16] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_19 
+ bl[17] br[17] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_20 
+ bl[18] br[18] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_21 
+ bl[19] br[19] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_22 
+ bl[20] br[20] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_23 
+ bl[21] br[21] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_24 
+ bl[22] br[22] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_25 
+ bl[23] br[23] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_26 
+ bl[24] br[24] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_27 
+ bl[25] br[25] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_28 
+ bl[26] br[26] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_29 
+ bl[27] br[27] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_30 
+ bl[28] br[28] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_31 
+ bl[29] br[29] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_32 
+ bl[30] br[30] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_33 
+ bl[31] br[31] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_34 
+ bl[32] br[32] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_35 
+ bl[33] br[33] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_36 
+ bl[34] br[34] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_37 
+ bl[35] br[35] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_38 
+ bl[36] br[36] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_39 
+ bl[37] br[37] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_40 
+ bl[38] br[38] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_41 
+ bl[39] br[39] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_42 
+ bl[40] br[40] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_43 
+ bl[41] br[41] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_44 
+ bl[42] br[42] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_45 
+ bl[43] br[43] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_46 
+ bl[44] br[44] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_47 
+ bl[45] br[45] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_48 
+ bl[46] br[46] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_49 
+ bl[47] br[47] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_50 
+ bl[48] br[48] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_51 
+ bl[49] br[49] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_52 
+ bl[50] br[50] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_53 
+ bl[51] br[51] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_54 
+ bl[52] br[52] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_55 
+ bl[53] br[53] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_56 
+ bl[54] br[54] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_57 
+ bl[55] br[55] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_58 
+ bl[56] br[56] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_59 
+ bl[57] br[57] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_60 
+ bl[58] br[58] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_61 
+ bl[59] br[59] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_62 
+ bl[60] br[60] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_63 
+ bl[61] br[61] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_64 
+ bl[62] br[62] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_65 
+ bl[63] br[63] vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_66 
+ vdd vdd vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_60_67 
+ vdd vdd vdd vss wl[58] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_0 
+ vdd vdd vss vdd vpb vnb wl[59] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_61_1 
+ rbl rbr vss vdd vpb vnb wl[59] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_61_2 
+ bl[0] br[0] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_3 
+ bl[1] br[1] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_4 
+ bl[2] br[2] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_5 
+ bl[3] br[3] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_6 
+ bl[4] br[4] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_7 
+ bl[5] br[5] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_8 
+ bl[6] br[6] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_9 
+ bl[7] br[7] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_10 
+ bl[8] br[8] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_11 
+ bl[9] br[9] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_12 
+ bl[10] br[10] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_13 
+ bl[11] br[11] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_14 
+ bl[12] br[12] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_15 
+ bl[13] br[13] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_16 
+ bl[14] br[14] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_17 
+ bl[15] br[15] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_18 
+ bl[16] br[16] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_19 
+ bl[17] br[17] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_20 
+ bl[18] br[18] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_21 
+ bl[19] br[19] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_22 
+ bl[20] br[20] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_23 
+ bl[21] br[21] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_24 
+ bl[22] br[22] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_25 
+ bl[23] br[23] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_26 
+ bl[24] br[24] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_27 
+ bl[25] br[25] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_28 
+ bl[26] br[26] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_29 
+ bl[27] br[27] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_30 
+ bl[28] br[28] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_31 
+ bl[29] br[29] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_32 
+ bl[30] br[30] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_33 
+ bl[31] br[31] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_34 
+ bl[32] br[32] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_35 
+ bl[33] br[33] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_36 
+ bl[34] br[34] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_37 
+ bl[35] br[35] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_38 
+ bl[36] br[36] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_39 
+ bl[37] br[37] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_40 
+ bl[38] br[38] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_41 
+ bl[39] br[39] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_42 
+ bl[40] br[40] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_43 
+ bl[41] br[41] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_44 
+ bl[42] br[42] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_45 
+ bl[43] br[43] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_46 
+ bl[44] br[44] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_47 
+ bl[45] br[45] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_48 
+ bl[46] br[46] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_49 
+ bl[47] br[47] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_50 
+ bl[48] br[48] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_51 
+ bl[49] br[49] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_52 
+ bl[50] br[50] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_53 
+ bl[51] br[51] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_54 
+ bl[52] br[52] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_55 
+ bl[53] br[53] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_56 
+ bl[54] br[54] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_57 
+ bl[55] br[55] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_58 
+ bl[56] br[56] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_59 
+ bl[57] br[57] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_60 
+ bl[58] br[58] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_61 
+ bl[59] br[59] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_62 
+ bl[60] br[60] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_63 
+ bl[61] br[61] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_64 
+ bl[62] br[62] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_65 
+ bl[63] br[63] vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_66 
+ vdd vdd vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_61_67 
+ vdd vdd vdd vss wl[59] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_0 
+ vdd vdd vss vdd vpb vnb wl[60] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_62_1 
+ rbl rbr vss vdd vpb vnb wl[60] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_62_2 
+ bl[0] br[0] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_3 
+ bl[1] br[1] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_4 
+ bl[2] br[2] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_5 
+ bl[3] br[3] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_6 
+ bl[4] br[4] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_7 
+ bl[5] br[5] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_8 
+ bl[6] br[6] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_9 
+ bl[7] br[7] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_10 
+ bl[8] br[8] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_11 
+ bl[9] br[9] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_12 
+ bl[10] br[10] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_13 
+ bl[11] br[11] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_14 
+ bl[12] br[12] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_15 
+ bl[13] br[13] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_16 
+ bl[14] br[14] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_17 
+ bl[15] br[15] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_18 
+ bl[16] br[16] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_19 
+ bl[17] br[17] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_20 
+ bl[18] br[18] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_21 
+ bl[19] br[19] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_22 
+ bl[20] br[20] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_23 
+ bl[21] br[21] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_24 
+ bl[22] br[22] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_25 
+ bl[23] br[23] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_26 
+ bl[24] br[24] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_27 
+ bl[25] br[25] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_28 
+ bl[26] br[26] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_29 
+ bl[27] br[27] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_30 
+ bl[28] br[28] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_31 
+ bl[29] br[29] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_32 
+ bl[30] br[30] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_33 
+ bl[31] br[31] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_34 
+ bl[32] br[32] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_35 
+ bl[33] br[33] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_36 
+ bl[34] br[34] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_37 
+ bl[35] br[35] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_38 
+ bl[36] br[36] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_39 
+ bl[37] br[37] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_40 
+ bl[38] br[38] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_41 
+ bl[39] br[39] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_42 
+ bl[40] br[40] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_43 
+ bl[41] br[41] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_44 
+ bl[42] br[42] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_45 
+ bl[43] br[43] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_46 
+ bl[44] br[44] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_47 
+ bl[45] br[45] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_48 
+ bl[46] br[46] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_49 
+ bl[47] br[47] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_50 
+ bl[48] br[48] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_51 
+ bl[49] br[49] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_52 
+ bl[50] br[50] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_53 
+ bl[51] br[51] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_54 
+ bl[52] br[52] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_55 
+ bl[53] br[53] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_56 
+ bl[54] br[54] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_57 
+ bl[55] br[55] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_58 
+ bl[56] br[56] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_59 
+ bl[57] br[57] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_60 
+ bl[58] br[58] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_61 
+ bl[59] br[59] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_62 
+ bl[60] br[60] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_63 
+ bl[61] br[61] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_64 
+ bl[62] br[62] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_65 
+ bl[63] br[63] vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_66 
+ vdd vdd vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_62_67 
+ vdd vdd vdd vss wl[60] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_0 
+ vdd vdd vss vdd vpb vnb wl[61] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_63_1 
+ rbl rbr vss vdd vpb vnb wl[61] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_63_2 
+ bl[0] br[0] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_3 
+ bl[1] br[1] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_4 
+ bl[2] br[2] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_5 
+ bl[3] br[3] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_6 
+ bl[4] br[4] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_7 
+ bl[5] br[5] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_8 
+ bl[6] br[6] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_9 
+ bl[7] br[7] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_10 
+ bl[8] br[8] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_11 
+ bl[9] br[9] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_12 
+ bl[10] br[10] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_13 
+ bl[11] br[11] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_14 
+ bl[12] br[12] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_15 
+ bl[13] br[13] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_16 
+ bl[14] br[14] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_17 
+ bl[15] br[15] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_18 
+ bl[16] br[16] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_19 
+ bl[17] br[17] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_20 
+ bl[18] br[18] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_21 
+ bl[19] br[19] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_22 
+ bl[20] br[20] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_23 
+ bl[21] br[21] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_24 
+ bl[22] br[22] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_25 
+ bl[23] br[23] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_26 
+ bl[24] br[24] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_27 
+ bl[25] br[25] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_28 
+ bl[26] br[26] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_29 
+ bl[27] br[27] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_30 
+ bl[28] br[28] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_31 
+ bl[29] br[29] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_32 
+ bl[30] br[30] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_33 
+ bl[31] br[31] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_34 
+ bl[32] br[32] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_35 
+ bl[33] br[33] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_36 
+ bl[34] br[34] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_37 
+ bl[35] br[35] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_38 
+ bl[36] br[36] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_39 
+ bl[37] br[37] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_40 
+ bl[38] br[38] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_41 
+ bl[39] br[39] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_42 
+ bl[40] br[40] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_43 
+ bl[41] br[41] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_44 
+ bl[42] br[42] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_45 
+ bl[43] br[43] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_46 
+ bl[44] br[44] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_47 
+ bl[45] br[45] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_48 
+ bl[46] br[46] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_49 
+ bl[47] br[47] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_50 
+ bl[48] br[48] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_51 
+ bl[49] br[49] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_52 
+ bl[50] br[50] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_53 
+ bl[51] br[51] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_54 
+ bl[52] br[52] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_55 
+ bl[53] br[53] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_56 
+ bl[54] br[54] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_57 
+ bl[55] br[55] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_58 
+ bl[56] br[56] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_59 
+ bl[57] br[57] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_60 
+ bl[58] br[58] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_61 
+ bl[59] br[59] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_62 
+ bl[60] br[60] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_63 
+ bl[61] br[61] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_64 
+ bl[62] br[62] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_65 
+ bl[63] br[63] vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_66 
+ vdd vdd vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_63_67 
+ vdd vdd vdd vss wl[61] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_0 
+ vdd vdd vss vdd vpb vnb wl[62] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_64_1 
+ rbl rbr vss vdd vpb vnb wl[62] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_64_2 
+ bl[0] br[0] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_3 
+ bl[1] br[1] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_4 
+ bl[2] br[2] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_5 
+ bl[3] br[3] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_6 
+ bl[4] br[4] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_7 
+ bl[5] br[5] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_8 
+ bl[6] br[6] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_9 
+ bl[7] br[7] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_10 
+ bl[8] br[8] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_11 
+ bl[9] br[9] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_12 
+ bl[10] br[10] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_13 
+ bl[11] br[11] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_14 
+ bl[12] br[12] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_15 
+ bl[13] br[13] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_16 
+ bl[14] br[14] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_17 
+ bl[15] br[15] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_18 
+ bl[16] br[16] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_19 
+ bl[17] br[17] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_20 
+ bl[18] br[18] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_21 
+ bl[19] br[19] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_22 
+ bl[20] br[20] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_23 
+ bl[21] br[21] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_24 
+ bl[22] br[22] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_25 
+ bl[23] br[23] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_26 
+ bl[24] br[24] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_27 
+ bl[25] br[25] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_28 
+ bl[26] br[26] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_29 
+ bl[27] br[27] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_30 
+ bl[28] br[28] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_31 
+ bl[29] br[29] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_32 
+ bl[30] br[30] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_33 
+ bl[31] br[31] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_34 
+ bl[32] br[32] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_35 
+ bl[33] br[33] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_36 
+ bl[34] br[34] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_37 
+ bl[35] br[35] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_38 
+ bl[36] br[36] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_39 
+ bl[37] br[37] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_40 
+ bl[38] br[38] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_41 
+ bl[39] br[39] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_42 
+ bl[40] br[40] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_43 
+ bl[41] br[41] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_44 
+ bl[42] br[42] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_45 
+ bl[43] br[43] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_46 
+ bl[44] br[44] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_47 
+ bl[45] br[45] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_48 
+ bl[46] br[46] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_49 
+ bl[47] br[47] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_50 
+ bl[48] br[48] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_51 
+ bl[49] br[49] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_52 
+ bl[50] br[50] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_53 
+ bl[51] br[51] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_54 
+ bl[52] br[52] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_55 
+ bl[53] br[53] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_56 
+ bl[54] br[54] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_57 
+ bl[55] br[55] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_58 
+ bl[56] br[56] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_59 
+ bl[57] br[57] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_60 
+ bl[58] br[58] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_61 
+ bl[59] br[59] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_62 
+ bl[60] br[60] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_63 
+ bl[61] br[61] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_64 
+ bl[62] br[62] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_65 
+ bl[63] br[63] vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_66 
+ vdd vdd vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_64_67 
+ vdd vdd vdd vss wl[62] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_0 
+ vdd vdd vss vdd vpb vnb wl[63] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_65_1 
+ rbl rbr vss vdd vpb vnb wl[63] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_65_2 
+ bl[0] br[0] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_3 
+ bl[1] br[1] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_4 
+ bl[2] br[2] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_5 
+ bl[3] br[3] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_6 
+ bl[4] br[4] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_7 
+ bl[5] br[5] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_8 
+ bl[6] br[6] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_9 
+ bl[7] br[7] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_10 
+ bl[8] br[8] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_11 
+ bl[9] br[9] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_12 
+ bl[10] br[10] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_13 
+ bl[11] br[11] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_14 
+ bl[12] br[12] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_15 
+ bl[13] br[13] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_16 
+ bl[14] br[14] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_17 
+ bl[15] br[15] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_18 
+ bl[16] br[16] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_19 
+ bl[17] br[17] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_20 
+ bl[18] br[18] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_21 
+ bl[19] br[19] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_22 
+ bl[20] br[20] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_23 
+ bl[21] br[21] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_24 
+ bl[22] br[22] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_25 
+ bl[23] br[23] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_26 
+ bl[24] br[24] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_27 
+ bl[25] br[25] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_28 
+ bl[26] br[26] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_29 
+ bl[27] br[27] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_30 
+ bl[28] br[28] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_31 
+ bl[29] br[29] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_32 
+ bl[30] br[30] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_33 
+ bl[31] br[31] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_34 
+ bl[32] br[32] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_35 
+ bl[33] br[33] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_36 
+ bl[34] br[34] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_37 
+ bl[35] br[35] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_38 
+ bl[36] br[36] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_39 
+ bl[37] br[37] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_40 
+ bl[38] br[38] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_41 
+ bl[39] br[39] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_42 
+ bl[40] br[40] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_43 
+ bl[41] br[41] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_44 
+ bl[42] br[42] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_45 
+ bl[43] br[43] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_46 
+ bl[44] br[44] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_47 
+ bl[45] br[45] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_48 
+ bl[46] br[46] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_49 
+ bl[47] br[47] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_50 
+ bl[48] br[48] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_51 
+ bl[49] br[49] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_52 
+ bl[50] br[50] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_53 
+ bl[51] br[51] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_54 
+ bl[52] br[52] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_55 
+ bl[53] br[53] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_56 
+ bl[54] br[54] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_57 
+ bl[55] br[55] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_58 
+ bl[56] br[56] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_59 
+ bl[57] br[57] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_60 
+ bl[58] br[58] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_61 
+ bl[59] br[59] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_62 
+ bl[60] br[60] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_63 
+ bl[61] br[61] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_64 
+ bl[62] br[62] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_65 
+ bl[63] br[63] vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_66 
+ vdd vdd vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_65_67 
+ vdd vdd vdd vss wl[63] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_0 
+ vdd vdd vss vdd vpb vnb wl[64] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_66_1 
+ rbl rbr vss vdd vpb vnb wl[64] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_66_2 
+ bl[0] br[0] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_3 
+ bl[1] br[1] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_4 
+ bl[2] br[2] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_5 
+ bl[3] br[3] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_6 
+ bl[4] br[4] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_7 
+ bl[5] br[5] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_8 
+ bl[6] br[6] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_9 
+ bl[7] br[7] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_10 
+ bl[8] br[8] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_11 
+ bl[9] br[9] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_12 
+ bl[10] br[10] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_13 
+ bl[11] br[11] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_14 
+ bl[12] br[12] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_15 
+ bl[13] br[13] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_16 
+ bl[14] br[14] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_17 
+ bl[15] br[15] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_18 
+ bl[16] br[16] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_19 
+ bl[17] br[17] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_20 
+ bl[18] br[18] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_21 
+ bl[19] br[19] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_22 
+ bl[20] br[20] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_23 
+ bl[21] br[21] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_24 
+ bl[22] br[22] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_25 
+ bl[23] br[23] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_26 
+ bl[24] br[24] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_27 
+ bl[25] br[25] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_28 
+ bl[26] br[26] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_29 
+ bl[27] br[27] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_30 
+ bl[28] br[28] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_31 
+ bl[29] br[29] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_32 
+ bl[30] br[30] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_33 
+ bl[31] br[31] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_34 
+ bl[32] br[32] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_35 
+ bl[33] br[33] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_36 
+ bl[34] br[34] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_37 
+ bl[35] br[35] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_38 
+ bl[36] br[36] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_39 
+ bl[37] br[37] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_40 
+ bl[38] br[38] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_41 
+ bl[39] br[39] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_42 
+ bl[40] br[40] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_43 
+ bl[41] br[41] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_44 
+ bl[42] br[42] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_45 
+ bl[43] br[43] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_46 
+ bl[44] br[44] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_47 
+ bl[45] br[45] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_48 
+ bl[46] br[46] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_49 
+ bl[47] br[47] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_50 
+ bl[48] br[48] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_51 
+ bl[49] br[49] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_52 
+ bl[50] br[50] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_53 
+ bl[51] br[51] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_54 
+ bl[52] br[52] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_55 
+ bl[53] br[53] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_56 
+ bl[54] br[54] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_57 
+ bl[55] br[55] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_58 
+ bl[56] br[56] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_59 
+ bl[57] br[57] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_60 
+ bl[58] br[58] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_61 
+ bl[59] br[59] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_62 
+ bl[60] br[60] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_63 
+ bl[61] br[61] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_64 
+ bl[62] br[62] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_65 
+ bl[63] br[63] vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_66 
+ vdd vdd vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_66_67 
+ vdd vdd vdd vss wl[64] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_0 
+ vdd vdd vss vdd vpb vnb wl[65] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_67_1 
+ rbl rbr vss vdd vpb vnb wl[65] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_67_2 
+ bl[0] br[0] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_3 
+ bl[1] br[1] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_4 
+ bl[2] br[2] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_5 
+ bl[3] br[3] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_6 
+ bl[4] br[4] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_7 
+ bl[5] br[5] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_8 
+ bl[6] br[6] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_9 
+ bl[7] br[7] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_10 
+ bl[8] br[8] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_11 
+ bl[9] br[9] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_12 
+ bl[10] br[10] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_13 
+ bl[11] br[11] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_14 
+ bl[12] br[12] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_15 
+ bl[13] br[13] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_16 
+ bl[14] br[14] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_17 
+ bl[15] br[15] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_18 
+ bl[16] br[16] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_19 
+ bl[17] br[17] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_20 
+ bl[18] br[18] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_21 
+ bl[19] br[19] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_22 
+ bl[20] br[20] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_23 
+ bl[21] br[21] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_24 
+ bl[22] br[22] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_25 
+ bl[23] br[23] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_26 
+ bl[24] br[24] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_27 
+ bl[25] br[25] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_28 
+ bl[26] br[26] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_29 
+ bl[27] br[27] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_30 
+ bl[28] br[28] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_31 
+ bl[29] br[29] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_32 
+ bl[30] br[30] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_33 
+ bl[31] br[31] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_34 
+ bl[32] br[32] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_35 
+ bl[33] br[33] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_36 
+ bl[34] br[34] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_37 
+ bl[35] br[35] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_38 
+ bl[36] br[36] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_39 
+ bl[37] br[37] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_40 
+ bl[38] br[38] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_41 
+ bl[39] br[39] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_42 
+ bl[40] br[40] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_43 
+ bl[41] br[41] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_44 
+ bl[42] br[42] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_45 
+ bl[43] br[43] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_46 
+ bl[44] br[44] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_47 
+ bl[45] br[45] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_48 
+ bl[46] br[46] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_49 
+ bl[47] br[47] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_50 
+ bl[48] br[48] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_51 
+ bl[49] br[49] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_52 
+ bl[50] br[50] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_53 
+ bl[51] br[51] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_54 
+ bl[52] br[52] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_55 
+ bl[53] br[53] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_56 
+ bl[54] br[54] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_57 
+ bl[55] br[55] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_58 
+ bl[56] br[56] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_59 
+ bl[57] br[57] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_60 
+ bl[58] br[58] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_61 
+ bl[59] br[59] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_62 
+ bl[60] br[60] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_63 
+ bl[61] br[61] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_64 
+ bl[62] br[62] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_65 
+ bl[63] br[63] vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_66 
+ vdd vdd vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_67_67 
+ vdd vdd vdd vss wl[65] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_0 
+ vdd vdd vss vdd vpb vnb wl[66] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_68_1 
+ rbl rbr vss vdd vpb vnb wl[66] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_68_2 
+ bl[0] br[0] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_3 
+ bl[1] br[1] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_4 
+ bl[2] br[2] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_5 
+ bl[3] br[3] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_6 
+ bl[4] br[4] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_7 
+ bl[5] br[5] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_8 
+ bl[6] br[6] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_9 
+ bl[7] br[7] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_10 
+ bl[8] br[8] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_11 
+ bl[9] br[9] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_12 
+ bl[10] br[10] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_13 
+ bl[11] br[11] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_14 
+ bl[12] br[12] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_15 
+ bl[13] br[13] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_16 
+ bl[14] br[14] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_17 
+ bl[15] br[15] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_18 
+ bl[16] br[16] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_19 
+ bl[17] br[17] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_20 
+ bl[18] br[18] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_21 
+ bl[19] br[19] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_22 
+ bl[20] br[20] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_23 
+ bl[21] br[21] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_24 
+ bl[22] br[22] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_25 
+ bl[23] br[23] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_26 
+ bl[24] br[24] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_27 
+ bl[25] br[25] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_28 
+ bl[26] br[26] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_29 
+ bl[27] br[27] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_30 
+ bl[28] br[28] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_31 
+ bl[29] br[29] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_32 
+ bl[30] br[30] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_33 
+ bl[31] br[31] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_34 
+ bl[32] br[32] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_35 
+ bl[33] br[33] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_36 
+ bl[34] br[34] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_37 
+ bl[35] br[35] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_38 
+ bl[36] br[36] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_39 
+ bl[37] br[37] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_40 
+ bl[38] br[38] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_41 
+ bl[39] br[39] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_42 
+ bl[40] br[40] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_43 
+ bl[41] br[41] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_44 
+ bl[42] br[42] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_45 
+ bl[43] br[43] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_46 
+ bl[44] br[44] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_47 
+ bl[45] br[45] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_48 
+ bl[46] br[46] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_49 
+ bl[47] br[47] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_50 
+ bl[48] br[48] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_51 
+ bl[49] br[49] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_52 
+ bl[50] br[50] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_53 
+ bl[51] br[51] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_54 
+ bl[52] br[52] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_55 
+ bl[53] br[53] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_56 
+ bl[54] br[54] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_57 
+ bl[55] br[55] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_58 
+ bl[56] br[56] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_59 
+ bl[57] br[57] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_60 
+ bl[58] br[58] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_61 
+ bl[59] br[59] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_62 
+ bl[60] br[60] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_63 
+ bl[61] br[61] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_64 
+ bl[62] br[62] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_65 
+ bl[63] br[63] vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_66 
+ vdd vdd vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_68_67 
+ vdd vdd vdd vss wl[66] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_0 
+ vdd vdd vss vdd vpb vnb wl[67] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_69_1 
+ rbl rbr vss vdd vpb vnb wl[67] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_69_2 
+ bl[0] br[0] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_3 
+ bl[1] br[1] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_4 
+ bl[2] br[2] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_5 
+ bl[3] br[3] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_6 
+ bl[4] br[4] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_7 
+ bl[5] br[5] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_8 
+ bl[6] br[6] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_9 
+ bl[7] br[7] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_10 
+ bl[8] br[8] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_11 
+ bl[9] br[9] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_12 
+ bl[10] br[10] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_13 
+ bl[11] br[11] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_14 
+ bl[12] br[12] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_15 
+ bl[13] br[13] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_16 
+ bl[14] br[14] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_17 
+ bl[15] br[15] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_18 
+ bl[16] br[16] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_19 
+ bl[17] br[17] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_20 
+ bl[18] br[18] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_21 
+ bl[19] br[19] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_22 
+ bl[20] br[20] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_23 
+ bl[21] br[21] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_24 
+ bl[22] br[22] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_25 
+ bl[23] br[23] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_26 
+ bl[24] br[24] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_27 
+ bl[25] br[25] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_28 
+ bl[26] br[26] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_29 
+ bl[27] br[27] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_30 
+ bl[28] br[28] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_31 
+ bl[29] br[29] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_32 
+ bl[30] br[30] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_33 
+ bl[31] br[31] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_34 
+ bl[32] br[32] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_35 
+ bl[33] br[33] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_36 
+ bl[34] br[34] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_37 
+ bl[35] br[35] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_38 
+ bl[36] br[36] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_39 
+ bl[37] br[37] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_40 
+ bl[38] br[38] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_41 
+ bl[39] br[39] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_42 
+ bl[40] br[40] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_43 
+ bl[41] br[41] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_44 
+ bl[42] br[42] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_45 
+ bl[43] br[43] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_46 
+ bl[44] br[44] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_47 
+ bl[45] br[45] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_48 
+ bl[46] br[46] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_49 
+ bl[47] br[47] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_50 
+ bl[48] br[48] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_51 
+ bl[49] br[49] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_52 
+ bl[50] br[50] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_53 
+ bl[51] br[51] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_54 
+ bl[52] br[52] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_55 
+ bl[53] br[53] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_56 
+ bl[54] br[54] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_57 
+ bl[55] br[55] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_58 
+ bl[56] br[56] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_59 
+ bl[57] br[57] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_60 
+ bl[58] br[58] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_61 
+ bl[59] br[59] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_62 
+ bl[60] br[60] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_63 
+ bl[61] br[61] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_64 
+ bl[62] br[62] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_65 
+ bl[63] br[63] vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_66 
+ vdd vdd vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_69_67 
+ vdd vdd vdd vss wl[67] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_0 
+ vdd vdd vss vdd vpb vnb wl[68] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_70_1 
+ rbl rbr vss vdd vpb vnb wl[68] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_70_2 
+ bl[0] br[0] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_3 
+ bl[1] br[1] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_4 
+ bl[2] br[2] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_5 
+ bl[3] br[3] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_6 
+ bl[4] br[4] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_7 
+ bl[5] br[5] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_8 
+ bl[6] br[6] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_9 
+ bl[7] br[7] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_10 
+ bl[8] br[8] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_11 
+ bl[9] br[9] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_12 
+ bl[10] br[10] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_13 
+ bl[11] br[11] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_14 
+ bl[12] br[12] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_15 
+ bl[13] br[13] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_16 
+ bl[14] br[14] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_17 
+ bl[15] br[15] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_18 
+ bl[16] br[16] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_19 
+ bl[17] br[17] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_20 
+ bl[18] br[18] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_21 
+ bl[19] br[19] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_22 
+ bl[20] br[20] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_23 
+ bl[21] br[21] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_24 
+ bl[22] br[22] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_25 
+ bl[23] br[23] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_26 
+ bl[24] br[24] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_27 
+ bl[25] br[25] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_28 
+ bl[26] br[26] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_29 
+ bl[27] br[27] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_30 
+ bl[28] br[28] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_31 
+ bl[29] br[29] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_32 
+ bl[30] br[30] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_33 
+ bl[31] br[31] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_34 
+ bl[32] br[32] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_35 
+ bl[33] br[33] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_36 
+ bl[34] br[34] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_37 
+ bl[35] br[35] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_38 
+ bl[36] br[36] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_39 
+ bl[37] br[37] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_40 
+ bl[38] br[38] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_41 
+ bl[39] br[39] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_42 
+ bl[40] br[40] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_43 
+ bl[41] br[41] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_44 
+ bl[42] br[42] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_45 
+ bl[43] br[43] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_46 
+ bl[44] br[44] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_47 
+ bl[45] br[45] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_48 
+ bl[46] br[46] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_49 
+ bl[47] br[47] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_50 
+ bl[48] br[48] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_51 
+ bl[49] br[49] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_52 
+ bl[50] br[50] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_53 
+ bl[51] br[51] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_54 
+ bl[52] br[52] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_55 
+ bl[53] br[53] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_56 
+ bl[54] br[54] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_57 
+ bl[55] br[55] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_58 
+ bl[56] br[56] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_59 
+ bl[57] br[57] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_60 
+ bl[58] br[58] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_61 
+ bl[59] br[59] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_62 
+ bl[60] br[60] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_63 
+ bl[61] br[61] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_64 
+ bl[62] br[62] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_65 
+ bl[63] br[63] vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_66 
+ vdd vdd vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_70_67 
+ vdd vdd vdd vss wl[68] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_0 
+ vdd vdd vss vdd vpb vnb wl[69] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_71_1 
+ rbl rbr vss vdd vpb vnb wl[69] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_71_2 
+ bl[0] br[0] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_3 
+ bl[1] br[1] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_4 
+ bl[2] br[2] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_5 
+ bl[3] br[3] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_6 
+ bl[4] br[4] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_7 
+ bl[5] br[5] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_8 
+ bl[6] br[6] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_9 
+ bl[7] br[7] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_10 
+ bl[8] br[8] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_11 
+ bl[9] br[9] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_12 
+ bl[10] br[10] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_13 
+ bl[11] br[11] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_14 
+ bl[12] br[12] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_15 
+ bl[13] br[13] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_16 
+ bl[14] br[14] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_17 
+ bl[15] br[15] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_18 
+ bl[16] br[16] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_19 
+ bl[17] br[17] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_20 
+ bl[18] br[18] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_21 
+ bl[19] br[19] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_22 
+ bl[20] br[20] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_23 
+ bl[21] br[21] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_24 
+ bl[22] br[22] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_25 
+ bl[23] br[23] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_26 
+ bl[24] br[24] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_27 
+ bl[25] br[25] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_28 
+ bl[26] br[26] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_29 
+ bl[27] br[27] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_30 
+ bl[28] br[28] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_31 
+ bl[29] br[29] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_32 
+ bl[30] br[30] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_33 
+ bl[31] br[31] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_34 
+ bl[32] br[32] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_35 
+ bl[33] br[33] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_36 
+ bl[34] br[34] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_37 
+ bl[35] br[35] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_38 
+ bl[36] br[36] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_39 
+ bl[37] br[37] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_40 
+ bl[38] br[38] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_41 
+ bl[39] br[39] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_42 
+ bl[40] br[40] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_43 
+ bl[41] br[41] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_44 
+ bl[42] br[42] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_45 
+ bl[43] br[43] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_46 
+ bl[44] br[44] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_47 
+ bl[45] br[45] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_48 
+ bl[46] br[46] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_49 
+ bl[47] br[47] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_50 
+ bl[48] br[48] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_51 
+ bl[49] br[49] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_52 
+ bl[50] br[50] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_53 
+ bl[51] br[51] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_54 
+ bl[52] br[52] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_55 
+ bl[53] br[53] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_56 
+ bl[54] br[54] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_57 
+ bl[55] br[55] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_58 
+ bl[56] br[56] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_59 
+ bl[57] br[57] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_60 
+ bl[58] br[58] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_61 
+ bl[59] br[59] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_62 
+ bl[60] br[60] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_63 
+ bl[61] br[61] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_64 
+ bl[62] br[62] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_65 
+ bl[63] br[63] vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_66 
+ vdd vdd vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_71_67 
+ vdd vdd vdd vss wl[69] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_0 
+ vdd vdd vss vdd vpb vnb wl[70] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_72_1 
+ rbl rbr vss vdd vpb vnb wl[70] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_72_2 
+ bl[0] br[0] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_3 
+ bl[1] br[1] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_4 
+ bl[2] br[2] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_5 
+ bl[3] br[3] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_6 
+ bl[4] br[4] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_7 
+ bl[5] br[5] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_8 
+ bl[6] br[6] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_9 
+ bl[7] br[7] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_10 
+ bl[8] br[8] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_11 
+ bl[9] br[9] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_12 
+ bl[10] br[10] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_13 
+ bl[11] br[11] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_14 
+ bl[12] br[12] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_15 
+ bl[13] br[13] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_16 
+ bl[14] br[14] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_17 
+ bl[15] br[15] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_18 
+ bl[16] br[16] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_19 
+ bl[17] br[17] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_20 
+ bl[18] br[18] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_21 
+ bl[19] br[19] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_22 
+ bl[20] br[20] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_23 
+ bl[21] br[21] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_24 
+ bl[22] br[22] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_25 
+ bl[23] br[23] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_26 
+ bl[24] br[24] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_27 
+ bl[25] br[25] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_28 
+ bl[26] br[26] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_29 
+ bl[27] br[27] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_30 
+ bl[28] br[28] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_31 
+ bl[29] br[29] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_32 
+ bl[30] br[30] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_33 
+ bl[31] br[31] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_34 
+ bl[32] br[32] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_35 
+ bl[33] br[33] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_36 
+ bl[34] br[34] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_37 
+ bl[35] br[35] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_38 
+ bl[36] br[36] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_39 
+ bl[37] br[37] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_40 
+ bl[38] br[38] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_41 
+ bl[39] br[39] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_42 
+ bl[40] br[40] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_43 
+ bl[41] br[41] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_44 
+ bl[42] br[42] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_45 
+ bl[43] br[43] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_46 
+ bl[44] br[44] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_47 
+ bl[45] br[45] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_48 
+ bl[46] br[46] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_49 
+ bl[47] br[47] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_50 
+ bl[48] br[48] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_51 
+ bl[49] br[49] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_52 
+ bl[50] br[50] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_53 
+ bl[51] br[51] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_54 
+ bl[52] br[52] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_55 
+ bl[53] br[53] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_56 
+ bl[54] br[54] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_57 
+ bl[55] br[55] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_58 
+ bl[56] br[56] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_59 
+ bl[57] br[57] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_60 
+ bl[58] br[58] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_61 
+ bl[59] br[59] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_62 
+ bl[60] br[60] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_63 
+ bl[61] br[61] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_64 
+ bl[62] br[62] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_65 
+ bl[63] br[63] vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_66 
+ vdd vdd vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_72_67 
+ vdd vdd vdd vss wl[70] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_0 
+ vdd vdd vss vdd vpb vnb wl[71] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_73_1 
+ rbl rbr vss vdd vpb vnb wl[71] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_73_2 
+ bl[0] br[0] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_3 
+ bl[1] br[1] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_4 
+ bl[2] br[2] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_5 
+ bl[3] br[3] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_6 
+ bl[4] br[4] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_7 
+ bl[5] br[5] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_8 
+ bl[6] br[6] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_9 
+ bl[7] br[7] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_10 
+ bl[8] br[8] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_11 
+ bl[9] br[9] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_12 
+ bl[10] br[10] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_13 
+ bl[11] br[11] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_14 
+ bl[12] br[12] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_15 
+ bl[13] br[13] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_16 
+ bl[14] br[14] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_17 
+ bl[15] br[15] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_18 
+ bl[16] br[16] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_19 
+ bl[17] br[17] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_20 
+ bl[18] br[18] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_21 
+ bl[19] br[19] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_22 
+ bl[20] br[20] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_23 
+ bl[21] br[21] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_24 
+ bl[22] br[22] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_25 
+ bl[23] br[23] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_26 
+ bl[24] br[24] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_27 
+ bl[25] br[25] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_28 
+ bl[26] br[26] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_29 
+ bl[27] br[27] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_30 
+ bl[28] br[28] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_31 
+ bl[29] br[29] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_32 
+ bl[30] br[30] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_33 
+ bl[31] br[31] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_34 
+ bl[32] br[32] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_35 
+ bl[33] br[33] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_36 
+ bl[34] br[34] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_37 
+ bl[35] br[35] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_38 
+ bl[36] br[36] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_39 
+ bl[37] br[37] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_40 
+ bl[38] br[38] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_41 
+ bl[39] br[39] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_42 
+ bl[40] br[40] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_43 
+ bl[41] br[41] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_44 
+ bl[42] br[42] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_45 
+ bl[43] br[43] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_46 
+ bl[44] br[44] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_47 
+ bl[45] br[45] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_48 
+ bl[46] br[46] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_49 
+ bl[47] br[47] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_50 
+ bl[48] br[48] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_51 
+ bl[49] br[49] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_52 
+ bl[50] br[50] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_53 
+ bl[51] br[51] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_54 
+ bl[52] br[52] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_55 
+ bl[53] br[53] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_56 
+ bl[54] br[54] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_57 
+ bl[55] br[55] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_58 
+ bl[56] br[56] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_59 
+ bl[57] br[57] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_60 
+ bl[58] br[58] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_61 
+ bl[59] br[59] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_62 
+ bl[60] br[60] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_63 
+ bl[61] br[61] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_64 
+ bl[62] br[62] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_65 
+ bl[63] br[63] vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_66 
+ vdd vdd vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_73_67 
+ vdd vdd vdd vss wl[71] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_0 
+ vdd vdd vss vdd vpb vnb wl[72] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_74_1 
+ rbl rbr vss vdd vpb vnb wl[72] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_74_2 
+ bl[0] br[0] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_3 
+ bl[1] br[1] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_4 
+ bl[2] br[2] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_5 
+ bl[3] br[3] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_6 
+ bl[4] br[4] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_7 
+ bl[5] br[5] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_8 
+ bl[6] br[6] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_9 
+ bl[7] br[7] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_10 
+ bl[8] br[8] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_11 
+ bl[9] br[9] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_12 
+ bl[10] br[10] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_13 
+ bl[11] br[11] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_14 
+ bl[12] br[12] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_15 
+ bl[13] br[13] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_16 
+ bl[14] br[14] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_17 
+ bl[15] br[15] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_18 
+ bl[16] br[16] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_19 
+ bl[17] br[17] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_20 
+ bl[18] br[18] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_21 
+ bl[19] br[19] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_22 
+ bl[20] br[20] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_23 
+ bl[21] br[21] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_24 
+ bl[22] br[22] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_25 
+ bl[23] br[23] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_26 
+ bl[24] br[24] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_27 
+ bl[25] br[25] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_28 
+ bl[26] br[26] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_29 
+ bl[27] br[27] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_30 
+ bl[28] br[28] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_31 
+ bl[29] br[29] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_32 
+ bl[30] br[30] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_33 
+ bl[31] br[31] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_34 
+ bl[32] br[32] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_35 
+ bl[33] br[33] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_36 
+ bl[34] br[34] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_37 
+ bl[35] br[35] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_38 
+ bl[36] br[36] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_39 
+ bl[37] br[37] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_40 
+ bl[38] br[38] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_41 
+ bl[39] br[39] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_42 
+ bl[40] br[40] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_43 
+ bl[41] br[41] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_44 
+ bl[42] br[42] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_45 
+ bl[43] br[43] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_46 
+ bl[44] br[44] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_47 
+ bl[45] br[45] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_48 
+ bl[46] br[46] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_49 
+ bl[47] br[47] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_50 
+ bl[48] br[48] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_51 
+ bl[49] br[49] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_52 
+ bl[50] br[50] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_53 
+ bl[51] br[51] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_54 
+ bl[52] br[52] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_55 
+ bl[53] br[53] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_56 
+ bl[54] br[54] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_57 
+ bl[55] br[55] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_58 
+ bl[56] br[56] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_59 
+ bl[57] br[57] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_60 
+ bl[58] br[58] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_61 
+ bl[59] br[59] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_62 
+ bl[60] br[60] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_63 
+ bl[61] br[61] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_64 
+ bl[62] br[62] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_65 
+ bl[63] br[63] vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_66 
+ vdd vdd vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_74_67 
+ vdd vdd vdd vss wl[72] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_0 
+ vdd vdd vss vdd vpb vnb wl[73] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_75_1 
+ rbl rbr vss vdd vpb vnb wl[73] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_75_2 
+ bl[0] br[0] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_3 
+ bl[1] br[1] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_4 
+ bl[2] br[2] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_5 
+ bl[3] br[3] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_6 
+ bl[4] br[4] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_7 
+ bl[5] br[5] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_8 
+ bl[6] br[6] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_9 
+ bl[7] br[7] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_10 
+ bl[8] br[8] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_11 
+ bl[9] br[9] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_12 
+ bl[10] br[10] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_13 
+ bl[11] br[11] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_14 
+ bl[12] br[12] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_15 
+ bl[13] br[13] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_16 
+ bl[14] br[14] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_17 
+ bl[15] br[15] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_18 
+ bl[16] br[16] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_19 
+ bl[17] br[17] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_20 
+ bl[18] br[18] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_21 
+ bl[19] br[19] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_22 
+ bl[20] br[20] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_23 
+ bl[21] br[21] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_24 
+ bl[22] br[22] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_25 
+ bl[23] br[23] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_26 
+ bl[24] br[24] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_27 
+ bl[25] br[25] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_28 
+ bl[26] br[26] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_29 
+ bl[27] br[27] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_30 
+ bl[28] br[28] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_31 
+ bl[29] br[29] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_32 
+ bl[30] br[30] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_33 
+ bl[31] br[31] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_34 
+ bl[32] br[32] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_35 
+ bl[33] br[33] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_36 
+ bl[34] br[34] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_37 
+ bl[35] br[35] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_38 
+ bl[36] br[36] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_39 
+ bl[37] br[37] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_40 
+ bl[38] br[38] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_41 
+ bl[39] br[39] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_42 
+ bl[40] br[40] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_43 
+ bl[41] br[41] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_44 
+ bl[42] br[42] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_45 
+ bl[43] br[43] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_46 
+ bl[44] br[44] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_47 
+ bl[45] br[45] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_48 
+ bl[46] br[46] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_49 
+ bl[47] br[47] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_50 
+ bl[48] br[48] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_51 
+ bl[49] br[49] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_52 
+ bl[50] br[50] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_53 
+ bl[51] br[51] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_54 
+ bl[52] br[52] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_55 
+ bl[53] br[53] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_56 
+ bl[54] br[54] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_57 
+ bl[55] br[55] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_58 
+ bl[56] br[56] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_59 
+ bl[57] br[57] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_60 
+ bl[58] br[58] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_61 
+ bl[59] br[59] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_62 
+ bl[60] br[60] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_63 
+ bl[61] br[61] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_64 
+ bl[62] br[62] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_65 
+ bl[63] br[63] vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_66 
+ vdd vdd vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_75_67 
+ vdd vdd vdd vss wl[73] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_0 
+ vdd vdd vss vdd vpb vnb wl[74] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_76_1 
+ rbl rbr vss vdd vpb vnb wl[74] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_76_2 
+ bl[0] br[0] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_3 
+ bl[1] br[1] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_4 
+ bl[2] br[2] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_5 
+ bl[3] br[3] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_6 
+ bl[4] br[4] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_7 
+ bl[5] br[5] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_8 
+ bl[6] br[6] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_9 
+ bl[7] br[7] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_10 
+ bl[8] br[8] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_11 
+ bl[9] br[9] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_12 
+ bl[10] br[10] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_13 
+ bl[11] br[11] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_14 
+ bl[12] br[12] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_15 
+ bl[13] br[13] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_16 
+ bl[14] br[14] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_17 
+ bl[15] br[15] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_18 
+ bl[16] br[16] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_19 
+ bl[17] br[17] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_20 
+ bl[18] br[18] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_21 
+ bl[19] br[19] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_22 
+ bl[20] br[20] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_23 
+ bl[21] br[21] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_24 
+ bl[22] br[22] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_25 
+ bl[23] br[23] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_26 
+ bl[24] br[24] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_27 
+ bl[25] br[25] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_28 
+ bl[26] br[26] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_29 
+ bl[27] br[27] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_30 
+ bl[28] br[28] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_31 
+ bl[29] br[29] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_32 
+ bl[30] br[30] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_33 
+ bl[31] br[31] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_34 
+ bl[32] br[32] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_35 
+ bl[33] br[33] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_36 
+ bl[34] br[34] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_37 
+ bl[35] br[35] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_38 
+ bl[36] br[36] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_39 
+ bl[37] br[37] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_40 
+ bl[38] br[38] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_41 
+ bl[39] br[39] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_42 
+ bl[40] br[40] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_43 
+ bl[41] br[41] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_44 
+ bl[42] br[42] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_45 
+ bl[43] br[43] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_46 
+ bl[44] br[44] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_47 
+ bl[45] br[45] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_48 
+ bl[46] br[46] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_49 
+ bl[47] br[47] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_50 
+ bl[48] br[48] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_51 
+ bl[49] br[49] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_52 
+ bl[50] br[50] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_53 
+ bl[51] br[51] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_54 
+ bl[52] br[52] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_55 
+ bl[53] br[53] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_56 
+ bl[54] br[54] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_57 
+ bl[55] br[55] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_58 
+ bl[56] br[56] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_59 
+ bl[57] br[57] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_60 
+ bl[58] br[58] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_61 
+ bl[59] br[59] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_62 
+ bl[60] br[60] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_63 
+ bl[61] br[61] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_64 
+ bl[62] br[62] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_65 
+ bl[63] br[63] vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_66 
+ vdd vdd vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_76_67 
+ vdd vdd vdd vss wl[74] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_0 
+ vdd vdd vss vdd vpb vnb wl[75] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_77_1 
+ rbl rbr vss vdd vpb vnb wl[75] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_77_2 
+ bl[0] br[0] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_3 
+ bl[1] br[1] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_4 
+ bl[2] br[2] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_5 
+ bl[3] br[3] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_6 
+ bl[4] br[4] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_7 
+ bl[5] br[5] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_8 
+ bl[6] br[6] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_9 
+ bl[7] br[7] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_10 
+ bl[8] br[8] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_11 
+ bl[9] br[9] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_12 
+ bl[10] br[10] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_13 
+ bl[11] br[11] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_14 
+ bl[12] br[12] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_15 
+ bl[13] br[13] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_16 
+ bl[14] br[14] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_17 
+ bl[15] br[15] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_18 
+ bl[16] br[16] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_19 
+ bl[17] br[17] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_20 
+ bl[18] br[18] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_21 
+ bl[19] br[19] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_22 
+ bl[20] br[20] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_23 
+ bl[21] br[21] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_24 
+ bl[22] br[22] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_25 
+ bl[23] br[23] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_26 
+ bl[24] br[24] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_27 
+ bl[25] br[25] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_28 
+ bl[26] br[26] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_29 
+ bl[27] br[27] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_30 
+ bl[28] br[28] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_31 
+ bl[29] br[29] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_32 
+ bl[30] br[30] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_33 
+ bl[31] br[31] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_34 
+ bl[32] br[32] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_35 
+ bl[33] br[33] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_36 
+ bl[34] br[34] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_37 
+ bl[35] br[35] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_38 
+ bl[36] br[36] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_39 
+ bl[37] br[37] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_40 
+ bl[38] br[38] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_41 
+ bl[39] br[39] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_42 
+ bl[40] br[40] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_43 
+ bl[41] br[41] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_44 
+ bl[42] br[42] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_45 
+ bl[43] br[43] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_46 
+ bl[44] br[44] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_47 
+ bl[45] br[45] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_48 
+ bl[46] br[46] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_49 
+ bl[47] br[47] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_50 
+ bl[48] br[48] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_51 
+ bl[49] br[49] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_52 
+ bl[50] br[50] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_53 
+ bl[51] br[51] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_54 
+ bl[52] br[52] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_55 
+ bl[53] br[53] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_56 
+ bl[54] br[54] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_57 
+ bl[55] br[55] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_58 
+ bl[56] br[56] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_59 
+ bl[57] br[57] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_60 
+ bl[58] br[58] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_61 
+ bl[59] br[59] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_62 
+ bl[60] br[60] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_63 
+ bl[61] br[61] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_64 
+ bl[62] br[62] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_65 
+ bl[63] br[63] vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_66 
+ vdd vdd vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_77_67 
+ vdd vdd vdd vss wl[75] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_0 
+ vdd vdd vss vdd vpb vnb wl[76] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_78_1 
+ rbl rbr vss vdd vpb vnb wl[76] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_78_2 
+ bl[0] br[0] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_3 
+ bl[1] br[1] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_4 
+ bl[2] br[2] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_5 
+ bl[3] br[3] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_6 
+ bl[4] br[4] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_7 
+ bl[5] br[5] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_8 
+ bl[6] br[6] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_9 
+ bl[7] br[7] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_10 
+ bl[8] br[8] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_11 
+ bl[9] br[9] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_12 
+ bl[10] br[10] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_13 
+ bl[11] br[11] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_14 
+ bl[12] br[12] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_15 
+ bl[13] br[13] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_16 
+ bl[14] br[14] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_17 
+ bl[15] br[15] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_18 
+ bl[16] br[16] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_19 
+ bl[17] br[17] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_20 
+ bl[18] br[18] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_21 
+ bl[19] br[19] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_22 
+ bl[20] br[20] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_23 
+ bl[21] br[21] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_24 
+ bl[22] br[22] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_25 
+ bl[23] br[23] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_26 
+ bl[24] br[24] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_27 
+ bl[25] br[25] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_28 
+ bl[26] br[26] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_29 
+ bl[27] br[27] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_30 
+ bl[28] br[28] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_31 
+ bl[29] br[29] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_32 
+ bl[30] br[30] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_33 
+ bl[31] br[31] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_34 
+ bl[32] br[32] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_35 
+ bl[33] br[33] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_36 
+ bl[34] br[34] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_37 
+ bl[35] br[35] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_38 
+ bl[36] br[36] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_39 
+ bl[37] br[37] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_40 
+ bl[38] br[38] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_41 
+ bl[39] br[39] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_42 
+ bl[40] br[40] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_43 
+ bl[41] br[41] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_44 
+ bl[42] br[42] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_45 
+ bl[43] br[43] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_46 
+ bl[44] br[44] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_47 
+ bl[45] br[45] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_48 
+ bl[46] br[46] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_49 
+ bl[47] br[47] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_50 
+ bl[48] br[48] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_51 
+ bl[49] br[49] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_52 
+ bl[50] br[50] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_53 
+ bl[51] br[51] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_54 
+ bl[52] br[52] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_55 
+ bl[53] br[53] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_56 
+ bl[54] br[54] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_57 
+ bl[55] br[55] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_58 
+ bl[56] br[56] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_59 
+ bl[57] br[57] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_60 
+ bl[58] br[58] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_61 
+ bl[59] br[59] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_62 
+ bl[60] br[60] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_63 
+ bl[61] br[61] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_64 
+ bl[62] br[62] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_65 
+ bl[63] br[63] vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_66 
+ vdd vdd vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_78_67 
+ vdd vdd vdd vss wl[76] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_0 
+ vdd vdd vss vdd vpb vnb wl[77] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_79_1 
+ rbl rbr vss vdd vpb vnb wl[77] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_79_2 
+ bl[0] br[0] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_3 
+ bl[1] br[1] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_4 
+ bl[2] br[2] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_5 
+ bl[3] br[3] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_6 
+ bl[4] br[4] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_7 
+ bl[5] br[5] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_8 
+ bl[6] br[6] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_9 
+ bl[7] br[7] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_10 
+ bl[8] br[8] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_11 
+ bl[9] br[9] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_12 
+ bl[10] br[10] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_13 
+ bl[11] br[11] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_14 
+ bl[12] br[12] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_15 
+ bl[13] br[13] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_16 
+ bl[14] br[14] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_17 
+ bl[15] br[15] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_18 
+ bl[16] br[16] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_19 
+ bl[17] br[17] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_20 
+ bl[18] br[18] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_21 
+ bl[19] br[19] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_22 
+ bl[20] br[20] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_23 
+ bl[21] br[21] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_24 
+ bl[22] br[22] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_25 
+ bl[23] br[23] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_26 
+ bl[24] br[24] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_27 
+ bl[25] br[25] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_28 
+ bl[26] br[26] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_29 
+ bl[27] br[27] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_30 
+ bl[28] br[28] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_31 
+ bl[29] br[29] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_32 
+ bl[30] br[30] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_33 
+ bl[31] br[31] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_34 
+ bl[32] br[32] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_35 
+ bl[33] br[33] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_36 
+ bl[34] br[34] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_37 
+ bl[35] br[35] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_38 
+ bl[36] br[36] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_39 
+ bl[37] br[37] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_40 
+ bl[38] br[38] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_41 
+ bl[39] br[39] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_42 
+ bl[40] br[40] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_43 
+ bl[41] br[41] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_44 
+ bl[42] br[42] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_45 
+ bl[43] br[43] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_46 
+ bl[44] br[44] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_47 
+ bl[45] br[45] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_48 
+ bl[46] br[46] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_49 
+ bl[47] br[47] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_50 
+ bl[48] br[48] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_51 
+ bl[49] br[49] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_52 
+ bl[50] br[50] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_53 
+ bl[51] br[51] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_54 
+ bl[52] br[52] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_55 
+ bl[53] br[53] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_56 
+ bl[54] br[54] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_57 
+ bl[55] br[55] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_58 
+ bl[56] br[56] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_59 
+ bl[57] br[57] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_60 
+ bl[58] br[58] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_61 
+ bl[59] br[59] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_62 
+ bl[60] br[60] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_63 
+ bl[61] br[61] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_64 
+ bl[62] br[62] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_65 
+ bl[63] br[63] vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_66 
+ vdd vdd vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_79_67 
+ vdd vdd vdd vss wl[77] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_0 
+ vdd vdd vss vdd vpb vnb wl[78] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_80_1 
+ rbl rbr vss vdd vpb vnb wl[78] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_80_2 
+ bl[0] br[0] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_3 
+ bl[1] br[1] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_4 
+ bl[2] br[2] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_5 
+ bl[3] br[3] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_6 
+ bl[4] br[4] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_7 
+ bl[5] br[5] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_8 
+ bl[6] br[6] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_9 
+ bl[7] br[7] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_10 
+ bl[8] br[8] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_11 
+ bl[9] br[9] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_12 
+ bl[10] br[10] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_13 
+ bl[11] br[11] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_14 
+ bl[12] br[12] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_15 
+ bl[13] br[13] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_16 
+ bl[14] br[14] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_17 
+ bl[15] br[15] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_18 
+ bl[16] br[16] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_19 
+ bl[17] br[17] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_20 
+ bl[18] br[18] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_21 
+ bl[19] br[19] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_22 
+ bl[20] br[20] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_23 
+ bl[21] br[21] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_24 
+ bl[22] br[22] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_25 
+ bl[23] br[23] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_26 
+ bl[24] br[24] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_27 
+ bl[25] br[25] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_28 
+ bl[26] br[26] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_29 
+ bl[27] br[27] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_30 
+ bl[28] br[28] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_31 
+ bl[29] br[29] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_32 
+ bl[30] br[30] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_33 
+ bl[31] br[31] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_34 
+ bl[32] br[32] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_35 
+ bl[33] br[33] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_36 
+ bl[34] br[34] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_37 
+ bl[35] br[35] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_38 
+ bl[36] br[36] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_39 
+ bl[37] br[37] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_40 
+ bl[38] br[38] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_41 
+ bl[39] br[39] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_42 
+ bl[40] br[40] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_43 
+ bl[41] br[41] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_44 
+ bl[42] br[42] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_45 
+ bl[43] br[43] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_46 
+ bl[44] br[44] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_47 
+ bl[45] br[45] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_48 
+ bl[46] br[46] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_49 
+ bl[47] br[47] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_50 
+ bl[48] br[48] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_51 
+ bl[49] br[49] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_52 
+ bl[50] br[50] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_53 
+ bl[51] br[51] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_54 
+ bl[52] br[52] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_55 
+ bl[53] br[53] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_56 
+ bl[54] br[54] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_57 
+ bl[55] br[55] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_58 
+ bl[56] br[56] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_59 
+ bl[57] br[57] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_60 
+ bl[58] br[58] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_61 
+ bl[59] br[59] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_62 
+ bl[60] br[60] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_63 
+ bl[61] br[61] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_64 
+ bl[62] br[62] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_65 
+ bl[63] br[63] vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_66 
+ vdd vdd vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_80_67 
+ vdd vdd vdd vss wl[78] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_0 
+ vdd vdd vss vdd vpb vnb wl[79] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_81_1 
+ rbl rbr vss vdd vpb vnb wl[79] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_81_2 
+ bl[0] br[0] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_3 
+ bl[1] br[1] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_4 
+ bl[2] br[2] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_5 
+ bl[3] br[3] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_6 
+ bl[4] br[4] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_7 
+ bl[5] br[5] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_8 
+ bl[6] br[6] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_9 
+ bl[7] br[7] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_10 
+ bl[8] br[8] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_11 
+ bl[9] br[9] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_12 
+ bl[10] br[10] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_13 
+ bl[11] br[11] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_14 
+ bl[12] br[12] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_15 
+ bl[13] br[13] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_16 
+ bl[14] br[14] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_17 
+ bl[15] br[15] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_18 
+ bl[16] br[16] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_19 
+ bl[17] br[17] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_20 
+ bl[18] br[18] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_21 
+ bl[19] br[19] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_22 
+ bl[20] br[20] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_23 
+ bl[21] br[21] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_24 
+ bl[22] br[22] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_25 
+ bl[23] br[23] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_26 
+ bl[24] br[24] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_27 
+ bl[25] br[25] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_28 
+ bl[26] br[26] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_29 
+ bl[27] br[27] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_30 
+ bl[28] br[28] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_31 
+ bl[29] br[29] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_32 
+ bl[30] br[30] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_33 
+ bl[31] br[31] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_34 
+ bl[32] br[32] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_35 
+ bl[33] br[33] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_36 
+ bl[34] br[34] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_37 
+ bl[35] br[35] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_38 
+ bl[36] br[36] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_39 
+ bl[37] br[37] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_40 
+ bl[38] br[38] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_41 
+ bl[39] br[39] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_42 
+ bl[40] br[40] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_43 
+ bl[41] br[41] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_44 
+ bl[42] br[42] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_45 
+ bl[43] br[43] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_46 
+ bl[44] br[44] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_47 
+ bl[45] br[45] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_48 
+ bl[46] br[46] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_49 
+ bl[47] br[47] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_50 
+ bl[48] br[48] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_51 
+ bl[49] br[49] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_52 
+ bl[50] br[50] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_53 
+ bl[51] br[51] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_54 
+ bl[52] br[52] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_55 
+ bl[53] br[53] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_56 
+ bl[54] br[54] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_57 
+ bl[55] br[55] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_58 
+ bl[56] br[56] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_59 
+ bl[57] br[57] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_60 
+ bl[58] br[58] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_61 
+ bl[59] br[59] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_62 
+ bl[60] br[60] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_63 
+ bl[61] br[61] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_64 
+ bl[62] br[62] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_65 
+ bl[63] br[63] vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_66 
+ vdd vdd vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_81_67 
+ vdd vdd vdd vss wl[79] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_0 
+ vdd vdd vss vdd vpb vnb wl[80] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_82_1 
+ rbl rbr vss vdd vpb vnb wl[80] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_82_2 
+ bl[0] br[0] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_3 
+ bl[1] br[1] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_4 
+ bl[2] br[2] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_5 
+ bl[3] br[3] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_6 
+ bl[4] br[4] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_7 
+ bl[5] br[5] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_8 
+ bl[6] br[6] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_9 
+ bl[7] br[7] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_10 
+ bl[8] br[8] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_11 
+ bl[9] br[9] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_12 
+ bl[10] br[10] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_13 
+ bl[11] br[11] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_14 
+ bl[12] br[12] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_15 
+ bl[13] br[13] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_16 
+ bl[14] br[14] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_17 
+ bl[15] br[15] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_18 
+ bl[16] br[16] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_19 
+ bl[17] br[17] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_20 
+ bl[18] br[18] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_21 
+ bl[19] br[19] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_22 
+ bl[20] br[20] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_23 
+ bl[21] br[21] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_24 
+ bl[22] br[22] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_25 
+ bl[23] br[23] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_26 
+ bl[24] br[24] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_27 
+ bl[25] br[25] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_28 
+ bl[26] br[26] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_29 
+ bl[27] br[27] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_30 
+ bl[28] br[28] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_31 
+ bl[29] br[29] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_32 
+ bl[30] br[30] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_33 
+ bl[31] br[31] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_34 
+ bl[32] br[32] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_35 
+ bl[33] br[33] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_36 
+ bl[34] br[34] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_37 
+ bl[35] br[35] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_38 
+ bl[36] br[36] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_39 
+ bl[37] br[37] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_40 
+ bl[38] br[38] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_41 
+ bl[39] br[39] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_42 
+ bl[40] br[40] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_43 
+ bl[41] br[41] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_44 
+ bl[42] br[42] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_45 
+ bl[43] br[43] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_46 
+ bl[44] br[44] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_47 
+ bl[45] br[45] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_48 
+ bl[46] br[46] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_49 
+ bl[47] br[47] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_50 
+ bl[48] br[48] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_51 
+ bl[49] br[49] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_52 
+ bl[50] br[50] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_53 
+ bl[51] br[51] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_54 
+ bl[52] br[52] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_55 
+ bl[53] br[53] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_56 
+ bl[54] br[54] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_57 
+ bl[55] br[55] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_58 
+ bl[56] br[56] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_59 
+ bl[57] br[57] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_60 
+ bl[58] br[58] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_61 
+ bl[59] br[59] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_62 
+ bl[60] br[60] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_63 
+ bl[61] br[61] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_64 
+ bl[62] br[62] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_65 
+ bl[63] br[63] vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_66 
+ vdd vdd vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_82_67 
+ vdd vdd vdd vss wl[80] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_0 
+ vdd vdd vss vdd vpb vnb wl[81] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_83_1 
+ rbl rbr vss vdd vpb vnb wl[81] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_83_2 
+ bl[0] br[0] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_3 
+ bl[1] br[1] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_4 
+ bl[2] br[2] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_5 
+ bl[3] br[3] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_6 
+ bl[4] br[4] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_7 
+ bl[5] br[5] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_8 
+ bl[6] br[6] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_9 
+ bl[7] br[7] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_10 
+ bl[8] br[8] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_11 
+ bl[9] br[9] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_12 
+ bl[10] br[10] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_13 
+ bl[11] br[11] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_14 
+ bl[12] br[12] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_15 
+ bl[13] br[13] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_16 
+ bl[14] br[14] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_17 
+ bl[15] br[15] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_18 
+ bl[16] br[16] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_19 
+ bl[17] br[17] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_20 
+ bl[18] br[18] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_21 
+ bl[19] br[19] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_22 
+ bl[20] br[20] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_23 
+ bl[21] br[21] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_24 
+ bl[22] br[22] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_25 
+ bl[23] br[23] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_26 
+ bl[24] br[24] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_27 
+ bl[25] br[25] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_28 
+ bl[26] br[26] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_29 
+ bl[27] br[27] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_30 
+ bl[28] br[28] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_31 
+ bl[29] br[29] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_32 
+ bl[30] br[30] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_33 
+ bl[31] br[31] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_34 
+ bl[32] br[32] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_35 
+ bl[33] br[33] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_36 
+ bl[34] br[34] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_37 
+ bl[35] br[35] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_38 
+ bl[36] br[36] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_39 
+ bl[37] br[37] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_40 
+ bl[38] br[38] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_41 
+ bl[39] br[39] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_42 
+ bl[40] br[40] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_43 
+ bl[41] br[41] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_44 
+ bl[42] br[42] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_45 
+ bl[43] br[43] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_46 
+ bl[44] br[44] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_47 
+ bl[45] br[45] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_48 
+ bl[46] br[46] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_49 
+ bl[47] br[47] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_50 
+ bl[48] br[48] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_51 
+ bl[49] br[49] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_52 
+ bl[50] br[50] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_53 
+ bl[51] br[51] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_54 
+ bl[52] br[52] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_55 
+ bl[53] br[53] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_56 
+ bl[54] br[54] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_57 
+ bl[55] br[55] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_58 
+ bl[56] br[56] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_59 
+ bl[57] br[57] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_60 
+ bl[58] br[58] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_61 
+ bl[59] br[59] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_62 
+ bl[60] br[60] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_63 
+ bl[61] br[61] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_64 
+ bl[62] br[62] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_65 
+ bl[63] br[63] vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_66 
+ vdd vdd vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_83_67 
+ vdd vdd vdd vss wl[81] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_0 
+ vdd vdd vss vdd vpb vnb wl[82] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_84_1 
+ rbl rbr vss vdd vpb vnb wl[82] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_84_2 
+ bl[0] br[0] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_3 
+ bl[1] br[1] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_4 
+ bl[2] br[2] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_5 
+ bl[3] br[3] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_6 
+ bl[4] br[4] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_7 
+ bl[5] br[5] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_8 
+ bl[6] br[6] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_9 
+ bl[7] br[7] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_10 
+ bl[8] br[8] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_11 
+ bl[9] br[9] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_12 
+ bl[10] br[10] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_13 
+ bl[11] br[11] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_14 
+ bl[12] br[12] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_15 
+ bl[13] br[13] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_16 
+ bl[14] br[14] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_17 
+ bl[15] br[15] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_18 
+ bl[16] br[16] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_19 
+ bl[17] br[17] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_20 
+ bl[18] br[18] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_21 
+ bl[19] br[19] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_22 
+ bl[20] br[20] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_23 
+ bl[21] br[21] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_24 
+ bl[22] br[22] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_25 
+ bl[23] br[23] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_26 
+ bl[24] br[24] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_27 
+ bl[25] br[25] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_28 
+ bl[26] br[26] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_29 
+ bl[27] br[27] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_30 
+ bl[28] br[28] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_31 
+ bl[29] br[29] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_32 
+ bl[30] br[30] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_33 
+ bl[31] br[31] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_34 
+ bl[32] br[32] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_35 
+ bl[33] br[33] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_36 
+ bl[34] br[34] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_37 
+ bl[35] br[35] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_38 
+ bl[36] br[36] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_39 
+ bl[37] br[37] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_40 
+ bl[38] br[38] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_41 
+ bl[39] br[39] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_42 
+ bl[40] br[40] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_43 
+ bl[41] br[41] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_44 
+ bl[42] br[42] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_45 
+ bl[43] br[43] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_46 
+ bl[44] br[44] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_47 
+ bl[45] br[45] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_48 
+ bl[46] br[46] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_49 
+ bl[47] br[47] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_50 
+ bl[48] br[48] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_51 
+ bl[49] br[49] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_52 
+ bl[50] br[50] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_53 
+ bl[51] br[51] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_54 
+ bl[52] br[52] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_55 
+ bl[53] br[53] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_56 
+ bl[54] br[54] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_57 
+ bl[55] br[55] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_58 
+ bl[56] br[56] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_59 
+ bl[57] br[57] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_60 
+ bl[58] br[58] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_61 
+ bl[59] br[59] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_62 
+ bl[60] br[60] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_63 
+ bl[61] br[61] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_64 
+ bl[62] br[62] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_65 
+ bl[63] br[63] vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_66 
+ vdd vdd vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_84_67 
+ vdd vdd vdd vss wl[82] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_0 
+ vdd vdd vss vdd vpb vnb wl[83] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_85_1 
+ rbl rbr vss vdd vpb vnb wl[83] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_85_2 
+ bl[0] br[0] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_3 
+ bl[1] br[1] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_4 
+ bl[2] br[2] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_5 
+ bl[3] br[3] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_6 
+ bl[4] br[4] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_7 
+ bl[5] br[5] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_8 
+ bl[6] br[6] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_9 
+ bl[7] br[7] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_10 
+ bl[8] br[8] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_11 
+ bl[9] br[9] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_12 
+ bl[10] br[10] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_13 
+ bl[11] br[11] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_14 
+ bl[12] br[12] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_15 
+ bl[13] br[13] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_16 
+ bl[14] br[14] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_17 
+ bl[15] br[15] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_18 
+ bl[16] br[16] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_19 
+ bl[17] br[17] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_20 
+ bl[18] br[18] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_21 
+ bl[19] br[19] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_22 
+ bl[20] br[20] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_23 
+ bl[21] br[21] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_24 
+ bl[22] br[22] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_25 
+ bl[23] br[23] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_26 
+ bl[24] br[24] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_27 
+ bl[25] br[25] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_28 
+ bl[26] br[26] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_29 
+ bl[27] br[27] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_30 
+ bl[28] br[28] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_31 
+ bl[29] br[29] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_32 
+ bl[30] br[30] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_33 
+ bl[31] br[31] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_34 
+ bl[32] br[32] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_35 
+ bl[33] br[33] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_36 
+ bl[34] br[34] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_37 
+ bl[35] br[35] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_38 
+ bl[36] br[36] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_39 
+ bl[37] br[37] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_40 
+ bl[38] br[38] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_41 
+ bl[39] br[39] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_42 
+ bl[40] br[40] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_43 
+ bl[41] br[41] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_44 
+ bl[42] br[42] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_45 
+ bl[43] br[43] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_46 
+ bl[44] br[44] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_47 
+ bl[45] br[45] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_48 
+ bl[46] br[46] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_49 
+ bl[47] br[47] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_50 
+ bl[48] br[48] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_51 
+ bl[49] br[49] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_52 
+ bl[50] br[50] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_53 
+ bl[51] br[51] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_54 
+ bl[52] br[52] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_55 
+ bl[53] br[53] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_56 
+ bl[54] br[54] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_57 
+ bl[55] br[55] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_58 
+ bl[56] br[56] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_59 
+ bl[57] br[57] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_60 
+ bl[58] br[58] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_61 
+ bl[59] br[59] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_62 
+ bl[60] br[60] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_63 
+ bl[61] br[61] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_64 
+ bl[62] br[62] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_65 
+ bl[63] br[63] vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_66 
+ vdd vdd vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_85_67 
+ vdd vdd vdd vss wl[83] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_0 
+ vdd vdd vss vdd vpb vnb wl[84] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_86_1 
+ rbl rbr vss vdd vpb vnb wl[84] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_86_2 
+ bl[0] br[0] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_3 
+ bl[1] br[1] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_4 
+ bl[2] br[2] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_5 
+ bl[3] br[3] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_6 
+ bl[4] br[4] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_7 
+ bl[5] br[5] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_8 
+ bl[6] br[6] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_9 
+ bl[7] br[7] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_10 
+ bl[8] br[8] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_11 
+ bl[9] br[9] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_12 
+ bl[10] br[10] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_13 
+ bl[11] br[11] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_14 
+ bl[12] br[12] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_15 
+ bl[13] br[13] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_16 
+ bl[14] br[14] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_17 
+ bl[15] br[15] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_18 
+ bl[16] br[16] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_19 
+ bl[17] br[17] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_20 
+ bl[18] br[18] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_21 
+ bl[19] br[19] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_22 
+ bl[20] br[20] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_23 
+ bl[21] br[21] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_24 
+ bl[22] br[22] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_25 
+ bl[23] br[23] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_26 
+ bl[24] br[24] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_27 
+ bl[25] br[25] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_28 
+ bl[26] br[26] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_29 
+ bl[27] br[27] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_30 
+ bl[28] br[28] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_31 
+ bl[29] br[29] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_32 
+ bl[30] br[30] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_33 
+ bl[31] br[31] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_34 
+ bl[32] br[32] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_35 
+ bl[33] br[33] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_36 
+ bl[34] br[34] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_37 
+ bl[35] br[35] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_38 
+ bl[36] br[36] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_39 
+ bl[37] br[37] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_40 
+ bl[38] br[38] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_41 
+ bl[39] br[39] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_42 
+ bl[40] br[40] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_43 
+ bl[41] br[41] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_44 
+ bl[42] br[42] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_45 
+ bl[43] br[43] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_46 
+ bl[44] br[44] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_47 
+ bl[45] br[45] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_48 
+ bl[46] br[46] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_49 
+ bl[47] br[47] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_50 
+ bl[48] br[48] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_51 
+ bl[49] br[49] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_52 
+ bl[50] br[50] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_53 
+ bl[51] br[51] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_54 
+ bl[52] br[52] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_55 
+ bl[53] br[53] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_56 
+ bl[54] br[54] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_57 
+ bl[55] br[55] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_58 
+ bl[56] br[56] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_59 
+ bl[57] br[57] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_60 
+ bl[58] br[58] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_61 
+ bl[59] br[59] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_62 
+ bl[60] br[60] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_63 
+ bl[61] br[61] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_64 
+ bl[62] br[62] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_65 
+ bl[63] br[63] vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_66 
+ vdd vdd vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_86_67 
+ vdd vdd vdd vss wl[84] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_0 
+ vdd vdd vss vdd vpb vnb wl[85] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_87_1 
+ rbl rbr vss vdd vpb vnb wl[85] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_87_2 
+ bl[0] br[0] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_3 
+ bl[1] br[1] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_4 
+ bl[2] br[2] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_5 
+ bl[3] br[3] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_6 
+ bl[4] br[4] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_7 
+ bl[5] br[5] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_8 
+ bl[6] br[6] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_9 
+ bl[7] br[7] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_10 
+ bl[8] br[8] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_11 
+ bl[9] br[9] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_12 
+ bl[10] br[10] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_13 
+ bl[11] br[11] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_14 
+ bl[12] br[12] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_15 
+ bl[13] br[13] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_16 
+ bl[14] br[14] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_17 
+ bl[15] br[15] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_18 
+ bl[16] br[16] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_19 
+ bl[17] br[17] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_20 
+ bl[18] br[18] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_21 
+ bl[19] br[19] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_22 
+ bl[20] br[20] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_23 
+ bl[21] br[21] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_24 
+ bl[22] br[22] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_25 
+ bl[23] br[23] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_26 
+ bl[24] br[24] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_27 
+ bl[25] br[25] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_28 
+ bl[26] br[26] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_29 
+ bl[27] br[27] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_30 
+ bl[28] br[28] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_31 
+ bl[29] br[29] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_32 
+ bl[30] br[30] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_33 
+ bl[31] br[31] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_34 
+ bl[32] br[32] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_35 
+ bl[33] br[33] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_36 
+ bl[34] br[34] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_37 
+ bl[35] br[35] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_38 
+ bl[36] br[36] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_39 
+ bl[37] br[37] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_40 
+ bl[38] br[38] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_41 
+ bl[39] br[39] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_42 
+ bl[40] br[40] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_43 
+ bl[41] br[41] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_44 
+ bl[42] br[42] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_45 
+ bl[43] br[43] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_46 
+ bl[44] br[44] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_47 
+ bl[45] br[45] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_48 
+ bl[46] br[46] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_49 
+ bl[47] br[47] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_50 
+ bl[48] br[48] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_51 
+ bl[49] br[49] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_52 
+ bl[50] br[50] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_53 
+ bl[51] br[51] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_54 
+ bl[52] br[52] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_55 
+ bl[53] br[53] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_56 
+ bl[54] br[54] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_57 
+ bl[55] br[55] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_58 
+ bl[56] br[56] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_59 
+ bl[57] br[57] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_60 
+ bl[58] br[58] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_61 
+ bl[59] br[59] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_62 
+ bl[60] br[60] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_63 
+ bl[61] br[61] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_64 
+ bl[62] br[62] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_65 
+ bl[63] br[63] vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_66 
+ vdd vdd vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_87_67 
+ vdd vdd vdd vss wl[85] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_0 
+ vdd vdd vss vdd vpb vnb wl[86] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_88_1 
+ rbl rbr vss vdd vpb vnb wl[86] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_88_2 
+ bl[0] br[0] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_3 
+ bl[1] br[1] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_4 
+ bl[2] br[2] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_5 
+ bl[3] br[3] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_6 
+ bl[4] br[4] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_7 
+ bl[5] br[5] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_8 
+ bl[6] br[6] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_9 
+ bl[7] br[7] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_10 
+ bl[8] br[8] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_11 
+ bl[9] br[9] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_12 
+ bl[10] br[10] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_13 
+ bl[11] br[11] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_14 
+ bl[12] br[12] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_15 
+ bl[13] br[13] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_16 
+ bl[14] br[14] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_17 
+ bl[15] br[15] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_18 
+ bl[16] br[16] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_19 
+ bl[17] br[17] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_20 
+ bl[18] br[18] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_21 
+ bl[19] br[19] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_22 
+ bl[20] br[20] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_23 
+ bl[21] br[21] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_24 
+ bl[22] br[22] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_25 
+ bl[23] br[23] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_26 
+ bl[24] br[24] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_27 
+ bl[25] br[25] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_28 
+ bl[26] br[26] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_29 
+ bl[27] br[27] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_30 
+ bl[28] br[28] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_31 
+ bl[29] br[29] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_32 
+ bl[30] br[30] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_33 
+ bl[31] br[31] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_34 
+ bl[32] br[32] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_35 
+ bl[33] br[33] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_36 
+ bl[34] br[34] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_37 
+ bl[35] br[35] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_38 
+ bl[36] br[36] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_39 
+ bl[37] br[37] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_40 
+ bl[38] br[38] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_41 
+ bl[39] br[39] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_42 
+ bl[40] br[40] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_43 
+ bl[41] br[41] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_44 
+ bl[42] br[42] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_45 
+ bl[43] br[43] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_46 
+ bl[44] br[44] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_47 
+ bl[45] br[45] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_48 
+ bl[46] br[46] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_49 
+ bl[47] br[47] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_50 
+ bl[48] br[48] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_51 
+ bl[49] br[49] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_52 
+ bl[50] br[50] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_53 
+ bl[51] br[51] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_54 
+ bl[52] br[52] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_55 
+ bl[53] br[53] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_56 
+ bl[54] br[54] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_57 
+ bl[55] br[55] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_58 
+ bl[56] br[56] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_59 
+ bl[57] br[57] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_60 
+ bl[58] br[58] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_61 
+ bl[59] br[59] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_62 
+ bl[60] br[60] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_63 
+ bl[61] br[61] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_64 
+ bl[62] br[62] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_65 
+ bl[63] br[63] vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_66 
+ vdd vdd vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_88_67 
+ vdd vdd vdd vss wl[86] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_0 
+ vdd vdd vss vdd vpb vnb wl[87] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_89_1 
+ rbl rbr vss vdd vpb vnb wl[87] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_89_2 
+ bl[0] br[0] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_3 
+ bl[1] br[1] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_4 
+ bl[2] br[2] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_5 
+ bl[3] br[3] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_6 
+ bl[4] br[4] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_7 
+ bl[5] br[5] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_8 
+ bl[6] br[6] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_9 
+ bl[7] br[7] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_10 
+ bl[8] br[8] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_11 
+ bl[9] br[9] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_12 
+ bl[10] br[10] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_13 
+ bl[11] br[11] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_14 
+ bl[12] br[12] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_15 
+ bl[13] br[13] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_16 
+ bl[14] br[14] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_17 
+ bl[15] br[15] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_18 
+ bl[16] br[16] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_19 
+ bl[17] br[17] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_20 
+ bl[18] br[18] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_21 
+ bl[19] br[19] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_22 
+ bl[20] br[20] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_23 
+ bl[21] br[21] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_24 
+ bl[22] br[22] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_25 
+ bl[23] br[23] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_26 
+ bl[24] br[24] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_27 
+ bl[25] br[25] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_28 
+ bl[26] br[26] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_29 
+ bl[27] br[27] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_30 
+ bl[28] br[28] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_31 
+ bl[29] br[29] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_32 
+ bl[30] br[30] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_33 
+ bl[31] br[31] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_34 
+ bl[32] br[32] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_35 
+ bl[33] br[33] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_36 
+ bl[34] br[34] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_37 
+ bl[35] br[35] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_38 
+ bl[36] br[36] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_39 
+ bl[37] br[37] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_40 
+ bl[38] br[38] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_41 
+ bl[39] br[39] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_42 
+ bl[40] br[40] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_43 
+ bl[41] br[41] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_44 
+ bl[42] br[42] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_45 
+ bl[43] br[43] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_46 
+ bl[44] br[44] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_47 
+ bl[45] br[45] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_48 
+ bl[46] br[46] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_49 
+ bl[47] br[47] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_50 
+ bl[48] br[48] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_51 
+ bl[49] br[49] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_52 
+ bl[50] br[50] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_53 
+ bl[51] br[51] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_54 
+ bl[52] br[52] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_55 
+ bl[53] br[53] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_56 
+ bl[54] br[54] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_57 
+ bl[55] br[55] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_58 
+ bl[56] br[56] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_59 
+ bl[57] br[57] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_60 
+ bl[58] br[58] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_61 
+ bl[59] br[59] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_62 
+ bl[60] br[60] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_63 
+ bl[61] br[61] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_64 
+ bl[62] br[62] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_65 
+ bl[63] br[63] vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_66 
+ vdd vdd vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_89_67 
+ vdd vdd vdd vss wl[87] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_0 
+ vdd vdd vss vdd vpb vnb wl[88] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_90_1 
+ rbl rbr vss vdd vpb vnb wl[88] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_90_2 
+ bl[0] br[0] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_3 
+ bl[1] br[1] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_4 
+ bl[2] br[2] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_5 
+ bl[3] br[3] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_6 
+ bl[4] br[4] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_7 
+ bl[5] br[5] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_8 
+ bl[6] br[6] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_9 
+ bl[7] br[7] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_10 
+ bl[8] br[8] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_11 
+ bl[9] br[9] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_12 
+ bl[10] br[10] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_13 
+ bl[11] br[11] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_14 
+ bl[12] br[12] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_15 
+ bl[13] br[13] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_16 
+ bl[14] br[14] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_17 
+ bl[15] br[15] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_18 
+ bl[16] br[16] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_19 
+ bl[17] br[17] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_20 
+ bl[18] br[18] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_21 
+ bl[19] br[19] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_22 
+ bl[20] br[20] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_23 
+ bl[21] br[21] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_24 
+ bl[22] br[22] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_25 
+ bl[23] br[23] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_26 
+ bl[24] br[24] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_27 
+ bl[25] br[25] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_28 
+ bl[26] br[26] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_29 
+ bl[27] br[27] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_30 
+ bl[28] br[28] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_31 
+ bl[29] br[29] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_32 
+ bl[30] br[30] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_33 
+ bl[31] br[31] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_34 
+ bl[32] br[32] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_35 
+ bl[33] br[33] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_36 
+ bl[34] br[34] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_37 
+ bl[35] br[35] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_38 
+ bl[36] br[36] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_39 
+ bl[37] br[37] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_40 
+ bl[38] br[38] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_41 
+ bl[39] br[39] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_42 
+ bl[40] br[40] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_43 
+ bl[41] br[41] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_44 
+ bl[42] br[42] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_45 
+ bl[43] br[43] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_46 
+ bl[44] br[44] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_47 
+ bl[45] br[45] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_48 
+ bl[46] br[46] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_49 
+ bl[47] br[47] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_50 
+ bl[48] br[48] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_51 
+ bl[49] br[49] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_52 
+ bl[50] br[50] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_53 
+ bl[51] br[51] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_54 
+ bl[52] br[52] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_55 
+ bl[53] br[53] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_56 
+ bl[54] br[54] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_57 
+ bl[55] br[55] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_58 
+ bl[56] br[56] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_59 
+ bl[57] br[57] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_60 
+ bl[58] br[58] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_61 
+ bl[59] br[59] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_62 
+ bl[60] br[60] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_63 
+ bl[61] br[61] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_64 
+ bl[62] br[62] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_65 
+ bl[63] br[63] vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_66 
+ vdd vdd vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_90_67 
+ vdd vdd vdd vss wl[88] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_0 
+ vdd vdd vss vdd vpb vnb wl[89] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_91_1 
+ rbl rbr vss vdd vpb vnb wl[89] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_91_2 
+ bl[0] br[0] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_3 
+ bl[1] br[1] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_4 
+ bl[2] br[2] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_5 
+ bl[3] br[3] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_6 
+ bl[4] br[4] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_7 
+ bl[5] br[5] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_8 
+ bl[6] br[6] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_9 
+ bl[7] br[7] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_10 
+ bl[8] br[8] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_11 
+ bl[9] br[9] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_12 
+ bl[10] br[10] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_13 
+ bl[11] br[11] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_14 
+ bl[12] br[12] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_15 
+ bl[13] br[13] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_16 
+ bl[14] br[14] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_17 
+ bl[15] br[15] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_18 
+ bl[16] br[16] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_19 
+ bl[17] br[17] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_20 
+ bl[18] br[18] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_21 
+ bl[19] br[19] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_22 
+ bl[20] br[20] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_23 
+ bl[21] br[21] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_24 
+ bl[22] br[22] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_25 
+ bl[23] br[23] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_26 
+ bl[24] br[24] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_27 
+ bl[25] br[25] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_28 
+ bl[26] br[26] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_29 
+ bl[27] br[27] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_30 
+ bl[28] br[28] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_31 
+ bl[29] br[29] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_32 
+ bl[30] br[30] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_33 
+ bl[31] br[31] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_34 
+ bl[32] br[32] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_35 
+ bl[33] br[33] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_36 
+ bl[34] br[34] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_37 
+ bl[35] br[35] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_38 
+ bl[36] br[36] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_39 
+ bl[37] br[37] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_40 
+ bl[38] br[38] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_41 
+ bl[39] br[39] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_42 
+ bl[40] br[40] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_43 
+ bl[41] br[41] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_44 
+ bl[42] br[42] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_45 
+ bl[43] br[43] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_46 
+ bl[44] br[44] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_47 
+ bl[45] br[45] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_48 
+ bl[46] br[46] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_49 
+ bl[47] br[47] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_50 
+ bl[48] br[48] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_51 
+ bl[49] br[49] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_52 
+ bl[50] br[50] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_53 
+ bl[51] br[51] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_54 
+ bl[52] br[52] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_55 
+ bl[53] br[53] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_56 
+ bl[54] br[54] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_57 
+ bl[55] br[55] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_58 
+ bl[56] br[56] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_59 
+ bl[57] br[57] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_60 
+ bl[58] br[58] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_61 
+ bl[59] br[59] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_62 
+ bl[60] br[60] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_63 
+ bl[61] br[61] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_64 
+ bl[62] br[62] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_65 
+ bl[63] br[63] vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_66 
+ vdd vdd vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_91_67 
+ vdd vdd vdd vss wl[89] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_0 
+ vdd vdd vss vdd vpb vnb wl[90] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_92_1 
+ rbl rbr vss vdd vpb vnb wl[90] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_92_2 
+ bl[0] br[0] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_3 
+ bl[1] br[1] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_4 
+ bl[2] br[2] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_5 
+ bl[3] br[3] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_6 
+ bl[4] br[4] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_7 
+ bl[5] br[5] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_8 
+ bl[6] br[6] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_9 
+ bl[7] br[7] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_10 
+ bl[8] br[8] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_11 
+ bl[9] br[9] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_12 
+ bl[10] br[10] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_13 
+ bl[11] br[11] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_14 
+ bl[12] br[12] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_15 
+ bl[13] br[13] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_16 
+ bl[14] br[14] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_17 
+ bl[15] br[15] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_18 
+ bl[16] br[16] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_19 
+ bl[17] br[17] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_20 
+ bl[18] br[18] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_21 
+ bl[19] br[19] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_22 
+ bl[20] br[20] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_23 
+ bl[21] br[21] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_24 
+ bl[22] br[22] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_25 
+ bl[23] br[23] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_26 
+ bl[24] br[24] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_27 
+ bl[25] br[25] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_28 
+ bl[26] br[26] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_29 
+ bl[27] br[27] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_30 
+ bl[28] br[28] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_31 
+ bl[29] br[29] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_32 
+ bl[30] br[30] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_33 
+ bl[31] br[31] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_34 
+ bl[32] br[32] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_35 
+ bl[33] br[33] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_36 
+ bl[34] br[34] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_37 
+ bl[35] br[35] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_38 
+ bl[36] br[36] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_39 
+ bl[37] br[37] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_40 
+ bl[38] br[38] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_41 
+ bl[39] br[39] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_42 
+ bl[40] br[40] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_43 
+ bl[41] br[41] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_44 
+ bl[42] br[42] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_45 
+ bl[43] br[43] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_46 
+ bl[44] br[44] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_47 
+ bl[45] br[45] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_48 
+ bl[46] br[46] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_49 
+ bl[47] br[47] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_50 
+ bl[48] br[48] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_51 
+ bl[49] br[49] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_52 
+ bl[50] br[50] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_53 
+ bl[51] br[51] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_54 
+ bl[52] br[52] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_55 
+ bl[53] br[53] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_56 
+ bl[54] br[54] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_57 
+ bl[55] br[55] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_58 
+ bl[56] br[56] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_59 
+ bl[57] br[57] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_60 
+ bl[58] br[58] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_61 
+ bl[59] br[59] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_62 
+ bl[60] br[60] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_63 
+ bl[61] br[61] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_64 
+ bl[62] br[62] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_65 
+ bl[63] br[63] vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_66 
+ vdd vdd vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_92_67 
+ vdd vdd vdd vss wl[90] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_0 
+ vdd vdd vss vdd vpb vnb wl[91] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_93_1 
+ rbl rbr vss vdd vpb vnb wl[91] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_93_2 
+ bl[0] br[0] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_3 
+ bl[1] br[1] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_4 
+ bl[2] br[2] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_5 
+ bl[3] br[3] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_6 
+ bl[4] br[4] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_7 
+ bl[5] br[5] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_8 
+ bl[6] br[6] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_9 
+ bl[7] br[7] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_10 
+ bl[8] br[8] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_11 
+ bl[9] br[9] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_12 
+ bl[10] br[10] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_13 
+ bl[11] br[11] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_14 
+ bl[12] br[12] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_15 
+ bl[13] br[13] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_16 
+ bl[14] br[14] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_17 
+ bl[15] br[15] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_18 
+ bl[16] br[16] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_19 
+ bl[17] br[17] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_20 
+ bl[18] br[18] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_21 
+ bl[19] br[19] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_22 
+ bl[20] br[20] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_23 
+ bl[21] br[21] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_24 
+ bl[22] br[22] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_25 
+ bl[23] br[23] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_26 
+ bl[24] br[24] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_27 
+ bl[25] br[25] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_28 
+ bl[26] br[26] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_29 
+ bl[27] br[27] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_30 
+ bl[28] br[28] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_31 
+ bl[29] br[29] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_32 
+ bl[30] br[30] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_33 
+ bl[31] br[31] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_34 
+ bl[32] br[32] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_35 
+ bl[33] br[33] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_36 
+ bl[34] br[34] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_37 
+ bl[35] br[35] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_38 
+ bl[36] br[36] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_39 
+ bl[37] br[37] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_40 
+ bl[38] br[38] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_41 
+ bl[39] br[39] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_42 
+ bl[40] br[40] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_43 
+ bl[41] br[41] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_44 
+ bl[42] br[42] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_45 
+ bl[43] br[43] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_46 
+ bl[44] br[44] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_47 
+ bl[45] br[45] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_48 
+ bl[46] br[46] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_49 
+ bl[47] br[47] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_50 
+ bl[48] br[48] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_51 
+ bl[49] br[49] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_52 
+ bl[50] br[50] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_53 
+ bl[51] br[51] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_54 
+ bl[52] br[52] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_55 
+ bl[53] br[53] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_56 
+ bl[54] br[54] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_57 
+ bl[55] br[55] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_58 
+ bl[56] br[56] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_59 
+ bl[57] br[57] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_60 
+ bl[58] br[58] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_61 
+ bl[59] br[59] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_62 
+ bl[60] br[60] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_63 
+ bl[61] br[61] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_64 
+ bl[62] br[62] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_65 
+ bl[63] br[63] vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_66 
+ vdd vdd vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_93_67 
+ vdd vdd vdd vss wl[91] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_0 
+ vdd vdd vss vdd vpb vnb wl[92] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_94_1 
+ rbl rbr vss vdd vpb vnb wl[92] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_94_2 
+ bl[0] br[0] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_3 
+ bl[1] br[1] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_4 
+ bl[2] br[2] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_5 
+ bl[3] br[3] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_6 
+ bl[4] br[4] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_7 
+ bl[5] br[5] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_8 
+ bl[6] br[6] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_9 
+ bl[7] br[7] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_10 
+ bl[8] br[8] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_11 
+ bl[9] br[9] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_12 
+ bl[10] br[10] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_13 
+ bl[11] br[11] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_14 
+ bl[12] br[12] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_15 
+ bl[13] br[13] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_16 
+ bl[14] br[14] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_17 
+ bl[15] br[15] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_18 
+ bl[16] br[16] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_19 
+ bl[17] br[17] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_20 
+ bl[18] br[18] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_21 
+ bl[19] br[19] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_22 
+ bl[20] br[20] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_23 
+ bl[21] br[21] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_24 
+ bl[22] br[22] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_25 
+ bl[23] br[23] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_26 
+ bl[24] br[24] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_27 
+ bl[25] br[25] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_28 
+ bl[26] br[26] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_29 
+ bl[27] br[27] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_30 
+ bl[28] br[28] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_31 
+ bl[29] br[29] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_32 
+ bl[30] br[30] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_33 
+ bl[31] br[31] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_34 
+ bl[32] br[32] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_35 
+ bl[33] br[33] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_36 
+ bl[34] br[34] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_37 
+ bl[35] br[35] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_38 
+ bl[36] br[36] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_39 
+ bl[37] br[37] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_40 
+ bl[38] br[38] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_41 
+ bl[39] br[39] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_42 
+ bl[40] br[40] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_43 
+ bl[41] br[41] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_44 
+ bl[42] br[42] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_45 
+ bl[43] br[43] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_46 
+ bl[44] br[44] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_47 
+ bl[45] br[45] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_48 
+ bl[46] br[46] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_49 
+ bl[47] br[47] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_50 
+ bl[48] br[48] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_51 
+ bl[49] br[49] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_52 
+ bl[50] br[50] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_53 
+ bl[51] br[51] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_54 
+ bl[52] br[52] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_55 
+ bl[53] br[53] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_56 
+ bl[54] br[54] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_57 
+ bl[55] br[55] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_58 
+ bl[56] br[56] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_59 
+ bl[57] br[57] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_60 
+ bl[58] br[58] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_61 
+ bl[59] br[59] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_62 
+ bl[60] br[60] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_63 
+ bl[61] br[61] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_64 
+ bl[62] br[62] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_65 
+ bl[63] br[63] vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_66 
+ vdd vdd vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_94_67 
+ vdd vdd vdd vss wl[92] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_0 
+ vdd vdd vss vdd vpb vnb wl[93] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_95_1 
+ rbl rbr vss vdd vpb vnb wl[93] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_95_2 
+ bl[0] br[0] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_3 
+ bl[1] br[1] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_4 
+ bl[2] br[2] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_5 
+ bl[3] br[3] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_6 
+ bl[4] br[4] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_7 
+ bl[5] br[5] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_8 
+ bl[6] br[6] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_9 
+ bl[7] br[7] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_10 
+ bl[8] br[8] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_11 
+ bl[9] br[9] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_12 
+ bl[10] br[10] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_13 
+ bl[11] br[11] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_14 
+ bl[12] br[12] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_15 
+ bl[13] br[13] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_16 
+ bl[14] br[14] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_17 
+ bl[15] br[15] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_18 
+ bl[16] br[16] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_19 
+ bl[17] br[17] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_20 
+ bl[18] br[18] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_21 
+ bl[19] br[19] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_22 
+ bl[20] br[20] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_23 
+ bl[21] br[21] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_24 
+ bl[22] br[22] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_25 
+ bl[23] br[23] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_26 
+ bl[24] br[24] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_27 
+ bl[25] br[25] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_28 
+ bl[26] br[26] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_29 
+ bl[27] br[27] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_30 
+ bl[28] br[28] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_31 
+ bl[29] br[29] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_32 
+ bl[30] br[30] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_33 
+ bl[31] br[31] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_34 
+ bl[32] br[32] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_35 
+ bl[33] br[33] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_36 
+ bl[34] br[34] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_37 
+ bl[35] br[35] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_38 
+ bl[36] br[36] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_39 
+ bl[37] br[37] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_40 
+ bl[38] br[38] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_41 
+ bl[39] br[39] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_42 
+ bl[40] br[40] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_43 
+ bl[41] br[41] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_44 
+ bl[42] br[42] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_45 
+ bl[43] br[43] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_46 
+ bl[44] br[44] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_47 
+ bl[45] br[45] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_48 
+ bl[46] br[46] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_49 
+ bl[47] br[47] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_50 
+ bl[48] br[48] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_51 
+ bl[49] br[49] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_52 
+ bl[50] br[50] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_53 
+ bl[51] br[51] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_54 
+ bl[52] br[52] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_55 
+ bl[53] br[53] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_56 
+ bl[54] br[54] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_57 
+ bl[55] br[55] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_58 
+ bl[56] br[56] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_59 
+ bl[57] br[57] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_60 
+ bl[58] br[58] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_61 
+ bl[59] br[59] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_62 
+ bl[60] br[60] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_63 
+ bl[61] br[61] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_64 
+ bl[62] br[62] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_65 
+ bl[63] br[63] vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_66 
+ vdd vdd vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_95_67 
+ vdd vdd vdd vss wl[93] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_0 
+ vdd vdd vss vdd vpb vnb wl[94] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_96_1 
+ rbl rbr vss vdd vpb vnb wl[94] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_96_2 
+ bl[0] br[0] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_3 
+ bl[1] br[1] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_4 
+ bl[2] br[2] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_5 
+ bl[3] br[3] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_6 
+ bl[4] br[4] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_7 
+ bl[5] br[5] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_8 
+ bl[6] br[6] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_9 
+ bl[7] br[7] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_10 
+ bl[8] br[8] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_11 
+ bl[9] br[9] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_12 
+ bl[10] br[10] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_13 
+ bl[11] br[11] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_14 
+ bl[12] br[12] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_15 
+ bl[13] br[13] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_16 
+ bl[14] br[14] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_17 
+ bl[15] br[15] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_18 
+ bl[16] br[16] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_19 
+ bl[17] br[17] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_20 
+ bl[18] br[18] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_21 
+ bl[19] br[19] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_22 
+ bl[20] br[20] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_23 
+ bl[21] br[21] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_24 
+ bl[22] br[22] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_25 
+ bl[23] br[23] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_26 
+ bl[24] br[24] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_27 
+ bl[25] br[25] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_28 
+ bl[26] br[26] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_29 
+ bl[27] br[27] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_30 
+ bl[28] br[28] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_31 
+ bl[29] br[29] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_32 
+ bl[30] br[30] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_33 
+ bl[31] br[31] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_34 
+ bl[32] br[32] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_35 
+ bl[33] br[33] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_36 
+ bl[34] br[34] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_37 
+ bl[35] br[35] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_38 
+ bl[36] br[36] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_39 
+ bl[37] br[37] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_40 
+ bl[38] br[38] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_41 
+ bl[39] br[39] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_42 
+ bl[40] br[40] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_43 
+ bl[41] br[41] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_44 
+ bl[42] br[42] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_45 
+ bl[43] br[43] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_46 
+ bl[44] br[44] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_47 
+ bl[45] br[45] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_48 
+ bl[46] br[46] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_49 
+ bl[47] br[47] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_50 
+ bl[48] br[48] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_51 
+ bl[49] br[49] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_52 
+ bl[50] br[50] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_53 
+ bl[51] br[51] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_54 
+ bl[52] br[52] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_55 
+ bl[53] br[53] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_56 
+ bl[54] br[54] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_57 
+ bl[55] br[55] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_58 
+ bl[56] br[56] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_59 
+ bl[57] br[57] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_60 
+ bl[58] br[58] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_61 
+ bl[59] br[59] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_62 
+ bl[60] br[60] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_63 
+ bl[61] br[61] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_64 
+ bl[62] br[62] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_65 
+ bl[63] br[63] vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_66 
+ vdd vdd vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_96_67 
+ vdd vdd vdd vss wl[94] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_0 
+ vdd vdd vss vdd vpb vnb wl[95] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_97_1 
+ rbl rbr vss vdd vpb vnb wl[95] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_97_2 
+ bl[0] br[0] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_3 
+ bl[1] br[1] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_4 
+ bl[2] br[2] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_5 
+ bl[3] br[3] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_6 
+ bl[4] br[4] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_7 
+ bl[5] br[5] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_8 
+ bl[6] br[6] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_9 
+ bl[7] br[7] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_10 
+ bl[8] br[8] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_11 
+ bl[9] br[9] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_12 
+ bl[10] br[10] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_13 
+ bl[11] br[11] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_14 
+ bl[12] br[12] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_15 
+ bl[13] br[13] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_16 
+ bl[14] br[14] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_17 
+ bl[15] br[15] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_18 
+ bl[16] br[16] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_19 
+ bl[17] br[17] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_20 
+ bl[18] br[18] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_21 
+ bl[19] br[19] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_22 
+ bl[20] br[20] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_23 
+ bl[21] br[21] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_24 
+ bl[22] br[22] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_25 
+ bl[23] br[23] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_26 
+ bl[24] br[24] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_27 
+ bl[25] br[25] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_28 
+ bl[26] br[26] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_29 
+ bl[27] br[27] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_30 
+ bl[28] br[28] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_31 
+ bl[29] br[29] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_32 
+ bl[30] br[30] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_33 
+ bl[31] br[31] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_34 
+ bl[32] br[32] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_35 
+ bl[33] br[33] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_36 
+ bl[34] br[34] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_37 
+ bl[35] br[35] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_38 
+ bl[36] br[36] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_39 
+ bl[37] br[37] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_40 
+ bl[38] br[38] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_41 
+ bl[39] br[39] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_42 
+ bl[40] br[40] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_43 
+ bl[41] br[41] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_44 
+ bl[42] br[42] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_45 
+ bl[43] br[43] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_46 
+ bl[44] br[44] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_47 
+ bl[45] br[45] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_48 
+ bl[46] br[46] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_49 
+ bl[47] br[47] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_50 
+ bl[48] br[48] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_51 
+ bl[49] br[49] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_52 
+ bl[50] br[50] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_53 
+ bl[51] br[51] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_54 
+ bl[52] br[52] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_55 
+ bl[53] br[53] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_56 
+ bl[54] br[54] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_57 
+ bl[55] br[55] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_58 
+ bl[56] br[56] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_59 
+ bl[57] br[57] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_60 
+ bl[58] br[58] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_61 
+ bl[59] br[59] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_62 
+ bl[60] br[60] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_63 
+ bl[61] br[61] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_64 
+ bl[62] br[62] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_65 
+ bl[63] br[63] vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_66 
+ vdd vdd vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_97_67 
+ vdd vdd vdd vss wl[95] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_0 
+ vdd vdd vss vdd vpb vnb wl[96] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_98_1 
+ rbl rbr vss vdd vpb vnb wl[96] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_98_2 
+ bl[0] br[0] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_3 
+ bl[1] br[1] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_4 
+ bl[2] br[2] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_5 
+ bl[3] br[3] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_6 
+ bl[4] br[4] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_7 
+ bl[5] br[5] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_8 
+ bl[6] br[6] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_9 
+ bl[7] br[7] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_10 
+ bl[8] br[8] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_11 
+ bl[9] br[9] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_12 
+ bl[10] br[10] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_13 
+ bl[11] br[11] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_14 
+ bl[12] br[12] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_15 
+ bl[13] br[13] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_16 
+ bl[14] br[14] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_17 
+ bl[15] br[15] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_18 
+ bl[16] br[16] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_19 
+ bl[17] br[17] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_20 
+ bl[18] br[18] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_21 
+ bl[19] br[19] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_22 
+ bl[20] br[20] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_23 
+ bl[21] br[21] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_24 
+ bl[22] br[22] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_25 
+ bl[23] br[23] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_26 
+ bl[24] br[24] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_27 
+ bl[25] br[25] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_28 
+ bl[26] br[26] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_29 
+ bl[27] br[27] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_30 
+ bl[28] br[28] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_31 
+ bl[29] br[29] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_32 
+ bl[30] br[30] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_33 
+ bl[31] br[31] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_34 
+ bl[32] br[32] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_35 
+ bl[33] br[33] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_36 
+ bl[34] br[34] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_37 
+ bl[35] br[35] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_38 
+ bl[36] br[36] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_39 
+ bl[37] br[37] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_40 
+ bl[38] br[38] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_41 
+ bl[39] br[39] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_42 
+ bl[40] br[40] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_43 
+ bl[41] br[41] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_44 
+ bl[42] br[42] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_45 
+ bl[43] br[43] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_46 
+ bl[44] br[44] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_47 
+ bl[45] br[45] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_48 
+ bl[46] br[46] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_49 
+ bl[47] br[47] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_50 
+ bl[48] br[48] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_51 
+ bl[49] br[49] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_52 
+ bl[50] br[50] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_53 
+ bl[51] br[51] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_54 
+ bl[52] br[52] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_55 
+ bl[53] br[53] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_56 
+ bl[54] br[54] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_57 
+ bl[55] br[55] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_58 
+ bl[56] br[56] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_59 
+ bl[57] br[57] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_60 
+ bl[58] br[58] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_61 
+ bl[59] br[59] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_62 
+ bl[60] br[60] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_63 
+ bl[61] br[61] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_64 
+ bl[62] br[62] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_65 
+ bl[63] br[63] vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_66 
+ vdd vdd vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_98_67 
+ vdd vdd vdd vss wl[96] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_0 
+ vdd vdd vss vdd vpb vnb wl[97] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_99_1 
+ rbl rbr vss vdd vpb vnb wl[97] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_99_2 
+ bl[0] br[0] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_3 
+ bl[1] br[1] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_4 
+ bl[2] br[2] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_5 
+ bl[3] br[3] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_6 
+ bl[4] br[4] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_7 
+ bl[5] br[5] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_8 
+ bl[6] br[6] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_9 
+ bl[7] br[7] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_10 
+ bl[8] br[8] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_11 
+ bl[9] br[9] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_12 
+ bl[10] br[10] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_13 
+ bl[11] br[11] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_14 
+ bl[12] br[12] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_15 
+ bl[13] br[13] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_16 
+ bl[14] br[14] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_17 
+ bl[15] br[15] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_18 
+ bl[16] br[16] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_19 
+ bl[17] br[17] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_20 
+ bl[18] br[18] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_21 
+ bl[19] br[19] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_22 
+ bl[20] br[20] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_23 
+ bl[21] br[21] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_24 
+ bl[22] br[22] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_25 
+ bl[23] br[23] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_26 
+ bl[24] br[24] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_27 
+ bl[25] br[25] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_28 
+ bl[26] br[26] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_29 
+ bl[27] br[27] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_30 
+ bl[28] br[28] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_31 
+ bl[29] br[29] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_32 
+ bl[30] br[30] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_33 
+ bl[31] br[31] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_34 
+ bl[32] br[32] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_35 
+ bl[33] br[33] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_36 
+ bl[34] br[34] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_37 
+ bl[35] br[35] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_38 
+ bl[36] br[36] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_39 
+ bl[37] br[37] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_40 
+ bl[38] br[38] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_41 
+ bl[39] br[39] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_42 
+ bl[40] br[40] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_43 
+ bl[41] br[41] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_44 
+ bl[42] br[42] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_45 
+ bl[43] br[43] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_46 
+ bl[44] br[44] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_47 
+ bl[45] br[45] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_48 
+ bl[46] br[46] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_49 
+ bl[47] br[47] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_50 
+ bl[48] br[48] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_51 
+ bl[49] br[49] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_52 
+ bl[50] br[50] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_53 
+ bl[51] br[51] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_54 
+ bl[52] br[52] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_55 
+ bl[53] br[53] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_56 
+ bl[54] br[54] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_57 
+ bl[55] br[55] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_58 
+ bl[56] br[56] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_59 
+ bl[57] br[57] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_60 
+ bl[58] br[58] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_61 
+ bl[59] br[59] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_62 
+ bl[60] br[60] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_63 
+ bl[61] br[61] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_64 
+ bl[62] br[62] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_65 
+ bl[63] br[63] vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_66 
+ vdd vdd vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_99_67 
+ vdd vdd vdd vss wl[97] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_0 
+ vdd vdd vss vdd vpb vnb wl[98] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_100_1 
+ rbl rbr vss vdd vpb vnb wl[98] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_100_2 
+ bl[0] br[0] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_3 
+ bl[1] br[1] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_4 
+ bl[2] br[2] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_5 
+ bl[3] br[3] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_6 
+ bl[4] br[4] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_7 
+ bl[5] br[5] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_8 
+ bl[6] br[6] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_9 
+ bl[7] br[7] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_10 
+ bl[8] br[8] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_11 
+ bl[9] br[9] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_12 
+ bl[10] br[10] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_13 
+ bl[11] br[11] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_14 
+ bl[12] br[12] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_15 
+ bl[13] br[13] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_16 
+ bl[14] br[14] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_17 
+ bl[15] br[15] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_18 
+ bl[16] br[16] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_19 
+ bl[17] br[17] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_20 
+ bl[18] br[18] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_21 
+ bl[19] br[19] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_22 
+ bl[20] br[20] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_23 
+ bl[21] br[21] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_24 
+ bl[22] br[22] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_25 
+ bl[23] br[23] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_26 
+ bl[24] br[24] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_27 
+ bl[25] br[25] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_28 
+ bl[26] br[26] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_29 
+ bl[27] br[27] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_30 
+ bl[28] br[28] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_31 
+ bl[29] br[29] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_32 
+ bl[30] br[30] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_33 
+ bl[31] br[31] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_34 
+ bl[32] br[32] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_35 
+ bl[33] br[33] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_36 
+ bl[34] br[34] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_37 
+ bl[35] br[35] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_38 
+ bl[36] br[36] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_39 
+ bl[37] br[37] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_40 
+ bl[38] br[38] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_41 
+ bl[39] br[39] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_42 
+ bl[40] br[40] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_43 
+ bl[41] br[41] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_44 
+ bl[42] br[42] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_45 
+ bl[43] br[43] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_46 
+ bl[44] br[44] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_47 
+ bl[45] br[45] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_48 
+ bl[46] br[46] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_49 
+ bl[47] br[47] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_50 
+ bl[48] br[48] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_51 
+ bl[49] br[49] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_52 
+ bl[50] br[50] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_53 
+ bl[51] br[51] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_54 
+ bl[52] br[52] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_55 
+ bl[53] br[53] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_56 
+ bl[54] br[54] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_57 
+ bl[55] br[55] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_58 
+ bl[56] br[56] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_59 
+ bl[57] br[57] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_60 
+ bl[58] br[58] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_61 
+ bl[59] br[59] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_62 
+ bl[60] br[60] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_63 
+ bl[61] br[61] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_64 
+ bl[62] br[62] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_65 
+ bl[63] br[63] vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_66 
+ vdd vdd vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_100_67 
+ vdd vdd vdd vss wl[98] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_0 
+ vdd vdd vss vdd vpb vnb wl[99] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_101_1 
+ rbl rbr vss vdd vpb vnb wl[99] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_101_2 
+ bl[0] br[0] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_3 
+ bl[1] br[1] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_4 
+ bl[2] br[2] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_5 
+ bl[3] br[3] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_6 
+ bl[4] br[4] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_7 
+ bl[5] br[5] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_8 
+ bl[6] br[6] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_9 
+ bl[7] br[7] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_10 
+ bl[8] br[8] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_11 
+ bl[9] br[9] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_12 
+ bl[10] br[10] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_13 
+ bl[11] br[11] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_14 
+ bl[12] br[12] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_15 
+ bl[13] br[13] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_16 
+ bl[14] br[14] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_17 
+ bl[15] br[15] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_18 
+ bl[16] br[16] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_19 
+ bl[17] br[17] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_20 
+ bl[18] br[18] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_21 
+ bl[19] br[19] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_22 
+ bl[20] br[20] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_23 
+ bl[21] br[21] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_24 
+ bl[22] br[22] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_25 
+ bl[23] br[23] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_26 
+ bl[24] br[24] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_27 
+ bl[25] br[25] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_28 
+ bl[26] br[26] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_29 
+ bl[27] br[27] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_30 
+ bl[28] br[28] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_31 
+ bl[29] br[29] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_32 
+ bl[30] br[30] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_33 
+ bl[31] br[31] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_34 
+ bl[32] br[32] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_35 
+ bl[33] br[33] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_36 
+ bl[34] br[34] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_37 
+ bl[35] br[35] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_38 
+ bl[36] br[36] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_39 
+ bl[37] br[37] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_40 
+ bl[38] br[38] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_41 
+ bl[39] br[39] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_42 
+ bl[40] br[40] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_43 
+ bl[41] br[41] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_44 
+ bl[42] br[42] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_45 
+ bl[43] br[43] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_46 
+ bl[44] br[44] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_47 
+ bl[45] br[45] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_48 
+ bl[46] br[46] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_49 
+ bl[47] br[47] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_50 
+ bl[48] br[48] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_51 
+ bl[49] br[49] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_52 
+ bl[50] br[50] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_53 
+ bl[51] br[51] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_54 
+ bl[52] br[52] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_55 
+ bl[53] br[53] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_56 
+ bl[54] br[54] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_57 
+ bl[55] br[55] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_58 
+ bl[56] br[56] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_59 
+ bl[57] br[57] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_60 
+ bl[58] br[58] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_61 
+ bl[59] br[59] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_62 
+ bl[60] br[60] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_63 
+ bl[61] br[61] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_64 
+ bl[62] br[62] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_65 
+ bl[63] br[63] vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_66 
+ vdd vdd vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_101_67 
+ vdd vdd vdd vss wl[99] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_0 
+ vdd vdd vss vdd vpb vnb wl[100] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_102_1 
+ rbl rbr vss vdd vpb vnb wl[100] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_102_2 
+ bl[0] br[0] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_3 
+ bl[1] br[1] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_4 
+ bl[2] br[2] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_5 
+ bl[3] br[3] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_6 
+ bl[4] br[4] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_7 
+ bl[5] br[5] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_8 
+ bl[6] br[6] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_9 
+ bl[7] br[7] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_10 
+ bl[8] br[8] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_11 
+ bl[9] br[9] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_12 
+ bl[10] br[10] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_13 
+ bl[11] br[11] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_14 
+ bl[12] br[12] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_15 
+ bl[13] br[13] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_16 
+ bl[14] br[14] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_17 
+ bl[15] br[15] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_18 
+ bl[16] br[16] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_19 
+ bl[17] br[17] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_20 
+ bl[18] br[18] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_21 
+ bl[19] br[19] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_22 
+ bl[20] br[20] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_23 
+ bl[21] br[21] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_24 
+ bl[22] br[22] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_25 
+ bl[23] br[23] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_26 
+ bl[24] br[24] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_27 
+ bl[25] br[25] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_28 
+ bl[26] br[26] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_29 
+ bl[27] br[27] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_30 
+ bl[28] br[28] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_31 
+ bl[29] br[29] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_32 
+ bl[30] br[30] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_33 
+ bl[31] br[31] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_34 
+ bl[32] br[32] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_35 
+ bl[33] br[33] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_36 
+ bl[34] br[34] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_37 
+ bl[35] br[35] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_38 
+ bl[36] br[36] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_39 
+ bl[37] br[37] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_40 
+ bl[38] br[38] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_41 
+ bl[39] br[39] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_42 
+ bl[40] br[40] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_43 
+ bl[41] br[41] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_44 
+ bl[42] br[42] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_45 
+ bl[43] br[43] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_46 
+ bl[44] br[44] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_47 
+ bl[45] br[45] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_48 
+ bl[46] br[46] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_49 
+ bl[47] br[47] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_50 
+ bl[48] br[48] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_51 
+ bl[49] br[49] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_52 
+ bl[50] br[50] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_53 
+ bl[51] br[51] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_54 
+ bl[52] br[52] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_55 
+ bl[53] br[53] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_56 
+ bl[54] br[54] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_57 
+ bl[55] br[55] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_58 
+ bl[56] br[56] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_59 
+ bl[57] br[57] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_60 
+ bl[58] br[58] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_61 
+ bl[59] br[59] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_62 
+ bl[60] br[60] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_63 
+ bl[61] br[61] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_64 
+ bl[62] br[62] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_65 
+ bl[63] br[63] vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_66 
+ vdd vdd vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_102_67 
+ vdd vdd vdd vss wl[100] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_0 
+ vdd vdd vss vdd vpb vnb wl[101] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_103_1 
+ rbl rbr vss vdd vpb vnb wl[101] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_103_2 
+ bl[0] br[0] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_3 
+ bl[1] br[1] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_4 
+ bl[2] br[2] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_5 
+ bl[3] br[3] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_6 
+ bl[4] br[4] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_7 
+ bl[5] br[5] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_8 
+ bl[6] br[6] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_9 
+ bl[7] br[7] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_10 
+ bl[8] br[8] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_11 
+ bl[9] br[9] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_12 
+ bl[10] br[10] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_13 
+ bl[11] br[11] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_14 
+ bl[12] br[12] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_15 
+ bl[13] br[13] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_16 
+ bl[14] br[14] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_17 
+ bl[15] br[15] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_18 
+ bl[16] br[16] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_19 
+ bl[17] br[17] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_20 
+ bl[18] br[18] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_21 
+ bl[19] br[19] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_22 
+ bl[20] br[20] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_23 
+ bl[21] br[21] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_24 
+ bl[22] br[22] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_25 
+ bl[23] br[23] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_26 
+ bl[24] br[24] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_27 
+ bl[25] br[25] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_28 
+ bl[26] br[26] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_29 
+ bl[27] br[27] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_30 
+ bl[28] br[28] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_31 
+ bl[29] br[29] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_32 
+ bl[30] br[30] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_33 
+ bl[31] br[31] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_34 
+ bl[32] br[32] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_35 
+ bl[33] br[33] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_36 
+ bl[34] br[34] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_37 
+ bl[35] br[35] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_38 
+ bl[36] br[36] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_39 
+ bl[37] br[37] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_40 
+ bl[38] br[38] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_41 
+ bl[39] br[39] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_42 
+ bl[40] br[40] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_43 
+ bl[41] br[41] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_44 
+ bl[42] br[42] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_45 
+ bl[43] br[43] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_46 
+ bl[44] br[44] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_47 
+ bl[45] br[45] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_48 
+ bl[46] br[46] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_49 
+ bl[47] br[47] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_50 
+ bl[48] br[48] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_51 
+ bl[49] br[49] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_52 
+ bl[50] br[50] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_53 
+ bl[51] br[51] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_54 
+ bl[52] br[52] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_55 
+ bl[53] br[53] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_56 
+ bl[54] br[54] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_57 
+ bl[55] br[55] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_58 
+ bl[56] br[56] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_59 
+ bl[57] br[57] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_60 
+ bl[58] br[58] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_61 
+ bl[59] br[59] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_62 
+ bl[60] br[60] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_63 
+ bl[61] br[61] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_64 
+ bl[62] br[62] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_65 
+ bl[63] br[63] vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_66 
+ vdd vdd vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_103_67 
+ vdd vdd vdd vss wl[101] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_0 
+ vdd vdd vss vdd vpb vnb wl[102] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_104_1 
+ rbl rbr vss vdd vpb vnb wl[102] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_104_2 
+ bl[0] br[0] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_3 
+ bl[1] br[1] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_4 
+ bl[2] br[2] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_5 
+ bl[3] br[3] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_6 
+ bl[4] br[4] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_7 
+ bl[5] br[5] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_8 
+ bl[6] br[6] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_9 
+ bl[7] br[7] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_10 
+ bl[8] br[8] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_11 
+ bl[9] br[9] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_12 
+ bl[10] br[10] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_13 
+ bl[11] br[11] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_14 
+ bl[12] br[12] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_15 
+ bl[13] br[13] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_16 
+ bl[14] br[14] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_17 
+ bl[15] br[15] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_18 
+ bl[16] br[16] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_19 
+ bl[17] br[17] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_20 
+ bl[18] br[18] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_21 
+ bl[19] br[19] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_22 
+ bl[20] br[20] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_23 
+ bl[21] br[21] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_24 
+ bl[22] br[22] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_25 
+ bl[23] br[23] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_26 
+ bl[24] br[24] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_27 
+ bl[25] br[25] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_28 
+ bl[26] br[26] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_29 
+ bl[27] br[27] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_30 
+ bl[28] br[28] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_31 
+ bl[29] br[29] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_32 
+ bl[30] br[30] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_33 
+ bl[31] br[31] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_34 
+ bl[32] br[32] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_35 
+ bl[33] br[33] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_36 
+ bl[34] br[34] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_37 
+ bl[35] br[35] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_38 
+ bl[36] br[36] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_39 
+ bl[37] br[37] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_40 
+ bl[38] br[38] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_41 
+ bl[39] br[39] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_42 
+ bl[40] br[40] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_43 
+ bl[41] br[41] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_44 
+ bl[42] br[42] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_45 
+ bl[43] br[43] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_46 
+ bl[44] br[44] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_47 
+ bl[45] br[45] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_48 
+ bl[46] br[46] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_49 
+ bl[47] br[47] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_50 
+ bl[48] br[48] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_51 
+ bl[49] br[49] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_52 
+ bl[50] br[50] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_53 
+ bl[51] br[51] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_54 
+ bl[52] br[52] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_55 
+ bl[53] br[53] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_56 
+ bl[54] br[54] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_57 
+ bl[55] br[55] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_58 
+ bl[56] br[56] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_59 
+ bl[57] br[57] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_60 
+ bl[58] br[58] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_61 
+ bl[59] br[59] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_62 
+ bl[60] br[60] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_63 
+ bl[61] br[61] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_64 
+ bl[62] br[62] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_65 
+ bl[63] br[63] vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_66 
+ vdd vdd vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_104_67 
+ vdd vdd vdd vss wl[102] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_0 
+ vdd vdd vss vdd vpb vnb wl[103] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_105_1 
+ rbl rbr vss vdd vpb vnb wl[103] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_105_2 
+ bl[0] br[0] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_3 
+ bl[1] br[1] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_4 
+ bl[2] br[2] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_5 
+ bl[3] br[3] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_6 
+ bl[4] br[4] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_7 
+ bl[5] br[5] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_8 
+ bl[6] br[6] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_9 
+ bl[7] br[7] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_10 
+ bl[8] br[8] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_11 
+ bl[9] br[9] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_12 
+ bl[10] br[10] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_13 
+ bl[11] br[11] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_14 
+ bl[12] br[12] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_15 
+ bl[13] br[13] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_16 
+ bl[14] br[14] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_17 
+ bl[15] br[15] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_18 
+ bl[16] br[16] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_19 
+ bl[17] br[17] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_20 
+ bl[18] br[18] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_21 
+ bl[19] br[19] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_22 
+ bl[20] br[20] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_23 
+ bl[21] br[21] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_24 
+ bl[22] br[22] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_25 
+ bl[23] br[23] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_26 
+ bl[24] br[24] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_27 
+ bl[25] br[25] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_28 
+ bl[26] br[26] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_29 
+ bl[27] br[27] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_30 
+ bl[28] br[28] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_31 
+ bl[29] br[29] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_32 
+ bl[30] br[30] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_33 
+ bl[31] br[31] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_34 
+ bl[32] br[32] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_35 
+ bl[33] br[33] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_36 
+ bl[34] br[34] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_37 
+ bl[35] br[35] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_38 
+ bl[36] br[36] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_39 
+ bl[37] br[37] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_40 
+ bl[38] br[38] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_41 
+ bl[39] br[39] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_42 
+ bl[40] br[40] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_43 
+ bl[41] br[41] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_44 
+ bl[42] br[42] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_45 
+ bl[43] br[43] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_46 
+ bl[44] br[44] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_47 
+ bl[45] br[45] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_48 
+ bl[46] br[46] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_49 
+ bl[47] br[47] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_50 
+ bl[48] br[48] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_51 
+ bl[49] br[49] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_52 
+ bl[50] br[50] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_53 
+ bl[51] br[51] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_54 
+ bl[52] br[52] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_55 
+ bl[53] br[53] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_56 
+ bl[54] br[54] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_57 
+ bl[55] br[55] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_58 
+ bl[56] br[56] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_59 
+ bl[57] br[57] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_60 
+ bl[58] br[58] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_61 
+ bl[59] br[59] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_62 
+ bl[60] br[60] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_63 
+ bl[61] br[61] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_64 
+ bl[62] br[62] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_65 
+ bl[63] br[63] vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_66 
+ vdd vdd vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_105_67 
+ vdd vdd vdd vss wl[103] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_0 
+ vdd vdd vss vdd vpb vnb wl[104] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_106_1 
+ rbl rbr vss vdd vpb vnb wl[104] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_106_2 
+ bl[0] br[0] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_3 
+ bl[1] br[1] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_4 
+ bl[2] br[2] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_5 
+ bl[3] br[3] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_6 
+ bl[4] br[4] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_7 
+ bl[5] br[5] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_8 
+ bl[6] br[6] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_9 
+ bl[7] br[7] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_10 
+ bl[8] br[8] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_11 
+ bl[9] br[9] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_12 
+ bl[10] br[10] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_13 
+ bl[11] br[11] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_14 
+ bl[12] br[12] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_15 
+ bl[13] br[13] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_16 
+ bl[14] br[14] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_17 
+ bl[15] br[15] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_18 
+ bl[16] br[16] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_19 
+ bl[17] br[17] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_20 
+ bl[18] br[18] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_21 
+ bl[19] br[19] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_22 
+ bl[20] br[20] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_23 
+ bl[21] br[21] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_24 
+ bl[22] br[22] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_25 
+ bl[23] br[23] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_26 
+ bl[24] br[24] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_27 
+ bl[25] br[25] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_28 
+ bl[26] br[26] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_29 
+ bl[27] br[27] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_30 
+ bl[28] br[28] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_31 
+ bl[29] br[29] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_32 
+ bl[30] br[30] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_33 
+ bl[31] br[31] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_34 
+ bl[32] br[32] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_35 
+ bl[33] br[33] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_36 
+ bl[34] br[34] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_37 
+ bl[35] br[35] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_38 
+ bl[36] br[36] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_39 
+ bl[37] br[37] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_40 
+ bl[38] br[38] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_41 
+ bl[39] br[39] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_42 
+ bl[40] br[40] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_43 
+ bl[41] br[41] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_44 
+ bl[42] br[42] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_45 
+ bl[43] br[43] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_46 
+ bl[44] br[44] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_47 
+ bl[45] br[45] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_48 
+ bl[46] br[46] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_49 
+ bl[47] br[47] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_50 
+ bl[48] br[48] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_51 
+ bl[49] br[49] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_52 
+ bl[50] br[50] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_53 
+ bl[51] br[51] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_54 
+ bl[52] br[52] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_55 
+ bl[53] br[53] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_56 
+ bl[54] br[54] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_57 
+ bl[55] br[55] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_58 
+ bl[56] br[56] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_59 
+ bl[57] br[57] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_60 
+ bl[58] br[58] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_61 
+ bl[59] br[59] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_62 
+ bl[60] br[60] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_63 
+ bl[61] br[61] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_64 
+ bl[62] br[62] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_65 
+ bl[63] br[63] vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_66 
+ vdd vdd vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_106_67 
+ vdd vdd vdd vss wl[104] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_0 
+ vdd vdd vss vdd vpb vnb wl[105] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_107_1 
+ rbl rbr vss vdd vpb vnb wl[105] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_107_2 
+ bl[0] br[0] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_3 
+ bl[1] br[1] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_4 
+ bl[2] br[2] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_5 
+ bl[3] br[3] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_6 
+ bl[4] br[4] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_7 
+ bl[5] br[5] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_8 
+ bl[6] br[6] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_9 
+ bl[7] br[7] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_10 
+ bl[8] br[8] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_11 
+ bl[9] br[9] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_12 
+ bl[10] br[10] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_13 
+ bl[11] br[11] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_14 
+ bl[12] br[12] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_15 
+ bl[13] br[13] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_16 
+ bl[14] br[14] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_17 
+ bl[15] br[15] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_18 
+ bl[16] br[16] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_19 
+ bl[17] br[17] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_20 
+ bl[18] br[18] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_21 
+ bl[19] br[19] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_22 
+ bl[20] br[20] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_23 
+ bl[21] br[21] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_24 
+ bl[22] br[22] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_25 
+ bl[23] br[23] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_26 
+ bl[24] br[24] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_27 
+ bl[25] br[25] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_28 
+ bl[26] br[26] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_29 
+ bl[27] br[27] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_30 
+ bl[28] br[28] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_31 
+ bl[29] br[29] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_32 
+ bl[30] br[30] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_33 
+ bl[31] br[31] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_34 
+ bl[32] br[32] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_35 
+ bl[33] br[33] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_36 
+ bl[34] br[34] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_37 
+ bl[35] br[35] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_38 
+ bl[36] br[36] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_39 
+ bl[37] br[37] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_40 
+ bl[38] br[38] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_41 
+ bl[39] br[39] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_42 
+ bl[40] br[40] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_43 
+ bl[41] br[41] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_44 
+ bl[42] br[42] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_45 
+ bl[43] br[43] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_46 
+ bl[44] br[44] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_47 
+ bl[45] br[45] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_48 
+ bl[46] br[46] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_49 
+ bl[47] br[47] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_50 
+ bl[48] br[48] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_51 
+ bl[49] br[49] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_52 
+ bl[50] br[50] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_53 
+ bl[51] br[51] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_54 
+ bl[52] br[52] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_55 
+ bl[53] br[53] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_56 
+ bl[54] br[54] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_57 
+ bl[55] br[55] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_58 
+ bl[56] br[56] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_59 
+ bl[57] br[57] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_60 
+ bl[58] br[58] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_61 
+ bl[59] br[59] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_62 
+ bl[60] br[60] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_63 
+ bl[61] br[61] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_64 
+ bl[62] br[62] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_65 
+ bl[63] br[63] vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_66 
+ vdd vdd vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_107_67 
+ vdd vdd vdd vss wl[105] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_0 
+ vdd vdd vss vdd vpb vnb wl[106] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_108_1 
+ rbl rbr vss vdd vpb vnb wl[106] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_108_2 
+ bl[0] br[0] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_3 
+ bl[1] br[1] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_4 
+ bl[2] br[2] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_5 
+ bl[3] br[3] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_6 
+ bl[4] br[4] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_7 
+ bl[5] br[5] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_8 
+ bl[6] br[6] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_9 
+ bl[7] br[7] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_10 
+ bl[8] br[8] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_11 
+ bl[9] br[9] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_12 
+ bl[10] br[10] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_13 
+ bl[11] br[11] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_14 
+ bl[12] br[12] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_15 
+ bl[13] br[13] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_16 
+ bl[14] br[14] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_17 
+ bl[15] br[15] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_18 
+ bl[16] br[16] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_19 
+ bl[17] br[17] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_20 
+ bl[18] br[18] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_21 
+ bl[19] br[19] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_22 
+ bl[20] br[20] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_23 
+ bl[21] br[21] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_24 
+ bl[22] br[22] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_25 
+ bl[23] br[23] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_26 
+ bl[24] br[24] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_27 
+ bl[25] br[25] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_28 
+ bl[26] br[26] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_29 
+ bl[27] br[27] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_30 
+ bl[28] br[28] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_31 
+ bl[29] br[29] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_32 
+ bl[30] br[30] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_33 
+ bl[31] br[31] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_34 
+ bl[32] br[32] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_35 
+ bl[33] br[33] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_36 
+ bl[34] br[34] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_37 
+ bl[35] br[35] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_38 
+ bl[36] br[36] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_39 
+ bl[37] br[37] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_40 
+ bl[38] br[38] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_41 
+ bl[39] br[39] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_42 
+ bl[40] br[40] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_43 
+ bl[41] br[41] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_44 
+ bl[42] br[42] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_45 
+ bl[43] br[43] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_46 
+ bl[44] br[44] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_47 
+ bl[45] br[45] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_48 
+ bl[46] br[46] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_49 
+ bl[47] br[47] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_50 
+ bl[48] br[48] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_51 
+ bl[49] br[49] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_52 
+ bl[50] br[50] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_53 
+ bl[51] br[51] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_54 
+ bl[52] br[52] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_55 
+ bl[53] br[53] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_56 
+ bl[54] br[54] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_57 
+ bl[55] br[55] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_58 
+ bl[56] br[56] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_59 
+ bl[57] br[57] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_60 
+ bl[58] br[58] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_61 
+ bl[59] br[59] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_62 
+ bl[60] br[60] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_63 
+ bl[61] br[61] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_64 
+ bl[62] br[62] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_65 
+ bl[63] br[63] vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_66 
+ vdd vdd vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_108_67 
+ vdd vdd vdd vss wl[106] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_0 
+ vdd vdd vss vdd vpb vnb wl[107] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_109_1 
+ rbl rbr vss vdd vpb vnb wl[107] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_109_2 
+ bl[0] br[0] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_3 
+ bl[1] br[1] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_4 
+ bl[2] br[2] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_5 
+ bl[3] br[3] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_6 
+ bl[4] br[4] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_7 
+ bl[5] br[5] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_8 
+ bl[6] br[6] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_9 
+ bl[7] br[7] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_10 
+ bl[8] br[8] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_11 
+ bl[9] br[9] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_12 
+ bl[10] br[10] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_13 
+ bl[11] br[11] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_14 
+ bl[12] br[12] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_15 
+ bl[13] br[13] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_16 
+ bl[14] br[14] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_17 
+ bl[15] br[15] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_18 
+ bl[16] br[16] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_19 
+ bl[17] br[17] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_20 
+ bl[18] br[18] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_21 
+ bl[19] br[19] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_22 
+ bl[20] br[20] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_23 
+ bl[21] br[21] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_24 
+ bl[22] br[22] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_25 
+ bl[23] br[23] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_26 
+ bl[24] br[24] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_27 
+ bl[25] br[25] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_28 
+ bl[26] br[26] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_29 
+ bl[27] br[27] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_30 
+ bl[28] br[28] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_31 
+ bl[29] br[29] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_32 
+ bl[30] br[30] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_33 
+ bl[31] br[31] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_34 
+ bl[32] br[32] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_35 
+ bl[33] br[33] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_36 
+ bl[34] br[34] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_37 
+ bl[35] br[35] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_38 
+ bl[36] br[36] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_39 
+ bl[37] br[37] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_40 
+ bl[38] br[38] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_41 
+ bl[39] br[39] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_42 
+ bl[40] br[40] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_43 
+ bl[41] br[41] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_44 
+ bl[42] br[42] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_45 
+ bl[43] br[43] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_46 
+ bl[44] br[44] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_47 
+ bl[45] br[45] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_48 
+ bl[46] br[46] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_49 
+ bl[47] br[47] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_50 
+ bl[48] br[48] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_51 
+ bl[49] br[49] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_52 
+ bl[50] br[50] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_53 
+ bl[51] br[51] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_54 
+ bl[52] br[52] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_55 
+ bl[53] br[53] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_56 
+ bl[54] br[54] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_57 
+ bl[55] br[55] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_58 
+ bl[56] br[56] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_59 
+ bl[57] br[57] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_60 
+ bl[58] br[58] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_61 
+ bl[59] br[59] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_62 
+ bl[60] br[60] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_63 
+ bl[61] br[61] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_64 
+ bl[62] br[62] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_65 
+ bl[63] br[63] vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_66 
+ vdd vdd vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_109_67 
+ vdd vdd vdd vss wl[107] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_0 
+ vdd vdd vss vdd vpb vnb wl[108] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_110_1 
+ rbl rbr vss vdd vpb vnb wl[108] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_110_2 
+ bl[0] br[0] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_3 
+ bl[1] br[1] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_4 
+ bl[2] br[2] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_5 
+ bl[3] br[3] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_6 
+ bl[4] br[4] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_7 
+ bl[5] br[5] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_8 
+ bl[6] br[6] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_9 
+ bl[7] br[7] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_10 
+ bl[8] br[8] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_11 
+ bl[9] br[9] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_12 
+ bl[10] br[10] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_13 
+ bl[11] br[11] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_14 
+ bl[12] br[12] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_15 
+ bl[13] br[13] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_16 
+ bl[14] br[14] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_17 
+ bl[15] br[15] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_18 
+ bl[16] br[16] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_19 
+ bl[17] br[17] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_20 
+ bl[18] br[18] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_21 
+ bl[19] br[19] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_22 
+ bl[20] br[20] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_23 
+ bl[21] br[21] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_24 
+ bl[22] br[22] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_25 
+ bl[23] br[23] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_26 
+ bl[24] br[24] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_27 
+ bl[25] br[25] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_28 
+ bl[26] br[26] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_29 
+ bl[27] br[27] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_30 
+ bl[28] br[28] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_31 
+ bl[29] br[29] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_32 
+ bl[30] br[30] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_33 
+ bl[31] br[31] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_34 
+ bl[32] br[32] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_35 
+ bl[33] br[33] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_36 
+ bl[34] br[34] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_37 
+ bl[35] br[35] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_38 
+ bl[36] br[36] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_39 
+ bl[37] br[37] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_40 
+ bl[38] br[38] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_41 
+ bl[39] br[39] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_42 
+ bl[40] br[40] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_43 
+ bl[41] br[41] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_44 
+ bl[42] br[42] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_45 
+ bl[43] br[43] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_46 
+ bl[44] br[44] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_47 
+ bl[45] br[45] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_48 
+ bl[46] br[46] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_49 
+ bl[47] br[47] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_50 
+ bl[48] br[48] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_51 
+ bl[49] br[49] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_52 
+ bl[50] br[50] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_53 
+ bl[51] br[51] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_54 
+ bl[52] br[52] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_55 
+ bl[53] br[53] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_56 
+ bl[54] br[54] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_57 
+ bl[55] br[55] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_58 
+ bl[56] br[56] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_59 
+ bl[57] br[57] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_60 
+ bl[58] br[58] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_61 
+ bl[59] br[59] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_62 
+ bl[60] br[60] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_63 
+ bl[61] br[61] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_64 
+ bl[62] br[62] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_65 
+ bl[63] br[63] vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_66 
+ vdd vdd vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_110_67 
+ vdd vdd vdd vss wl[108] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_0 
+ vdd vdd vss vdd vpb vnb wl[109] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_111_1 
+ rbl rbr vss vdd vpb vnb wl[109] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_111_2 
+ bl[0] br[0] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_3 
+ bl[1] br[1] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_4 
+ bl[2] br[2] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_5 
+ bl[3] br[3] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_6 
+ bl[4] br[4] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_7 
+ bl[5] br[5] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_8 
+ bl[6] br[6] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_9 
+ bl[7] br[7] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_10 
+ bl[8] br[8] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_11 
+ bl[9] br[9] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_12 
+ bl[10] br[10] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_13 
+ bl[11] br[11] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_14 
+ bl[12] br[12] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_15 
+ bl[13] br[13] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_16 
+ bl[14] br[14] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_17 
+ bl[15] br[15] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_18 
+ bl[16] br[16] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_19 
+ bl[17] br[17] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_20 
+ bl[18] br[18] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_21 
+ bl[19] br[19] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_22 
+ bl[20] br[20] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_23 
+ bl[21] br[21] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_24 
+ bl[22] br[22] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_25 
+ bl[23] br[23] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_26 
+ bl[24] br[24] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_27 
+ bl[25] br[25] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_28 
+ bl[26] br[26] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_29 
+ bl[27] br[27] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_30 
+ bl[28] br[28] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_31 
+ bl[29] br[29] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_32 
+ bl[30] br[30] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_33 
+ bl[31] br[31] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_34 
+ bl[32] br[32] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_35 
+ bl[33] br[33] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_36 
+ bl[34] br[34] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_37 
+ bl[35] br[35] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_38 
+ bl[36] br[36] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_39 
+ bl[37] br[37] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_40 
+ bl[38] br[38] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_41 
+ bl[39] br[39] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_42 
+ bl[40] br[40] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_43 
+ bl[41] br[41] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_44 
+ bl[42] br[42] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_45 
+ bl[43] br[43] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_46 
+ bl[44] br[44] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_47 
+ bl[45] br[45] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_48 
+ bl[46] br[46] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_49 
+ bl[47] br[47] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_50 
+ bl[48] br[48] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_51 
+ bl[49] br[49] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_52 
+ bl[50] br[50] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_53 
+ bl[51] br[51] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_54 
+ bl[52] br[52] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_55 
+ bl[53] br[53] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_56 
+ bl[54] br[54] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_57 
+ bl[55] br[55] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_58 
+ bl[56] br[56] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_59 
+ bl[57] br[57] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_60 
+ bl[58] br[58] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_61 
+ bl[59] br[59] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_62 
+ bl[60] br[60] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_63 
+ bl[61] br[61] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_64 
+ bl[62] br[62] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_65 
+ bl[63] br[63] vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_66 
+ vdd vdd vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_111_67 
+ vdd vdd vdd vss wl[109] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_0 
+ vdd vdd vss vdd vpb vnb wl[110] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_112_1 
+ rbl rbr vss vdd vpb vnb wl[110] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_112_2 
+ bl[0] br[0] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_3 
+ bl[1] br[1] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_4 
+ bl[2] br[2] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_5 
+ bl[3] br[3] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_6 
+ bl[4] br[4] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_7 
+ bl[5] br[5] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_8 
+ bl[6] br[6] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_9 
+ bl[7] br[7] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_10 
+ bl[8] br[8] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_11 
+ bl[9] br[9] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_12 
+ bl[10] br[10] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_13 
+ bl[11] br[11] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_14 
+ bl[12] br[12] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_15 
+ bl[13] br[13] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_16 
+ bl[14] br[14] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_17 
+ bl[15] br[15] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_18 
+ bl[16] br[16] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_19 
+ bl[17] br[17] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_20 
+ bl[18] br[18] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_21 
+ bl[19] br[19] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_22 
+ bl[20] br[20] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_23 
+ bl[21] br[21] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_24 
+ bl[22] br[22] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_25 
+ bl[23] br[23] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_26 
+ bl[24] br[24] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_27 
+ bl[25] br[25] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_28 
+ bl[26] br[26] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_29 
+ bl[27] br[27] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_30 
+ bl[28] br[28] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_31 
+ bl[29] br[29] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_32 
+ bl[30] br[30] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_33 
+ bl[31] br[31] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_34 
+ bl[32] br[32] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_35 
+ bl[33] br[33] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_36 
+ bl[34] br[34] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_37 
+ bl[35] br[35] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_38 
+ bl[36] br[36] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_39 
+ bl[37] br[37] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_40 
+ bl[38] br[38] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_41 
+ bl[39] br[39] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_42 
+ bl[40] br[40] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_43 
+ bl[41] br[41] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_44 
+ bl[42] br[42] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_45 
+ bl[43] br[43] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_46 
+ bl[44] br[44] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_47 
+ bl[45] br[45] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_48 
+ bl[46] br[46] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_49 
+ bl[47] br[47] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_50 
+ bl[48] br[48] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_51 
+ bl[49] br[49] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_52 
+ bl[50] br[50] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_53 
+ bl[51] br[51] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_54 
+ bl[52] br[52] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_55 
+ bl[53] br[53] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_56 
+ bl[54] br[54] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_57 
+ bl[55] br[55] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_58 
+ bl[56] br[56] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_59 
+ bl[57] br[57] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_60 
+ bl[58] br[58] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_61 
+ bl[59] br[59] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_62 
+ bl[60] br[60] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_63 
+ bl[61] br[61] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_64 
+ bl[62] br[62] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_65 
+ bl[63] br[63] vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_66 
+ vdd vdd vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_112_67 
+ vdd vdd vdd vss wl[110] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_0 
+ vdd vdd vss vdd vpb vnb wl[111] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_113_1 
+ rbl rbr vss vdd vpb vnb wl[111] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_113_2 
+ bl[0] br[0] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_3 
+ bl[1] br[1] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_4 
+ bl[2] br[2] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_5 
+ bl[3] br[3] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_6 
+ bl[4] br[4] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_7 
+ bl[5] br[5] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_8 
+ bl[6] br[6] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_9 
+ bl[7] br[7] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_10 
+ bl[8] br[8] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_11 
+ bl[9] br[9] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_12 
+ bl[10] br[10] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_13 
+ bl[11] br[11] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_14 
+ bl[12] br[12] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_15 
+ bl[13] br[13] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_16 
+ bl[14] br[14] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_17 
+ bl[15] br[15] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_18 
+ bl[16] br[16] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_19 
+ bl[17] br[17] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_20 
+ bl[18] br[18] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_21 
+ bl[19] br[19] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_22 
+ bl[20] br[20] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_23 
+ bl[21] br[21] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_24 
+ bl[22] br[22] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_25 
+ bl[23] br[23] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_26 
+ bl[24] br[24] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_27 
+ bl[25] br[25] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_28 
+ bl[26] br[26] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_29 
+ bl[27] br[27] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_30 
+ bl[28] br[28] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_31 
+ bl[29] br[29] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_32 
+ bl[30] br[30] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_33 
+ bl[31] br[31] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_34 
+ bl[32] br[32] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_35 
+ bl[33] br[33] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_36 
+ bl[34] br[34] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_37 
+ bl[35] br[35] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_38 
+ bl[36] br[36] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_39 
+ bl[37] br[37] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_40 
+ bl[38] br[38] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_41 
+ bl[39] br[39] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_42 
+ bl[40] br[40] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_43 
+ bl[41] br[41] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_44 
+ bl[42] br[42] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_45 
+ bl[43] br[43] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_46 
+ bl[44] br[44] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_47 
+ bl[45] br[45] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_48 
+ bl[46] br[46] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_49 
+ bl[47] br[47] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_50 
+ bl[48] br[48] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_51 
+ bl[49] br[49] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_52 
+ bl[50] br[50] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_53 
+ bl[51] br[51] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_54 
+ bl[52] br[52] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_55 
+ bl[53] br[53] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_56 
+ bl[54] br[54] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_57 
+ bl[55] br[55] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_58 
+ bl[56] br[56] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_59 
+ bl[57] br[57] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_60 
+ bl[58] br[58] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_61 
+ bl[59] br[59] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_62 
+ bl[60] br[60] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_63 
+ bl[61] br[61] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_64 
+ bl[62] br[62] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_65 
+ bl[63] br[63] vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_66 
+ vdd vdd vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_113_67 
+ vdd vdd vdd vss wl[111] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_0 
+ vdd vdd vss vdd vpb vnb wl[112] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_114_1 
+ rbl rbr vss vdd vpb vnb wl[112] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_114_2 
+ bl[0] br[0] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_3 
+ bl[1] br[1] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_4 
+ bl[2] br[2] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_5 
+ bl[3] br[3] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_6 
+ bl[4] br[4] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_7 
+ bl[5] br[5] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_8 
+ bl[6] br[6] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_9 
+ bl[7] br[7] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_10 
+ bl[8] br[8] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_11 
+ bl[9] br[9] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_12 
+ bl[10] br[10] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_13 
+ bl[11] br[11] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_14 
+ bl[12] br[12] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_15 
+ bl[13] br[13] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_16 
+ bl[14] br[14] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_17 
+ bl[15] br[15] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_18 
+ bl[16] br[16] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_19 
+ bl[17] br[17] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_20 
+ bl[18] br[18] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_21 
+ bl[19] br[19] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_22 
+ bl[20] br[20] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_23 
+ bl[21] br[21] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_24 
+ bl[22] br[22] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_25 
+ bl[23] br[23] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_26 
+ bl[24] br[24] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_27 
+ bl[25] br[25] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_28 
+ bl[26] br[26] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_29 
+ bl[27] br[27] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_30 
+ bl[28] br[28] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_31 
+ bl[29] br[29] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_32 
+ bl[30] br[30] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_33 
+ bl[31] br[31] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_34 
+ bl[32] br[32] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_35 
+ bl[33] br[33] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_36 
+ bl[34] br[34] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_37 
+ bl[35] br[35] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_38 
+ bl[36] br[36] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_39 
+ bl[37] br[37] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_40 
+ bl[38] br[38] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_41 
+ bl[39] br[39] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_42 
+ bl[40] br[40] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_43 
+ bl[41] br[41] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_44 
+ bl[42] br[42] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_45 
+ bl[43] br[43] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_46 
+ bl[44] br[44] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_47 
+ bl[45] br[45] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_48 
+ bl[46] br[46] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_49 
+ bl[47] br[47] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_50 
+ bl[48] br[48] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_51 
+ bl[49] br[49] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_52 
+ bl[50] br[50] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_53 
+ bl[51] br[51] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_54 
+ bl[52] br[52] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_55 
+ bl[53] br[53] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_56 
+ bl[54] br[54] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_57 
+ bl[55] br[55] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_58 
+ bl[56] br[56] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_59 
+ bl[57] br[57] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_60 
+ bl[58] br[58] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_61 
+ bl[59] br[59] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_62 
+ bl[60] br[60] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_63 
+ bl[61] br[61] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_64 
+ bl[62] br[62] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_65 
+ bl[63] br[63] vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_66 
+ vdd vdd vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_114_67 
+ vdd vdd vdd vss wl[112] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_0 
+ vdd vdd vss vdd vpb vnb wl[113] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_115_1 
+ rbl rbr vss vdd vpb vnb wl[113] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_115_2 
+ bl[0] br[0] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_3 
+ bl[1] br[1] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_4 
+ bl[2] br[2] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_5 
+ bl[3] br[3] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_6 
+ bl[4] br[4] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_7 
+ bl[5] br[5] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_8 
+ bl[6] br[6] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_9 
+ bl[7] br[7] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_10 
+ bl[8] br[8] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_11 
+ bl[9] br[9] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_12 
+ bl[10] br[10] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_13 
+ bl[11] br[11] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_14 
+ bl[12] br[12] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_15 
+ bl[13] br[13] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_16 
+ bl[14] br[14] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_17 
+ bl[15] br[15] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_18 
+ bl[16] br[16] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_19 
+ bl[17] br[17] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_20 
+ bl[18] br[18] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_21 
+ bl[19] br[19] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_22 
+ bl[20] br[20] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_23 
+ bl[21] br[21] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_24 
+ bl[22] br[22] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_25 
+ bl[23] br[23] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_26 
+ bl[24] br[24] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_27 
+ bl[25] br[25] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_28 
+ bl[26] br[26] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_29 
+ bl[27] br[27] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_30 
+ bl[28] br[28] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_31 
+ bl[29] br[29] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_32 
+ bl[30] br[30] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_33 
+ bl[31] br[31] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_34 
+ bl[32] br[32] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_35 
+ bl[33] br[33] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_36 
+ bl[34] br[34] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_37 
+ bl[35] br[35] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_38 
+ bl[36] br[36] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_39 
+ bl[37] br[37] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_40 
+ bl[38] br[38] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_41 
+ bl[39] br[39] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_42 
+ bl[40] br[40] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_43 
+ bl[41] br[41] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_44 
+ bl[42] br[42] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_45 
+ bl[43] br[43] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_46 
+ bl[44] br[44] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_47 
+ bl[45] br[45] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_48 
+ bl[46] br[46] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_49 
+ bl[47] br[47] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_50 
+ bl[48] br[48] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_51 
+ bl[49] br[49] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_52 
+ bl[50] br[50] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_53 
+ bl[51] br[51] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_54 
+ bl[52] br[52] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_55 
+ bl[53] br[53] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_56 
+ bl[54] br[54] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_57 
+ bl[55] br[55] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_58 
+ bl[56] br[56] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_59 
+ bl[57] br[57] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_60 
+ bl[58] br[58] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_61 
+ bl[59] br[59] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_62 
+ bl[60] br[60] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_63 
+ bl[61] br[61] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_64 
+ bl[62] br[62] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_65 
+ bl[63] br[63] vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_66 
+ vdd vdd vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_115_67 
+ vdd vdd vdd vss wl[113] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_0 
+ vdd vdd vss vdd vpb vnb wl[114] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_116_1 
+ rbl rbr vss vdd vpb vnb wl[114] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_116_2 
+ bl[0] br[0] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_3 
+ bl[1] br[1] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_4 
+ bl[2] br[2] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_5 
+ bl[3] br[3] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_6 
+ bl[4] br[4] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_7 
+ bl[5] br[5] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_8 
+ bl[6] br[6] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_9 
+ bl[7] br[7] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_10 
+ bl[8] br[8] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_11 
+ bl[9] br[9] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_12 
+ bl[10] br[10] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_13 
+ bl[11] br[11] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_14 
+ bl[12] br[12] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_15 
+ bl[13] br[13] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_16 
+ bl[14] br[14] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_17 
+ bl[15] br[15] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_18 
+ bl[16] br[16] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_19 
+ bl[17] br[17] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_20 
+ bl[18] br[18] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_21 
+ bl[19] br[19] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_22 
+ bl[20] br[20] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_23 
+ bl[21] br[21] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_24 
+ bl[22] br[22] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_25 
+ bl[23] br[23] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_26 
+ bl[24] br[24] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_27 
+ bl[25] br[25] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_28 
+ bl[26] br[26] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_29 
+ bl[27] br[27] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_30 
+ bl[28] br[28] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_31 
+ bl[29] br[29] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_32 
+ bl[30] br[30] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_33 
+ bl[31] br[31] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_34 
+ bl[32] br[32] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_35 
+ bl[33] br[33] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_36 
+ bl[34] br[34] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_37 
+ bl[35] br[35] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_38 
+ bl[36] br[36] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_39 
+ bl[37] br[37] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_40 
+ bl[38] br[38] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_41 
+ bl[39] br[39] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_42 
+ bl[40] br[40] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_43 
+ bl[41] br[41] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_44 
+ bl[42] br[42] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_45 
+ bl[43] br[43] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_46 
+ bl[44] br[44] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_47 
+ bl[45] br[45] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_48 
+ bl[46] br[46] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_49 
+ bl[47] br[47] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_50 
+ bl[48] br[48] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_51 
+ bl[49] br[49] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_52 
+ bl[50] br[50] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_53 
+ bl[51] br[51] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_54 
+ bl[52] br[52] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_55 
+ bl[53] br[53] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_56 
+ bl[54] br[54] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_57 
+ bl[55] br[55] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_58 
+ bl[56] br[56] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_59 
+ bl[57] br[57] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_60 
+ bl[58] br[58] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_61 
+ bl[59] br[59] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_62 
+ bl[60] br[60] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_63 
+ bl[61] br[61] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_64 
+ bl[62] br[62] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_65 
+ bl[63] br[63] vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_66 
+ vdd vdd vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_116_67 
+ vdd vdd vdd vss wl[114] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_0 
+ vdd vdd vss vdd vpb vnb wl[115] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_117_1 
+ rbl rbr vss vdd vpb vnb wl[115] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_117_2 
+ bl[0] br[0] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_3 
+ bl[1] br[1] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_4 
+ bl[2] br[2] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_5 
+ bl[3] br[3] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_6 
+ bl[4] br[4] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_7 
+ bl[5] br[5] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_8 
+ bl[6] br[6] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_9 
+ bl[7] br[7] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_10 
+ bl[8] br[8] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_11 
+ bl[9] br[9] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_12 
+ bl[10] br[10] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_13 
+ bl[11] br[11] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_14 
+ bl[12] br[12] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_15 
+ bl[13] br[13] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_16 
+ bl[14] br[14] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_17 
+ bl[15] br[15] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_18 
+ bl[16] br[16] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_19 
+ bl[17] br[17] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_20 
+ bl[18] br[18] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_21 
+ bl[19] br[19] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_22 
+ bl[20] br[20] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_23 
+ bl[21] br[21] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_24 
+ bl[22] br[22] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_25 
+ bl[23] br[23] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_26 
+ bl[24] br[24] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_27 
+ bl[25] br[25] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_28 
+ bl[26] br[26] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_29 
+ bl[27] br[27] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_30 
+ bl[28] br[28] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_31 
+ bl[29] br[29] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_32 
+ bl[30] br[30] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_33 
+ bl[31] br[31] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_34 
+ bl[32] br[32] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_35 
+ bl[33] br[33] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_36 
+ bl[34] br[34] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_37 
+ bl[35] br[35] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_38 
+ bl[36] br[36] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_39 
+ bl[37] br[37] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_40 
+ bl[38] br[38] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_41 
+ bl[39] br[39] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_42 
+ bl[40] br[40] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_43 
+ bl[41] br[41] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_44 
+ bl[42] br[42] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_45 
+ bl[43] br[43] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_46 
+ bl[44] br[44] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_47 
+ bl[45] br[45] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_48 
+ bl[46] br[46] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_49 
+ bl[47] br[47] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_50 
+ bl[48] br[48] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_51 
+ bl[49] br[49] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_52 
+ bl[50] br[50] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_53 
+ bl[51] br[51] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_54 
+ bl[52] br[52] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_55 
+ bl[53] br[53] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_56 
+ bl[54] br[54] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_57 
+ bl[55] br[55] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_58 
+ bl[56] br[56] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_59 
+ bl[57] br[57] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_60 
+ bl[58] br[58] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_61 
+ bl[59] br[59] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_62 
+ bl[60] br[60] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_63 
+ bl[61] br[61] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_64 
+ bl[62] br[62] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_65 
+ bl[63] br[63] vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_66 
+ vdd vdd vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_117_67 
+ vdd vdd vdd vss wl[115] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_0 
+ vdd vdd vss vdd vpb vnb wl[116] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_118_1 
+ rbl rbr vss vdd vpb vnb wl[116] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_118_2 
+ bl[0] br[0] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_3 
+ bl[1] br[1] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_4 
+ bl[2] br[2] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_5 
+ bl[3] br[3] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_6 
+ bl[4] br[4] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_7 
+ bl[5] br[5] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_8 
+ bl[6] br[6] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_9 
+ bl[7] br[7] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_10 
+ bl[8] br[8] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_11 
+ bl[9] br[9] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_12 
+ bl[10] br[10] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_13 
+ bl[11] br[11] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_14 
+ bl[12] br[12] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_15 
+ bl[13] br[13] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_16 
+ bl[14] br[14] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_17 
+ bl[15] br[15] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_18 
+ bl[16] br[16] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_19 
+ bl[17] br[17] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_20 
+ bl[18] br[18] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_21 
+ bl[19] br[19] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_22 
+ bl[20] br[20] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_23 
+ bl[21] br[21] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_24 
+ bl[22] br[22] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_25 
+ bl[23] br[23] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_26 
+ bl[24] br[24] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_27 
+ bl[25] br[25] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_28 
+ bl[26] br[26] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_29 
+ bl[27] br[27] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_30 
+ bl[28] br[28] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_31 
+ bl[29] br[29] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_32 
+ bl[30] br[30] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_33 
+ bl[31] br[31] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_34 
+ bl[32] br[32] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_35 
+ bl[33] br[33] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_36 
+ bl[34] br[34] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_37 
+ bl[35] br[35] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_38 
+ bl[36] br[36] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_39 
+ bl[37] br[37] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_40 
+ bl[38] br[38] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_41 
+ bl[39] br[39] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_42 
+ bl[40] br[40] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_43 
+ bl[41] br[41] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_44 
+ bl[42] br[42] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_45 
+ bl[43] br[43] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_46 
+ bl[44] br[44] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_47 
+ bl[45] br[45] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_48 
+ bl[46] br[46] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_49 
+ bl[47] br[47] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_50 
+ bl[48] br[48] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_51 
+ bl[49] br[49] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_52 
+ bl[50] br[50] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_53 
+ bl[51] br[51] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_54 
+ bl[52] br[52] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_55 
+ bl[53] br[53] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_56 
+ bl[54] br[54] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_57 
+ bl[55] br[55] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_58 
+ bl[56] br[56] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_59 
+ bl[57] br[57] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_60 
+ bl[58] br[58] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_61 
+ bl[59] br[59] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_62 
+ bl[60] br[60] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_63 
+ bl[61] br[61] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_64 
+ bl[62] br[62] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_65 
+ bl[63] br[63] vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_66 
+ vdd vdd vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_118_67 
+ vdd vdd vdd vss wl[116] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_0 
+ vdd vdd vss vdd vpb vnb wl[117] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_119_1 
+ rbl rbr vss vdd vpb vnb wl[117] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_119_2 
+ bl[0] br[0] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_3 
+ bl[1] br[1] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_4 
+ bl[2] br[2] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_5 
+ bl[3] br[3] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_6 
+ bl[4] br[4] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_7 
+ bl[5] br[5] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_8 
+ bl[6] br[6] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_9 
+ bl[7] br[7] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_10 
+ bl[8] br[8] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_11 
+ bl[9] br[9] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_12 
+ bl[10] br[10] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_13 
+ bl[11] br[11] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_14 
+ bl[12] br[12] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_15 
+ bl[13] br[13] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_16 
+ bl[14] br[14] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_17 
+ bl[15] br[15] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_18 
+ bl[16] br[16] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_19 
+ bl[17] br[17] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_20 
+ bl[18] br[18] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_21 
+ bl[19] br[19] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_22 
+ bl[20] br[20] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_23 
+ bl[21] br[21] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_24 
+ bl[22] br[22] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_25 
+ bl[23] br[23] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_26 
+ bl[24] br[24] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_27 
+ bl[25] br[25] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_28 
+ bl[26] br[26] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_29 
+ bl[27] br[27] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_30 
+ bl[28] br[28] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_31 
+ bl[29] br[29] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_32 
+ bl[30] br[30] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_33 
+ bl[31] br[31] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_34 
+ bl[32] br[32] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_35 
+ bl[33] br[33] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_36 
+ bl[34] br[34] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_37 
+ bl[35] br[35] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_38 
+ bl[36] br[36] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_39 
+ bl[37] br[37] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_40 
+ bl[38] br[38] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_41 
+ bl[39] br[39] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_42 
+ bl[40] br[40] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_43 
+ bl[41] br[41] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_44 
+ bl[42] br[42] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_45 
+ bl[43] br[43] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_46 
+ bl[44] br[44] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_47 
+ bl[45] br[45] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_48 
+ bl[46] br[46] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_49 
+ bl[47] br[47] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_50 
+ bl[48] br[48] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_51 
+ bl[49] br[49] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_52 
+ bl[50] br[50] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_53 
+ bl[51] br[51] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_54 
+ bl[52] br[52] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_55 
+ bl[53] br[53] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_56 
+ bl[54] br[54] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_57 
+ bl[55] br[55] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_58 
+ bl[56] br[56] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_59 
+ bl[57] br[57] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_60 
+ bl[58] br[58] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_61 
+ bl[59] br[59] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_62 
+ bl[60] br[60] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_63 
+ bl[61] br[61] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_64 
+ bl[62] br[62] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_65 
+ bl[63] br[63] vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_66 
+ vdd vdd vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_119_67 
+ vdd vdd vdd vss wl[117] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_0 
+ vdd vdd vss vdd vpb vnb wl[118] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_120_1 
+ rbl rbr vss vdd vpb vnb wl[118] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_120_2 
+ bl[0] br[0] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_3 
+ bl[1] br[1] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_4 
+ bl[2] br[2] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_5 
+ bl[3] br[3] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_6 
+ bl[4] br[4] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_7 
+ bl[5] br[5] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_8 
+ bl[6] br[6] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_9 
+ bl[7] br[7] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_10 
+ bl[8] br[8] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_11 
+ bl[9] br[9] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_12 
+ bl[10] br[10] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_13 
+ bl[11] br[11] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_14 
+ bl[12] br[12] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_15 
+ bl[13] br[13] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_16 
+ bl[14] br[14] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_17 
+ bl[15] br[15] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_18 
+ bl[16] br[16] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_19 
+ bl[17] br[17] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_20 
+ bl[18] br[18] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_21 
+ bl[19] br[19] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_22 
+ bl[20] br[20] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_23 
+ bl[21] br[21] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_24 
+ bl[22] br[22] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_25 
+ bl[23] br[23] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_26 
+ bl[24] br[24] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_27 
+ bl[25] br[25] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_28 
+ bl[26] br[26] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_29 
+ bl[27] br[27] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_30 
+ bl[28] br[28] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_31 
+ bl[29] br[29] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_32 
+ bl[30] br[30] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_33 
+ bl[31] br[31] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_34 
+ bl[32] br[32] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_35 
+ bl[33] br[33] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_36 
+ bl[34] br[34] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_37 
+ bl[35] br[35] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_38 
+ bl[36] br[36] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_39 
+ bl[37] br[37] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_40 
+ bl[38] br[38] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_41 
+ bl[39] br[39] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_42 
+ bl[40] br[40] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_43 
+ bl[41] br[41] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_44 
+ bl[42] br[42] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_45 
+ bl[43] br[43] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_46 
+ bl[44] br[44] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_47 
+ bl[45] br[45] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_48 
+ bl[46] br[46] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_49 
+ bl[47] br[47] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_50 
+ bl[48] br[48] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_51 
+ bl[49] br[49] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_52 
+ bl[50] br[50] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_53 
+ bl[51] br[51] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_54 
+ bl[52] br[52] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_55 
+ bl[53] br[53] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_56 
+ bl[54] br[54] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_57 
+ bl[55] br[55] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_58 
+ bl[56] br[56] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_59 
+ bl[57] br[57] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_60 
+ bl[58] br[58] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_61 
+ bl[59] br[59] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_62 
+ bl[60] br[60] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_63 
+ bl[61] br[61] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_64 
+ bl[62] br[62] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_65 
+ bl[63] br[63] vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_66 
+ vdd vdd vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_120_67 
+ vdd vdd vdd vss wl[118] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_0 
+ vdd vdd vss vdd vpb vnb wl[119] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_121_1 
+ rbl rbr vss vdd vpb vnb wl[119] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_121_2 
+ bl[0] br[0] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_3 
+ bl[1] br[1] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_4 
+ bl[2] br[2] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_5 
+ bl[3] br[3] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_6 
+ bl[4] br[4] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_7 
+ bl[5] br[5] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_8 
+ bl[6] br[6] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_9 
+ bl[7] br[7] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_10 
+ bl[8] br[8] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_11 
+ bl[9] br[9] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_12 
+ bl[10] br[10] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_13 
+ bl[11] br[11] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_14 
+ bl[12] br[12] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_15 
+ bl[13] br[13] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_16 
+ bl[14] br[14] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_17 
+ bl[15] br[15] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_18 
+ bl[16] br[16] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_19 
+ bl[17] br[17] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_20 
+ bl[18] br[18] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_21 
+ bl[19] br[19] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_22 
+ bl[20] br[20] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_23 
+ bl[21] br[21] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_24 
+ bl[22] br[22] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_25 
+ bl[23] br[23] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_26 
+ bl[24] br[24] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_27 
+ bl[25] br[25] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_28 
+ bl[26] br[26] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_29 
+ bl[27] br[27] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_30 
+ bl[28] br[28] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_31 
+ bl[29] br[29] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_32 
+ bl[30] br[30] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_33 
+ bl[31] br[31] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_34 
+ bl[32] br[32] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_35 
+ bl[33] br[33] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_36 
+ bl[34] br[34] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_37 
+ bl[35] br[35] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_38 
+ bl[36] br[36] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_39 
+ bl[37] br[37] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_40 
+ bl[38] br[38] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_41 
+ bl[39] br[39] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_42 
+ bl[40] br[40] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_43 
+ bl[41] br[41] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_44 
+ bl[42] br[42] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_45 
+ bl[43] br[43] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_46 
+ bl[44] br[44] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_47 
+ bl[45] br[45] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_48 
+ bl[46] br[46] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_49 
+ bl[47] br[47] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_50 
+ bl[48] br[48] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_51 
+ bl[49] br[49] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_52 
+ bl[50] br[50] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_53 
+ bl[51] br[51] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_54 
+ bl[52] br[52] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_55 
+ bl[53] br[53] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_56 
+ bl[54] br[54] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_57 
+ bl[55] br[55] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_58 
+ bl[56] br[56] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_59 
+ bl[57] br[57] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_60 
+ bl[58] br[58] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_61 
+ bl[59] br[59] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_62 
+ bl[60] br[60] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_63 
+ bl[61] br[61] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_64 
+ bl[62] br[62] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_65 
+ bl[63] br[63] vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_66 
+ vdd vdd vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_121_67 
+ vdd vdd vdd vss wl[119] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_0 
+ vdd vdd vss vdd vpb vnb wl[120] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_122_1 
+ rbl rbr vss vdd vpb vnb wl[120] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_122_2 
+ bl[0] br[0] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_3 
+ bl[1] br[1] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_4 
+ bl[2] br[2] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_5 
+ bl[3] br[3] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_6 
+ bl[4] br[4] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_7 
+ bl[5] br[5] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_8 
+ bl[6] br[6] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_9 
+ bl[7] br[7] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_10 
+ bl[8] br[8] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_11 
+ bl[9] br[9] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_12 
+ bl[10] br[10] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_13 
+ bl[11] br[11] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_14 
+ bl[12] br[12] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_15 
+ bl[13] br[13] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_16 
+ bl[14] br[14] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_17 
+ bl[15] br[15] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_18 
+ bl[16] br[16] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_19 
+ bl[17] br[17] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_20 
+ bl[18] br[18] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_21 
+ bl[19] br[19] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_22 
+ bl[20] br[20] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_23 
+ bl[21] br[21] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_24 
+ bl[22] br[22] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_25 
+ bl[23] br[23] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_26 
+ bl[24] br[24] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_27 
+ bl[25] br[25] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_28 
+ bl[26] br[26] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_29 
+ bl[27] br[27] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_30 
+ bl[28] br[28] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_31 
+ bl[29] br[29] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_32 
+ bl[30] br[30] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_33 
+ bl[31] br[31] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_34 
+ bl[32] br[32] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_35 
+ bl[33] br[33] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_36 
+ bl[34] br[34] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_37 
+ bl[35] br[35] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_38 
+ bl[36] br[36] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_39 
+ bl[37] br[37] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_40 
+ bl[38] br[38] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_41 
+ bl[39] br[39] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_42 
+ bl[40] br[40] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_43 
+ bl[41] br[41] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_44 
+ bl[42] br[42] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_45 
+ bl[43] br[43] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_46 
+ bl[44] br[44] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_47 
+ bl[45] br[45] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_48 
+ bl[46] br[46] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_49 
+ bl[47] br[47] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_50 
+ bl[48] br[48] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_51 
+ bl[49] br[49] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_52 
+ bl[50] br[50] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_53 
+ bl[51] br[51] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_54 
+ bl[52] br[52] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_55 
+ bl[53] br[53] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_56 
+ bl[54] br[54] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_57 
+ bl[55] br[55] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_58 
+ bl[56] br[56] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_59 
+ bl[57] br[57] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_60 
+ bl[58] br[58] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_61 
+ bl[59] br[59] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_62 
+ bl[60] br[60] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_63 
+ bl[61] br[61] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_64 
+ bl[62] br[62] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_65 
+ bl[63] br[63] vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_66 
+ vdd vdd vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_122_67 
+ vdd vdd vdd vss wl[120] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_0 
+ vdd vdd vss vdd vpb vnb wl[121] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_123_1 
+ rbl rbr vss vdd vpb vnb wl[121] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_123_2 
+ bl[0] br[0] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_3 
+ bl[1] br[1] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_4 
+ bl[2] br[2] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_5 
+ bl[3] br[3] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_6 
+ bl[4] br[4] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_7 
+ bl[5] br[5] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_8 
+ bl[6] br[6] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_9 
+ bl[7] br[7] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_10 
+ bl[8] br[8] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_11 
+ bl[9] br[9] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_12 
+ bl[10] br[10] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_13 
+ bl[11] br[11] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_14 
+ bl[12] br[12] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_15 
+ bl[13] br[13] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_16 
+ bl[14] br[14] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_17 
+ bl[15] br[15] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_18 
+ bl[16] br[16] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_19 
+ bl[17] br[17] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_20 
+ bl[18] br[18] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_21 
+ bl[19] br[19] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_22 
+ bl[20] br[20] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_23 
+ bl[21] br[21] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_24 
+ bl[22] br[22] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_25 
+ bl[23] br[23] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_26 
+ bl[24] br[24] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_27 
+ bl[25] br[25] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_28 
+ bl[26] br[26] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_29 
+ bl[27] br[27] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_30 
+ bl[28] br[28] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_31 
+ bl[29] br[29] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_32 
+ bl[30] br[30] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_33 
+ bl[31] br[31] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_34 
+ bl[32] br[32] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_35 
+ bl[33] br[33] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_36 
+ bl[34] br[34] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_37 
+ bl[35] br[35] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_38 
+ bl[36] br[36] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_39 
+ bl[37] br[37] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_40 
+ bl[38] br[38] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_41 
+ bl[39] br[39] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_42 
+ bl[40] br[40] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_43 
+ bl[41] br[41] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_44 
+ bl[42] br[42] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_45 
+ bl[43] br[43] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_46 
+ bl[44] br[44] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_47 
+ bl[45] br[45] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_48 
+ bl[46] br[46] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_49 
+ bl[47] br[47] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_50 
+ bl[48] br[48] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_51 
+ bl[49] br[49] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_52 
+ bl[50] br[50] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_53 
+ bl[51] br[51] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_54 
+ bl[52] br[52] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_55 
+ bl[53] br[53] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_56 
+ bl[54] br[54] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_57 
+ bl[55] br[55] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_58 
+ bl[56] br[56] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_59 
+ bl[57] br[57] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_60 
+ bl[58] br[58] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_61 
+ bl[59] br[59] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_62 
+ bl[60] br[60] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_63 
+ bl[61] br[61] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_64 
+ bl[62] br[62] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_65 
+ bl[63] br[63] vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_66 
+ vdd vdd vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_123_67 
+ vdd vdd vdd vss wl[121] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_0 
+ vdd vdd vss vdd vpb vnb wl[122] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_124_1 
+ rbl rbr vss vdd vpb vnb wl[122] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_124_2 
+ bl[0] br[0] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_3 
+ bl[1] br[1] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_4 
+ bl[2] br[2] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_5 
+ bl[3] br[3] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_6 
+ bl[4] br[4] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_7 
+ bl[5] br[5] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_8 
+ bl[6] br[6] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_9 
+ bl[7] br[7] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_10 
+ bl[8] br[8] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_11 
+ bl[9] br[9] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_12 
+ bl[10] br[10] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_13 
+ bl[11] br[11] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_14 
+ bl[12] br[12] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_15 
+ bl[13] br[13] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_16 
+ bl[14] br[14] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_17 
+ bl[15] br[15] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_18 
+ bl[16] br[16] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_19 
+ bl[17] br[17] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_20 
+ bl[18] br[18] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_21 
+ bl[19] br[19] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_22 
+ bl[20] br[20] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_23 
+ bl[21] br[21] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_24 
+ bl[22] br[22] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_25 
+ bl[23] br[23] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_26 
+ bl[24] br[24] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_27 
+ bl[25] br[25] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_28 
+ bl[26] br[26] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_29 
+ bl[27] br[27] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_30 
+ bl[28] br[28] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_31 
+ bl[29] br[29] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_32 
+ bl[30] br[30] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_33 
+ bl[31] br[31] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_34 
+ bl[32] br[32] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_35 
+ bl[33] br[33] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_36 
+ bl[34] br[34] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_37 
+ bl[35] br[35] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_38 
+ bl[36] br[36] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_39 
+ bl[37] br[37] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_40 
+ bl[38] br[38] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_41 
+ bl[39] br[39] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_42 
+ bl[40] br[40] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_43 
+ bl[41] br[41] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_44 
+ bl[42] br[42] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_45 
+ bl[43] br[43] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_46 
+ bl[44] br[44] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_47 
+ bl[45] br[45] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_48 
+ bl[46] br[46] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_49 
+ bl[47] br[47] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_50 
+ bl[48] br[48] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_51 
+ bl[49] br[49] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_52 
+ bl[50] br[50] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_53 
+ bl[51] br[51] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_54 
+ bl[52] br[52] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_55 
+ bl[53] br[53] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_56 
+ bl[54] br[54] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_57 
+ bl[55] br[55] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_58 
+ bl[56] br[56] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_59 
+ bl[57] br[57] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_60 
+ bl[58] br[58] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_61 
+ bl[59] br[59] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_62 
+ bl[60] br[60] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_63 
+ bl[61] br[61] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_64 
+ bl[62] br[62] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_65 
+ bl[63] br[63] vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_66 
+ vdd vdd vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_124_67 
+ vdd vdd vdd vss wl[122] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_0 
+ vdd vdd vss vdd vpb vnb wl[123] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_125_1 
+ rbl rbr vss vdd vpb vnb wl[123] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_125_2 
+ bl[0] br[0] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_3 
+ bl[1] br[1] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_4 
+ bl[2] br[2] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_5 
+ bl[3] br[3] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_6 
+ bl[4] br[4] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_7 
+ bl[5] br[5] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_8 
+ bl[6] br[6] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_9 
+ bl[7] br[7] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_10 
+ bl[8] br[8] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_11 
+ bl[9] br[9] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_12 
+ bl[10] br[10] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_13 
+ bl[11] br[11] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_14 
+ bl[12] br[12] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_15 
+ bl[13] br[13] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_16 
+ bl[14] br[14] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_17 
+ bl[15] br[15] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_18 
+ bl[16] br[16] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_19 
+ bl[17] br[17] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_20 
+ bl[18] br[18] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_21 
+ bl[19] br[19] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_22 
+ bl[20] br[20] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_23 
+ bl[21] br[21] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_24 
+ bl[22] br[22] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_25 
+ bl[23] br[23] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_26 
+ bl[24] br[24] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_27 
+ bl[25] br[25] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_28 
+ bl[26] br[26] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_29 
+ bl[27] br[27] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_30 
+ bl[28] br[28] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_31 
+ bl[29] br[29] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_32 
+ bl[30] br[30] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_33 
+ bl[31] br[31] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_34 
+ bl[32] br[32] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_35 
+ bl[33] br[33] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_36 
+ bl[34] br[34] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_37 
+ bl[35] br[35] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_38 
+ bl[36] br[36] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_39 
+ bl[37] br[37] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_40 
+ bl[38] br[38] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_41 
+ bl[39] br[39] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_42 
+ bl[40] br[40] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_43 
+ bl[41] br[41] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_44 
+ bl[42] br[42] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_45 
+ bl[43] br[43] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_46 
+ bl[44] br[44] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_47 
+ bl[45] br[45] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_48 
+ bl[46] br[46] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_49 
+ bl[47] br[47] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_50 
+ bl[48] br[48] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_51 
+ bl[49] br[49] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_52 
+ bl[50] br[50] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_53 
+ bl[51] br[51] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_54 
+ bl[52] br[52] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_55 
+ bl[53] br[53] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_56 
+ bl[54] br[54] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_57 
+ bl[55] br[55] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_58 
+ bl[56] br[56] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_59 
+ bl[57] br[57] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_60 
+ bl[58] br[58] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_61 
+ bl[59] br[59] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_62 
+ bl[60] br[60] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_63 
+ bl[61] br[61] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_64 
+ bl[62] br[62] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_65 
+ bl[63] br[63] vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_66 
+ vdd vdd vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_125_67 
+ vdd vdd vdd vss wl[123] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_0 
+ vdd vdd vss vdd vpb vnb wl[124] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_126_1 
+ rbl rbr vss vdd vpb vnb wl[124] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_126_2 
+ bl[0] br[0] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_3 
+ bl[1] br[1] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_4 
+ bl[2] br[2] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_5 
+ bl[3] br[3] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_6 
+ bl[4] br[4] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_7 
+ bl[5] br[5] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_8 
+ bl[6] br[6] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_9 
+ bl[7] br[7] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_10 
+ bl[8] br[8] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_11 
+ bl[9] br[9] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_12 
+ bl[10] br[10] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_13 
+ bl[11] br[11] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_14 
+ bl[12] br[12] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_15 
+ bl[13] br[13] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_16 
+ bl[14] br[14] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_17 
+ bl[15] br[15] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_18 
+ bl[16] br[16] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_19 
+ bl[17] br[17] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_20 
+ bl[18] br[18] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_21 
+ bl[19] br[19] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_22 
+ bl[20] br[20] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_23 
+ bl[21] br[21] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_24 
+ bl[22] br[22] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_25 
+ bl[23] br[23] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_26 
+ bl[24] br[24] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_27 
+ bl[25] br[25] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_28 
+ bl[26] br[26] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_29 
+ bl[27] br[27] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_30 
+ bl[28] br[28] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_31 
+ bl[29] br[29] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_32 
+ bl[30] br[30] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_33 
+ bl[31] br[31] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_34 
+ bl[32] br[32] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_35 
+ bl[33] br[33] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_36 
+ bl[34] br[34] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_37 
+ bl[35] br[35] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_38 
+ bl[36] br[36] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_39 
+ bl[37] br[37] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_40 
+ bl[38] br[38] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_41 
+ bl[39] br[39] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_42 
+ bl[40] br[40] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_43 
+ bl[41] br[41] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_44 
+ bl[42] br[42] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_45 
+ bl[43] br[43] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_46 
+ bl[44] br[44] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_47 
+ bl[45] br[45] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_48 
+ bl[46] br[46] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_49 
+ bl[47] br[47] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_50 
+ bl[48] br[48] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_51 
+ bl[49] br[49] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_52 
+ bl[50] br[50] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_53 
+ bl[51] br[51] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_54 
+ bl[52] br[52] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_55 
+ bl[53] br[53] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_56 
+ bl[54] br[54] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_57 
+ bl[55] br[55] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_58 
+ bl[56] br[56] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_59 
+ bl[57] br[57] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_60 
+ bl[58] br[58] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_61 
+ bl[59] br[59] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_62 
+ bl[60] br[60] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_63 
+ bl[61] br[61] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_64 
+ bl[62] br[62] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_65 
+ bl[63] br[63] vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_66 
+ vdd vdd vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_126_67 
+ vdd vdd vdd vss wl[124] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_0 
+ vdd vdd vss vdd vpb vnb wl[125] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_127_1 
+ rbl rbr vss vdd vpb vnb wl[125] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_127_2 
+ bl[0] br[0] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_3 
+ bl[1] br[1] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_4 
+ bl[2] br[2] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_5 
+ bl[3] br[3] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_6 
+ bl[4] br[4] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_7 
+ bl[5] br[5] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_8 
+ bl[6] br[6] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_9 
+ bl[7] br[7] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_10 
+ bl[8] br[8] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_11 
+ bl[9] br[9] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_12 
+ bl[10] br[10] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_13 
+ bl[11] br[11] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_14 
+ bl[12] br[12] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_15 
+ bl[13] br[13] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_16 
+ bl[14] br[14] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_17 
+ bl[15] br[15] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_18 
+ bl[16] br[16] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_19 
+ bl[17] br[17] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_20 
+ bl[18] br[18] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_21 
+ bl[19] br[19] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_22 
+ bl[20] br[20] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_23 
+ bl[21] br[21] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_24 
+ bl[22] br[22] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_25 
+ bl[23] br[23] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_26 
+ bl[24] br[24] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_27 
+ bl[25] br[25] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_28 
+ bl[26] br[26] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_29 
+ bl[27] br[27] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_30 
+ bl[28] br[28] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_31 
+ bl[29] br[29] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_32 
+ bl[30] br[30] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_33 
+ bl[31] br[31] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_34 
+ bl[32] br[32] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_35 
+ bl[33] br[33] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_36 
+ bl[34] br[34] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_37 
+ bl[35] br[35] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_38 
+ bl[36] br[36] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_39 
+ bl[37] br[37] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_40 
+ bl[38] br[38] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_41 
+ bl[39] br[39] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_42 
+ bl[40] br[40] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_43 
+ bl[41] br[41] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_44 
+ bl[42] br[42] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_45 
+ bl[43] br[43] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_46 
+ bl[44] br[44] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_47 
+ bl[45] br[45] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_48 
+ bl[46] br[46] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_49 
+ bl[47] br[47] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_50 
+ bl[48] br[48] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_51 
+ bl[49] br[49] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_52 
+ bl[50] br[50] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_53 
+ bl[51] br[51] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_54 
+ bl[52] br[52] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_55 
+ bl[53] br[53] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_56 
+ bl[54] br[54] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_57 
+ bl[55] br[55] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_58 
+ bl[56] br[56] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_59 
+ bl[57] br[57] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_60 
+ bl[58] br[58] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_61 
+ bl[59] br[59] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_62 
+ bl[60] br[60] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_63 
+ bl[61] br[61] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_64 
+ bl[62] br[62] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_65 
+ bl[63] br[63] vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_66 
+ vdd vdd vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_127_67 
+ vdd vdd vdd vss wl[125] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_0 
+ vdd vdd vss vdd vpb vnb wl[126] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_128_1 
+ rbl rbr vss vdd vpb vnb wl[126] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_128_2 
+ bl[0] br[0] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_3 
+ bl[1] br[1] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_4 
+ bl[2] br[2] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_5 
+ bl[3] br[3] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_6 
+ bl[4] br[4] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_7 
+ bl[5] br[5] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_8 
+ bl[6] br[6] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_9 
+ bl[7] br[7] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_10 
+ bl[8] br[8] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_11 
+ bl[9] br[9] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_12 
+ bl[10] br[10] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_13 
+ bl[11] br[11] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_14 
+ bl[12] br[12] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_15 
+ bl[13] br[13] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_16 
+ bl[14] br[14] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_17 
+ bl[15] br[15] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_18 
+ bl[16] br[16] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_19 
+ bl[17] br[17] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_20 
+ bl[18] br[18] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_21 
+ bl[19] br[19] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_22 
+ bl[20] br[20] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_23 
+ bl[21] br[21] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_24 
+ bl[22] br[22] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_25 
+ bl[23] br[23] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_26 
+ bl[24] br[24] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_27 
+ bl[25] br[25] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_28 
+ bl[26] br[26] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_29 
+ bl[27] br[27] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_30 
+ bl[28] br[28] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_31 
+ bl[29] br[29] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_32 
+ bl[30] br[30] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_33 
+ bl[31] br[31] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_34 
+ bl[32] br[32] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_35 
+ bl[33] br[33] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_36 
+ bl[34] br[34] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_37 
+ bl[35] br[35] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_38 
+ bl[36] br[36] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_39 
+ bl[37] br[37] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_40 
+ bl[38] br[38] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_41 
+ bl[39] br[39] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_42 
+ bl[40] br[40] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_43 
+ bl[41] br[41] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_44 
+ bl[42] br[42] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_45 
+ bl[43] br[43] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_46 
+ bl[44] br[44] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_47 
+ bl[45] br[45] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_48 
+ bl[46] br[46] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_49 
+ bl[47] br[47] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_50 
+ bl[48] br[48] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_51 
+ bl[49] br[49] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_52 
+ bl[50] br[50] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_53 
+ bl[51] br[51] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_54 
+ bl[52] br[52] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_55 
+ bl[53] br[53] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_56 
+ bl[54] br[54] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_57 
+ bl[55] br[55] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_58 
+ bl[56] br[56] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_59 
+ bl[57] br[57] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_60 
+ bl[58] br[58] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_61 
+ bl[59] br[59] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_62 
+ bl[60] br[60] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_63 
+ bl[61] br[61] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_64 
+ bl[62] br[62] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_65 
+ bl[63] br[63] vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_66 
+ vdd vdd vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_128_67 
+ vdd vdd vdd vss wl[126] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_0 
+ vdd vdd vss vdd vpb vnb wl[127] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_129_1 
+ rbl rbr vss vdd vpb vnb wl[127] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_129_2 
+ bl[0] br[0] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_3 
+ bl[1] br[1] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_4 
+ bl[2] br[2] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_5 
+ bl[3] br[3] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_6 
+ bl[4] br[4] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_7 
+ bl[5] br[5] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_8 
+ bl[6] br[6] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_9 
+ bl[7] br[7] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_10 
+ bl[8] br[8] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_11 
+ bl[9] br[9] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_12 
+ bl[10] br[10] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_13 
+ bl[11] br[11] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_14 
+ bl[12] br[12] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_15 
+ bl[13] br[13] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_16 
+ bl[14] br[14] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_17 
+ bl[15] br[15] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_18 
+ bl[16] br[16] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_19 
+ bl[17] br[17] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_20 
+ bl[18] br[18] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_21 
+ bl[19] br[19] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_22 
+ bl[20] br[20] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_23 
+ bl[21] br[21] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_24 
+ bl[22] br[22] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_25 
+ bl[23] br[23] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_26 
+ bl[24] br[24] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_27 
+ bl[25] br[25] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_28 
+ bl[26] br[26] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_29 
+ bl[27] br[27] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_30 
+ bl[28] br[28] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_31 
+ bl[29] br[29] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_32 
+ bl[30] br[30] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_33 
+ bl[31] br[31] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_34 
+ bl[32] br[32] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_35 
+ bl[33] br[33] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_36 
+ bl[34] br[34] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_37 
+ bl[35] br[35] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_38 
+ bl[36] br[36] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_39 
+ bl[37] br[37] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_40 
+ bl[38] br[38] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_41 
+ bl[39] br[39] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_42 
+ bl[40] br[40] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_43 
+ bl[41] br[41] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_44 
+ bl[42] br[42] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_45 
+ bl[43] br[43] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_46 
+ bl[44] br[44] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_47 
+ bl[45] br[45] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_48 
+ bl[46] br[46] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_49 
+ bl[47] br[47] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_50 
+ bl[48] br[48] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_51 
+ bl[49] br[49] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_52 
+ bl[50] br[50] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_53 
+ bl[51] br[51] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_54 
+ bl[52] br[52] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_55 
+ bl[53] br[53] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_56 
+ bl[54] br[54] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_57 
+ bl[55] br[55] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_58 
+ bl[56] br[56] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_59 
+ bl[57] br[57] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_60 
+ bl[58] br[58] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_61 
+ bl[59] br[59] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_62 
+ bl[60] br[60] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_63 
+ bl[61] br[61] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_64 
+ bl[62] br[62] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_65 
+ bl[63] br[63] vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_66 
+ vdd vdd vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_129_67 
+ vdd vdd vdd vss wl[127] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_0 
+ vdd vdd vss vdd vpb vnb wl[128] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_130_1 
+ rbl rbr vss vdd vpb vnb wl[128] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_130_2 
+ bl[0] br[0] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_3 
+ bl[1] br[1] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_4 
+ bl[2] br[2] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_5 
+ bl[3] br[3] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_6 
+ bl[4] br[4] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_7 
+ bl[5] br[5] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_8 
+ bl[6] br[6] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_9 
+ bl[7] br[7] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_10 
+ bl[8] br[8] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_11 
+ bl[9] br[9] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_12 
+ bl[10] br[10] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_13 
+ bl[11] br[11] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_14 
+ bl[12] br[12] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_15 
+ bl[13] br[13] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_16 
+ bl[14] br[14] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_17 
+ bl[15] br[15] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_18 
+ bl[16] br[16] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_19 
+ bl[17] br[17] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_20 
+ bl[18] br[18] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_21 
+ bl[19] br[19] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_22 
+ bl[20] br[20] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_23 
+ bl[21] br[21] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_24 
+ bl[22] br[22] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_25 
+ bl[23] br[23] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_26 
+ bl[24] br[24] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_27 
+ bl[25] br[25] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_28 
+ bl[26] br[26] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_29 
+ bl[27] br[27] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_30 
+ bl[28] br[28] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_31 
+ bl[29] br[29] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_32 
+ bl[30] br[30] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_33 
+ bl[31] br[31] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_34 
+ bl[32] br[32] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_35 
+ bl[33] br[33] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_36 
+ bl[34] br[34] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_37 
+ bl[35] br[35] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_38 
+ bl[36] br[36] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_39 
+ bl[37] br[37] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_40 
+ bl[38] br[38] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_41 
+ bl[39] br[39] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_42 
+ bl[40] br[40] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_43 
+ bl[41] br[41] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_44 
+ bl[42] br[42] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_45 
+ bl[43] br[43] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_46 
+ bl[44] br[44] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_47 
+ bl[45] br[45] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_48 
+ bl[46] br[46] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_49 
+ bl[47] br[47] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_50 
+ bl[48] br[48] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_51 
+ bl[49] br[49] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_52 
+ bl[50] br[50] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_53 
+ bl[51] br[51] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_54 
+ bl[52] br[52] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_55 
+ bl[53] br[53] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_56 
+ bl[54] br[54] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_57 
+ bl[55] br[55] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_58 
+ bl[56] br[56] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_59 
+ bl[57] br[57] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_60 
+ bl[58] br[58] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_61 
+ bl[59] br[59] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_62 
+ bl[60] br[60] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_63 
+ bl[61] br[61] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_64 
+ bl[62] br[62] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_65 
+ bl[63] br[63] vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_66 
+ vdd vdd vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_130_67 
+ vdd vdd vdd vss wl[128] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_0 
+ vdd vdd vss vdd vpb vnb wl[129] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_131_1 
+ rbl rbr vss vdd vpb vnb wl[129] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_131_2 
+ bl[0] br[0] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_3 
+ bl[1] br[1] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_4 
+ bl[2] br[2] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_5 
+ bl[3] br[3] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_6 
+ bl[4] br[4] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_7 
+ bl[5] br[5] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_8 
+ bl[6] br[6] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_9 
+ bl[7] br[7] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_10 
+ bl[8] br[8] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_11 
+ bl[9] br[9] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_12 
+ bl[10] br[10] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_13 
+ bl[11] br[11] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_14 
+ bl[12] br[12] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_15 
+ bl[13] br[13] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_16 
+ bl[14] br[14] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_17 
+ bl[15] br[15] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_18 
+ bl[16] br[16] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_19 
+ bl[17] br[17] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_20 
+ bl[18] br[18] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_21 
+ bl[19] br[19] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_22 
+ bl[20] br[20] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_23 
+ bl[21] br[21] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_24 
+ bl[22] br[22] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_25 
+ bl[23] br[23] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_26 
+ bl[24] br[24] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_27 
+ bl[25] br[25] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_28 
+ bl[26] br[26] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_29 
+ bl[27] br[27] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_30 
+ bl[28] br[28] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_31 
+ bl[29] br[29] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_32 
+ bl[30] br[30] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_33 
+ bl[31] br[31] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_34 
+ bl[32] br[32] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_35 
+ bl[33] br[33] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_36 
+ bl[34] br[34] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_37 
+ bl[35] br[35] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_38 
+ bl[36] br[36] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_39 
+ bl[37] br[37] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_40 
+ bl[38] br[38] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_41 
+ bl[39] br[39] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_42 
+ bl[40] br[40] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_43 
+ bl[41] br[41] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_44 
+ bl[42] br[42] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_45 
+ bl[43] br[43] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_46 
+ bl[44] br[44] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_47 
+ bl[45] br[45] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_48 
+ bl[46] br[46] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_49 
+ bl[47] br[47] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_50 
+ bl[48] br[48] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_51 
+ bl[49] br[49] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_52 
+ bl[50] br[50] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_53 
+ bl[51] br[51] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_54 
+ bl[52] br[52] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_55 
+ bl[53] br[53] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_56 
+ bl[54] br[54] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_57 
+ bl[55] br[55] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_58 
+ bl[56] br[56] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_59 
+ bl[57] br[57] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_60 
+ bl[58] br[58] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_61 
+ bl[59] br[59] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_62 
+ bl[60] br[60] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_63 
+ bl[61] br[61] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_64 
+ bl[62] br[62] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_65 
+ bl[63] br[63] vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_66 
+ vdd vdd vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_131_67 
+ vdd vdd vdd vss wl[129] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_0 
+ vdd vdd vss vdd vpb vnb wl[130] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_132_1 
+ rbl rbr vss vdd vpb vnb wl[130] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_132_2 
+ bl[0] br[0] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_3 
+ bl[1] br[1] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_4 
+ bl[2] br[2] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_5 
+ bl[3] br[3] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_6 
+ bl[4] br[4] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_7 
+ bl[5] br[5] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_8 
+ bl[6] br[6] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_9 
+ bl[7] br[7] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_10 
+ bl[8] br[8] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_11 
+ bl[9] br[9] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_12 
+ bl[10] br[10] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_13 
+ bl[11] br[11] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_14 
+ bl[12] br[12] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_15 
+ bl[13] br[13] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_16 
+ bl[14] br[14] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_17 
+ bl[15] br[15] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_18 
+ bl[16] br[16] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_19 
+ bl[17] br[17] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_20 
+ bl[18] br[18] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_21 
+ bl[19] br[19] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_22 
+ bl[20] br[20] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_23 
+ bl[21] br[21] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_24 
+ bl[22] br[22] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_25 
+ bl[23] br[23] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_26 
+ bl[24] br[24] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_27 
+ bl[25] br[25] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_28 
+ bl[26] br[26] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_29 
+ bl[27] br[27] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_30 
+ bl[28] br[28] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_31 
+ bl[29] br[29] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_32 
+ bl[30] br[30] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_33 
+ bl[31] br[31] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_34 
+ bl[32] br[32] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_35 
+ bl[33] br[33] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_36 
+ bl[34] br[34] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_37 
+ bl[35] br[35] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_38 
+ bl[36] br[36] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_39 
+ bl[37] br[37] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_40 
+ bl[38] br[38] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_41 
+ bl[39] br[39] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_42 
+ bl[40] br[40] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_43 
+ bl[41] br[41] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_44 
+ bl[42] br[42] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_45 
+ bl[43] br[43] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_46 
+ bl[44] br[44] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_47 
+ bl[45] br[45] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_48 
+ bl[46] br[46] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_49 
+ bl[47] br[47] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_50 
+ bl[48] br[48] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_51 
+ bl[49] br[49] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_52 
+ bl[50] br[50] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_53 
+ bl[51] br[51] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_54 
+ bl[52] br[52] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_55 
+ bl[53] br[53] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_56 
+ bl[54] br[54] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_57 
+ bl[55] br[55] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_58 
+ bl[56] br[56] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_59 
+ bl[57] br[57] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_60 
+ bl[58] br[58] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_61 
+ bl[59] br[59] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_62 
+ bl[60] br[60] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_63 
+ bl[61] br[61] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_64 
+ bl[62] br[62] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_65 
+ bl[63] br[63] vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_66 
+ vdd vdd vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_132_67 
+ vdd vdd vdd vss wl[130] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_0 
+ vdd vdd vss vdd vpb vnb wl[131] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_133_1 
+ rbl rbr vss vdd vpb vnb wl[131] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_133_2 
+ bl[0] br[0] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_3 
+ bl[1] br[1] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_4 
+ bl[2] br[2] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_5 
+ bl[3] br[3] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_6 
+ bl[4] br[4] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_7 
+ bl[5] br[5] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_8 
+ bl[6] br[6] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_9 
+ bl[7] br[7] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_10 
+ bl[8] br[8] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_11 
+ bl[9] br[9] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_12 
+ bl[10] br[10] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_13 
+ bl[11] br[11] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_14 
+ bl[12] br[12] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_15 
+ bl[13] br[13] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_16 
+ bl[14] br[14] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_17 
+ bl[15] br[15] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_18 
+ bl[16] br[16] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_19 
+ bl[17] br[17] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_20 
+ bl[18] br[18] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_21 
+ bl[19] br[19] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_22 
+ bl[20] br[20] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_23 
+ bl[21] br[21] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_24 
+ bl[22] br[22] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_25 
+ bl[23] br[23] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_26 
+ bl[24] br[24] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_27 
+ bl[25] br[25] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_28 
+ bl[26] br[26] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_29 
+ bl[27] br[27] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_30 
+ bl[28] br[28] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_31 
+ bl[29] br[29] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_32 
+ bl[30] br[30] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_33 
+ bl[31] br[31] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_34 
+ bl[32] br[32] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_35 
+ bl[33] br[33] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_36 
+ bl[34] br[34] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_37 
+ bl[35] br[35] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_38 
+ bl[36] br[36] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_39 
+ bl[37] br[37] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_40 
+ bl[38] br[38] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_41 
+ bl[39] br[39] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_42 
+ bl[40] br[40] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_43 
+ bl[41] br[41] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_44 
+ bl[42] br[42] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_45 
+ bl[43] br[43] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_46 
+ bl[44] br[44] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_47 
+ bl[45] br[45] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_48 
+ bl[46] br[46] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_49 
+ bl[47] br[47] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_50 
+ bl[48] br[48] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_51 
+ bl[49] br[49] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_52 
+ bl[50] br[50] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_53 
+ bl[51] br[51] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_54 
+ bl[52] br[52] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_55 
+ bl[53] br[53] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_56 
+ bl[54] br[54] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_57 
+ bl[55] br[55] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_58 
+ bl[56] br[56] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_59 
+ bl[57] br[57] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_60 
+ bl[58] br[58] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_61 
+ bl[59] br[59] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_62 
+ bl[60] br[60] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_63 
+ bl[61] br[61] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_64 
+ bl[62] br[62] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_65 
+ bl[63] br[63] vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_66 
+ vdd vdd vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_133_67 
+ vdd vdd vdd vss wl[131] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_0 
+ vdd vdd vss vdd vpb vnb wl[132] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_134_1 
+ rbl rbr vss vdd vpb vnb wl[132] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_134_2 
+ bl[0] br[0] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_3 
+ bl[1] br[1] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_4 
+ bl[2] br[2] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_5 
+ bl[3] br[3] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_6 
+ bl[4] br[4] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_7 
+ bl[5] br[5] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_8 
+ bl[6] br[6] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_9 
+ bl[7] br[7] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_10 
+ bl[8] br[8] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_11 
+ bl[9] br[9] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_12 
+ bl[10] br[10] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_13 
+ bl[11] br[11] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_14 
+ bl[12] br[12] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_15 
+ bl[13] br[13] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_16 
+ bl[14] br[14] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_17 
+ bl[15] br[15] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_18 
+ bl[16] br[16] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_19 
+ bl[17] br[17] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_20 
+ bl[18] br[18] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_21 
+ bl[19] br[19] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_22 
+ bl[20] br[20] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_23 
+ bl[21] br[21] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_24 
+ bl[22] br[22] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_25 
+ bl[23] br[23] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_26 
+ bl[24] br[24] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_27 
+ bl[25] br[25] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_28 
+ bl[26] br[26] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_29 
+ bl[27] br[27] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_30 
+ bl[28] br[28] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_31 
+ bl[29] br[29] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_32 
+ bl[30] br[30] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_33 
+ bl[31] br[31] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_34 
+ bl[32] br[32] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_35 
+ bl[33] br[33] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_36 
+ bl[34] br[34] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_37 
+ bl[35] br[35] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_38 
+ bl[36] br[36] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_39 
+ bl[37] br[37] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_40 
+ bl[38] br[38] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_41 
+ bl[39] br[39] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_42 
+ bl[40] br[40] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_43 
+ bl[41] br[41] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_44 
+ bl[42] br[42] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_45 
+ bl[43] br[43] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_46 
+ bl[44] br[44] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_47 
+ bl[45] br[45] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_48 
+ bl[46] br[46] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_49 
+ bl[47] br[47] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_50 
+ bl[48] br[48] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_51 
+ bl[49] br[49] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_52 
+ bl[50] br[50] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_53 
+ bl[51] br[51] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_54 
+ bl[52] br[52] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_55 
+ bl[53] br[53] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_56 
+ bl[54] br[54] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_57 
+ bl[55] br[55] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_58 
+ bl[56] br[56] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_59 
+ bl[57] br[57] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_60 
+ bl[58] br[58] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_61 
+ bl[59] br[59] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_62 
+ bl[60] br[60] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_63 
+ bl[61] br[61] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_64 
+ bl[62] br[62] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_65 
+ bl[63] br[63] vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_66 
+ vdd vdd vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_134_67 
+ vdd vdd vdd vss wl[132] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_0 
+ vdd vdd vss vdd vpb vnb wl[133] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_135_1 
+ rbl rbr vss vdd vpb vnb wl[133] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_135_2 
+ bl[0] br[0] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_3 
+ bl[1] br[1] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_4 
+ bl[2] br[2] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_5 
+ bl[3] br[3] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_6 
+ bl[4] br[4] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_7 
+ bl[5] br[5] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_8 
+ bl[6] br[6] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_9 
+ bl[7] br[7] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_10 
+ bl[8] br[8] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_11 
+ bl[9] br[9] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_12 
+ bl[10] br[10] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_13 
+ bl[11] br[11] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_14 
+ bl[12] br[12] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_15 
+ bl[13] br[13] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_16 
+ bl[14] br[14] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_17 
+ bl[15] br[15] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_18 
+ bl[16] br[16] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_19 
+ bl[17] br[17] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_20 
+ bl[18] br[18] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_21 
+ bl[19] br[19] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_22 
+ bl[20] br[20] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_23 
+ bl[21] br[21] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_24 
+ bl[22] br[22] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_25 
+ bl[23] br[23] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_26 
+ bl[24] br[24] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_27 
+ bl[25] br[25] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_28 
+ bl[26] br[26] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_29 
+ bl[27] br[27] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_30 
+ bl[28] br[28] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_31 
+ bl[29] br[29] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_32 
+ bl[30] br[30] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_33 
+ bl[31] br[31] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_34 
+ bl[32] br[32] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_35 
+ bl[33] br[33] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_36 
+ bl[34] br[34] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_37 
+ bl[35] br[35] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_38 
+ bl[36] br[36] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_39 
+ bl[37] br[37] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_40 
+ bl[38] br[38] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_41 
+ bl[39] br[39] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_42 
+ bl[40] br[40] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_43 
+ bl[41] br[41] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_44 
+ bl[42] br[42] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_45 
+ bl[43] br[43] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_46 
+ bl[44] br[44] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_47 
+ bl[45] br[45] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_48 
+ bl[46] br[46] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_49 
+ bl[47] br[47] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_50 
+ bl[48] br[48] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_51 
+ bl[49] br[49] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_52 
+ bl[50] br[50] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_53 
+ bl[51] br[51] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_54 
+ bl[52] br[52] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_55 
+ bl[53] br[53] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_56 
+ bl[54] br[54] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_57 
+ bl[55] br[55] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_58 
+ bl[56] br[56] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_59 
+ bl[57] br[57] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_60 
+ bl[58] br[58] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_61 
+ bl[59] br[59] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_62 
+ bl[60] br[60] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_63 
+ bl[61] br[61] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_64 
+ bl[62] br[62] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_65 
+ bl[63] br[63] vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_66 
+ vdd vdd vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_135_67 
+ vdd vdd vdd vss wl[133] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_0 
+ vdd vdd vss vdd vpb vnb wl[134] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_136_1 
+ rbl rbr vss vdd vpb vnb wl[134] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_136_2 
+ bl[0] br[0] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_3 
+ bl[1] br[1] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_4 
+ bl[2] br[2] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_5 
+ bl[3] br[3] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_6 
+ bl[4] br[4] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_7 
+ bl[5] br[5] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_8 
+ bl[6] br[6] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_9 
+ bl[7] br[7] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_10 
+ bl[8] br[8] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_11 
+ bl[9] br[9] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_12 
+ bl[10] br[10] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_13 
+ bl[11] br[11] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_14 
+ bl[12] br[12] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_15 
+ bl[13] br[13] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_16 
+ bl[14] br[14] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_17 
+ bl[15] br[15] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_18 
+ bl[16] br[16] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_19 
+ bl[17] br[17] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_20 
+ bl[18] br[18] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_21 
+ bl[19] br[19] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_22 
+ bl[20] br[20] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_23 
+ bl[21] br[21] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_24 
+ bl[22] br[22] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_25 
+ bl[23] br[23] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_26 
+ bl[24] br[24] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_27 
+ bl[25] br[25] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_28 
+ bl[26] br[26] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_29 
+ bl[27] br[27] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_30 
+ bl[28] br[28] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_31 
+ bl[29] br[29] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_32 
+ bl[30] br[30] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_33 
+ bl[31] br[31] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_34 
+ bl[32] br[32] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_35 
+ bl[33] br[33] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_36 
+ bl[34] br[34] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_37 
+ bl[35] br[35] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_38 
+ bl[36] br[36] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_39 
+ bl[37] br[37] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_40 
+ bl[38] br[38] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_41 
+ bl[39] br[39] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_42 
+ bl[40] br[40] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_43 
+ bl[41] br[41] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_44 
+ bl[42] br[42] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_45 
+ bl[43] br[43] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_46 
+ bl[44] br[44] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_47 
+ bl[45] br[45] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_48 
+ bl[46] br[46] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_49 
+ bl[47] br[47] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_50 
+ bl[48] br[48] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_51 
+ bl[49] br[49] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_52 
+ bl[50] br[50] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_53 
+ bl[51] br[51] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_54 
+ bl[52] br[52] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_55 
+ bl[53] br[53] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_56 
+ bl[54] br[54] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_57 
+ bl[55] br[55] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_58 
+ bl[56] br[56] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_59 
+ bl[57] br[57] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_60 
+ bl[58] br[58] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_61 
+ bl[59] br[59] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_62 
+ bl[60] br[60] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_63 
+ bl[61] br[61] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_64 
+ bl[62] br[62] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_65 
+ bl[63] br[63] vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_66 
+ vdd vdd vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_136_67 
+ vdd vdd vdd vss wl[134] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_0 
+ vdd vdd vss vdd vpb vnb wl[135] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_137_1 
+ rbl rbr vss vdd vpb vnb wl[135] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_137_2 
+ bl[0] br[0] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_3 
+ bl[1] br[1] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_4 
+ bl[2] br[2] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_5 
+ bl[3] br[3] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_6 
+ bl[4] br[4] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_7 
+ bl[5] br[5] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_8 
+ bl[6] br[6] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_9 
+ bl[7] br[7] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_10 
+ bl[8] br[8] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_11 
+ bl[9] br[9] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_12 
+ bl[10] br[10] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_13 
+ bl[11] br[11] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_14 
+ bl[12] br[12] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_15 
+ bl[13] br[13] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_16 
+ bl[14] br[14] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_17 
+ bl[15] br[15] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_18 
+ bl[16] br[16] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_19 
+ bl[17] br[17] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_20 
+ bl[18] br[18] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_21 
+ bl[19] br[19] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_22 
+ bl[20] br[20] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_23 
+ bl[21] br[21] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_24 
+ bl[22] br[22] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_25 
+ bl[23] br[23] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_26 
+ bl[24] br[24] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_27 
+ bl[25] br[25] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_28 
+ bl[26] br[26] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_29 
+ bl[27] br[27] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_30 
+ bl[28] br[28] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_31 
+ bl[29] br[29] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_32 
+ bl[30] br[30] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_33 
+ bl[31] br[31] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_34 
+ bl[32] br[32] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_35 
+ bl[33] br[33] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_36 
+ bl[34] br[34] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_37 
+ bl[35] br[35] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_38 
+ bl[36] br[36] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_39 
+ bl[37] br[37] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_40 
+ bl[38] br[38] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_41 
+ bl[39] br[39] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_42 
+ bl[40] br[40] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_43 
+ bl[41] br[41] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_44 
+ bl[42] br[42] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_45 
+ bl[43] br[43] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_46 
+ bl[44] br[44] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_47 
+ bl[45] br[45] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_48 
+ bl[46] br[46] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_49 
+ bl[47] br[47] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_50 
+ bl[48] br[48] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_51 
+ bl[49] br[49] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_52 
+ bl[50] br[50] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_53 
+ bl[51] br[51] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_54 
+ bl[52] br[52] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_55 
+ bl[53] br[53] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_56 
+ bl[54] br[54] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_57 
+ bl[55] br[55] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_58 
+ bl[56] br[56] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_59 
+ bl[57] br[57] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_60 
+ bl[58] br[58] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_61 
+ bl[59] br[59] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_62 
+ bl[60] br[60] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_63 
+ bl[61] br[61] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_64 
+ bl[62] br[62] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_65 
+ bl[63] br[63] vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_66 
+ vdd vdd vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_137_67 
+ vdd vdd vdd vss wl[135] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_0 
+ vdd vdd vss vdd vpb vnb wl[136] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_138_1 
+ rbl rbr vss vdd vpb vnb wl[136] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_138_2 
+ bl[0] br[0] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_3 
+ bl[1] br[1] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_4 
+ bl[2] br[2] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_5 
+ bl[3] br[3] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_6 
+ bl[4] br[4] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_7 
+ bl[5] br[5] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_8 
+ bl[6] br[6] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_9 
+ bl[7] br[7] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_10 
+ bl[8] br[8] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_11 
+ bl[9] br[9] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_12 
+ bl[10] br[10] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_13 
+ bl[11] br[11] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_14 
+ bl[12] br[12] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_15 
+ bl[13] br[13] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_16 
+ bl[14] br[14] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_17 
+ bl[15] br[15] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_18 
+ bl[16] br[16] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_19 
+ bl[17] br[17] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_20 
+ bl[18] br[18] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_21 
+ bl[19] br[19] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_22 
+ bl[20] br[20] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_23 
+ bl[21] br[21] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_24 
+ bl[22] br[22] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_25 
+ bl[23] br[23] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_26 
+ bl[24] br[24] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_27 
+ bl[25] br[25] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_28 
+ bl[26] br[26] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_29 
+ bl[27] br[27] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_30 
+ bl[28] br[28] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_31 
+ bl[29] br[29] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_32 
+ bl[30] br[30] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_33 
+ bl[31] br[31] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_34 
+ bl[32] br[32] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_35 
+ bl[33] br[33] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_36 
+ bl[34] br[34] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_37 
+ bl[35] br[35] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_38 
+ bl[36] br[36] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_39 
+ bl[37] br[37] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_40 
+ bl[38] br[38] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_41 
+ bl[39] br[39] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_42 
+ bl[40] br[40] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_43 
+ bl[41] br[41] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_44 
+ bl[42] br[42] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_45 
+ bl[43] br[43] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_46 
+ bl[44] br[44] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_47 
+ bl[45] br[45] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_48 
+ bl[46] br[46] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_49 
+ bl[47] br[47] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_50 
+ bl[48] br[48] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_51 
+ bl[49] br[49] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_52 
+ bl[50] br[50] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_53 
+ bl[51] br[51] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_54 
+ bl[52] br[52] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_55 
+ bl[53] br[53] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_56 
+ bl[54] br[54] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_57 
+ bl[55] br[55] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_58 
+ bl[56] br[56] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_59 
+ bl[57] br[57] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_60 
+ bl[58] br[58] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_61 
+ bl[59] br[59] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_62 
+ bl[60] br[60] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_63 
+ bl[61] br[61] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_64 
+ bl[62] br[62] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_65 
+ bl[63] br[63] vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_66 
+ vdd vdd vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_138_67 
+ vdd vdd vdd vss wl[136] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_0 
+ vdd vdd vss vdd vpb vnb wl[137] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_139_1 
+ rbl rbr vss vdd vpb vnb wl[137] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_139_2 
+ bl[0] br[0] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_3 
+ bl[1] br[1] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_4 
+ bl[2] br[2] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_5 
+ bl[3] br[3] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_6 
+ bl[4] br[4] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_7 
+ bl[5] br[5] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_8 
+ bl[6] br[6] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_9 
+ bl[7] br[7] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_10 
+ bl[8] br[8] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_11 
+ bl[9] br[9] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_12 
+ bl[10] br[10] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_13 
+ bl[11] br[11] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_14 
+ bl[12] br[12] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_15 
+ bl[13] br[13] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_16 
+ bl[14] br[14] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_17 
+ bl[15] br[15] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_18 
+ bl[16] br[16] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_19 
+ bl[17] br[17] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_20 
+ bl[18] br[18] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_21 
+ bl[19] br[19] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_22 
+ bl[20] br[20] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_23 
+ bl[21] br[21] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_24 
+ bl[22] br[22] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_25 
+ bl[23] br[23] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_26 
+ bl[24] br[24] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_27 
+ bl[25] br[25] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_28 
+ bl[26] br[26] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_29 
+ bl[27] br[27] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_30 
+ bl[28] br[28] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_31 
+ bl[29] br[29] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_32 
+ bl[30] br[30] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_33 
+ bl[31] br[31] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_34 
+ bl[32] br[32] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_35 
+ bl[33] br[33] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_36 
+ bl[34] br[34] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_37 
+ bl[35] br[35] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_38 
+ bl[36] br[36] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_39 
+ bl[37] br[37] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_40 
+ bl[38] br[38] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_41 
+ bl[39] br[39] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_42 
+ bl[40] br[40] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_43 
+ bl[41] br[41] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_44 
+ bl[42] br[42] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_45 
+ bl[43] br[43] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_46 
+ bl[44] br[44] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_47 
+ bl[45] br[45] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_48 
+ bl[46] br[46] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_49 
+ bl[47] br[47] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_50 
+ bl[48] br[48] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_51 
+ bl[49] br[49] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_52 
+ bl[50] br[50] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_53 
+ bl[51] br[51] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_54 
+ bl[52] br[52] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_55 
+ bl[53] br[53] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_56 
+ bl[54] br[54] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_57 
+ bl[55] br[55] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_58 
+ bl[56] br[56] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_59 
+ bl[57] br[57] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_60 
+ bl[58] br[58] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_61 
+ bl[59] br[59] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_62 
+ bl[60] br[60] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_63 
+ bl[61] br[61] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_64 
+ bl[62] br[62] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_65 
+ bl[63] br[63] vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_66 
+ vdd vdd vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_139_67 
+ vdd vdd vdd vss wl[137] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_0 
+ vdd vdd vss vdd vpb vnb wl[138] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_140_1 
+ rbl rbr vss vdd vpb vnb wl[138] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_140_2 
+ bl[0] br[0] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_3 
+ bl[1] br[1] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_4 
+ bl[2] br[2] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_5 
+ bl[3] br[3] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_6 
+ bl[4] br[4] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_7 
+ bl[5] br[5] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_8 
+ bl[6] br[6] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_9 
+ bl[7] br[7] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_10 
+ bl[8] br[8] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_11 
+ bl[9] br[9] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_12 
+ bl[10] br[10] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_13 
+ bl[11] br[11] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_14 
+ bl[12] br[12] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_15 
+ bl[13] br[13] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_16 
+ bl[14] br[14] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_17 
+ bl[15] br[15] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_18 
+ bl[16] br[16] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_19 
+ bl[17] br[17] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_20 
+ bl[18] br[18] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_21 
+ bl[19] br[19] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_22 
+ bl[20] br[20] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_23 
+ bl[21] br[21] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_24 
+ bl[22] br[22] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_25 
+ bl[23] br[23] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_26 
+ bl[24] br[24] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_27 
+ bl[25] br[25] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_28 
+ bl[26] br[26] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_29 
+ bl[27] br[27] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_30 
+ bl[28] br[28] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_31 
+ bl[29] br[29] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_32 
+ bl[30] br[30] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_33 
+ bl[31] br[31] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_34 
+ bl[32] br[32] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_35 
+ bl[33] br[33] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_36 
+ bl[34] br[34] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_37 
+ bl[35] br[35] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_38 
+ bl[36] br[36] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_39 
+ bl[37] br[37] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_40 
+ bl[38] br[38] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_41 
+ bl[39] br[39] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_42 
+ bl[40] br[40] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_43 
+ bl[41] br[41] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_44 
+ bl[42] br[42] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_45 
+ bl[43] br[43] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_46 
+ bl[44] br[44] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_47 
+ bl[45] br[45] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_48 
+ bl[46] br[46] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_49 
+ bl[47] br[47] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_50 
+ bl[48] br[48] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_51 
+ bl[49] br[49] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_52 
+ bl[50] br[50] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_53 
+ bl[51] br[51] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_54 
+ bl[52] br[52] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_55 
+ bl[53] br[53] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_56 
+ bl[54] br[54] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_57 
+ bl[55] br[55] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_58 
+ bl[56] br[56] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_59 
+ bl[57] br[57] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_60 
+ bl[58] br[58] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_61 
+ bl[59] br[59] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_62 
+ bl[60] br[60] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_63 
+ bl[61] br[61] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_64 
+ bl[62] br[62] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_65 
+ bl[63] br[63] vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_66 
+ vdd vdd vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_140_67 
+ vdd vdd vdd vss wl[138] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_0 
+ vdd vdd vss vdd vpb vnb wl[139] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_141_1 
+ rbl rbr vss vdd vpb vnb wl[139] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_141_2 
+ bl[0] br[0] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_3 
+ bl[1] br[1] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_4 
+ bl[2] br[2] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_5 
+ bl[3] br[3] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_6 
+ bl[4] br[4] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_7 
+ bl[5] br[5] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_8 
+ bl[6] br[6] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_9 
+ bl[7] br[7] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_10 
+ bl[8] br[8] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_11 
+ bl[9] br[9] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_12 
+ bl[10] br[10] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_13 
+ bl[11] br[11] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_14 
+ bl[12] br[12] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_15 
+ bl[13] br[13] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_16 
+ bl[14] br[14] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_17 
+ bl[15] br[15] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_18 
+ bl[16] br[16] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_19 
+ bl[17] br[17] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_20 
+ bl[18] br[18] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_21 
+ bl[19] br[19] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_22 
+ bl[20] br[20] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_23 
+ bl[21] br[21] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_24 
+ bl[22] br[22] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_25 
+ bl[23] br[23] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_26 
+ bl[24] br[24] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_27 
+ bl[25] br[25] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_28 
+ bl[26] br[26] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_29 
+ bl[27] br[27] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_30 
+ bl[28] br[28] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_31 
+ bl[29] br[29] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_32 
+ bl[30] br[30] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_33 
+ bl[31] br[31] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_34 
+ bl[32] br[32] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_35 
+ bl[33] br[33] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_36 
+ bl[34] br[34] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_37 
+ bl[35] br[35] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_38 
+ bl[36] br[36] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_39 
+ bl[37] br[37] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_40 
+ bl[38] br[38] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_41 
+ bl[39] br[39] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_42 
+ bl[40] br[40] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_43 
+ bl[41] br[41] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_44 
+ bl[42] br[42] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_45 
+ bl[43] br[43] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_46 
+ bl[44] br[44] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_47 
+ bl[45] br[45] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_48 
+ bl[46] br[46] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_49 
+ bl[47] br[47] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_50 
+ bl[48] br[48] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_51 
+ bl[49] br[49] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_52 
+ bl[50] br[50] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_53 
+ bl[51] br[51] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_54 
+ bl[52] br[52] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_55 
+ bl[53] br[53] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_56 
+ bl[54] br[54] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_57 
+ bl[55] br[55] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_58 
+ bl[56] br[56] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_59 
+ bl[57] br[57] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_60 
+ bl[58] br[58] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_61 
+ bl[59] br[59] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_62 
+ bl[60] br[60] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_63 
+ bl[61] br[61] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_64 
+ bl[62] br[62] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_65 
+ bl[63] br[63] vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_66 
+ vdd vdd vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_141_67 
+ vdd vdd vdd vss wl[139] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_0 
+ vdd vdd vss vdd vpb vnb wl[140] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_142_1 
+ rbl rbr vss vdd vpb vnb wl[140] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_142_2 
+ bl[0] br[0] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_3 
+ bl[1] br[1] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_4 
+ bl[2] br[2] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_5 
+ bl[3] br[3] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_6 
+ bl[4] br[4] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_7 
+ bl[5] br[5] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_8 
+ bl[6] br[6] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_9 
+ bl[7] br[7] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_10 
+ bl[8] br[8] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_11 
+ bl[9] br[9] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_12 
+ bl[10] br[10] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_13 
+ bl[11] br[11] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_14 
+ bl[12] br[12] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_15 
+ bl[13] br[13] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_16 
+ bl[14] br[14] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_17 
+ bl[15] br[15] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_18 
+ bl[16] br[16] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_19 
+ bl[17] br[17] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_20 
+ bl[18] br[18] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_21 
+ bl[19] br[19] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_22 
+ bl[20] br[20] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_23 
+ bl[21] br[21] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_24 
+ bl[22] br[22] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_25 
+ bl[23] br[23] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_26 
+ bl[24] br[24] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_27 
+ bl[25] br[25] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_28 
+ bl[26] br[26] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_29 
+ bl[27] br[27] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_30 
+ bl[28] br[28] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_31 
+ bl[29] br[29] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_32 
+ bl[30] br[30] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_33 
+ bl[31] br[31] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_34 
+ bl[32] br[32] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_35 
+ bl[33] br[33] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_36 
+ bl[34] br[34] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_37 
+ bl[35] br[35] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_38 
+ bl[36] br[36] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_39 
+ bl[37] br[37] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_40 
+ bl[38] br[38] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_41 
+ bl[39] br[39] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_42 
+ bl[40] br[40] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_43 
+ bl[41] br[41] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_44 
+ bl[42] br[42] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_45 
+ bl[43] br[43] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_46 
+ bl[44] br[44] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_47 
+ bl[45] br[45] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_48 
+ bl[46] br[46] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_49 
+ bl[47] br[47] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_50 
+ bl[48] br[48] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_51 
+ bl[49] br[49] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_52 
+ bl[50] br[50] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_53 
+ bl[51] br[51] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_54 
+ bl[52] br[52] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_55 
+ bl[53] br[53] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_56 
+ bl[54] br[54] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_57 
+ bl[55] br[55] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_58 
+ bl[56] br[56] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_59 
+ bl[57] br[57] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_60 
+ bl[58] br[58] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_61 
+ bl[59] br[59] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_62 
+ bl[60] br[60] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_63 
+ bl[61] br[61] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_64 
+ bl[62] br[62] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_65 
+ bl[63] br[63] vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_66 
+ vdd vdd vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_142_67 
+ vdd vdd vdd vss wl[140] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_0 
+ vdd vdd vss vdd vpb vnb wl[141] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_143_1 
+ rbl rbr vss vdd vpb vnb wl[141] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_143_2 
+ bl[0] br[0] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_3 
+ bl[1] br[1] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_4 
+ bl[2] br[2] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_5 
+ bl[3] br[3] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_6 
+ bl[4] br[4] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_7 
+ bl[5] br[5] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_8 
+ bl[6] br[6] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_9 
+ bl[7] br[7] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_10 
+ bl[8] br[8] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_11 
+ bl[9] br[9] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_12 
+ bl[10] br[10] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_13 
+ bl[11] br[11] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_14 
+ bl[12] br[12] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_15 
+ bl[13] br[13] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_16 
+ bl[14] br[14] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_17 
+ bl[15] br[15] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_18 
+ bl[16] br[16] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_19 
+ bl[17] br[17] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_20 
+ bl[18] br[18] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_21 
+ bl[19] br[19] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_22 
+ bl[20] br[20] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_23 
+ bl[21] br[21] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_24 
+ bl[22] br[22] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_25 
+ bl[23] br[23] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_26 
+ bl[24] br[24] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_27 
+ bl[25] br[25] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_28 
+ bl[26] br[26] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_29 
+ bl[27] br[27] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_30 
+ bl[28] br[28] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_31 
+ bl[29] br[29] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_32 
+ bl[30] br[30] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_33 
+ bl[31] br[31] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_34 
+ bl[32] br[32] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_35 
+ bl[33] br[33] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_36 
+ bl[34] br[34] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_37 
+ bl[35] br[35] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_38 
+ bl[36] br[36] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_39 
+ bl[37] br[37] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_40 
+ bl[38] br[38] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_41 
+ bl[39] br[39] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_42 
+ bl[40] br[40] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_43 
+ bl[41] br[41] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_44 
+ bl[42] br[42] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_45 
+ bl[43] br[43] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_46 
+ bl[44] br[44] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_47 
+ bl[45] br[45] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_48 
+ bl[46] br[46] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_49 
+ bl[47] br[47] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_50 
+ bl[48] br[48] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_51 
+ bl[49] br[49] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_52 
+ bl[50] br[50] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_53 
+ bl[51] br[51] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_54 
+ bl[52] br[52] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_55 
+ bl[53] br[53] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_56 
+ bl[54] br[54] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_57 
+ bl[55] br[55] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_58 
+ bl[56] br[56] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_59 
+ bl[57] br[57] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_60 
+ bl[58] br[58] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_61 
+ bl[59] br[59] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_62 
+ bl[60] br[60] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_63 
+ bl[61] br[61] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_64 
+ bl[62] br[62] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_65 
+ bl[63] br[63] vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_66 
+ vdd vdd vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_143_67 
+ vdd vdd vdd vss wl[141] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_0 
+ vdd vdd vss vdd vpb vnb wl[142] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_144_1 
+ rbl rbr vss vdd vpb vnb wl[142] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_144_2 
+ bl[0] br[0] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_3 
+ bl[1] br[1] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_4 
+ bl[2] br[2] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_5 
+ bl[3] br[3] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_6 
+ bl[4] br[4] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_7 
+ bl[5] br[5] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_8 
+ bl[6] br[6] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_9 
+ bl[7] br[7] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_10 
+ bl[8] br[8] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_11 
+ bl[9] br[9] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_12 
+ bl[10] br[10] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_13 
+ bl[11] br[11] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_14 
+ bl[12] br[12] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_15 
+ bl[13] br[13] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_16 
+ bl[14] br[14] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_17 
+ bl[15] br[15] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_18 
+ bl[16] br[16] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_19 
+ bl[17] br[17] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_20 
+ bl[18] br[18] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_21 
+ bl[19] br[19] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_22 
+ bl[20] br[20] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_23 
+ bl[21] br[21] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_24 
+ bl[22] br[22] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_25 
+ bl[23] br[23] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_26 
+ bl[24] br[24] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_27 
+ bl[25] br[25] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_28 
+ bl[26] br[26] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_29 
+ bl[27] br[27] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_30 
+ bl[28] br[28] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_31 
+ bl[29] br[29] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_32 
+ bl[30] br[30] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_33 
+ bl[31] br[31] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_34 
+ bl[32] br[32] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_35 
+ bl[33] br[33] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_36 
+ bl[34] br[34] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_37 
+ bl[35] br[35] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_38 
+ bl[36] br[36] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_39 
+ bl[37] br[37] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_40 
+ bl[38] br[38] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_41 
+ bl[39] br[39] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_42 
+ bl[40] br[40] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_43 
+ bl[41] br[41] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_44 
+ bl[42] br[42] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_45 
+ bl[43] br[43] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_46 
+ bl[44] br[44] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_47 
+ bl[45] br[45] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_48 
+ bl[46] br[46] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_49 
+ bl[47] br[47] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_50 
+ bl[48] br[48] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_51 
+ bl[49] br[49] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_52 
+ bl[50] br[50] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_53 
+ bl[51] br[51] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_54 
+ bl[52] br[52] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_55 
+ bl[53] br[53] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_56 
+ bl[54] br[54] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_57 
+ bl[55] br[55] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_58 
+ bl[56] br[56] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_59 
+ bl[57] br[57] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_60 
+ bl[58] br[58] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_61 
+ bl[59] br[59] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_62 
+ bl[60] br[60] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_63 
+ bl[61] br[61] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_64 
+ bl[62] br[62] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_65 
+ bl[63] br[63] vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_66 
+ vdd vdd vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_144_67 
+ vdd vdd vdd vss wl[142] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_0 
+ vdd vdd vss vdd vpb vnb wl[143] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_145_1 
+ rbl rbr vss vdd vpb vnb wl[143] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_145_2 
+ bl[0] br[0] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_3 
+ bl[1] br[1] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_4 
+ bl[2] br[2] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_5 
+ bl[3] br[3] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_6 
+ bl[4] br[4] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_7 
+ bl[5] br[5] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_8 
+ bl[6] br[6] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_9 
+ bl[7] br[7] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_10 
+ bl[8] br[8] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_11 
+ bl[9] br[9] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_12 
+ bl[10] br[10] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_13 
+ bl[11] br[11] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_14 
+ bl[12] br[12] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_15 
+ bl[13] br[13] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_16 
+ bl[14] br[14] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_17 
+ bl[15] br[15] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_18 
+ bl[16] br[16] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_19 
+ bl[17] br[17] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_20 
+ bl[18] br[18] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_21 
+ bl[19] br[19] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_22 
+ bl[20] br[20] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_23 
+ bl[21] br[21] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_24 
+ bl[22] br[22] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_25 
+ bl[23] br[23] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_26 
+ bl[24] br[24] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_27 
+ bl[25] br[25] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_28 
+ bl[26] br[26] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_29 
+ bl[27] br[27] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_30 
+ bl[28] br[28] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_31 
+ bl[29] br[29] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_32 
+ bl[30] br[30] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_33 
+ bl[31] br[31] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_34 
+ bl[32] br[32] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_35 
+ bl[33] br[33] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_36 
+ bl[34] br[34] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_37 
+ bl[35] br[35] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_38 
+ bl[36] br[36] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_39 
+ bl[37] br[37] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_40 
+ bl[38] br[38] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_41 
+ bl[39] br[39] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_42 
+ bl[40] br[40] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_43 
+ bl[41] br[41] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_44 
+ bl[42] br[42] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_45 
+ bl[43] br[43] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_46 
+ bl[44] br[44] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_47 
+ bl[45] br[45] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_48 
+ bl[46] br[46] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_49 
+ bl[47] br[47] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_50 
+ bl[48] br[48] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_51 
+ bl[49] br[49] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_52 
+ bl[50] br[50] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_53 
+ bl[51] br[51] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_54 
+ bl[52] br[52] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_55 
+ bl[53] br[53] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_56 
+ bl[54] br[54] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_57 
+ bl[55] br[55] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_58 
+ bl[56] br[56] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_59 
+ bl[57] br[57] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_60 
+ bl[58] br[58] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_61 
+ bl[59] br[59] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_62 
+ bl[60] br[60] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_63 
+ bl[61] br[61] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_64 
+ bl[62] br[62] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_65 
+ bl[63] br[63] vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_66 
+ vdd vdd vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_145_67 
+ vdd vdd vdd vss wl[143] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_0 
+ vdd vdd vss vdd vpb vnb wl[144] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_146_1 
+ rbl rbr vss vdd vpb vnb wl[144] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_146_2 
+ bl[0] br[0] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_3 
+ bl[1] br[1] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_4 
+ bl[2] br[2] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_5 
+ bl[3] br[3] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_6 
+ bl[4] br[4] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_7 
+ bl[5] br[5] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_8 
+ bl[6] br[6] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_9 
+ bl[7] br[7] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_10 
+ bl[8] br[8] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_11 
+ bl[9] br[9] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_12 
+ bl[10] br[10] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_13 
+ bl[11] br[11] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_14 
+ bl[12] br[12] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_15 
+ bl[13] br[13] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_16 
+ bl[14] br[14] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_17 
+ bl[15] br[15] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_18 
+ bl[16] br[16] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_19 
+ bl[17] br[17] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_20 
+ bl[18] br[18] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_21 
+ bl[19] br[19] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_22 
+ bl[20] br[20] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_23 
+ bl[21] br[21] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_24 
+ bl[22] br[22] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_25 
+ bl[23] br[23] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_26 
+ bl[24] br[24] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_27 
+ bl[25] br[25] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_28 
+ bl[26] br[26] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_29 
+ bl[27] br[27] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_30 
+ bl[28] br[28] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_31 
+ bl[29] br[29] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_32 
+ bl[30] br[30] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_33 
+ bl[31] br[31] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_34 
+ bl[32] br[32] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_35 
+ bl[33] br[33] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_36 
+ bl[34] br[34] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_37 
+ bl[35] br[35] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_38 
+ bl[36] br[36] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_39 
+ bl[37] br[37] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_40 
+ bl[38] br[38] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_41 
+ bl[39] br[39] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_42 
+ bl[40] br[40] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_43 
+ bl[41] br[41] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_44 
+ bl[42] br[42] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_45 
+ bl[43] br[43] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_46 
+ bl[44] br[44] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_47 
+ bl[45] br[45] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_48 
+ bl[46] br[46] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_49 
+ bl[47] br[47] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_50 
+ bl[48] br[48] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_51 
+ bl[49] br[49] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_52 
+ bl[50] br[50] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_53 
+ bl[51] br[51] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_54 
+ bl[52] br[52] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_55 
+ bl[53] br[53] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_56 
+ bl[54] br[54] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_57 
+ bl[55] br[55] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_58 
+ bl[56] br[56] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_59 
+ bl[57] br[57] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_60 
+ bl[58] br[58] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_61 
+ bl[59] br[59] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_62 
+ bl[60] br[60] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_63 
+ bl[61] br[61] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_64 
+ bl[62] br[62] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_65 
+ bl[63] br[63] vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_66 
+ vdd vdd vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_146_67 
+ vdd vdd vdd vss wl[144] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_0 
+ vdd vdd vss vdd vpb vnb wl[145] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_147_1 
+ rbl rbr vss vdd vpb vnb wl[145] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_147_2 
+ bl[0] br[0] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_3 
+ bl[1] br[1] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_4 
+ bl[2] br[2] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_5 
+ bl[3] br[3] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_6 
+ bl[4] br[4] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_7 
+ bl[5] br[5] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_8 
+ bl[6] br[6] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_9 
+ bl[7] br[7] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_10 
+ bl[8] br[8] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_11 
+ bl[9] br[9] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_12 
+ bl[10] br[10] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_13 
+ bl[11] br[11] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_14 
+ bl[12] br[12] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_15 
+ bl[13] br[13] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_16 
+ bl[14] br[14] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_17 
+ bl[15] br[15] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_18 
+ bl[16] br[16] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_19 
+ bl[17] br[17] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_20 
+ bl[18] br[18] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_21 
+ bl[19] br[19] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_22 
+ bl[20] br[20] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_23 
+ bl[21] br[21] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_24 
+ bl[22] br[22] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_25 
+ bl[23] br[23] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_26 
+ bl[24] br[24] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_27 
+ bl[25] br[25] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_28 
+ bl[26] br[26] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_29 
+ bl[27] br[27] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_30 
+ bl[28] br[28] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_31 
+ bl[29] br[29] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_32 
+ bl[30] br[30] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_33 
+ bl[31] br[31] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_34 
+ bl[32] br[32] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_35 
+ bl[33] br[33] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_36 
+ bl[34] br[34] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_37 
+ bl[35] br[35] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_38 
+ bl[36] br[36] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_39 
+ bl[37] br[37] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_40 
+ bl[38] br[38] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_41 
+ bl[39] br[39] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_42 
+ bl[40] br[40] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_43 
+ bl[41] br[41] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_44 
+ bl[42] br[42] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_45 
+ bl[43] br[43] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_46 
+ bl[44] br[44] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_47 
+ bl[45] br[45] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_48 
+ bl[46] br[46] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_49 
+ bl[47] br[47] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_50 
+ bl[48] br[48] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_51 
+ bl[49] br[49] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_52 
+ bl[50] br[50] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_53 
+ bl[51] br[51] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_54 
+ bl[52] br[52] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_55 
+ bl[53] br[53] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_56 
+ bl[54] br[54] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_57 
+ bl[55] br[55] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_58 
+ bl[56] br[56] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_59 
+ bl[57] br[57] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_60 
+ bl[58] br[58] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_61 
+ bl[59] br[59] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_62 
+ bl[60] br[60] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_63 
+ bl[61] br[61] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_64 
+ bl[62] br[62] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_65 
+ bl[63] br[63] vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_66 
+ vdd vdd vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_147_67 
+ vdd vdd vdd vss wl[145] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_0 
+ vdd vdd vss vdd vpb vnb wl[146] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_148_1 
+ rbl rbr vss vdd vpb vnb wl[146] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_148_2 
+ bl[0] br[0] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_3 
+ bl[1] br[1] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_4 
+ bl[2] br[2] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_5 
+ bl[3] br[3] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_6 
+ bl[4] br[4] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_7 
+ bl[5] br[5] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_8 
+ bl[6] br[6] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_9 
+ bl[7] br[7] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_10 
+ bl[8] br[8] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_11 
+ bl[9] br[9] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_12 
+ bl[10] br[10] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_13 
+ bl[11] br[11] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_14 
+ bl[12] br[12] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_15 
+ bl[13] br[13] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_16 
+ bl[14] br[14] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_17 
+ bl[15] br[15] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_18 
+ bl[16] br[16] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_19 
+ bl[17] br[17] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_20 
+ bl[18] br[18] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_21 
+ bl[19] br[19] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_22 
+ bl[20] br[20] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_23 
+ bl[21] br[21] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_24 
+ bl[22] br[22] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_25 
+ bl[23] br[23] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_26 
+ bl[24] br[24] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_27 
+ bl[25] br[25] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_28 
+ bl[26] br[26] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_29 
+ bl[27] br[27] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_30 
+ bl[28] br[28] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_31 
+ bl[29] br[29] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_32 
+ bl[30] br[30] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_33 
+ bl[31] br[31] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_34 
+ bl[32] br[32] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_35 
+ bl[33] br[33] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_36 
+ bl[34] br[34] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_37 
+ bl[35] br[35] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_38 
+ bl[36] br[36] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_39 
+ bl[37] br[37] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_40 
+ bl[38] br[38] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_41 
+ bl[39] br[39] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_42 
+ bl[40] br[40] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_43 
+ bl[41] br[41] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_44 
+ bl[42] br[42] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_45 
+ bl[43] br[43] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_46 
+ bl[44] br[44] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_47 
+ bl[45] br[45] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_48 
+ bl[46] br[46] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_49 
+ bl[47] br[47] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_50 
+ bl[48] br[48] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_51 
+ bl[49] br[49] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_52 
+ bl[50] br[50] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_53 
+ bl[51] br[51] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_54 
+ bl[52] br[52] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_55 
+ bl[53] br[53] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_56 
+ bl[54] br[54] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_57 
+ bl[55] br[55] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_58 
+ bl[56] br[56] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_59 
+ bl[57] br[57] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_60 
+ bl[58] br[58] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_61 
+ bl[59] br[59] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_62 
+ bl[60] br[60] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_63 
+ bl[61] br[61] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_64 
+ bl[62] br[62] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_65 
+ bl[63] br[63] vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_66 
+ vdd vdd vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_148_67 
+ vdd vdd vdd vss wl[146] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_0 
+ vdd vdd vss vdd vpb vnb wl[147] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_149_1 
+ rbl rbr vss vdd vpb vnb wl[147] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_149_2 
+ bl[0] br[0] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_3 
+ bl[1] br[1] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_4 
+ bl[2] br[2] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_5 
+ bl[3] br[3] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_6 
+ bl[4] br[4] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_7 
+ bl[5] br[5] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_8 
+ bl[6] br[6] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_9 
+ bl[7] br[7] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_10 
+ bl[8] br[8] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_11 
+ bl[9] br[9] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_12 
+ bl[10] br[10] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_13 
+ bl[11] br[11] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_14 
+ bl[12] br[12] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_15 
+ bl[13] br[13] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_16 
+ bl[14] br[14] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_17 
+ bl[15] br[15] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_18 
+ bl[16] br[16] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_19 
+ bl[17] br[17] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_20 
+ bl[18] br[18] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_21 
+ bl[19] br[19] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_22 
+ bl[20] br[20] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_23 
+ bl[21] br[21] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_24 
+ bl[22] br[22] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_25 
+ bl[23] br[23] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_26 
+ bl[24] br[24] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_27 
+ bl[25] br[25] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_28 
+ bl[26] br[26] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_29 
+ bl[27] br[27] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_30 
+ bl[28] br[28] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_31 
+ bl[29] br[29] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_32 
+ bl[30] br[30] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_33 
+ bl[31] br[31] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_34 
+ bl[32] br[32] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_35 
+ bl[33] br[33] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_36 
+ bl[34] br[34] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_37 
+ bl[35] br[35] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_38 
+ bl[36] br[36] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_39 
+ bl[37] br[37] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_40 
+ bl[38] br[38] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_41 
+ bl[39] br[39] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_42 
+ bl[40] br[40] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_43 
+ bl[41] br[41] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_44 
+ bl[42] br[42] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_45 
+ bl[43] br[43] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_46 
+ bl[44] br[44] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_47 
+ bl[45] br[45] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_48 
+ bl[46] br[46] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_49 
+ bl[47] br[47] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_50 
+ bl[48] br[48] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_51 
+ bl[49] br[49] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_52 
+ bl[50] br[50] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_53 
+ bl[51] br[51] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_54 
+ bl[52] br[52] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_55 
+ bl[53] br[53] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_56 
+ bl[54] br[54] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_57 
+ bl[55] br[55] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_58 
+ bl[56] br[56] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_59 
+ bl[57] br[57] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_60 
+ bl[58] br[58] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_61 
+ bl[59] br[59] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_62 
+ bl[60] br[60] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_63 
+ bl[61] br[61] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_64 
+ bl[62] br[62] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_65 
+ bl[63] br[63] vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_66 
+ vdd vdd vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_149_67 
+ vdd vdd vdd vss wl[147] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_0 
+ vdd vdd vss vdd vpb vnb wl[148] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_150_1 
+ rbl rbr vss vdd vpb vnb wl[148] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_150_2 
+ bl[0] br[0] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_3 
+ bl[1] br[1] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_4 
+ bl[2] br[2] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_5 
+ bl[3] br[3] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_6 
+ bl[4] br[4] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_7 
+ bl[5] br[5] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_8 
+ bl[6] br[6] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_9 
+ bl[7] br[7] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_10 
+ bl[8] br[8] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_11 
+ bl[9] br[9] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_12 
+ bl[10] br[10] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_13 
+ bl[11] br[11] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_14 
+ bl[12] br[12] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_15 
+ bl[13] br[13] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_16 
+ bl[14] br[14] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_17 
+ bl[15] br[15] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_18 
+ bl[16] br[16] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_19 
+ bl[17] br[17] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_20 
+ bl[18] br[18] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_21 
+ bl[19] br[19] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_22 
+ bl[20] br[20] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_23 
+ bl[21] br[21] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_24 
+ bl[22] br[22] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_25 
+ bl[23] br[23] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_26 
+ bl[24] br[24] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_27 
+ bl[25] br[25] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_28 
+ bl[26] br[26] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_29 
+ bl[27] br[27] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_30 
+ bl[28] br[28] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_31 
+ bl[29] br[29] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_32 
+ bl[30] br[30] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_33 
+ bl[31] br[31] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_34 
+ bl[32] br[32] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_35 
+ bl[33] br[33] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_36 
+ bl[34] br[34] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_37 
+ bl[35] br[35] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_38 
+ bl[36] br[36] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_39 
+ bl[37] br[37] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_40 
+ bl[38] br[38] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_41 
+ bl[39] br[39] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_42 
+ bl[40] br[40] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_43 
+ bl[41] br[41] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_44 
+ bl[42] br[42] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_45 
+ bl[43] br[43] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_46 
+ bl[44] br[44] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_47 
+ bl[45] br[45] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_48 
+ bl[46] br[46] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_49 
+ bl[47] br[47] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_50 
+ bl[48] br[48] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_51 
+ bl[49] br[49] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_52 
+ bl[50] br[50] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_53 
+ bl[51] br[51] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_54 
+ bl[52] br[52] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_55 
+ bl[53] br[53] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_56 
+ bl[54] br[54] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_57 
+ bl[55] br[55] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_58 
+ bl[56] br[56] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_59 
+ bl[57] br[57] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_60 
+ bl[58] br[58] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_61 
+ bl[59] br[59] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_62 
+ bl[60] br[60] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_63 
+ bl[61] br[61] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_64 
+ bl[62] br[62] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_65 
+ bl[63] br[63] vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_66 
+ vdd vdd vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_150_67 
+ vdd vdd vdd vss wl[148] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_0 
+ vdd vdd vss vdd vpb vnb wl[149] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_151_1 
+ rbl rbr vss vdd vpb vnb wl[149] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_151_2 
+ bl[0] br[0] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_3 
+ bl[1] br[1] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_4 
+ bl[2] br[2] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_5 
+ bl[3] br[3] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_6 
+ bl[4] br[4] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_7 
+ bl[5] br[5] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_8 
+ bl[6] br[6] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_9 
+ bl[7] br[7] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_10 
+ bl[8] br[8] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_11 
+ bl[9] br[9] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_12 
+ bl[10] br[10] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_13 
+ bl[11] br[11] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_14 
+ bl[12] br[12] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_15 
+ bl[13] br[13] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_16 
+ bl[14] br[14] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_17 
+ bl[15] br[15] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_18 
+ bl[16] br[16] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_19 
+ bl[17] br[17] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_20 
+ bl[18] br[18] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_21 
+ bl[19] br[19] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_22 
+ bl[20] br[20] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_23 
+ bl[21] br[21] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_24 
+ bl[22] br[22] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_25 
+ bl[23] br[23] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_26 
+ bl[24] br[24] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_27 
+ bl[25] br[25] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_28 
+ bl[26] br[26] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_29 
+ bl[27] br[27] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_30 
+ bl[28] br[28] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_31 
+ bl[29] br[29] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_32 
+ bl[30] br[30] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_33 
+ bl[31] br[31] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_34 
+ bl[32] br[32] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_35 
+ bl[33] br[33] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_36 
+ bl[34] br[34] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_37 
+ bl[35] br[35] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_38 
+ bl[36] br[36] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_39 
+ bl[37] br[37] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_40 
+ bl[38] br[38] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_41 
+ bl[39] br[39] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_42 
+ bl[40] br[40] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_43 
+ bl[41] br[41] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_44 
+ bl[42] br[42] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_45 
+ bl[43] br[43] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_46 
+ bl[44] br[44] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_47 
+ bl[45] br[45] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_48 
+ bl[46] br[46] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_49 
+ bl[47] br[47] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_50 
+ bl[48] br[48] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_51 
+ bl[49] br[49] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_52 
+ bl[50] br[50] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_53 
+ bl[51] br[51] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_54 
+ bl[52] br[52] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_55 
+ bl[53] br[53] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_56 
+ bl[54] br[54] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_57 
+ bl[55] br[55] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_58 
+ bl[56] br[56] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_59 
+ bl[57] br[57] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_60 
+ bl[58] br[58] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_61 
+ bl[59] br[59] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_62 
+ bl[60] br[60] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_63 
+ bl[61] br[61] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_64 
+ bl[62] br[62] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_65 
+ bl[63] br[63] vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_66 
+ vdd vdd vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_151_67 
+ vdd vdd vdd vss wl[149] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_0 
+ vdd vdd vss vdd vpb vnb wl[150] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_152_1 
+ rbl rbr vss vdd vpb vnb wl[150] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_152_2 
+ bl[0] br[0] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_3 
+ bl[1] br[1] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_4 
+ bl[2] br[2] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_5 
+ bl[3] br[3] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_6 
+ bl[4] br[4] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_7 
+ bl[5] br[5] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_8 
+ bl[6] br[6] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_9 
+ bl[7] br[7] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_10 
+ bl[8] br[8] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_11 
+ bl[9] br[9] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_12 
+ bl[10] br[10] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_13 
+ bl[11] br[11] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_14 
+ bl[12] br[12] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_15 
+ bl[13] br[13] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_16 
+ bl[14] br[14] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_17 
+ bl[15] br[15] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_18 
+ bl[16] br[16] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_19 
+ bl[17] br[17] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_20 
+ bl[18] br[18] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_21 
+ bl[19] br[19] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_22 
+ bl[20] br[20] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_23 
+ bl[21] br[21] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_24 
+ bl[22] br[22] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_25 
+ bl[23] br[23] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_26 
+ bl[24] br[24] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_27 
+ bl[25] br[25] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_28 
+ bl[26] br[26] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_29 
+ bl[27] br[27] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_30 
+ bl[28] br[28] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_31 
+ bl[29] br[29] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_32 
+ bl[30] br[30] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_33 
+ bl[31] br[31] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_34 
+ bl[32] br[32] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_35 
+ bl[33] br[33] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_36 
+ bl[34] br[34] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_37 
+ bl[35] br[35] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_38 
+ bl[36] br[36] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_39 
+ bl[37] br[37] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_40 
+ bl[38] br[38] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_41 
+ bl[39] br[39] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_42 
+ bl[40] br[40] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_43 
+ bl[41] br[41] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_44 
+ bl[42] br[42] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_45 
+ bl[43] br[43] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_46 
+ bl[44] br[44] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_47 
+ bl[45] br[45] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_48 
+ bl[46] br[46] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_49 
+ bl[47] br[47] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_50 
+ bl[48] br[48] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_51 
+ bl[49] br[49] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_52 
+ bl[50] br[50] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_53 
+ bl[51] br[51] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_54 
+ bl[52] br[52] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_55 
+ bl[53] br[53] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_56 
+ bl[54] br[54] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_57 
+ bl[55] br[55] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_58 
+ bl[56] br[56] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_59 
+ bl[57] br[57] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_60 
+ bl[58] br[58] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_61 
+ bl[59] br[59] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_62 
+ bl[60] br[60] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_63 
+ bl[61] br[61] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_64 
+ bl[62] br[62] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_65 
+ bl[63] br[63] vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_66 
+ vdd vdd vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_152_67 
+ vdd vdd vdd vss wl[150] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_0 
+ vdd vdd vss vdd vpb vnb wl[151] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_153_1 
+ rbl rbr vss vdd vpb vnb wl[151] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_153_2 
+ bl[0] br[0] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_3 
+ bl[1] br[1] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_4 
+ bl[2] br[2] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_5 
+ bl[3] br[3] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_6 
+ bl[4] br[4] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_7 
+ bl[5] br[5] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_8 
+ bl[6] br[6] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_9 
+ bl[7] br[7] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_10 
+ bl[8] br[8] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_11 
+ bl[9] br[9] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_12 
+ bl[10] br[10] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_13 
+ bl[11] br[11] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_14 
+ bl[12] br[12] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_15 
+ bl[13] br[13] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_16 
+ bl[14] br[14] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_17 
+ bl[15] br[15] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_18 
+ bl[16] br[16] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_19 
+ bl[17] br[17] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_20 
+ bl[18] br[18] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_21 
+ bl[19] br[19] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_22 
+ bl[20] br[20] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_23 
+ bl[21] br[21] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_24 
+ bl[22] br[22] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_25 
+ bl[23] br[23] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_26 
+ bl[24] br[24] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_27 
+ bl[25] br[25] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_28 
+ bl[26] br[26] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_29 
+ bl[27] br[27] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_30 
+ bl[28] br[28] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_31 
+ bl[29] br[29] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_32 
+ bl[30] br[30] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_33 
+ bl[31] br[31] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_34 
+ bl[32] br[32] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_35 
+ bl[33] br[33] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_36 
+ bl[34] br[34] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_37 
+ bl[35] br[35] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_38 
+ bl[36] br[36] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_39 
+ bl[37] br[37] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_40 
+ bl[38] br[38] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_41 
+ bl[39] br[39] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_42 
+ bl[40] br[40] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_43 
+ bl[41] br[41] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_44 
+ bl[42] br[42] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_45 
+ bl[43] br[43] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_46 
+ bl[44] br[44] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_47 
+ bl[45] br[45] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_48 
+ bl[46] br[46] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_49 
+ bl[47] br[47] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_50 
+ bl[48] br[48] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_51 
+ bl[49] br[49] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_52 
+ bl[50] br[50] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_53 
+ bl[51] br[51] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_54 
+ bl[52] br[52] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_55 
+ bl[53] br[53] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_56 
+ bl[54] br[54] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_57 
+ bl[55] br[55] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_58 
+ bl[56] br[56] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_59 
+ bl[57] br[57] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_60 
+ bl[58] br[58] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_61 
+ bl[59] br[59] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_62 
+ bl[60] br[60] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_63 
+ bl[61] br[61] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_64 
+ bl[62] br[62] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_65 
+ bl[63] br[63] vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_66 
+ vdd vdd vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_153_67 
+ vdd vdd vdd vss wl[151] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_0 
+ vdd vdd vss vdd vpb vnb wl[152] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_154_1 
+ rbl rbr vss vdd vpb vnb wl[152] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_154_2 
+ bl[0] br[0] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_3 
+ bl[1] br[1] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_4 
+ bl[2] br[2] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_5 
+ bl[3] br[3] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_6 
+ bl[4] br[4] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_7 
+ bl[5] br[5] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_8 
+ bl[6] br[6] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_9 
+ bl[7] br[7] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_10 
+ bl[8] br[8] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_11 
+ bl[9] br[9] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_12 
+ bl[10] br[10] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_13 
+ bl[11] br[11] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_14 
+ bl[12] br[12] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_15 
+ bl[13] br[13] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_16 
+ bl[14] br[14] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_17 
+ bl[15] br[15] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_18 
+ bl[16] br[16] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_19 
+ bl[17] br[17] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_20 
+ bl[18] br[18] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_21 
+ bl[19] br[19] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_22 
+ bl[20] br[20] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_23 
+ bl[21] br[21] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_24 
+ bl[22] br[22] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_25 
+ bl[23] br[23] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_26 
+ bl[24] br[24] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_27 
+ bl[25] br[25] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_28 
+ bl[26] br[26] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_29 
+ bl[27] br[27] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_30 
+ bl[28] br[28] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_31 
+ bl[29] br[29] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_32 
+ bl[30] br[30] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_33 
+ bl[31] br[31] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_34 
+ bl[32] br[32] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_35 
+ bl[33] br[33] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_36 
+ bl[34] br[34] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_37 
+ bl[35] br[35] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_38 
+ bl[36] br[36] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_39 
+ bl[37] br[37] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_40 
+ bl[38] br[38] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_41 
+ bl[39] br[39] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_42 
+ bl[40] br[40] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_43 
+ bl[41] br[41] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_44 
+ bl[42] br[42] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_45 
+ bl[43] br[43] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_46 
+ bl[44] br[44] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_47 
+ bl[45] br[45] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_48 
+ bl[46] br[46] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_49 
+ bl[47] br[47] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_50 
+ bl[48] br[48] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_51 
+ bl[49] br[49] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_52 
+ bl[50] br[50] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_53 
+ bl[51] br[51] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_54 
+ bl[52] br[52] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_55 
+ bl[53] br[53] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_56 
+ bl[54] br[54] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_57 
+ bl[55] br[55] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_58 
+ bl[56] br[56] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_59 
+ bl[57] br[57] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_60 
+ bl[58] br[58] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_61 
+ bl[59] br[59] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_62 
+ bl[60] br[60] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_63 
+ bl[61] br[61] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_64 
+ bl[62] br[62] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_65 
+ bl[63] br[63] vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_66 
+ vdd vdd vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_154_67 
+ vdd vdd vdd vss wl[152] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_0 
+ vdd vdd vss vdd vpb vnb wl[153] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_155_1 
+ rbl rbr vss vdd vpb vnb wl[153] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_155_2 
+ bl[0] br[0] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_3 
+ bl[1] br[1] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_4 
+ bl[2] br[2] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_5 
+ bl[3] br[3] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_6 
+ bl[4] br[4] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_7 
+ bl[5] br[5] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_8 
+ bl[6] br[6] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_9 
+ bl[7] br[7] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_10 
+ bl[8] br[8] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_11 
+ bl[9] br[9] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_12 
+ bl[10] br[10] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_13 
+ bl[11] br[11] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_14 
+ bl[12] br[12] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_15 
+ bl[13] br[13] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_16 
+ bl[14] br[14] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_17 
+ bl[15] br[15] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_18 
+ bl[16] br[16] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_19 
+ bl[17] br[17] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_20 
+ bl[18] br[18] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_21 
+ bl[19] br[19] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_22 
+ bl[20] br[20] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_23 
+ bl[21] br[21] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_24 
+ bl[22] br[22] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_25 
+ bl[23] br[23] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_26 
+ bl[24] br[24] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_27 
+ bl[25] br[25] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_28 
+ bl[26] br[26] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_29 
+ bl[27] br[27] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_30 
+ bl[28] br[28] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_31 
+ bl[29] br[29] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_32 
+ bl[30] br[30] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_33 
+ bl[31] br[31] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_34 
+ bl[32] br[32] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_35 
+ bl[33] br[33] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_36 
+ bl[34] br[34] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_37 
+ bl[35] br[35] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_38 
+ bl[36] br[36] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_39 
+ bl[37] br[37] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_40 
+ bl[38] br[38] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_41 
+ bl[39] br[39] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_42 
+ bl[40] br[40] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_43 
+ bl[41] br[41] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_44 
+ bl[42] br[42] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_45 
+ bl[43] br[43] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_46 
+ bl[44] br[44] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_47 
+ bl[45] br[45] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_48 
+ bl[46] br[46] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_49 
+ bl[47] br[47] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_50 
+ bl[48] br[48] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_51 
+ bl[49] br[49] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_52 
+ bl[50] br[50] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_53 
+ bl[51] br[51] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_54 
+ bl[52] br[52] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_55 
+ bl[53] br[53] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_56 
+ bl[54] br[54] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_57 
+ bl[55] br[55] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_58 
+ bl[56] br[56] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_59 
+ bl[57] br[57] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_60 
+ bl[58] br[58] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_61 
+ bl[59] br[59] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_62 
+ bl[60] br[60] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_63 
+ bl[61] br[61] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_64 
+ bl[62] br[62] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_65 
+ bl[63] br[63] vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_66 
+ vdd vdd vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_155_67 
+ vdd vdd vdd vss wl[153] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_0 
+ vdd vdd vss vdd vpb vnb wl[154] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_156_1 
+ rbl rbr vss vdd vpb vnb wl[154] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_156_2 
+ bl[0] br[0] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_3 
+ bl[1] br[1] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_4 
+ bl[2] br[2] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_5 
+ bl[3] br[3] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_6 
+ bl[4] br[4] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_7 
+ bl[5] br[5] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_8 
+ bl[6] br[6] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_9 
+ bl[7] br[7] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_10 
+ bl[8] br[8] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_11 
+ bl[9] br[9] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_12 
+ bl[10] br[10] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_13 
+ bl[11] br[11] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_14 
+ bl[12] br[12] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_15 
+ bl[13] br[13] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_16 
+ bl[14] br[14] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_17 
+ bl[15] br[15] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_18 
+ bl[16] br[16] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_19 
+ bl[17] br[17] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_20 
+ bl[18] br[18] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_21 
+ bl[19] br[19] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_22 
+ bl[20] br[20] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_23 
+ bl[21] br[21] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_24 
+ bl[22] br[22] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_25 
+ bl[23] br[23] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_26 
+ bl[24] br[24] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_27 
+ bl[25] br[25] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_28 
+ bl[26] br[26] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_29 
+ bl[27] br[27] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_30 
+ bl[28] br[28] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_31 
+ bl[29] br[29] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_32 
+ bl[30] br[30] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_33 
+ bl[31] br[31] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_34 
+ bl[32] br[32] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_35 
+ bl[33] br[33] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_36 
+ bl[34] br[34] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_37 
+ bl[35] br[35] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_38 
+ bl[36] br[36] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_39 
+ bl[37] br[37] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_40 
+ bl[38] br[38] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_41 
+ bl[39] br[39] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_42 
+ bl[40] br[40] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_43 
+ bl[41] br[41] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_44 
+ bl[42] br[42] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_45 
+ bl[43] br[43] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_46 
+ bl[44] br[44] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_47 
+ bl[45] br[45] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_48 
+ bl[46] br[46] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_49 
+ bl[47] br[47] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_50 
+ bl[48] br[48] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_51 
+ bl[49] br[49] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_52 
+ bl[50] br[50] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_53 
+ bl[51] br[51] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_54 
+ bl[52] br[52] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_55 
+ bl[53] br[53] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_56 
+ bl[54] br[54] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_57 
+ bl[55] br[55] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_58 
+ bl[56] br[56] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_59 
+ bl[57] br[57] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_60 
+ bl[58] br[58] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_61 
+ bl[59] br[59] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_62 
+ bl[60] br[60] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_63 
+ bl[61] br[61] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_64 
+ bl[62] br[62] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_65 
+ bl[63] br[63] vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_66 
+ vdd vdd vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_156_67 
+ vdd vdd vdd vss wl[154] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_0 
+ vdd vdd vss vdd vpb vnb wl[155] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_157_1 
+ rbl rbr vss vdd vpb vnb wl[155] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_157_2 
+ bl[0] br[0] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_3 
+ bl[1] br[1] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_4 
+ bl[2] br[2] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_5 
+ bl[3] br[3] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_6 
+ bl[4] br[4] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_7 
+ bl[5] br[5] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_8 
+ bl[6] br[6] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_9 
+ bl[7] br[7] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_10 
+ bl[8] br[8] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_11 
+ bl[9] br[9] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_12 
+ bl[10] br[10] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_13 
+ bl[11] br[11] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_14 
+ bl[12] br[12] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_15 
+ bl[13] br[13] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_16 
+ bl[14] br[14] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_17 
+ bl[15] br[15] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_18 
+ bl[16] br[16] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_19 
+ bl[17] br[17] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_20 
+ bl[18] br[18] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_21 
+ bl[19] br[19] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_22 
+ bl[20] br[20] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_23 
+ bl[21] br[21] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_24 
+ bl[22] br[22] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_25 
+ bl[23] br[23] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_26 
+ bl[24] br[24] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_27 
+ bl[25] br[25] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_28 
+ bl[26] br[26] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_29 
+ bl[27] br[27] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_30 
+ bl[28] br[28] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_31 
+ bl[29] br[29] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_32 
+ bl[30] br[30] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_33 
+ bl[31] br[31] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_34 
+ bl[32] br[32] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_35 
+ bl[33] br[33] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_36 
+ bl[34] br[34] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_37 
+ bl[35] br[35] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_38 
+ bl[36] br[36] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_39 
+ bl[37] br[37] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_40 
+ bl[38] br[38] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_41 
+ bl[39] br[39] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_42 
+ bl[40] br[40] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_43 
+ bl[41] br[41] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_44 
+ bl[42] br[42] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_45 
+ bl[43] br[43] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_46 
+ bl[44] br[44] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_47 
+ bl[45] br[45] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_48 
+ bl[46] br[46] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_49 
+ bl[47] br[47] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_50 
+ bl[48] br[48] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_51 
+ bl[49] br[49] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_52 
+ bl[50] br[50] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_53 
+ bl[51] br[51] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_54 
+ bl[52] br[52] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_55 
+ bl[53] br[53] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_56 
+ bl[54] br[54] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_57 
+ bl[55] br[55] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_58 
+ bl[56] br[56] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_59 
+ bl[57] br[57] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_60 
+ bl[58] br[58] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_61 
+ bl[59] br[59] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_62 
+ bl[60] br[60] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_63 
+ bl[61] br[61] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_64 
+ bl[62] br[62] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_65 
+ bl[63] br[63] vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_66 
+ vdd vdd vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_157_67 
+ vdd vdd vdd vss wl[155] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_0 
+ vdd vdd vss vdd vpb vnb wl[156] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_158_1 
+ rbl rbr vss vdd vpb vnb wl[156] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_158_2 
+ bl[0] br[0] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_3 
+ bl[1] br[1] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_4 
+ bl[2] br[2] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_5 
+ bl[3] br[3] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_6 
+ bl[4] br[4] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_7 
+ bl[5] br[5] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_8 
+ bl[6] br[6] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_9 
+ bl[7] br[7] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_10 
+ bl[8] br[8] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_11 
+ bl[9] br[9] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_12 
+ bl[10] br[10] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_13 
+ bl[11] br[11] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_14 
+ bl[12] br[12] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_15 
+ bl[13] br[13] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_16 
+ bl[14] br[14] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_17 
+ bl[15] br[15] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_18 
+ bl[16] br[16] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_19 
+ bl[17] br[17] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_20 
+ bl[18] br[18] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_21 
+ bl[19] br[19] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_22 
+ bl[20] br[20] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_23 
+ bl[21] br[21] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_24 
+ bl[22] br[22] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_25 
+ bl[23] br[23] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_26 
+ bl[24] br[24] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_27 
+ bl[25] br[25] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_28 
+ bl[26] br[26] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_29 
+ bl[27] br[27] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_30 
+ bl[28] br[28] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_31 
+ bl[29] br[29] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_32 
+ bl[30] br[30] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_33 
+ bl[31] br[31] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_34 
+ bl[32] br[32] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_35 
+ bl[33] br[33] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_36 
+ bl[34] br[34] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_37 
+ bl[35] br[35] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_38 
+ bl[36] br[36] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_39 
+ bl[37] br[37] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_40 
+ bl[38] br[38] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_41 
+ bl[39] br[39] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_42 
+ bl[40] br[40] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_43 
+ bl[41] br[41] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_44 
+ bl[42] br[42] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_45 
+ bl[43] br[43] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_46 
+ bl[44] br[44] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_47 
+ bl[45] br[45] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_48 
+ bl[46] br[46] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_49 
+ bl[47] br[47] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_50 
+ bl[48] br[48] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_51 
+ bl[49] br[49] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_52 
+ bl[50] br[50] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_53 
+ bl[51] br[51] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_54 
+ bl[52] br[52] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_55 
+ bl[53] br[53] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_56 
+ bl[54] br[54] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_57 
+ bl[55] br[55] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_58 
+ bl[56] br[56] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_59 
+ bl[57] br[57] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_60 
+ bl[58] br[58] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_61 
+ bl[59] br[59] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_62 
+ bl[60] br[60] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_63 
+ bl[61] br[61] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_64 
+ bl[62] br[62] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_65 
+ bl[63] br[63] vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_66 
+ vdd vdd vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_158_67 
+ vdd vdd vdd vss wl[156] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_0 
+ vdd vdd vss vdd vpb vnb wl[157] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_159_1 
+ rbl rbr vss vdd vpb vnb wl[157] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_159_2 
+ bl[0] br[0] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_3 
+ bl[1] br[1] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_4 
+ bl[2] br[2] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_5 
+ bl[3] br[3] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_6 
+ bl[4] br[4] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_7 
+ bl[5] br[5] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_8 
+ bl[6] br[6] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_9 
+ bl[7] br[7] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_10 
+ bl[8] br[8] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_11 
+ bl[9] br[9] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_12 
+ bl[10] br[10] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_13 
+ bl[11] br[11] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_14 
+ bl[12] br[12] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_15 
+ bl[13] br[13] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_16 
+ bl[14] br[14] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_17 
+ bl[15] br[15] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_18 
+ bl[16] br[16] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_19 
+ bl[17] br[17] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_20 
+ bl[18] br[18] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_21 
+ bl[19] br[19] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_22 
+ bl[20] br[20] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_23 
+ bl[21] br[21] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_24 
+ bl[22] br[22] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_25 
+ bl[23] br[23] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_26 
+ bl[24] br[24] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_27 
+ bl[25] br[25] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_28 
+ bl[26] br[26] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_29 
+ bl[27] br[27] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_30 
+ bl[28] br[28] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_31 
+ bl[29] br[29] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_32 
+ bl[30] br[30] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_33 
+ bl[31] br[31] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_34 
+ bl[32] br[32] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_35 
+ bl[33] br[33] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_36 
+ bl[34] br[34] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_37 
+ bl[35] br[35] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_38 
+ bl[36] br[36] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_39 
+ bl[37] br[37] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_40 
+ bl[38] br[38] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_41 
+ bl[39] br[39] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_42 
+ bl[40] br[40] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_43 
+ bl[41] br[41] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_44 
+ bl[42] br[42] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_45 
+ bl[43] br[43] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_46 
+ bl[44] br[44] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_47 
+ bl[45] br[45] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_48 
+ bl[46] br[46] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_49 
+ bl[47] br[47] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_50 
+ bl[48] br[48] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_51 
+ bl[49] br[49] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_52 
+ bl[50] br[50] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_53 
+ bl[51] br[51] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_54 
+ bl[52] br[52] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_55 
+ bl[53] br[53] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_56 
+ bl[54] br[54] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_57 
+ bl[55] br[55] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_58 
+ bl[56] br[56] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_59 
+ bl[57] br[57] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_60 
+ bl[58] br[58] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_61 
+ bl[59] br[59] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_62 
+ bl[60] br[60] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_63 
+ bl[61] br[61] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_64 
+ bl[62] br[62] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_65 
+ bl[63] br[63] vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_66 
+ vdd vdd vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_159_67 
+ vdd vdd vdd vss wl[157] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_0 
+ vdd vdd vss vdd vpb vnb wl[158] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_160_1 
+ rbl rbr vss vdd vpb vnb wl[158] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_160_2 
+ bl[0] br[0] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_3 
+ bl[1] br[1] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_4 
+ bl[2] br[2] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_5 
+ bl[3] br[3] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_6 
+ bl[4] br[4] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_7 
+ bl[5] br[5] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_8 
+ bl[6] br[6] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_9 
+ bl[7] br[7] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_10 
+ bl[8] br[8] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_11 
+ bl[9] br[9] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_12 
+ bl[10] br[10] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_13 
+ bl[11] br[11] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_14 
+ bl[12] br[12] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_15 
+ bl[13] br[13] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_16 
+ bl[14] br[14] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_17 
+ bl[15] br[15] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_18 
+ bl[16] br[16] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_19 
+ bl[17] br[17] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_20 
+ bl[18] br[18] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_21 
+ bl[19] br[19] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_22 
+ bl[20] br[20] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_23 
+ bl[21] br[21] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_24 
+ bl[22] br[22] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_25 
+ bl[23] br[23] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_26 
+ bl[24] br[24] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_27 
+ bl[25] br[25] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_28 
+ bl[26] br[26] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_29 
+ bl[27] br[27] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_30 
+ bl[28] br[28] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_31 
+ bl[29] br[29] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_32 
+ bl[30] br[30] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_33 
+ bl[31] br[31] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_34 
+ bl[32] br[32] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_35 
+ bl[33] br[33] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_36 
+ bl[34] br[34] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_37 
+ bl[35] br[35] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_38 
+ bl[36] br[36] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_39 
+ bl[37] br[37] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_40 
+ bl[38] br[38] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_41 
+ bl[39] br[39] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_42 
+ bl[40] br[40] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_43 
+ bl[41] br[41] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_44 
+ bl[42] br[42] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_45 
+ bl[43] br[43] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_46 
+ bl[44] br[44] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_47 
+ bl[45] br[45] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_48 
+ bl[46] br[46] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_49 
+ bl[47] br[47] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_50 
+ bl[48] br[48] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_51 
+ bl[49] br[49] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_52 
+ bl[50] br[50] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_53 
+ bl[51] br[51] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_54 
+ bl[52] br[52] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_55 
+ bl[53] br[53] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_56 
+ bl[54] br[54] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_57 
+ bl[55] br[55] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_58 
+ bl[56] br[56] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_59 
+ bl[57] br[57] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_60 
+ bl[58] br[58] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_61 
+ bl[59] br[59] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_62 
+ bl[60] br[60] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_63 
+ bl[61] br[61] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_64 
+ bl[62] br[62] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_65 
+ bl[63] br[63] vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_66 
+ vdd vdd vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_160_67 
+ vdd vdd vdd vss wl[158] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_0 
+ vdd vdd vss vdd vpb vnb wl[159] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_161_1 
+ rbl rbr vss vdd vpb vnb wl[159] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_161_2 
+ bl[0] br[0] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_3 
+ bl[1] br[1] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_4 
+ bl[2] br[2] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_5 
+ bl[3] br[3] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_6 
+ bl[4] br[4] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_7 
+ bl[5] br[5] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_8 
+ bl[6] br[6] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_9 
+ bl[7] br[7] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_10 
+ bl[8] br[8] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_11 
+ bl[9] br[9] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_12 
+ bl[10] br[10] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_13 
+ bl[11] br[11] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_14 
+ bl[12] br[12] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_15 
+ bl[13] br[13] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_16 
+ bl[14] br[14] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_17 
+ bl[15] br[15] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_18 
+ bl[16] br[16] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_19 
+ bl[17] br[17] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_20 
+ bl[18] br[18] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_21 
+ bl[19] br[19] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_22 
+ bl[20] br[20] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_23 
+ bl[21] br[21] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_24 
+ bl[22] br[22] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_25 
+ bl[23] br[23] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_26 
+ bl[24] br[24] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_27 
+ bl[25] br[25] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_28 
+ bl[26] br[26] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_29 
+ bl[27] br[27] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_30 
+ bl[28] br[28] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_31 
+ bl[29] br[29] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_32 
+ bl[30] br[30] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_33 
+ bl[31] br[31] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_34 
+ bl[32] br[32] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_35 
+ bl[33] br[33] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_36 
+ bl[34] br[34] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_37 
+ bl[35] br[35] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_38 
+ bl[36] br[36] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_39 
+ bl[37] br[37] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_40 
+ bl[38] br[38] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_41 
+ bl[39] br[39] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_42 
+ bl[40] br[40] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_43 
+ bl[41] br[41] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_44 
+ bl[42] br[42] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_45 
+ bl[43] br[43] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_46 
+ bl[44] br[44] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_47 
+ bl[45] br[45] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_48 
+ bl[46] br[46] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_49 
+ bl[47] br[47] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_50 
+ bl[48] br[48] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_51 
+ bl[49] br[49] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_52 
+ bl[50] br[50] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_53 
+ bl[51] br[51] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_54 
+ bl[52] br[52] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_55 
+ bl[53] br[53] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_56 
+ bl[54] br[54] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_57 
+ bl[55] br[55] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_58 
+ bl[56] br[56] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_59 
+ bl[57] br[57] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_60 
+ bl[58] br[58] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_61 
+ bl[59] br[59] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_62 
+ bl[60] br[60] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_63 
+ bl[61] br[61] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_64 
+ bl[62] br[62] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_65 
+ bl[63] br[63] vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_66 
+ vdd vdd vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_161_67 
+ vdd vdd vdd vss wl[159] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_0 
+ vdd vdd vss vdd vpb vnb wl[160] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_162_1 
+ rbl rbr vss vdd vpb vnb wl[160] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_162_2 
+ bl[0] br[0] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_3 
+ bl[1] br[1] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_4 
+ bl[2] br[2] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_5 
+ bl[3] br[3] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_6 
+ bl[4] br[4] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_7 
+ bl[5] br[5] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_8 
+ bl[6] br[6] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_9 
+ bl[7] br[7] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_10 
+ bl[8] br[8] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_11 
+ bl[9] br[9] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_12 
+ bl[10] br[10] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_13 
+ bl[11] br[11] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_14 
+ bl[12] br[12] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_15 
+ bl[13] br[13] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_16 
+ bl[14] br[14] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_17 
+ bl[15] br[15] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_18 
+ bl[16] br[16] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_19 
+ bl[17] br[17] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_20 
+ bl[18] br[18] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_21 
+ bl[19] br[19] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_22 
+ bl[20] br[20] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_23 
+ bl[21] br[21] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_24 
+ bl[22] br[22] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_25 
+ bl[23] br[23] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_26 
+ bl[24] br[24] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_27 
+ bl[25] br[25] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_28 
+ bl[26] br[26] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_29 
+ bl[27] br[27] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_30 
+ bl[28] br[28] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_31 
+ bl[29] br[29] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_32 
+ bl[30] br[30] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_33 
+ bl[31] br[31] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_34 
+ bl[32] br[32] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_35 
+ bl[33] br[33] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_36 
+ bl[34] br[34] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_37 
+ bl[35] br[35] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_38 
+ bl[36] br[36] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_39 
+ bl[37] br[37] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_40 
+ bl[38] br[38] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_41 
+ bl[39] br[39] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_42 
+ bl[40] br[40] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_43 
+ bl[41] br[41] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_44 
+ bl[42] br[42] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_45 
+ bl[43] br[43] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_46 
+ bl[44] br[44] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_47 
+ bl[45] br[45] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_48 
+ bl[46] br[46] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_49 
+ bl[47] br[47] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_50 
+ bl[48] br[48] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_51 
+ bl[49] br[49] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_52 
+ bl[50] br[50] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_53 
+ bl[51] br[51] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_54 
+ bl[52] br[52] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_55 
+ bl[53] br[53] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_56 
+ bl[54] br[54] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_57 
+ bl[55] br[55] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_58 
+ bl[56] br[56] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_59 
+ bl[57] br[57] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_60 
+ bl[58] br[58] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_61 
+ bl[59] br[59] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_62 
+ bl[60] br[60] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_63 
+ bl[61] br[61] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_64 
+ bl[62] br[62] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_65 
+ bl[63] br[63] vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_66 
+ vdd vdd vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_162_67 
+ vdd vdd vdd vss wl[160] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_0 
+ vdd vdd vss vdd vpb vnb wl[161] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_163_1 
+ rbl rbr vss vdd vpb vnb wl[161] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_163_2 
+ bl[0] br[0] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_3 
+ bl[1] br[1] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_4 
+ bl[2] br[2] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_5 
+ bl[3] br[3] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_6 
+ bl[4] br[4] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_7 
+ bl[5] br[5] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_8 
+ bl[6] br[6] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_9 
+ bl[7] br[7] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_10 
+ bl[8] br[8] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_11 
+ bl[9] br[9] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_12 
+ bl[10] br[10] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_13 
+ bl[11] br[11] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_14 
+ bl[12] br[12] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_15 
+ bl[13] br[13] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_16 
+ bl[14] br[14] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_17 
+ bl[15] br[15] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_18 
+ bl[16] br[16] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_19 
+ bl[17] br[17] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_20 
+ bl[18] br[18] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_21 
+ bl[19] br[19] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_22 
+ bl[20] br[20] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_23 
+ bl[21] br[21] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_24 
+ bl[22] br[22] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_25 
+ bl[23] br[23] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_26 
+ bl[24] br[24] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_27 
+ bl[25] br[25] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_28 
+ bl[26] br[26] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_29 
+ bl[27] br[27] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_30 
+ bl[28] br[28] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_31 
+ bl[29] br[29] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_32 
+ bl[30] br[30] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_33 
+ bl[31] br[31] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_34 
+ bl[32] br[32] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_35 
+ bl[33] br[33] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_36 
+ bl[34] br[34] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_37 
+ bl[35] br[35] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_38 
+ bl[36] br[36] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_39 
+ bl[37] br[37] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_40 
+ bl[38] br[38] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_41 
+ bl[39] br[39] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_42 
+ bl[40] br[40] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_43 
+ bl[41] br[41] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_44 
+ bl[42] br[42] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_45 
+ bl[43] br[43] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_46 
+ bl[44] br[44] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_47 
+ bl[45] br[45] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_48 
+ bl[46] br[46] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_49 
+ bl[47] br[47] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_50 
+ bl[48] br[48] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_51 
+ bl[49] br[49] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_52 
+ bl[50] br[50] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_53 
+ bl[51] br[51] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_54 
+ bl[52] br[52] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_55 
+ bl[53] br[53] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_56 
+ bl[54] br[54] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_57 
+ bl[55] br[55] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_58 
+ bl[56] br[56] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_59 
+ bl[57] br[57] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_60 
+ bl[58] br[58] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_61 
+ bl[59] br[59] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_62 
+ bl[60] br[60] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_63 
+ bl[61] br[61] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_64 
+ bl[62] br[62] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_65 
+ bl[63] br[63] vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_66 
+ vdd vdd vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_163_67 
+ vdd vdd vdd vss wl[161] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_0 
+ vdd vdd vss vdd vpb vnb wl[162] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_164_1 
+ rbl rbr vss vdd vpb vnb wl[162] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_164_2 
+ bl[0] br[0] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_3 
+ bl[1] br[1] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_4 
+ bl[2] br[2] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_5 
+ bl[3] br[3] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_6 
+ bl[4] br[4] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_7 
+ bl[5] br[5] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_8 
+ bl[6] br[6] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_9 
+ bl[7] br[7] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_10 
+ bl[8] br[8] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_11 
+ bl[9] br[9] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_12 
+ bl[10] br[10] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_13 
+ bl[11] br[11] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_14 
+ bl[12] br[12] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_15 
+ bl[13] br[13] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_16 
+ bl[14] br[14] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_17 
+ bl[15] br[15] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_18 
+ bl[16] br[16] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_19 
+ bl[17] br[17] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_20 
+ bl[18] br[18] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_21 
+ bl[19] br[19] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_22 
+ bl[20] br[20] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_23 
+ bl[21] br[21] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_24 
+ bl[22] br[22] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_25 
+ bl[23] br[23] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_26 
+ bl[24] br[24] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_27 
+ bl[25] br[25] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_28 
+ bl[26] br[26] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_29 
+ bl[27] br[27] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_30 
+ bl[28] br[28] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_31 
+ bl[29] br[29] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_32 
+ bl[30] br[30] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_33 
+ bl[31] br[31] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_34 
+ bl[32] br[32] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_35 
+ bl[33] br[33] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_36 
+ bl[34] br[34] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_37 
+ bl[35] br[35] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_38 
+ bl[36] br[36] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_39 
+ bl[37] br[37] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_40 
+ bl[38] br[38] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_41 
+ bl[39] br[39] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_42 
+ bl[40] br[40] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_43 
+ bl[41] br[41] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_44 
+ bl[42] br[42] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_45 
+ bl[43] br[43] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_46 
+ bl[44] br[44] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_47 
+ bl[45] br[45] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_48 
+ bl[46] br[46] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_49 
+ bl[47] br[47] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_50 
+ bl[48] br[48] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_51 
+ bl[49] br[49] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_52 
+ bl[50] br[50] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_53 
+ bl[51] br[51] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_54 
+ bl[52] br[52] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_55 
+ bl[53] br[53] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_56 
+ bl[54] br[54] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_57 
+ bl[55] br[55] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_58 
+ bl[56] br[56] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_59 
+ bl[57] br[57] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_60 
+ bl[58] br[58] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_61 
+ bl[59] br[59] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_62 
+ bl[60] br[60] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_63 
+ bl[61] br[61] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_64 
+ bl[62] br[62] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_65 
+ bl[63] br[63] vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_66 
+ vdd vdd vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_164_67 
+ vdd vdd vdd vss wl[162] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_0 
+ vdd vdd vss vdd vpb vnb wl[163] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_165_1 
+ rbl rbr vss vdd vpb vnb wl[163] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_165_2 
+ bl[0] br[0] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_3 
+ bl[1] br[1] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_4 
+ bl[2] br[2] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_5 
+ bl[3] br[3] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_6 
+ bl[4] br[4] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_7 
+ bl[5] br[5] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_8 
+ bl[6] br[6] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_9 
+ bl[7] br[7] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_10 
+ bl[8] br[8] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_11 
+ bl[9] br[9] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_12 
+ bl[10] br[10] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_13 
+ bl[11] br[11] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_14 
+ bl[12] br[12] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_15 
+ bl[13] br[13] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_16 
+ bl[14] br[14] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_17 
+ bl[15] br[15] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_18 
+ bl[16] br[16] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_19 
+ bl[17] br[17] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_20 
+ bl[18] br[18] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_21 
+ bl[19] br[19] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_22 
+ bl[20] br[20] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_23 
+ bl[21] br[21] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_24 
+ bl[22] br[22] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_25 
+ bl[23] br[23] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_26 
+ bl[24] br[24] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_27 
+ bl[25] br[25] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_28 
+ bl[26] br[26] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_29 
+ bl[27] br[27] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_30 
+ bl[28] br[28] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_31 
+ bl[29] br[29] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_32 
+ bl[30] br[30] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_33 
+ bl[31] br[31] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_34 
+ bl[32] br[32] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_35 
+ bl[33] br[33] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_36 
+ bl[34] br[34] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_37 
+ bl[35] br[35] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_38 
+ bl[36] br[36] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_39 
+ bl[37] br[37] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_40 
+ bl[38] br[38] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_41 
+ bl[39] br[39] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_42 
+ bl[40] br[40] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_43 
+ bl[41] br[41] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_44 
+ bl[42] br[42] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_45 
+ bl[43] br[43] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_46 
+ bl[44] br[44] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_47 
+ bl[45] br[45] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_48 
+ bl[46] br[46] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_49 
+ bl[47] br[47] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_50 
+ bl[48] br[48] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_51 
+ bl[49] br[49] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_52 
+ bl[50] br[50] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_53 
+ bl[51] br[51] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_54 
+ bl[52] br[52] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_55 
+ bl[53] br[53] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_56 
+ bl[54] br[54] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_57 
+ bl[55] br[55] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_58 
+ bl[56] br[56] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_59 
+ bl[57] br[57] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_60 
+ bl[58] br[58] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_61 
+ bl[59] br[59] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_62 
+ bl[60] br[60] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_63 
+ bl[61] br[61] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_64 
+ bl[62] br[62] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_65 
+ bl[63] br[63] vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_66 
+ vdd vdd vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_165_67 
+ vdd vdd vdd vss wl[163] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_0 
+ vdd vdd vss vdd vpb vnb wl[164] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_166_1 
+ rbl rbr vss vdd vpb vnb wl[164] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_166_2 
+ bl[0] br[0] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_3 
+ bl[1] br[1] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_4 
+ bl[2] br[2] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_5 
+ bl[3] br[3] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_6 
+ bl[4] br[4] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_7 
+ bl[5] br[5] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_8 
+ bl[6] br[6] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_9 
+ bl[7] br[7] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_10 
+ bl[8] br[8] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_11 
+ bl[9] br[9] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_12 
+ bl[10] br[10] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_13 
+ bl[11] br[11] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_14 
+ bl[12] br[12] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_15 
+ bl[13] br[13] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_16 
+ bl[14] br[14] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_17 
+ bl[15] br[15] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_18 
+ bl[16] br[16] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_19 
+ bl[17] br[17] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_20 
+ bl[18] br[18] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_21 
+ bl[19] br[19] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_22 
+ bl[20] br[20] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_23 
+ bl[21] br[21] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_24 
+ bl[22] br[22] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_25 
+ bl[23] br[23] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_26 
+ bl[24] br[24] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_27 
+ bl[25] br[25] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_28 
+ bl[26] br[26] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_29 
+ bl[27] br[27] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_30 
+ bl[28] br[28] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_31 
+ bl[29] br[29] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_32 
+ bl[30] br[30] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_33 
+ bl[31] br[31] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_34 
+ bl[32] br[32] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_35 
+ bl[33] br[33] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_36 
+ bl[34] br[34] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_37 
+ bl[35] br[35] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_38 
+ bl[36] br[36] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_39 
+ bl[37] br[37] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_40 
+ bl[38] br[38] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_41 
+ bl[39] br[39] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_42 
+ bl[40] br[40] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_43 
+ bl[41] br[41] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_44 
+ bl[42] br[42] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_45 
+ bl[43] br[43] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_46 
+ bl[44] br[44] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_47 
+ bl[45] br[45] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_48 
+ bl[46] br[46] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_49 
+ bl[47] br[47] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_50 
+ bl[48] br[48] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_51 
+ bl[49] br[49] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_52 
+ bl[50] br[50] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_53 
+ bl[51] br[51] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_54 
+ bl[52] br[52] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_55 
+ bl[53] br[53] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_56 
+ bl[54] br[54] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_57 
+ bl[55] br[55] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_58 
+ bl[56] br[56] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_59 
+ bl[57] br[57] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_60 
+ bl[58] br[58] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_61 
+ bl[59] br[59] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_62 
+ bl[60] br[60] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_63 
+ bl[61] br[61] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_64 
+ bl[62] br[62] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_65 
+ bl[63] br[63] vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_66 
+ vdd vdd vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_166_67 
+ vdd vdd vdd vss wl[164] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_0 
+ vdd vdd vss vdd vpb vnb wl[165] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_167_1 
+ rbl rbr vss vdd vpb vnb wl[165] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_167_2 
+ bl[0] br[0] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_3 
+ bl[1] br[1] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_4 
+ bl[2] br[2] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_5 
+ bl[3] br[3] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_6 
+ bl[4] br[4] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_7 
+ bl[5] br[5] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_8 
+ bl[6] br[6] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_9 
+ bl[7] br[7] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_10 
+ bl[8] br[8] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_11 
+ bl[9] br[9] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_12 
+ bl[10] br[10] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_13 
+ bl[11] br[11] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_14 
+ bl[12] br[12] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_15 
+ bl[13] br[13] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_16 
+ bl[14] br[14] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_17 
+ bl[15] br[15] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_18 
+ bl[16] br[16] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_19 
+ bl[17] br[17] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_20 
+ bl[18] br[18] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_21 
+ bl[19] br[19] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_22 
+ bl[20] br[20] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_23 
+ bl[21] br[21] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_24 
+ bl[22] br[22] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_25 
+ bl[23] br[23] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_26 
+ bl[24] br[24] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_27 
+ bl[25] br[25] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_28 
+ bl[26] br[26] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_29 
+ bl[27] br[27] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_30 
+ bl[28] br[28] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_31 
+ bl[29] br[29] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_32 
+ bl[30] br[30] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_33 
+ bl[31] br[31] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_34 
+ bl[32] br[32] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_35 
+ bl[33] br[33] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_36 
+ bl[34] br[34] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_37 
+ bl[35] br[35] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_38 
+ bl[36] br[36] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_39 
+ bl[37] br[37] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_40 
+ bl[38] br[38] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_41 
+ bl[39] br[39] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_42 
+ bl[40] br[40] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_43 
+ bl[41] br[41] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_44 
+ bl[42] br[42] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_45 
+ bl[43] br[43] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_46 
+ bl[44] br[44] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_47 
+ bl[45] br[45] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_48 
+ bl[46] br[46] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_49 
+ bl[47] br[47] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_50 
+ bl[48] br[48] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_51 
+ bl[49] br[49] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_52 
+ bl[50] br[50] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_53 
+ bl[51] br[51] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_54 
+ bl[52] br[52] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_55 
+ bl[53] br[53] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_56 
+ bl[54] br[54] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_57 
+ bl[55] br[55] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_58 
+ bl[56] br[56] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_59 
+ bl[57] br[57] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_60 
+ bl[58] br[58] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_61 
+ bl[59] br[59] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_62 
+ bl[60] br[60] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_63 
+ bl[61] br[61] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_64 
+ bl[62] br[62] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_65 
+ bl[63] br[63] vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_66 
+ vdd vdd vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_167_67 
+ vdd vdd vdd vss wl[165] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_0 
+ vdd vdd vss vdd vpb vnb wl[166] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_168_1 
+ rbl rbr vss vdd vpb vnb wl[166] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_168_2 
+ bl[0] br[0] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_3 
+ bl[1] br[1] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_4 
+ bl[2] br[2] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_5 
+ bl[3] br[3] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_6 
+ bl[4] br[4] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_7 
+ bl[5] br[5] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_8 
+ bl[6] br[6] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_9 
+ bl[7] br[7] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_10 
+ bl[8] br[8] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_11 
+ bl[9] br[9] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_12 
+ bl[10] br[10] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_13 
+ bl[11] br[11] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_14 
+ bl[12] br[12] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_15 
+ bl[13] br[13] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_16 
+ bl[14] br[14] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_17 
+ bl[15] br[15] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_18 
+ bl[16] br[16] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_19 
+ bl[17] br[17] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_20 
+ bl[18] br[18] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_21 
+ bl[19] br[19] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_22 
+ bl[20] br[20] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_23 
+ bl[21] br[21] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_24 
+ bl[22] br[22] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_25 
+ bl[23] br[23] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_26 
+ bl[24] br[24] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_27 
+ bl[25] br[25] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_28 
+ bl[26] br[26] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_29 
+ bl[27] br[27] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_30 
+ bl[28] br[28] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_31 
+ bl[29] br[29] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_32 
+ bl[30] br[30] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_33 
+ bl[31] br[31] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_34 
+ bl[32] br[32] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_35 
+ bl[33] br[33] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_36 
+ bl[34] br[34] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_37 
+ bl[35] br[35] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_38 
+ bl[36] br[36] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_39 
+ bl[37] br[37] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_40 
+ bl[38] br[38] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_41 
+ bl[39] br[39] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_42 
+ bl[40] br[40] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_43 
+ bl[41] br[41] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_44 
+ bl[42] br[42] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_45 
+ bl[43] br[43] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_46 
+ bl[44] br[44] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_47 
+ bl[45] br[45] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_48 
+ bl[46] br[46] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_49 
+ bl[47] br[47] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_50 
+ bl[48] br[48] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_51 
+ bl[49] br[49] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_52 
+ bl[50] br[50] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_53 
+ bl[51] br[51] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_54 
+ bl[52] br[52] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_55 
+ bl[53] br[53] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_56 
+ bl[54] br[54] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_57 
+ bl[55] br[55] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_58 
+ bl[56] br[56] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_59 
+ bl[57] br[57] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_60 
+ bl[58] br[58] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_61 
+ bl[59] br[59] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_62 
+ bl[60] br[60] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_63 
+ bl[61] br[61] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_64 
+ bl[62] br[62] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_65 
+ bl[63] br[63] vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_66 
+ vdd vdd vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_168_67 
+ vdd vdd vdd vss wl[166] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_0 
+ vdd vdd vss vdd vpb vnb wl[167] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_169_1 
+ rbl rbr vss vdd vpb vnb wl[167] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_169_2 
+ bl[0] br[0] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_3 
+ bl[1] br[1] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_4 
+ bl[2] br[2] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_5 
+ bl[3] br[3] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_6 
+ bl[4] br[4] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_7 
+ bl[5] br[5] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_8 
+ bl[6] br[6] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_9 
+ bl[7] br[7] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_10 
+ bl[8] br[8] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_11 
+ bl[9] br[9] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_12 
+ bl[10] br[10] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_13 
+ bl[11] br[11] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_14 
+ bl[12] br[12] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_15 
+ bl[13] br[13] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_16 
+ bl[14] br[14] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_17 
+ bl[15] br[15] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_18 
+ bl[16] br[16] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_19 
+ bl[17] br[17] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_20 
+ bl[18] br[18] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_21 
+ bl[19] br[19] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_22 
+ bl[20] br[20] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_23 
+ bl[21] br[21] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_24 
+ bl[22] br[22] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_25 
+ bl[23] br[23] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_26 
+ bl[24] br[24] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_27 
+ bl[25] br[25] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_28 
+ bl[26] br[26] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_29 
+ bl[27] br[27] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_30 
+ bl[28] br[28] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_31 
+ bl[29] br[29] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_32 
+ bl[30] br[30] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_33 
+ bl[31] br[31] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_34 
+ bl[32] br[32] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_35 
+ bl[33] br[33] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_36 
+ bl[34] br[34] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_37 
+ bl[35] br[35] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_38 
+ bl[36] br[36] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_39 
+ bl[37] br[37] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_40 
+ bl[38] br[38] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_41 
+ bl[39] br[39] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_42 
+ bl[40] br[40] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_43 
+ bl[41] br[41] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_44 
+ bl[42] br[42] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_45 
+ bl[43] br[43] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_46 
+ bl[44] br[44] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_47 
+ bl[45] br[45] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_48 
+ bl[46] br[46] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_49 
+ bl[47] br[47] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_50 
+ bl[48] br[48] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_51 
+ bl[49] br[49] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_52 
+ bl[50] br[50] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_53 
+ bl[51] br[51] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_54 
+ bl[52] br[52] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_55 
+ bl[53] br[53] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_56 
+ bl[54] br[54] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_57 
+ bl[55] br[55] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_58 
+ bl[56] br[56] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_59 
+ bl[57] br[57] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_60 
+ bl[58] br[58] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_61 
+ bl[59] br[59] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_62 
+ bl[60] br[60] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_63 
+ bl[61] br[61] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_64 
+ bl[62] br[62] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_65 
+ bl[63] br[63] vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_66 
+ vdd vdd vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_169_67 
+ vdd vdd vdd vss wl[167] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_0 
+ vdd vdd vss vdd vpb vnb wl[168] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_170_1 
+ rbl rbr vss vdd vpb vnb wl[168] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_170_2 
+ bl[0] br[0] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_3 
+ bl[1] br[1] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_4 
+ bl[2] br[2] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_5 
+ bl[3] br[3] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_6 
+ bl[4] br[4] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_7 
+ bl[5] br[5] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_8 
+ bl[6] br[6] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_9 
+ bl[7] br[7] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_10 
+ bl[8] br[8] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_11 
+ bl[9] br[9] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_12 
+ bl[10] br[10] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_13 
+ bl[11] br[11] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_14 
+ bl[12] br[12] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_15 
+ bl[13] br[13] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_16 
+ bl[14] br[14] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_17 
+ bl[15] br[15] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_18 
+ bl[16] br[16] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_19 
+ bl[17] br[17] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_20 
+ bl[18] br[18] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_21 
+ bl[19] br[19] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_22 
+ bl[20] br[20] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_23 
+ bl[21] br[21] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_24 
+ bl[22] br[22] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_25 
+ bl[23] br[23] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_26 
+ bl[24] br[24] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_27 
+ bl[25] br[25] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_28 
+ bl[26] br[26] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_29 
+ bl[27] br[27] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_30 
+ bl[28] br[28] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_31 
+ bl[29] br[29] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_32 
+ bl[30] br[30] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_33 
+ bl[31] br[31] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_34 
+ bl[32] br[32] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_35 
+ bl[33] br[33] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_36 
+ bl[34] br[34] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_37 
+ bl[35] br[35] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_38 
+ bl[36] br[36] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_39 
+ bl[37] br[37] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_40 
+ bl[38] br[38] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_41 
+ bl[39] br[39] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_42 
+ bl[40] br[40] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_43 
+ bl[41] br[41] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_44 
+ bl[42] br[42] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_45 
+ bl[43] br[43] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_46 
+ bl[44] br[44] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_47 
+ bl[45] br[45] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_48 
+ bl[46] br[46] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_49 
+ bl[47] br[47] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_50 
+ bl[48] br[48] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_51 
+ bl[49] br[49] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_52 
+ bl[50] br[50] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_53 
+ bl[51] br[51] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_54 
+ bl[52] br[52] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_55 
+ bl[53] br[53] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_56 
+ bl[54] br[54] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_57 
+ bl[55] br[55] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_58 
+ bl[56] br[56] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_59 
+ bl[57] br[57] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_60 
+ bl[58] br[58] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_61 
+ bl[59] br[59] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_62 
+ bl[60] br[60] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_63 
+ bl[61] br[61] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_64 
+ bl[62] br[62] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_65 
+ bl[63] br[63] vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_66 
+ vdd vdd vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_170_67 
+ vdd vdd vdd vss wl[168] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_0 
+ vdd vdd vss vdd vpb vnb wl[169] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_171_1 
+ rbl rbr vss vdd vpb vnb wl[169] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_171_2 
+ bl[0] br[0] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_3 
+ bl[1] br[1] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_4 
+ bl[2] br[2] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_5 
+ bl[3] br[3] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_6 
+ bl[4] br[4] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_7 
+ bl[5] br[5] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_8 
+ bl[6] br[6] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_9 
+ bl[7] br[7] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_10 
+ bl[8] br[8] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_11 
+ bl[9] br[9] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_12 
+ bl[10] br[10] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_13 
+ bl[11] br[11] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_14 
+ bl[12] br[12] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_15 
+ bl[13] br[13] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_16 
+ bl[14] br[14] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_17 
+ bl[15] br[15] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_18 
+ bl[16] br[16] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_19 
+ bl[17] br[17] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_20 
+ bl[18] br[18] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_21 
+ bl[19] br[19] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_22 
+ bl[20] br[20] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_23 
+ bl[21] br[21] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_24 
+ bl[22] br[22] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_25 
+ bl[23] br[23] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_26 
+ bl[24] br[24] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_27 
+ bl[25] br[25] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_28 
+ bl[26] br[26] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_29 
+ bl[27] br[27] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_30 
+ bl[28] br[28] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_31 
+ bl[29] br[29] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_32 
+ bl[30] br[30] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_33 
+ bl[31] br[31] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_34 
+ bl[32] br[32] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_35 
+ bl[33] br[33] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_36 
+ bl[34] br[34] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_37 
+ bl[35] br[35] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_38 
+ bl[36] br[36] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_39 
+ bl[37] br[37] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_40 
+ bl[38] br[38] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_41 
+ bl[39] br[39] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_42 
+ bl[40] br[40] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_43 
+ bl[41] br[41] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_44 
+ bl[42] br[42] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_45 
+ bl[43] br[43] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_46 
+ bl[44] br[44] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_47 
+ bl[45] br[45] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_48 
+ bl[46] br[46] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_49 
+ bl[47] br[47] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_50 
+ bl[48] br[48] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_51 
+ bl[49] br[49] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_52 
+ bl[50] br[50] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_53 
+ bl[51] br[51] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_54 
+ bl[52] br[52] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_55 
+ bl[53] br[53] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_56 
+ bl[54] br[54] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_57 
+ bl[55] br[55] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_58 
+ bl[56] br[56] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_59 
+ bl[57] br[57] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_60 
+ bl[58] br[58] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_61 
+ bl[59] br[59] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_62 
+ bl[60] br[60] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_63 
+ bl[61] br[61] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_64 
+ bl[62] br[62] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_65 
+ bl[63] br[63] vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_66 
+ vdd vdd vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_171_67 
+ vdd vdd vdd vss wl[169] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_0 
+ vdd vdd vss vdd vpb vnb wl[170] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_172_1 
+ rbl rbr vss vdd vpb vnb wl[170] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_172_2 
+ bl[0] br[0] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_3 
+ bl[1] br[1] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_4 
+ bl[2] br[2] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_5 
+ bl[3] br[3] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_6 
+ bl[4] br[4] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_7 
+ bl[5] br[5] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_8 
+ bl[6] br[6] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_9 
+ bl[7] br[7] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_10 
+ bl[8] br[8] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_11 
+ bl[9] br[9] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_12 
+ bl[10] br[10] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_13 
+ bl[11] br[11] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_14 
+ bl[12] br[12] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_15 
+ bl[13] br[13] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_16 
+ bl[14] br[14] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_17 
+ bl[15] br[15] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_18 
+ bl[16] br[16] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_19 
+ bl[17] br[17] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_20 
+ bl[18] br[18] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_21 
+ bl[19] br[19] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_22 
+ bl[20] br[20] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_23 
+ bl[21] br[21] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_24 
+ bl[22] br[22] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_25 
+ bl[23] br[23] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_26 
+ bl[24] br[24] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_27 
+ bl[25] br[25] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_28 
+ bl[26] br[26] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_29 
+ bl[27] br[27] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_30 
+ bl[28] br[28] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_31 
+ bl[29] br[29] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_32 
+ bl[30] br[30] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_33 
+ bl[31] br[31] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_34 
+ bl[32] br[32] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_35 
+ bl[33] br[33] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_36 
+ bl[34] br[34] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_37 
+ bl[35] br[35] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_38 
+ bl[36] br[36] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_39 
+ bl[37] br[37] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_40 
+ bl[38] br[38] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_41 
+ bl[39] br[39] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_42 
+ bl[40] br[40] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_43 
+ bl[41] br[41] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_44 
+ bl[42] br[42] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_45 
+ bl[43] br[43] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_46 
+ bl[44] br[44] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_47 
+ bl[45] br[45] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_48 
+ bl[46] br[46] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_49 
+ bl[47] br[47] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_50 
+ bl[48] br[48] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_51 
+ bl[49] br[49] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_52 
+ bl[50] br[50] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_53 
+ bl[51] br[51] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_54 
+ bl[52] br[52] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_55 
+ bl[53] br[53] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_56 
+ bl[54] br[54] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_57 
+ bl[55] br[55] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_58 
+ bl[56] br[56] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_59 
+ bl[57] br[57] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_60 
+ bl[58] br[58] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_61 
+ bl[59] br[59] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_62 
+ bl[60] br[60] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_63 
+ bl[61] br[61] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_64 
+ bl[62] br[62] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_65 
+ bl[63] br[63] vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_66 
+ vdd vdd vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_172_67 
+ vdd vdd vdd vss wl[170] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_0 
+ vdd vdd vss vdd vpb vnb wl[171] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_173_1 
+ rbl rbr vss vdd vpb vnb wl[171] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_173_2 
+ bl[0] br[0] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_3 
+ bl[1] br[1] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_4 
+ bl[2] br[2] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_5 
+ bl[3] br[3] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_6 
+ bl[4] br[4] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_7 
+ bl[5] br[5] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_8 
+ bl[6] br[6] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_9 
+ bl[7] br[7] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_10 
+ bl[8] br[8] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_11 
+ bl[9] br[9] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_12 
+ bl[10] br[10] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_13 
+ bl[11] br[11] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_14 
+ bl[12] br[12] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_15 
+ bl[13] br[13] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_16 
+ bl[14] br[14] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_17 
+ bl[15] br[15] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_18 
+ bl[16] br[16] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_19 
+ bl[17] br[17] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_20 
+ bl[18] br[18] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_21 
+ bl[19] br[19] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_22 
+ bl[20] br[20] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_23 
+ bl[21] br[21] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_24 
+ bl[22] br[22] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_25 
+ bl[23] br[23] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_26 
+ bl[24] br[24] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_27 
+ bl[25] br[25] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_28 
+ bl[26] br[26] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_29 
+ bl[27] br[27] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_30 
+ bl[28] br[28] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_31 
+ bl[29] br[29] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_32 
+ bl[30] br[30] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_33 
+ bl[31] br[31] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_34 
+ bl[32] br[32] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_35 
+ bl[33] br[33] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_36 
+ bl[34] br[34] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_37 
+ bl[35] br[35] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_38 
+ bl[36] br[36] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_39 
+ bl[37] br[37] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_40 
+ bl[38] br[38] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_41 
+ bl[39] br[39] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_42 
+ bl[40] br[40] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_43 
+ bl[41] br[41] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_44 
+ bl[42] br[42] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_45 
+ bl[43] br[43] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_46 
+ bl[44] br[44] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_47 
+ bl[45] br[45] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_48 
+ bl[46] br[46] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_49 
+ bl[47] br[47] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_50 
+ bl[48] br[48] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_51 
+ bl[49] br[49] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_52 
+ bl[50] br[50] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_53 
+ bl[51] br[51] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_54 
+ bl[52] br[52] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_55 
+ bl[53] br[53] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_56 
+ bl[54] br[54] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_57 
+ bl[55] br[55] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_58 
+ bl[56] br[56] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_59 
+ bl[57] br[57] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_60 
+ bl[58] br[58] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_61 
+ bl[59] br[59] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_62 
+ bl[60] br[60] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_63 
+ bl[61] br[61] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_64 
+ bl[62] br[62] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_65 
+ bl[63] br[63] vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_66 
+ vdd vdd vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_173_67 
+ vdd vdd vdd vss wl[171] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_0 
+ vdd vdd vss vdd vpb vnb wl[172] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_174_1 
+ rbl rbr vss vdd vpb vnb wl[172] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_174_2 
+ bl[0] br[0] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_3 
+ bl[1] br[1] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_4 
+ bl[2] br[2] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_5 
+ bl[3] br[3] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_6 
+ bl[4] br[4] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_7 
+ bl[5] br[5] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_8 
+ bl[6] br[6] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_9 
+ bl[7] br[7] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_10 
+ bl[8] br[8] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_11 
+ bl[9] br[9] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_12 
+ bl[10] br[10] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_13 
+ bl[11] br[11] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_14 
+ bl[12] br[12] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_15 
+ bl[13] br[13] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_16 
+ bl[14] br[14] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_17 
+ bl[15] br[15] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_18 
+ bl[16] br[16] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_19 
+ bl[17] br[17] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_20 
+ bl[18] br[18] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_21 
+ bl[19] br[19] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_22 
+ bl[20] br[20] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_23 
+ bl[21] br[21] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_24 
+ bl[22] br[22] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_25 
+ bl[23] br[23] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_26 
+ bl[24] br[24] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_27 
+ bl[25] br[25] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_28 
+ bl[26] br[26] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_29 
+ bl[27] br[27] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_30 
+ bl[28] br[28] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_31 
+ bl[29] br[29] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_32 
+ bl[30] br[30] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_33 
+ bl[31] br[31] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_34 
+ bl[32] br[32] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_35 
+ bl[33] br[33] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_36 
+ bl[34] br[34] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_37 
+ bl[35] br[35] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_38 
+ bl[36] br[36] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_39 
+ bl[37] br[37] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_40 
+ bl[38] br[38] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_41 
+ bl[39] br[39] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_42 
+ bl[40] br[40] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_43 
+ bl[41] br[41] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_44 
+ bl[42] br[42] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_45 
+ bl[43] br[43] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_46 
+ bl[44] br[44] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_47 
+ bl[45] br[45] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_48 
+ bl[46] br[46] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_49 
+ bl[47] br[47] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_50 
+ bl[48] br[48] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_51 
+ bl[49] br[49] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_52 
+ bl[50] br[50] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_53 
+ bl[51] br[51] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_54 
+ bl[52] br[52] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_55 
+ bl[53] br[53] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_56 
+ bl[54] br[54] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_57 
+ bl[55] br[55] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_58 
+ bl[56] br[56] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_59 
+ bl[57] br[57] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_60 
+ bl[58] br[58] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_61 
+ bl[59] br[59] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_62 
+ bl[60] br[60] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_63 
+ bl[61] br[61] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_64 
+ bl[62] br[62] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_65 
+ bl[63] br[63] vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_66 
+ vdd vdd vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_174_67 
+ vdd vdd vdd vss wl[172] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_0 
+ vdd vdd vss vdd vpb vnb wl[173] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_175_1 
+ rbl rbr vss vdd vpb vnb wl[173] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_175_2 
+ bl[0] br[0] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_3 
+ bl[1] br[1] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_4 
+ bl[2] br[2] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_5 
+ bl[3] br[3] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_6 
+ bl[4] br[4] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_7 
+ bl[5] br[5] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_8 
+ bl[6] br[6] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_9 
+ bl[7] br[7] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_10 
+ bl[8] br[8] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_11 
+ bl[9] br[9] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_12 
+ bl[10] br[10] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_13 
+ bl[11] br[11] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_14 
+ bl[12] br[12] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_15 
+ bl[13] br[13] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_16 
+ bl[14] br[14] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_17 
+ bl[15] br[15] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_18 
+ bl[16] br[16] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_19 
+ bl[17] br[17] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_20 
+ bl[18] br[18] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_21 
+ bl[19] br[19] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_22 
+ bl[20] br[20] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_23 
+ bl[21] br[21] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_24 
+ bl[22] br[22] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_25 
+ bl[23] br[23] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_26 
+ bl[24] br[24] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_27 
+ bl[25] br[25] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_28 
+ bl[26] br[26] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_29 
+ bl[27] br[27] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_30 
+ bl[28] br[28] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_31 
+ bl[29] br[29] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_32 
+ bl[30] br[30] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_33 
+ bl[31] br[31] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_34 
+ bl[32] br[32] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_35 
+ bl[33] br[33] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_36 
+ bl[34] br[34] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_37 
+ bl[35] br[35] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_38 
+ bl[36] br[36] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_39 
+ bl[37] br[37] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_40 
+ bl[38] br[38] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_41 
+ bl[39] br[39] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_42 
+ bl[40] br[40] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_43 
+ bl[41] br[41] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_44 
+ bl[42] br[42] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_45 
+ bl[43] br[43] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_46 
+ bl[44] br[44] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_47 
+ bl[45] br[45] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_48 
+ bl[46] br[46] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_49 
+ bl[47] br[47] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_50 
+ bl[48] br[48] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_51 
+ bl[49] br[49] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_52 
+ bl[50] br[50] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_53 
+ bl[51] br[51] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_54 
+ bl[52] br[52] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_55 
+ bl[53] br[53] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_56 
+ bl[54] br[54] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_57 
+ bl[55] br[55] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_58 
+ bl[56] br[56] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_59 
+ bl[57] br[57] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_60 
+ bl[58] br[58] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_61 
+ bl[59] br[59] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_62 
+ bl[60] br[60] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_63 
+ bl[61] br[61] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_64 
+ bl[62] br[62] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_65 
+ bl[63] br[63] vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_66 
+ vdd vdd vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_175_67 
+ vdd vdd vdd vss wl[173] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_0 
+ vdd vdd vss vdd vpb vnb wl[174] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_176_1 
+ rbl rbr vss vdd vpb vnb wl[174] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_176_2 
+ bl[0] br[0] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_3 
+ bl[1] br[1] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_4 
+ bl[2] br[2] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_5 
+ bl[3] br[3] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_6 
+ bl[4] br[4] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_7 
+ bl[5] br[5] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_8 
+ bl[6] br[6] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_9 
+ bl[7] br[7] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_10 
+ bl[8] br[8] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_11 
+ bl[9] br[9] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_12 
+ bl[10] br[10] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_13 
+ bl[11] br[11] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_14 
+ bl[12] br[12] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_15 
+ bl[13] br[13] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_16 
+ bl[14] br[14] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_17 
+ bl[15] br[15] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_18 
+ bl[16] br[16] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_19 
+ bl[17] br[17] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_20 
+ bl[18] br[18] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_21 
+ bl[19] br[19] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_22 
+ bl[20] br[20] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_23 
+ bl[21] br[21] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_24 
+ bl[22] br[22] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_25 
+ bl[23] br[23] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_26 
+ bl[24] br[24] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_27 
+ bl[25] br[25] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_28 
+ bl[26] br[26] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_29 
+ bl[27] br[27] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_30 
+ bl[28] br[28] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_31 
+ bl[29] br[29] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_32 
+ bl[30] br[30] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_33 
+ bl[31] br[31] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_34 
+ bl[32] br[32] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_35 
+ bl[33] br[33] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_36 
+ bl[34] br[34] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_37 
+ bl[35] br[35] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_38 
+ bl[36] br[36] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_39 
+ bl[37] br[37] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_40 
+ bl[38] br[38] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_41 
+ bl[39] br[39] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_42 
+ bl[40] br[40] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_43 
+ bl[41] br[41] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_44 
+ bl[42] br[42] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_45 
+ bl[43] br[43] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_46 
+ bl[44] br[44] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_47 
+ bl[45] br[45] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_48 
+ bl[46] br[46] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_49 
+ bl[47] br[47] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_50 
+ bl[48] br[48] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_51 
+ bl[49] br[49] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_52 
+ bl[50] br[50] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_53 
+ bl[51] br[51] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_54 
+ bl[52] br[52] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_55 
+ bl[53] br[53] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_56 
+ bl[54] br[54] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_57 
+ bl[55] br[55] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_58 
+ bl[56] br[56] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_59 
+ bl[57] br[57] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_60 
+ bl[58] br[58] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_61 
+ bl[59] br[59] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_62 
+ bl[60] br[60] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_63 
+ bl[61] br[61] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_64 
+ bl[62] br[62] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_65 
+ bl[63] br[63] vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_66 
+ vdd vdd vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_176_67 
+ vdd vdd vdd vss wl[174] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_0 
+ vdd vdd vss vdd vpb vnb wl[175] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_177_1 
+ rbl rbr vss vdd vpb vnb wl[175] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_177_2 
+ bl[0] br[0] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_3 
+ bl[1] br[1] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_4 
+ bl[2] br[2] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_5 
+ bl[3] br[3] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_6 
+ bl[4] br[4] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_7 
+ bl[5] br[5] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_8 
+ bl[6] br[6] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_9 
+ bl[7] br[7] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_10 
+ bl[8] br[8] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_11 
+ bl[9] br[9] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_12 
+ bl[10] br[10] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_13 
+ bl[11] br[11] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_14 
+ bl[12] br[12] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_15 
+ bl[13] br[13] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_16 
+ bl[14] br[14] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_17 
+ bl[15] br[15] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_18 
+ bl[16] br[16] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_19 
+ bl[17] br[17] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_20 
+ bl[18] br[18] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_21 
+ bl[19] br[19] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_22 
+ bl[20] br[20] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_23 
+ bl[21] br[21] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_24 
+ bl[22] br[22] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_25 
+ bl[23] br[23] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_26 
+ bl[24] br[24] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_27 
+ bl[25] br[25] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_28 
+ bl[26] br[26] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_29 
+ bl[27] br[27] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_30 
+ bl[28] br[28] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_31 
+ bl[29] br[29] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_32 
+ bl[30] br[30] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_33 
+ bl[31] br[31] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_34 
+ bl[32] br[32] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_35 
+ bl[33] br[33] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_36 
+ bl[34] br[34] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_37 
+ bl[35] br[35] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_38 
+ bl[36] br[36] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_39 
+ bl[37] br[37] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_40 
+ bl[38] br[38] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_41 
+ bl[39] br[39] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_42 
+ bl[40] br[40] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_43 
+ bl[41] br[41] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_44 
+ bl[42] br[42] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_45 
+ bl[43] br[43] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_46 
+ bl[44] br[44] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_47 
+ bl[45] br[45] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_48 
+ bl[46] br[46] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_49 
+ bl[47] br[47] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_50 
+ bl[48] br[48] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_51 
+ bl[49] br[49] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_52 
+ bl[50] br[50] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_53 
+ bl[51] br[51] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_54 
+ bl[52] br[52] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_55 
+ bl[53] br[53] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_56 
+ bl[54] br[54] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_57 
+ bl[55] br[55] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_58 
+ bl[56] br[56] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_59 
+ bl[57] br[57] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_60 
+ bl[58] br[58] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_61 
+ bl[59] br[59] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_62 
+ bl[60] br[60] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_63 
+ bl[61] br[61] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_64 
+ bl[62] br[62] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_65 
+ bl[63] br[63] vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_66 
+ vdd vdd vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_177_67 
+ vdd vdd vdd vss wl[175] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_0 
+ vdd vdd vss vdd vpb vnb wl[176] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_178_1 
+ rbl rbr vss vdd vpb vnb wl[176] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_178_2 
+ bl[0] br[0] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_3 
+ bl[1] br[1] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_4 
+ bl[2] br[2] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_5 
+ bl[3] br[3] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_6 
+ bl[4] br[4] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_7 
+ bl[5] br[5] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_8 
+ bl[6] br[6] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_9 
+ bl[7] br[7] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_10 
+ bl[8] br[8] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_11 
+ bl[9] br[9] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_12 
+ bl[10] br[10] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_13 
+ bl[11] br[11] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_14 
+ bl[12] br[12] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_15 
+ bl[13] br[13] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_16 
+ bl[14] br[14] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_17 
+ bl[15] br[15] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_18 
+ bl[16] br[16] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_19 
+ bl[17] br[17] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_20 
+ bl[18] br[18] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_21 
+ bl[19] br[19] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_22 
+ bl[20] br[20] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_23 
+ bl[21] br[21] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_24 
+ bl[22] br[22] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_25 
+ bl[23] br[23] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_26 
+ bl[24] br[24] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_27 
+ bl[25] br[25] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_28 
+ bl[26] br[26] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_29 
+ bl[27] br[27] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_30 
+ bl[28] br[28] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_31 
+ bl[29] br[29] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_32 
+ bl[30] br[30] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_33 
+ bl[31] br[31] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_34 
+ bl[32] br[32] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_35 
+ bl[33] br[33] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_36 
+ bl[34] br[34] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_37 
+ bl[35] br[35] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_38 
+ bl[36] br[36] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_39 
+ bl[37] br[37] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_40 
+ bl[38] br[38] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_41 
+ bl[39] br[39] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_42 
+ bl[40] br[40] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_43 
+ bl[41] br[41] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_44 
+ bl[42] br[42] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_45 
+ bl[43] br[43] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_46 
+ bl[44] br[44] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_47 
+ bl[45] br[45] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_48 
+ bl[46] br[46] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_49 
+ bl[47] br[47] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_50 
+ bl[48] br[48] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_51 
+ bl[49] br[49] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_52 
+ bl[50] br[50] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_53 
+ bl[51] br[51] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_54 
+ bl[52] br[52] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_55 
+ bl[53] br[53] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_56 
+ bl[54] br[54] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_57 
+ bl[55] br[55] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_58 
+ bl[56] br[56] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_59 
+ bl[57] br[57] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_60 
+ bl[58] br[58] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_61 
+ bl[59] br[59] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_62 
+ bl[60] br[60] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_63 
+ bl[61] br[61] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_64 
+ bl[62] br[62] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_65 
+ bl[63] br[63] vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_66 
+ vdd vdd vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_178_67 
+ vdd vdd vdd vss wl[176] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_0 
+ vdd vdd vss vdd vpb vnb wl[177] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_179_1 
+ rbl rbr vss vdd vpb vnb wl[177] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_179_2 
+ bl[0] br[0] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_3 
+ bl[1] br[1] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_4 
+ bl[2] br[2] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_5 
+ bl[3] br[3] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_6 
+ bl[4] br[4] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_7 
+ bl[5] br[5] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_8 
+ bl[6] br[6] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_9 
+ bl[7] br[7] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_10 
+ bl[8] br[8] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_11 
+ bl[9] br[9] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_12 
+ bl[10] br[10] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_13 
+ bl[11] br[11] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_14 
+ bl[12] br[12] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_15 
+ bl[13] br[13] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_16 
+ bl[14] br[14] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_17 
+ bl[15] br[15] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_18 
+ bl[16] br[16] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_19 
+ bl[17] br[17] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_20 
+ bl[18] br[18] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_21 
+ bl[19] br[19] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_22 
+ bl[20] br[20] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_23 
+ bl[21] br[21] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_24 
+ bl[22] br[22] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_25 
+ bl[23] br[23] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_26 
+ bl[24] br[24] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_27 
+ bl[25] br[25] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_28 
+ bl[26] br[26] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_29 
+ bl[27] br[27] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_30 
+ bl[28] br[28] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_31 
+ bl[29] br[29] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_32 
+ bl[30] br[30] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_33 
+ bl[31] br[31] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_34 
+ bl[32] br[32] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_35 
+ bl[33] br[33] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_36 
+ bl[34] br[34] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_37 
+ bl[35] br[35] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_38 
+ bl[36] br[36] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_39 
+ bl[37] br[37] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_40 
+ bl[38] br[38] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_41 
+ bl[39] br[39] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_42 
+ bl[40] br[40] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_43 
+ bl[41] br[41] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_44 
+ bl[42] br[42] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_45 
+ bl[43] br[43] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_46 
+ bl[44] br[44] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_47 
+ bl[45] br[45] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_48 
+ bl[46] br[46] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_49 
+ bl[47] br[47] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_50 
+ bl[48] br[48] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_51 
+ bl[49] br[49] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_52 
+ bl[50] br[50] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_53 
+ bl[51] br[51] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_54 
+ bl[52] br[52] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_55 
+ bl[53] br[53] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_56 
+ bl[54] br[54] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_57 
+ bl[55] br[55] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_58 
+ bl[56] br[56] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_59 
+ bl[57] br[57] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_60 
+ bl[58] br[58] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_61 
+ bl[59] br[59] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_62 
+ bl[60] br[60] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_63 
+ bl[61] br[61] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_64 
+ bl[62] br[62] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_65 
+ bl[63] br[63] vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_66 
+ vdd vdd vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_179_67 
+ vdd vdd vdd vss wl[177] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_0 
+ vdd vdd vss vdd vpb vnb wl[178] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_180_1 
+ rbl rbr vss vdd vpb vnb wl[178] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_180_2 
+ bl[0] br[0] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_3 
+ bl[1] br[1] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_4 
+ bl[2] br[2] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_5 
+ bl[3] br[3] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_6 
+ bl[4] br[4] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_7 
+ bl[5] br[5] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_8 
+ bl[6] br[6] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_9 
+ bl[7] br[7] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_10 
+ bl[8] br[8] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_11 
+ bl[9] br[9] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_12 
+ bl[10] br[10] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_13 
+ bl[11] br[11] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_14 
+ bl[12] br[12] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_15 
+ bl[13] br[13] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_16 
+ bl[14] br[14] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_17 
+ bl[15] br[15] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_18 
+ bl[16] br[16] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_19 
+ bl[17] br[17] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_20 
+ bl[18] br[18] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_21 
+ bl[19] br[19] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_22 
+ bl[20] br[20] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_23 
+ bl[21] br[21] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_24 
+ bl[22] br[22] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_25 
+ bl[23] br[23] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_26 
+ bl[24] br[24] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_27 
+ bl[25] br[25] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_28 
+ bl[26] br[26] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_29 
+ bl[27] br[27] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_30 
+ bl[28] br[28] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_31 
+ bl[29] br[29] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_32 
+ bl[30] br[30] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_33 
+ bl[31] br[31] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_34 
+ bl[32] br[32] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_35 
+ bl[33] br[33] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_36 
+ bl[34] br[34] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_37 
+ bl[35] br[35] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_38 
+ bl[36] br[36] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_39 
+ bl[37] br[37] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_40 
+ bl[38] br[38] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_41 
+ bl[39] br[39] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_42 
+ bl[40] br[40] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_43 
+ bl[41] br[41] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_44 
+ bl[42] br[42] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_45 
+ bl[43] br[43] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_46 
+ bl[44] br[44] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_47 
+ bl[45] br[45] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_48 
+ bl[46] br[46] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_49 
+ bl[47] br[47] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_50 
+ bl[48] br[48] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_51 
+ bl[49] br[49] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_52 
+ bl[50] br[50] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_53 
+ bl[51] br[51] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_54 
+ bl[52] br[52] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_55 
+ bl[53] br[53] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_56 
+ bl[54] br[54] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_57 
+ bl[55] br[55] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_58 
+ bl[56] br[56] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_59 
+ bl[57] br[57] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_60 
+ bl[58] br[58] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_61 
+ bl[59] br[59] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_62 
+ bl[60] br[60] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_63 
+ bl[61] br[61] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_64 
+ bl[62] br[62] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_65 
+ bl[63] br[63] vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_66 
+ vdd vdd vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_180_67 
+ vdd vdd vdd vss wl[178] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_0 
+ vdd vdd vss vdd vpb vnb wl[179] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_181_1 
+ rbl rbr vss vdd vpb vnb wl[179] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_181_2 
+ bl[0] br[0] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_3 
+ bl[1] br[1] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_4 
+ bl[2] br[2] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_5 
+ bl[3] br[3] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_6 
+ bl[4] br[4] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_7 
+ bl[5] br[5] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_8 
+ bl[6] br[6] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_9 
+ bl[7] br[7] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_10 
+ bl[8] br[8] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_11 
+ bl[9] br[9] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_12 
+ bl[10] br[10] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_13 
+ bl[11] br[11] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_14 
+ bl[12] br[12] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_15 
+ bl[13] br[13] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_16 
+ bl[14] br[14] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_17 
+ bl[15] br[15] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_18 
+ bl[16] br[16] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_19 
+ bl[17] br[17] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_20 
+ bl[18] br[18] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_21 
+ bl[19] br[19] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_22 
+ bl[20] br[20] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_23 
+ bl[21] br[21] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_24 
+ bl[22] br[22] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_25 
+ bl[23] br[23] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_26 
+ bl[24] br[24] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_27 
+ bl[25] br[25] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_28 
+ bl[26] br[26] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_29 
+ bl[27] br[27] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_30 
+ bl[28] br[28] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_31 
+ bl[29] br[29] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_32 
+ bl[30] br[30] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_33 
+ bl[31] br[31] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_34 
+ bl[32] br[32] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_35 
+ bl[33] br[33] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_36 
+ bl[34] br[34] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_37 
+ bl[35] br[35] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_38 
+ bl[36] br[36] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_39 
+ bl[37] br[37] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_40 
+ bl[38] br[38] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_41 
+ bl[39] br[39] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_42 
+ bl[40] br[40] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_43 
+ bl[41] br[41] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_44 
+ bl[42] br[42] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_45 
+ bl[43] br[43] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_46 
+ bl[44] br[44] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_47 
+ bl[45] br[45] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_48 
+ bl[46] br[46] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_49 
+ bl[47] br[47] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_50 
+ bl[48] br[48] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_51 
+ bl[49] br[49] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_52 
+ bl[50] br[50] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_53 
+ bl[51] br[51] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_54 
+ bl[52] br[52] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_55 
+ bl[53] br[53] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_56 
+ bl[54] br[54] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_57 
+ bl[55] br[55] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_58 
+ bl[56] br[56] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_59 
+ bl[57] br[57] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_60 
+ bl[58] br[58] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_61 
+ bl[59] br[59] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_62 
+ bl[60] br[60] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_63 
+ bl[61] br[61] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_64 
+ bl[62] br[62] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_65 
+ bl[63] br[63] vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_66 
+ vdd vdd vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_181_67 
+ vdd vdd vdd vss wl[179] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_0 
+ vdd vdd vss vdd vpb vnb wl[180] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_182_1 
+ rbl rbr vss vdd vpb vnb wl[180] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_182_2 
+ bl[0] br[0] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_3 
+ bl[1] br[1] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_4 
+ bl[2] br[2] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_5 
+ bl[3] br[3] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_6 
+ bl[4] br[4] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_7 
+ bl[5] br[5] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_8 
+ bl[6] br[6] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_9 
+ bl[7] br[7] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_10 
+ bl[8] br[8] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_11 
+ bl[9] br[9] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_12 
+ bl[10] br[10] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_13 
+ bl[11] br[11] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_14 
+ bl[12] br[12] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_15 
+ bl[13] br[13] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_16 
+ bl[14] br[14] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_17 
+ bl[15] br[15] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_18 
+ bl[16] br[16] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_19 
+ bl[17] br[17] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_20 
+ bl[18] br[18] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_21 
+ bl[19] br[19] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_22 
+ bl[20] br[20] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_23 
+ bl[21] br[21] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_24 
+ bl[22] br[22] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_25 
+ bl[23] br[23] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_26 
+ bl[24] br[24] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_27 
+ bl[25] br[25] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_28 
+ bl[26] br[26] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_29 
+ bl[27] br[27] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_30 
+ bl[28] br[28] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_31 
+ bl[29] br[29] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_32 
+ bl[30] br[30] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_33 
+ bl[31] br[31] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_34 
+ bl[32] br[32] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_35 
+ bl[33] br[33] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_36 
+ bl[34] br[34] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_37 
+ bl[35] br[35] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_38 
+ bl[36] br[36] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_39 
+ bl[37] br[37] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_40 
+ bl[38] br[38] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_41 
+ bl[39] br[39] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_42 
+ bl[40] br[40] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_43 
+ bl[41] br[41] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_44 
+ bl[42] br[42] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_45 
+ bl[43] br[43] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_46 
+ bl[44] br[44] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_47 
+ bl[45] br[45] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_48 
+ bl[46] br[46] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_49 
+ bl[47] br[47] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_50 
+ bl[48] br[48] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_51 
+ bl[49] br[49] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_52 
+ bl[50] br[50] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_53 
+ bl[51] br[51] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_54 
+ bl[52] br[52] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_55 
+ bl[53] br[53] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_56 
+ bl[54] br[54] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_57 
+ bl[55] br[55] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_58 
+ bl[56] br[56] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_59 
+ bl[57] br[57] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_60 
+ bl[58] br[58] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_61 
+ bl[59] br[59] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_62 
+ bl[60] br[60] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_63 
+ bl[61] br[61] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_64 
+ bl[62] br[62] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_65 
+ bl[63] br[63] vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_66 
+ vdd vdd vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_182_67 
+ vdd vdd vdd vss wl[180] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_0 
+ vdd vdd vss vdd vpb vnb wl[181] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_183_1 
+ rbl rbr vss vdd vpb vnb wl[181] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_183_2 
+ bl[0] br[0] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_3 
+ bl[1] br[1] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_4 
+ bl[2] br[2] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_5 
+ bl[3] br[3] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_6 
+ bl[4] br[4] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_7 
+ bl[5] br[5] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_8 
+ bl[6] br[6] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_9 
+ bl[7] br[7] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_10 
+ bl[8] br[8] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_11 
+ bl[9] br[9] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_12 
+ bl[10] br[10] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_13 
+ bl[11] br[11] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_14 
+ bl[12] br[12] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_15 
+ bl[13] br[13] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_16 
+ bl[14] br[14] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_17 
+ bl[15] br[15] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_18 
+ bl[16] br[16] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_19 
+ bl[17] br[17] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_20 
+ bl[18] br[18] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_21 
+ bl[19] br[19] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_22 
+ bl[20] br[20] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_23 
+ bl[21] br[21] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_24 
+ bl[22] br[22] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_25 
+ bl[23] br[23] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_26 
+ bl[24] br[24] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_27 
+ bl[25] br[25] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_28 
+ bl[26] br[26] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_29 
+ bl[27] br[27] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_30 
+ bl[28] br[28] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_31 
+ bl[29] br[29] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_32 
+ bl[30] br[30] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_33 
+ bl[31] br[31] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_34 
+ bl[32] br[32] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_35 
+ bl[33] br[33] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_36 
+ bl[34] br[34] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_37 
+ bl[35] br[35] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_38 
+ bl[36] br[36] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_39 
+ bl[37] br[37] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_40 
+ bl[38] br[38] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_41 
+ bl[39] br[39] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_42 
+ bl[40] br[40] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_43 
+ bl[41] br[41] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_44 
+ bl[42] br[42] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_45 
+ bl[43] br[43] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_46 
+ bl[44] br[44] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_47 
+ bl[45] br[45] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_48 
+ bl[46] br[46] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_49 
+ bl[47] br[47] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_50 
+ bl[48] br[48] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_51 
+ bl[49] br[49] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_52 
+ bl[50] br[50] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_53 
+ bl[51] br[51] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_54 
+ bl[52] br[52] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_55 
+ bl[53] br[53] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_56 
+ bl[54] br[54] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_57 
+ bl[55] br[55] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_58 
+ bl[56] br[56] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_59 
+ bl[57] br[57] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_60 
+ bl[58] br[58] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_61 
+ bl[59] br[59] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_62 
+ bl[60] br[60] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_63 
+ bl[61] br[61] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_64 
+ bl[62] br[62] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_65 
+ bl[63] br[63] vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_66 
+ vdd vdd vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_183_67 
+ vdd vdd vdd vss wl[181] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_0 
+ vdd vdd vss vdd vpb vnb wl[182] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_184_1 
+ rbl rbr vss vdd vpb vnb wl[182] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_184_2 
+ bl[0] br[0] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_3 
+ bl[1] br[1] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_4 
+ bl[2] br[2] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_5 
+ bl[3] br[3] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_6 
+ bl[4] br[4] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_7 
+ bl[5] br[5] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_8 
+ bl[6] br[6] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_9 
+ bl[7] br[7] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_10 
+ bl[8] br[8] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_11 
+ bl[9] br[9] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_12 
+ bl[10] br[10] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_13 
+ bl[11] br[11] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_14 
+ bl[12] br[12] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_15 
+ bl[13] br[13] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_16 
+ bl[14] br[14] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_17 
+ bl[15] br[15] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_18 
+ bl[16] br[16] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_19 
+ bl[17] br[17] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_20 
+ bl[18] br[18] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_21 
+ bl[19] br[19] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_22 
+ bl[20] br[20] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_23 
+ bl[21] br[21] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_24 
+ bl[22] br[22] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_25 
+ bl[23] br[23] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_26 
+ bl[24] br[24] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_27 
+ bl[25] br[25] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_28 
+ bl[26] br[26] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_29 
+ bl[27] br[27] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_30 
+ bl[28] br[28] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_31 
+ bl[29] br[29] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_32 
+ bl[30] br[30] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_33 
+ bl[31] br[31] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_34 
+ bl[32] br[32] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_35 
+ bl[33] br[33] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_36 
+ bl[34] br[34] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_37 
+ bl[35] br[35] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_38 
+ bl[36] br[36] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_39 
+ bl[37] br[37] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_40 
+ bl[38] br[38] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_41 
+ bl[39] br[39] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_42 
+ bl[40] br[40] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_43 
+ bl[41] br[41] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_44 
+ bl[42] br[42] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_45 
+ bl[43] br[43] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_46 
+ bl[44] br[44] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_47 
+ bl[45] br[45] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_48 
+ bl[46] br[46] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_49 
+ bl[47] br[47] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_50 
+ bl[48] br[48] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_51 
+ bl[49] br[49] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_52 
+ bl[50] br[50] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_53 
+ bl[51] br[51] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_54 
+ bl[52] br[52] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_55 
+ bl[53] br[53] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_56 
+ bl[54] br[54] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_57 
+ bl[55] br[55] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_58 
+ bl[56] br[56] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_59 
+ bl[57] br[57] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_60 
+ bl[58] br[58] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_61 
+ bl[59] br[59] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_62 
+ bl[60] br[60] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_63 
+ bl[61] br[61] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_64 
+ bl[62] br[62] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_65 
+ bl[63] br[63] vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_66 
+ vdd vdd vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_184_67 
+ vdd vdd vdd vss wl[182] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_0 
+ vdd vdd vss vdd vpb vnb wl[183] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_185_1 
+ rbl rbr vss vdd vpb vnb wl[183] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_185_2 
+ bl[0] br[0] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_3 
+ bl[1] br[1] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_4 
+ bl[2] br[2] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_5 
+ bl[3] br[3] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_6 
+ bl[4] br[4] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_7 
+ bl[5] br[5] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_8 
+ bl[6] br[6] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_9 
+ bl[7] br[7] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_10 
+ bl[8] br[8] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_11 
+ bl[9] br[9] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_12 
+ bl[10] br[10] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_13 
+ bl[11] br[11] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_14 
+ bl[12] br[12] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_15 
+ bl[13] br[13] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_16 
+ bl[14] br[14] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_17 
+ bl[15] br[15] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_18 
+ bl[16] br[16] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_19 
+ bl[17] br[17] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_20 
+ bl[18] br[18] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_21 
+ bl[19] br[19] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_22 
+ bl[20] br[20] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_23 
+ bl[21] br[21] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_24 
+ bl[22] br[22] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_25 
+ bl[23] br[23] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_26 
+ bl[24] br[24] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_27 
+ bl[25] br[25] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_28 
+ bl[26] br[26] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_29 
+ bl[27] br[27] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_30 
+ bl[28] br[28] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_31 
+ bl[29] br[29] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_32 
+ bl[30] br[30] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_33 
+ bl[31] br[31] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_34 
+ bl[32] br[32] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_35 
+ bl[33] br[33] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_36 
+ bl[34] br[34] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_37 
+ bl[35] br[35] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_38 
+ bl[36] br[36] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_39 
+ bl[37] br[37] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_40 
+ bl[38] br[38] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_41 
+ bl[39] br[39] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_42 
+ bl[40] br[40] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_43 
+ bl[41] br[41] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_44 
+ bl[42] br[42] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_45 
+ bl[43] br[43] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_46 
+ bl[44] br[44] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_47 
+ bl[45] br[45] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_48 
+ bl[46] br[46] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_49 
+ bl[47] br[47] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_50 
+ bl[48] br[48] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_51 
+ bl[49] br[49] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_52 
+ bl[50] br[50] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_53 
+ bl[51] br[51] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_54 
+ bl[52] br[52] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_55 
+ bl[53] br[53] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_56 
+ bl[54] br[54] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_57 
+ bl[55] br[55] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_58 
+ bl[56] br[56] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_59 
+ bl[57] br[57] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_60 
+ bl[58] br[58] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_61 
+ bl[59] br[59] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_62 
+ bl[60] br[60] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_63 
+ bl[61] br[61] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_64 
+ bl[62] br[62] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_65 
+ bl[63] br[63] vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_66 
+ vdd vdd vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_185_67 
+ vdd vdd vdd vss wl[183] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_0 
+ vdd vdd vss vdd vpb vnb wl[184] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_186_1 
+ rbl rbr vss vdd vpb vnb wl[184] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_186_2 
+ bl[0] br[0] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_3 
+ bl[1] br[1] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_4 
+ bl[2] br[2] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_5 
+ bl[3] br[3] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_6 
+ bl[4] br[4] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_7 
+ bl[5] br[5] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_8 
+ bl[6] br[6] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_9 
+ bl[7] br[7] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_10 
+ bl[8] br[8] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_11 
+ bl[9] br[9] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_12 
+ bl[10] br[10] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_13 
+ bl[11] br[11] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_14 
+ bl[12] br[12] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_15 
+ bl[13] br[13] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_16 
+ bl[14] br[14] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_17 
+ bl[15] br[15] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_18 
+ bl[16] br[16] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_19 
+ bl[17] br[17] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_20 
+ bl[18] br[18] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_21 
+ bl[19] br[19] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_22 
+ bl[20] br[20] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_23 
+ bl[21] br[21] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_24 
+ bl[22] br[22] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_25 
+ bl[23] br[23] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_26 
+ bl[24] br[24] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_27 
+ bl[25] br[25] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_28 
+ bl[26] br[26] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_29 
+ bl[27] br[27] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_30 
+ bl[28] br[28] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_31 
+ bl[29] br[29] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_32 
+ bl[30] br[30] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_33 
+ bl[31] br[31] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_34 
+ bl[32] br[32] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_35 
+ bl[33] br[33] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_36 
+ bl[34] br[34] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_37 
+ bl[35] br[35] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_38 
+ bl[36] br[36] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_39 
+ bl[37] br[37] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_40 
+ bl[38] br[38] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_41 
+ bl[39] br[39] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_42 
+ bl[40] br[40] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_43 
+ bl[41] br[41] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_44 
+ bl[42] br[42] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_45 
+ bl[43] br[43] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_46 
+ bl[44] br[44] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_47 
+ bl[45] br[45] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_48 
+ bl[46] br[46] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_49 
+ bl[47] br[47] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_50 
+ bl[48] br[48] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_51 
+ bl[49] br[49] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_52 
+ bl[50] br[50] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_53 
+ bl[51] br[51] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_54 
+ bl[52] br[52] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_55 
+ bl[53] br[53] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_56 
+ bl[54] br[54] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_57 
+ bl[55] br[55] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_58 
+ bl[56] br[56] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_59 
+ bl[57] br[57] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_60 
+ bl[58] br[58] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_61 
+ bl[59] br[59] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_62 
+ bl[60] br[60] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_63 
+ bl[61] br[61] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_64 
+ bl[62] br[62] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_65 
+ bl[63] br[63] vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_66 
+ vdd vdd vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_186_67 
+ vdd vdd vdd vss wl[184] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_0 
+ vdd vdd vss vdd vpb vnb wl[185] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_187_1 
+ rbl rbr vss vdd vpb vnb wl[185] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_187_2 
+ bl[0] br[0] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_3 
+ bl[1] br[1] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_4 
+ bl[2] br[2] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_5 
+ bl[3] br[3] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_6 
+ bl[4] br[4] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_7 
+ bl[5] br[5] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_8 
+ bl[6] br[6] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_9 
+ bl[7] br[7] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_10 
+ bl[8] br[8] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_11 
+ bl[9] br[9] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_12 
+ bl[10] br[10] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_13 
+ bl[11] br[11] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_14 
+ bl[12] br[12] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_15 
+ bl[13] br[13] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_16 
+ bl[14] br[14] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_17 
+ bl[15] br[15] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_18 
+ bl[16] br[16] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_19 
+ bl[17] br[17] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_20 
+ bl[18] br[18] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_21 
+ bl[19] br[19] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_22 
+ bl[20] br[20] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_23 
+ bl[21] br[21] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_24 
+ bl[22] br[22] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_25 
+ bl[23] br[23] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_26 
+ bl[24] br[24] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_27 
+ bl[25] br[25] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_28 
+ bl[26] br[26] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_29 
+ bl[27] br[27] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_30 
+ bl[28] br[28] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_31 
+ bl[29] br[29] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_32 
+ bl[30] br[30] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_33 
+ bl[31] br[31] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_34 
+ bl[32] br[32] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_35 
+ bl[33] br[33] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_36 
+ bl[34] br[34] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_37 
+ bl[35] br[35] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_38 
+ bl[36] br[36] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_39 
+ bl[37] br[37] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_40 
+ bl[38] br[38] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_41 
+ bl[39] br[39] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_42 
+ bl[40] br[40] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_43 
+ bl[41] br[41] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_44 
+ bl[42] br[42] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_45 
+ bl[43] br[43] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_46 
+ bl[44] br[44] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_47 
+ bl[45] br[45] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_48 
+ bl[46] br[46] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_49 
+ bl[47] br[47] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_50 
+ bl[48] br[48] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_51 
+ bl[49] br[49] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_52 
+ bl[50] br[50] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_53 
+ bl[51] br[51] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_54 
+ bl[52] br[52] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_55 
+ bl[53] br[53] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_56 
+ bl[54] br[54] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_57 
+ bl[55] br[55] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_58 
+ bl[56] br[56] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_59 
+ bl[57] br[57] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_60 
+ bl[58] br[58] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_61 
+ bl[59] br[59] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_62 
+ bl[60] br[60] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_63 
+ bl[61] br[61] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_64 
+ bl[62] br[62] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_65 
+ bl[63] br[63] vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_66 
+ vdd vdd vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_187_67 
+ vdd vdd vdd vss wl[185] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_0 
+ vdd vdd vss vdd vpb vnb wl[186] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_188_1 
+ rbl rbr vss vdd vpb vnb wl[186] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_188_2 
+ bl[0] br[0] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_3 
+ bl[1] br[1] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_4 
+ bl[2] br[2] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_5 
+ bl[3] br[3] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_6 
+ bl[4] br[4] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_7 
+ bl[5] br[5] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_8 
+ bl[6] br[6] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_9 
+ bl[7] br[7] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_10 
+ bl[8] br[8] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_11 
+ bl[9] br[9] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_12 
+ bl[10] br[10] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_13 
+ bl[11] br[11] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_14 
+ bl[12] br[12] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_15 
+ bl[13] br[13] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_16 
+ bl[14] br[14] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_17 
+ bl[15] br[15] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_18 
+ bl[16] br[16] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_19 
+ bl[17] br[17] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_20 
+ bl[18] br[18] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_21 
+ bl[19] br[19] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_22 
+ bl[20] br[20] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_23 
+ bl[21] br[21] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_24 
+ bl[22] br[22] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_25 
+ bl[23] br[23] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_26 
+ bl[24] br[24] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_27 
+ bl[25] br[25] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_28 
+ bl[26] br[26] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_29 
+ bl[27] br[27] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_30 
+ bl[28] br[28] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_31 
+ bl[29] br[29] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_32 
+ bl[30] br[30] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_33 
+ bl[31] br[31] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_34 
+ bl[32] br[32] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_35 
+ bl[33] br[33] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_36 
+ bl[34] br[34] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_37 
+ bl[35] br[35] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_38 
+ bl[36] br[36] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_39 
+ bl[37] br[37] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_40 
+ bl[38] br[38] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_41 
+ bl[39] br[39] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_42 
+ bl[40] br[40] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_43 
+ bl[41] br[41] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_44 
+ bl[42] br[42] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_45 
+ bl[43] br[43] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_46 
+ bl[44] br[44] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_47 
+ bl[45] br[45] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_48 
+ bl[46] br[46] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_49 
+ bl[47] br[47] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_50 
+ bl[48] br[48] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_51 
+ bl[49] br[49] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_52 
+ bl[50] br[50] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_53 
+ bl[51] br[51] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_54 
+ bl[52] br[52] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_55 
+ bl[53] br[53] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_56 
+ bl[54] br[54] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_57 
+ bl[55] br[55] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_58 
+ bl[56] br[56] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_59 
+ bl[57] br[57] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_60 
+ bl[58] br[58] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_61 
+ bl[59] br[59] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_62 
+ bl[60] br[60] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_63 
+ bl[61] br[61] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_64 
+ bl[62] br[62] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_65 
+ bl[63] br[63] vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_66 
+ vdd vdd vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_188_67 
+ vdd vdd vdd vss wl[186] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_0 
+ vdd vdd vss vdd vpb vnb wl[187] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_189_1 
+ rbl rbr vss vdd vpb vnb wl[187] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_189_2 
+ bl[0] br[0] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_3 
+ bl[1] br[1] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_4 
+ bl[2] br[2] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_5 
+ bl[3] br[3] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_6 
+ bl[4] br[4] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_7 
+ bl[5] br[5] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_8 
+ bl[6] br[6] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_9 
+ bl[7] br[7] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_10 
+ bl[8] br[8] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_11 
+ bl[9] br[9] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_12 
+ bl[10] br[10] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_13 
+ bl[11] br[11] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_14 
+ bl[12] br[12] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_15 
+ bl[13] br[13] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_16 
+ bl[14] br[14] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_17 
+ bl[15] br[15] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_18 
+ bl[16] br[16] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_19 
+ bl[17] br[17] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_20 
+ bl[18] br[18] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_21 
+ bl[19] br[19] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_22 
+ bl[20] br[20] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_23 
+ bl[21] br[21] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_24 
+ bl[22] br[22] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_25 
+ bl[23] br[23] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_26 
+ bl[24] br[24] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_27 
+ bl[25] br[25] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_28 
+ bl[26] br[26] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_29 
+ bl[27] br[27] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_30 
+ bl[28] br[28] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_31 
+ bl[29] br[29] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_32 
+ bl[30] br[30] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_33 
+ bl[31] br[31] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_34 
+ bl[32] br[32] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_35 
+ bl[33] br[33] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_36 
+ bl[34] br[34] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_37 
+ bl[35] br[35] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_38 
+ bl[36] br[36] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_39 
+ bl[37] br[37] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_40 
+ bl[38] br[38] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_41 
+ bl[39] br[39] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_42 
+ bl[40] br[40] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_43 
+ bl[41] br[41] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_44 
+ bl[42] br[42] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_45 
+ bl[43] br[43] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_46 
+ bl[44] br[44] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_47 
+ bl[45] br[45] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_48 
+ bl[46] br[46] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_49 
+ bl[47] br[47] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_50 
+ bl[48] br[48] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_51 
+ bl[49] br[49] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_52 
+ bl[50] br[50] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_53 
+ bl[51] br[51] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_54 
+ bl[52] br[52] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_55 
+ bl[53] br[53] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_56 
+ bl[54] br[54] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_57 
+ bl[55] br[55] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_58 
+ bl[56] br[56] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_59 
+ bl[57] br[57] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_60 
+ bl[58] br[58] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_61 
+ bl[59] br[59] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_62 
+ bl[60] br[60] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_63 
+ bl[61] br[61] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_64 
+ bl[62] br[62] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_65 
+ bl[63] br[63] vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_66 
+ vdd vdd vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_189_67 
+ vdd vdd vdd vss wl[187] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_0 
+ vdd vdd vss vdd vpb vnb wl[188] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_190_1 
+ rbl rbr vss vdd vpb vnb wl[188] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_190_2 
+ bl[0] br[0] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_3 
+ bl[1] br[1] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_4 
+ bl[2] br[2] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_5 
+ bl[3] br[3] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_6 
+ bl[4] br[4] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_7 
+ bl[5] br[5] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_8 
+ bl[6] br[6] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_9 
+ bl[7] br[7] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_10 
+ bl[8] br[8] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_11 
+ bl[9] br[9] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_12 
+ bl[10] br[10] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_13 
+ bl[11] br[11] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_14 
+ bl[12] br[12] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_15 
+ bl[13] br[13] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_16 
+ bl[14] br[14] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_17 
+ bl[15] br[15] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_18 
+ bl[16] br[16] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_19 
+ bl[17] br[17] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_20 
+ bl[18] br[18] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_21 
+ bl[19] br[19] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_22 
+ bl[20] br[20] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_23 
+ bl[21] br[21] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_24 
+ bl[22] br[22] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_25 
+ bl[23] br[23] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_26 
+ bl[24] br[24] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_27 
+ bl[25] br[25] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_28 
+ bl[26] br[26] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_29 
+ bl[27] br[27] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_30 
+ bl[28] br[28] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_31 
+ bl[29] br[29] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_32 
+ bl[30] br[30] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_33 
+ bl[31] br[31] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_34 
+ bl[32] br[32] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_35 
+ bl[33] br[33] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_36 
+ bl[34] br[34] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_37 
+ bl[35] br[35] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_38 
+ bl[36] br[36] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_39 
+ bl[37] br[37] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_40 
+ bl[38] br[38] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_41 
+ bl[39] br[39] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_42 
+ bl[40] br[40] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_43 
+ bl[41] br[41] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_44 
+ bl[42] br[42] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_45 
+ bl[43] br[43] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_46 
+ bl[44] br[44] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_47 
+ bl[45] br[45] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_48 
+ bl[46] br[46] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_49 
+ bl[47] br[47] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_50 
+ bl[48] br[48] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_51 
+ bl[49] br[49] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_52 
+ bl[50] br[50] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_53 
+ bl[51] br[51] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_54 
+ bl[52] br[52] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_55 
+ bl[53] br[53] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_56 
+ bl[54] br[54] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_57 
+ bl[55] br[55] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_58 
+ bl[56] br[56] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_59 
+ bl[57] br[57] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_60 
+ bl[58] br[58] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_61 
+ bl[59] br[59] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_62 
+ bl[60] br[60] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_63 
+ bl[61] br[61] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_64 
+ bl[62] br[62] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_65 
+ bl[63] br[63] vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_66 
+ vdd vdd vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_190_67 
+ vdd vdd vdd vss wl[188] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_0 
+ vdd vdd vss vdd vpb vnb wl[189] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_191_1 
+ rbl rbr vss vdd vpb vnb wl[189] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_191_2 
+ bl[0] br[0] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_3 
+ bl[1] br[1] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_4 
+ bl[2] br[2] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_5 
+ bl[3] br[3] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_6 
+ bl[4] br[4] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_7 
+ bl[5] br[5] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_8 
+ bl[6] br[6] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_9 
+ bl[7] br[7] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_10 
+ bl[8] br[8] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_11 
+ bl[9] br[9] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_12 
+ bl[10] br[10] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_13 
+ bl[11] br[11] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_14 
+ bl[12] br[12] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_15 
+ bl[13] br[13] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_16 
+ bl[14] br[14] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_17 
+ bl[15] br[15] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_18 
+ bl[16] br[16] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_19 
+ bl[17] br[17] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_20 
+ bl[18] br[18] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_21 
+ bl[19] br[19] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_22 
+ bl[20] br[20] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_23 
+ bl[21] br[21] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_24 
+ bl[22] br[22] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_25 
+ bl[23] br[23] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_26 
+ bl[24] br[24] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_27 
+ bl[25] br[25] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_28 
+ bl[26] br[26] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_29 
+ bl[27] br[27] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_30 
+ bl[28] br[28] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_31 
+ bl[29] br[29] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_32 
+ bl[30] br[30] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_33 
+ bl[31] br[31] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_34 
+ bl[32] br[32] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_35 
+ bl[33] br[33] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_36 
+ bl[34] br[34] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_37 
+ bl[35] br[35] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_38 
+ bl[36] br[36] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_39 
+ bl[37] br[37] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_40 
+ bl[38] br[38] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_41 
+ bl[39] br[39] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_42 
+ bl[40] br[40] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_43 
+ bl[41] br[41] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_44 
+ bl[42] br[42] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_45 
+ bl[43] br[43] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_46 
+ bl[44] br[44] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_47 
+ bl[45] br[45] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_48 
+ bl[46] br[46] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_49 
+ bl[47] br[47] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_50 
+ bl[48] br[48] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_51 
+ bl[49] br[49] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_52 
+ bl[50] br[50] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_53 
+ bl[51] br[51] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_54 
+ bl[52] br[52] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_55 
+ bl[53] br[53] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_56 
+ bl[54] br[54] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_57 
+ bl[55] br[55] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_58 
+ bl[56] br[56] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_59 
+ bl[57] br[57] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_60 
+ bl[58] br[58] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_61 
+ bl[59] br[59] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_62 
+ bl[60] br[60] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_63 
+ bl[61] br[61] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_64 
+ bl[62] br[62] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_65 
+ bl[63] br[63] vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_66 
+ vdd vdd vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_191_67 
+ vdd vdd vdd vss wl[189] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_0 
+ vdd vdd vss vdd vpb vnb wl[190] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_192_1 
+ rbl rbr vss vdd vpb vnb wl[190] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_192_2 
+ bl[0] br[0] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_3 
+ bl[1] br[1] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_4 
+ bl[2] br[2] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_5 
+ bl[3] br[3] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_6 
+ bl[4] br[4] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_7 
+ bl[5] br[5] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_8 
+ bl[6] br[6] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_9 
+ bl[7] br[7] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_10 
+ bl[8] br[8] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_11 
+ bl[9] br[9] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_12 
+ bl[10] br[10] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_13 
+ bl[11] br[11] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_14 
+ bl[12] br[12] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_15 
+ bl[13] br[13] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_16 
+ bl[14] br[14] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_17 
+ bl[15] br[15] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_18 
+ bl[16] br[16] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_19 
+ bl[17] br[17] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_20 
+ bl[18] br[18] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_21 
+ bl[19] br[19] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_22 
+ bl[20] br[20] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_23 
+ bl[21] br[21] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_24 
+ bl[22] br[22] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_25 
+ bl[23] br[23] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_26 
+ bl[24] br[24] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_27 
+ bl[25] br[25] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_28 
+ bl[26] br[26] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_29 
+ bl[27] br[27] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_30 
+ bl[28] br[28] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_31 
+ bl[29] br[29] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_32 
+ bl[30] br[30] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_33 
+ bl[31] br[31] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_34 
+ bl[32] br[32] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_35 
+ bl[33] br[33] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_36 
+ bl[34] br[34] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_37 
+ bl[35] br[35] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_38 
+ bl[36] br[36] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_39 
+ bl[37] br[37] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_40 
+ bl[38] br[38] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_41 
+ bl[39] br[39] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_42 
+ bl[40] br[40] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_43 
+ bl[41] br[41] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_44 
+ bl[42] br[42] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_45 
+ bl[43] br[43] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_46 
+ bl[44] br[44] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_47 
+ bl[45] br[45] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_48 
+ bl[46] br[46] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_49 
+ bl[47] br[47] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_50 
+ bl[48] br[48] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_51 
+ bl[49] br[49] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_52 
+ bl[50] br[50] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_53 
+ bl[51] br[51] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_54 
+ bl[52] br[52] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_55 
+ bl[53] br[53] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_56 
+ bl[54] br[54] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_57 
+ bl[55] br[55] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_58 
+ bl[56] br[56] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_59 
+ bl[57] br[57] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_60 
+ bl[58] br[58] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_61 
+ bl[59] br[59] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_62 
+ bl[60] br[60] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_63 
+ bl[61] br[61] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_64 
+ bl[62] br[62] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_65 
+ bl[63] br[63] vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_66 
+ vdd vdd vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_192_67 
+ vdd vdd vdd vss wl[190] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_0 
+ vdd vdd vss vdd vpb vnb wl[191] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_193_1 
+ rbl rbr vss vdd vpb vnb wl[191] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_193_2 
+ bl[0] br[0] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_3 
+ bl[1] br[1] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_4 
+ bl[2] br[2] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_5 
+ bl[3] br[3] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_6 
+ bl[4] br[4] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_7 
+ bl[5] br[5] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_8 
+ bl[6] br[6] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_9 
+ bl[7] br[7] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_10 
+ bl[8] br[8] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_11 
+ bl[9] br[9] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_12 
+ bl[10] br[10] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_13 
+ bl[11] br[11] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_14 
+ bl[12] br[12] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_15 
+ bl[13] br[13] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_16 
+ bl[14] br[14] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_17 
+ bl[15] br[15] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_18 
+ bl[16] br[16] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_19 
+ bl[17] br[17] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_20 
+ bl[18] br[18] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_21 
+ bl[19] br[19] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_22 
+ bl[20] br[20] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_23 
+ bl[21] br[21] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_24 
+ bl[22] br[22] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_25 
+ bl[23] br[23] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_26 
+ bl[24] br[24] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_27 
+ bl[25] br[25] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_28 
+ bl[26] br[26] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_29 
+ bl[27] br[27] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_30 
+ bl[28] br[28] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_31 
+ bl[29] br[29] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_32 
+ bl[30] br[30] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_33 
+ bl[31] br[31] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_34 
+ bl[32] br[32] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_35 
+ bl[33] br[33] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_36 
+ bl[34] br[34] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_37 
+ bl[35] br[35] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_38 
+ bl[36] br[36] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_39 
+ bl[37] br[37] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_40 
+ bl[38] br[38] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_41 
+ bl[39] br[39] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_42 
+ bl[40] br[40] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_43 
+ bl[41] br[41] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_44 
+ bl[42] br[42] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_45 
+ bl[43] br[43] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_46 
+ bl[44] br[44] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_47 
+ bl[45] br[45] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_48 
+ bl[46] br[46] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_49 
+ bl[47] br[47] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_50 
+ bl[48] br[48] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_51 
+ bl[49] br[49] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_52 
+ bl[50] br[50] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_53 
+ bl[51] br[51] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_54 
+ bl[52] br[52] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_55 
+ bl[53] br[53] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_56 
+ bl[54] br[54] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_57 
+ bl[55] br[55] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_58 
+ bl[56] br[56] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_59 
+ bl[57] br[57] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_60 
+ bl[58] br[58] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_61 
+ bl[59] br[59] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_62 
+ bl[60] br[60] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_63 
+ bl[61] br[61] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_64 
+ bl[62] br[62] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_65 
+ bl[63] br[63] vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_66 
+ vdd vdd vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_193_67 
+ vdd vdd vdd vss wl[191] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_0 
+ vdd vdd vss vdd vpb vnb wl[192] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_194_1 
+ rbl rbr vss vdd vpb vnb wl[192] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_194_2 
+ bl[0] br[0] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_3 
+ bl[1] br[1] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_4 
+ bl[2] br[2] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_5 
+ bl[3] br[3] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_6 
+ bl[4] br[4] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_7 
+ bl[5] br[5] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_8 
+ bl[6] br[6] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_9 
+ bl[7] br[7] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_10 
+ bl[8] br[8] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_11 
+ bl[9] br[9] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_12 
+ bl[10] br[10] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_13 
+ bl[11] br[11] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_14 
+ bl[12] br[12] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_15 
+ bl[13] br[13] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_16 
+ bl[14] br[14] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_17 
+ bl[15] br[15] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_18 
+ bl[16] br[16] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_19 
+ bl[17] br[17] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_20 
+ bl[18] br[18] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_21 
+ bl[19] br[19] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_22 
+ bl[20] br[20] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_23 
+ bl[21] br[21] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_24 
+ bl[22] br[22] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_25 
+ bl[23] br[23] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_26 
+ bl[24] br[24] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_27 
+ bl[25] br[25] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_28 
+ bl[26] br[26] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_29 
+ bl[27] br[27] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_30 
+ bl[28] br[28] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_31 
+ bl[29] br[29] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_32 
+ bl[30] br[30] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_33 
+ bl[31] br[31] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_34 
+ bl[32] br[32] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_35 
+ bl[33] br[33] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_36 
+ bl[34] br[34] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_37 
+ bl[35] br[35] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_38 
+ bl[36] br[36] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_39 
+ bl[37] br[37] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_40 
+ bl[38] br[38] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_41 
+ bl[39] br[39] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_42 
+ bl[40] br[40] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_43 
+ bl[41] br[41] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_44 
+ bl[42] br[42] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_45 
+ bl[43] br[43] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_46 
+ bl[44] br[44] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_47 
+ bl[45] br[45] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_48 
+ bl[46] br[46] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_49 
+ bl[47] br[47] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_50 
+ bl[48] br[48] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_51 
+ bl[49] br[49] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_52 
+ bl[50] br[50] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_53 
+ bl[51] br[51] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_54 
+ bl[52] br[52] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_55 
+ bl[53] br[53] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_56 
+ bl[54] br[54] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_57 
+ bl[55] br[55] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_58 
+ bl[56] br[56] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_59 
+ bl[57] br[57] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_60 
+ bl[58] br[58] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_61 
+ bl[59] br[59] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_62 
+ bl[60] br[60] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_63 
+ bl[61] br[61] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_64 
+ bl[62] br[62] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_65 
+ bl[63] br[63] vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_66 
+ vdd vdd vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_194_67 
+ vdd vdd vdd vss wl[192] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_0 
+ vdd vdd vss vdd vpb vnb wl[193] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_195_1 
+ rbl rbr vss vdd vpb vnb wl[193] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_195_2 
+ bl[0] br[0] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_3 
+ bl[1] br[1] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_4 
+ bl[2] br[2] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_5 
+ bl[3] br[3] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_6 
+ bl[4] br[4] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_7 
+ bl[5] br[5] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_8 
+ bl[6] br[6] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_9 
+ bl[7] br[7] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_10 
+ bl[8] br[8] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_11 
+ bl[9] br[9] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_12 
+ bl[10] br[10] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_13 
+ bl[11] br[11] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_14 
+ bl[12] br[12] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_15 
+ bl[13] br[13] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_16 
+ bl[14] br[14] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_17 
+ bl[15] br[15] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_18 
+ bl[16] br[16] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_19 
+ bl[17] br[17] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_20 
+ bl[18] br[18] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_21 
+ bl[19] br[19] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_22 
+ bl[20] br[20] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_23 
+ bl[21] br[21] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_24 
+ bl[22] br[22] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_25 
+ bl[23] br[23] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_26 
+ bl[24] br[24] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_27 
+ bl[25] br[25] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_28 
+ bl[26] br[26] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_29 
+ bl[27] br[27] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_30 
+ bl[28] br[28] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_31 
+ bl[29] br[29] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_32 
+ bl[30] br[30] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_33 
+ bl[31] br[31] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_34 
+ bl[32] br[32] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_35 
+ bl[33] br[33] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_36 
+ bl[34] br[34] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_37 
+ bl[35] br[35] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_38 
+ bl[36] br[36] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_39 
+ bl[37] br[37] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_40 
+ bl[38] br[38] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_41 
+ bl[39] br[39] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_42 
+ bl[40] br[40] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_43 
+ bl[41] br[41] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_44 
+ bl[42] br[42] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_45 
+ bl[43] br[43] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_46 
+ bl[44] br[44] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_47 
+ bl[45] br[45] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_48 
+ bl[46] br[46] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_49 
+ bl[47] br[47] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_50 
+ bl[48] br[48] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_51 
+ bl[49] br[49] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_52 
+ bl[50] br[50] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_53 
+ bl[51] br[51] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_54 
+ bl[52] br[52] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_55 
+ bl[53] br[53] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_56 
+ bl[54] br[54] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_57 
+ bl[55] br[55] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_58 
+ bl[56] br[56] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_59 
+ bl[57] br[57] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_60 
+ bl[58] br[58] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_61 
+ bl[59] br[59] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_62 
+ bl[60] br[60] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_63 
+ bl[61] br[61] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_64 
+ bl[62] br[62] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_65 
+ bl[63] br[63] vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_66 
+ vdd vdd vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_195_67 
+ vdd vdd vdd vss wl[193] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_0 
+ vdd vdd vss vdd vpb vnb wl[194] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_196_1 
+ rbl rbr vss vdd vpb vnb wl[194] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_196_2 
+ bl[0] br[0] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_3 
+ bl[1] br[1] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_4 
+ bl[2] br[2] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_5 
+ bl[3] br[3] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_6 
+ bl[4] br[4] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_7 
+ bl[5] br[5] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_8 
+ bl[6] br[6] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_9 
+ bl[7] br[7] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_10 
+ bl[8] br[8] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_11 
+ bl[9] br[9] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_12 
+ bl[10] br[10] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_13 
+ bl[11] br[11] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_14 
+ bl[12] br[12] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_15 
+ bl[13] br[13] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_16 
+ bl[14] br[14] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_17 
+ bl[15] br[15] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_18 
+ bl[16] br[16] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_19 
+ bl[17] br[17] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_20 
+ bl[18] br[18] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_21 
+ bl[19] br[19] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_22 
+ bl[20] br[20] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_23 
+ bl[21] br[21] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_24 
+ bl[22] br[22] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_25 
+ bl[23] br[23] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_26 
+ bl[24] br[24] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_27 
+ bl[25] br[25] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_28 
+ bl[26] br[26] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_29 
+ bl[27] br[27] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_30 
+ bl[28] br[28] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_31 
+ bl[29] br[29] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_32 
+ bl[30] br[30] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_33 
+ bl[31] br[31] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_34 
+ bl[32] br[32] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_35 
+ bl[33] br[33] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_36 
+ bl[34] br[34] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_37 
+ bl[35] br[35] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_38 
+ bl[36] br[36] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_39 
+ bl[37] br[37] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_40 
+ bl[38] br[38] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_41 
+ bl[39] br[39] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_42 
+ bl[40] br[40] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_43 
+ bl[41] br[41] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_44 
+ bl[42] br[42] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_45 
+ bl[43] br[43] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_46 
+ bl[44] br[44] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_47 
+ bl[45] br[45] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_48 
+ bl[46] br[46] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_49 
+ bl[47] br[47] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_50 
+ bl[48] br[48] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_51 
+ bl[49] br[49] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_52 
+ bl[50] br[50] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_53 
+ bl[51] br[51] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_54 
+ bl[52] br[52] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_55 
+ bl[53] br[53] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_56 
+ bl[54] br[54] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_57 
+ bl[55] br[55] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_58 
+ bl[56] br[56] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_59 
+ bl[57] br[57] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_60 
+ bl[58] br[58] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_61 
+ bl[59] br[59] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_62 
+ bl[60] br[60] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_63 
+ bl[61] br[61] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_64 
+ bl[62] br[62] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_65 
+ bl[63] br[63] vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_66 
+ vdd vdd vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_196_67 
+ vdd vdd vdd vss wl[194] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_0 
+ vdd vdd vss vdd vpb vnb wl[195] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_197_1 
+ rbl rbr vss vdd vpb vnb wl[195] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_197_2 
+ bl[0] br[0] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_3 
+ bl[1] br[1] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_4 
+ bl[2] br[2] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_5 
+ bl[3] br[3] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_6 
+ bl[4] br[4] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_7 
+ bl[5] br[5] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_8 
+ bl[6] br[6] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_9 
+ bl[7] br[7] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_10 
+ bl[8] br[8] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_11 
+ bl[9] br[9] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_12 
+ bl[10] br[10] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_13 
+ bl[11] br[11] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_14 
+ bl[12] br[12] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_15 
+ bl[13] br[13] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_16 
+ bl[14] br[14] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_17 
+ bl[15] br[15] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_18 
+ bl[16] br[16] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_19 
+ bl[17] br[17] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_20 
+ bl[18] br[18] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_21 
+ bl[19] br[19] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_22 
+ bl[20] br[20] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_23 
+ bl[21] br[21] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_24 
+ bl[22] br[22] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_25 
+ bl[23] br[23] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_26 
+ bl[24] br[24] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_27 
+ bl[25] br[25] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_28 
+ bl[26] br[26] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_29 
+ bl[27] br[27] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_30 
+ bl[28] br[28] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_31 
+ bl[29] br[29] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_32 
+ bl[30] br[30] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_33 
+ bl[31] br[31] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_34 
+ bl[32] br[32] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_35 
+ bl[33] br[33] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_36 
+ bl[34] br[34] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_37 
+ bl[35] br[35] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_38 
+ bl[36] br[36] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_39 
+ bl[37] br[37] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_40 
+ bl[38] br[38] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_41 
+ bl[39] br[39] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_42 
+ bl[40] br[40] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_43 
+ bl[41] br[41] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_44 
+ bl[42] br[42] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_45 
+ bl[43] br[43] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_46 
+ bl[44] br[44] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_47 
+ bl[45] br[45] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_48 
+ bl[46] br[46] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_49 
+ bl[47] br[47] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_50 
+ bl[48] br[48] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_51 
+ bl[49] br[49] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_52 
+ bl[50] br[50] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_53 
+ bl[51] br[51] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_54 
+ bl[52] br[52] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_55 
+ bl[53] br[53] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_56 
+ bl[54] br[54] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_57 
+ bl[55] br[55] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_58 
+ bl[56] br[56] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_59 
+ bl[57] br[57] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_60 
+ bl[58] br[58] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_61 
+ bl[59] br[59] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_62 
+ bl[60] br[60] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_63 
+ bl[61] br[61] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_64 
+ bl[62] br[62] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_65 
+ bl[63] br[63] vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_66 
+ vdd vdd vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_197_67 
+ vdd vdd vdd vss wl[195] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_0 
+ vdd vdd vss vdd vpb vnb wl[196] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_198_1 
+ rbl rbr vss vdd vpb vnb wl[196] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_198_2 
+ bl[0] br[0] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_3 
+ bl[1] br[1] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_4 
+ bl[2] br[2] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_5 
+ bl[3] br[3] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_6 
+ bl[4] br[4] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_7 
+ bl[5] br[5] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_8 
+ bl[6] br[6] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_9 
+ bl[7] br[7] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_10 
+ bl[8] br[8] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_11 
+ bl[9] br[9] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_12 
+ bl[10] br[10] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_13 
+ bl[11] br[11] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_14 
+ bl[12] br[12] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_15 
+ bl[13] br[13] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_16 
+ bl[14] br[14] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_17 
+ bl[15] br[15] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_18 
+ bl[16] br[16] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_19 
+ bl[17] br[17] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_20 
+ bl[18] br[18] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_21 
+ bl[19] br[19] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_22 
+ bl[20] br[20] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_23 
+ bl[21] br[21] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_24 
+ bl[22] br[22] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_25 
+ bl[23] br[23] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_26 
+ bl[24] br[24] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_27 
+ bl[25] br[25] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_28 
+ bl[26] br[26] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_29 
+ bl[27] br[27] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_30 
+ bl[28] br[28] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_31 
+ bl[29] br[29] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_32 
+ bl[30] br[30] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_33 
+ bl[31] br[31] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_34 
+ bl[32] br[32] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_35 
+ bl[33] br[33] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_36 
+ bl[34] br[34] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_37 
+ bl[35] br[35] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_38 
+ bl[36] br[36] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_39 
+ bl[37] br[37] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_40 
+ bl[38] br[38] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_41 
+ bl[39] br[39] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_42 
+ bl[40] br[40] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_43 
+ bl[41] br[41] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_44 
+ bl[42] br[42] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_45 
+ bl[43] br[43] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_46 
+ bl[44] br[44] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_47 
+ bl[45] br[45] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_48 
+ bl[46] br[46] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_49 
+ bl[47] br[47] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_50 
+ bl[48] br[48] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_51 
+ bl[49] br[49] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_52 
+ bl[50] br[50] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_53 
+ bl[51] br[51] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_54 
+ bl[52] br[52] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_55 
+ bl[53] br[53] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_56 
+ bl[54] br[54] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_57 
+ bl[55] br[55] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_58 
+ bl[56] br[56] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_59 
+ bl[57] br[57] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_60 
+ bl[58] br[58] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_61 
+ bl[59] br[59] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_62 
+ bl[60] br[60] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_63 
+ bl[61] br[61] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_64 
+ bl[62] br[62] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_65 
+ bl[63] br[63] vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_66 
+ vdd vdd vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_198_67 
+ vdd vdd vdd vss wl[196] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_0 
+ vdd vdd vss vdd vpb vnb wl[197] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_199_1 
+ rbl rbr vss vdd vpb vnb wl[197] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_199_2 
+ bl[0] br[0] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_3 
+ bl[1] br[1] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_4 
+ bl[2] br[2] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_5 
+ bl[3] br[3] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_6 
+ bl[4] br[4] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_7 
+ bl[5] br[5] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_8 
+ bl[6] br[6] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_9 
+ bl[7] br[7] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_10 
+ bl[8] br[8] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_11 
+ bl[9] br[9] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_12 
+ bl[10] br[10] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_13 
+ bl[11] br[11] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_14 
+ bl[12] br[12] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_15 
+ bl[13] br[13] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_16 
+ bl[14] br[14] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_17 
+ bl[15] br[15] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_18 
+ bl[16] br[16] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_19 
+ bl[17] br[17] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_20 
+ bl[18] br[18] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_21 
+ bl[19] br[19] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_22 
+ bl[20] br[20] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_23 
+ bl[21] br[21] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_24 
+ bl[22] br[22] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_25 
+ bl[23] br[23] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_26 
+ bl[24] br[24] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_27 
+ bl[25] br[25] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_28 
+ bl[26] br[26] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_29 
+ bl[27] br[27] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_30 
+ bl[28] br[28] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_31 
+ bl[29] br[29] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_32 
+ bl[30] br[30] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_33 
+ bl[31] br[31] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_34 
+ bl[32] br[32] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_35 
+ bl[33] br[33] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_36 
+ bl[34] br[34] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_37 
+ bl[35] br[35] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_38 
+ bl[36] br[36] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_39 
+ bl[37] br[37] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_40 
+ bl[38] br[38] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_41 
+ bl[39] br[39] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_42 
+ bl[40] br[40] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_43 
+ bl[41] br[41] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_44 
+ bl[42] br[42] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_45 
+ bl[43] br[43] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_46 
+ bl[44] br[44] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_47 
+ bl[45] br[45] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_48 
+ bl[46] br[46] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_49 
+ bl[47] br[47] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_50 
+ bl[48] br[48] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_51 
+ bl[49] br[49] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_52 
+ bl[50] br[50] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_53 
+ bl[51] br[51] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_54 
+ bl[52] br[52] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_55 
+ bl[53] br[53] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_56 
+ bl[54] br[54] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_57 
+ bl[55] br[55] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_58 
+ bl[56] br[56] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_59 
+ bl[57] br[57] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_60 
+ bl[58] br[58] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_61 
+ bl[59] br[59] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_62 
+ bl[60] br[60] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_63 
+ bl[61] br[61] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_64 
+ bl[62] br[62] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_65 
+ bl[63] br[63] vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_66 
+ vdd vdd vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_199_67 
+ vdd vdd vdd vss wl[197] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_0 
+ vdd vdd vss vdd vpb vnb wl[198] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_200_1 
+ rbl rbr vss vdd vpb vnb wl[198] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_200_2 
+ bl[0] br[0] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_3 
+ bl[1] br[1] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_4 
+ bl[2] br[2] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_5 
+ bl[3] br[3] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_6 
+ bl[4] br[4] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_7 
+ bl[5] br[5] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_8 
+ bl[6] br[6] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_9 
+ bl[7] br[7] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_10 
+ bl[8] br[8] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_11 
+ bl[9] br[9] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_12 
+ bl[10] br[10] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_13 
+ bl[11] br[11] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_14 
+ bl[12] br[12] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_15 
+ bl[13] br[13] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_16 
+ bl[14] br[14] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_17 
+ bl[15] br[15] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_18 
+ bl[16] br[16] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_19 
+ bl[17] br[17] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_20 
+ bl[18] br[18] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_21 
+ bl[19] br[19] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_22 
+ bl[20] br[20] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_23 
+ bl[21] br[21] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_24 
+ bl[22] br[22] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_25 
+ bl[23] br[23] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_26 
+ bl[24] br[24] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_27 
+ bl[25] br[25] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_28 
+ bl[26] br[26] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_29 
+ bl[27] br[27] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_30 
+ bl[28] br[28] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_31 
+ bl[29] br[29] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_32 
+ bl[30] br[30] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_33 
+ bl[31] br[31] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_34 
+ bl[32] br[32] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_35 
+ bl[33] br[33] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_36 
+ bl[34] br[34] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_37 
+ bl[35] br[35] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_38 
+ bl[36] br[36] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_39 
+ bl[37] br[37] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_40 
+ bl[38] br[38] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_41 
+ bl[39] br[39] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_42 
+ bl[40] br[40] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_43 
+ bl[41] br[41] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_44 
+ bl[42] br[42] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_45 
+ bl[43] br[43] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_46 
+ bl[44] br[44] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_47 
+ bl[45] br[45] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_48 
+ bl[46] br[46] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_49 
+ bl[47] br[47] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_50 
+ bl[48] br[48] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_51 
+ bl[49] br[49] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_52 
+ bl[50] br[50] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_53 
+ bl[51] br[51] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_54 
+ bl[52] br[52] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_55 
+ bl[53] br[53] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_56 
+ bl[54] br[54] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_57 
+ bl[55] br[55] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_58 
+ bl[56] br[56] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_59 
+ bl[57] br[57] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_60 
+ bl[58] br[58] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_61 
+ bl[59] br[59] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_62 
+ bl[60] br[60] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_63 
+ bl[61] br[61] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_64 
+ bl[62] br[62] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_65 
+ bl[63] br[63] vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_66 
+ vdd vdd vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_200_67 
+ vdd vdd vdd vss wl[198] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_0 
+ vdd vdd vss vdd vpb vnb wl[199] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_201_1 
+ rbl rbr vss vdd vpb vnb wl[199] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_201_2 
+ bl[0] br[0] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_3 
+ bl[1] br[1] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_4 
+ bl[2] br[2] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_5 
+ bl[3] br[3] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_6 
+ bl[4] br[4] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_7 
+ bl[5] br[5] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_8 
+ bl[6] br[6] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_9 
+ bl[7] br[7] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_10 
+ bl[8] br[8] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_11 
+ bl[9] br[9] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_12 
+ bl[10] br[10] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_13 
+ bl[11] br[11] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_14 
+ bl[12] br[12] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_15 
+ bl[13] br[13] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_16 
+ bl[14] br[14] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_17 
+ bl[15] br[15] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_18 
+ bl[16] br[16] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_19 
+ bl[17] br[17] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_20 
+ bl[18] br[18] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_21 
+ bl[19] br[19] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_22 
+ bl[20] br[20] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_23 
+ bl[21] br[21] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_24 
+ bl[22] br[22] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_25 
+ bl[23] br[23] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_26 
+ bl[24] br[24] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_27 
+ bl[25] br[25] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_28 
+ bl[26] br[26] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_29 
+ bl[27] br[27] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_30 
+ bl[28] br[28] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_31 
+ bl[29] br[29] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_32 
+ bl[30] br[30] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_33 
+ bl[31] br[31] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_34 
+ bl[32] br[32] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_35 
+ bl[33] br[33] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_36 
+ bl[34] br[34] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_37 
+ bl[35] br[35] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_38 
+ bl[36] br[36] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_39 
+ bl[37] br[37] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_40 
+ bl[38] br[38] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_41 
+ bl[39] br[39] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_42 
+ bl[40] br[40] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_43 
+ bl[41] br[41] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_44 
+ bl[42] br[42] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_45 
+ bl[43] br[43] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_46 
+ bl[44] br[44] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_47 
+ bl[45] br[45] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_48 
+ bl[46] br[46] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_49 
+ bl[47] br[47] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_50 
+ bl[48] br[48] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_51 
+ bl[49] br[49] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_52 
+ bl[50] br[50] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_53 
+ bl[51] br[51] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_54 
+ bl[52] br[52] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_55 
+ bl[53] br[53] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_56 
+ bl[54] br[54] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_57 
+ bl[55] br[55] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_58 
+ bl[56] br[56] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_59 
+ bl[57] br[57] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_60 
+ bl[58] br[58] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_61 
+ bl[59] br[59] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_62 
+ bl[60] br[60] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_63 
+ bl[61] br[61] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_64 
+ bl[62] br[62] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_65 
+ bl[63] br[63] vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_66 
+ vdd vdd vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_201_67 
+ vdd vdd vdd vss wl[199] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_0 
+ vdd vdd vss vdd vpb vnb wl[200] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_202_1 
+ rbl rbr vss vdd vpb vnb wl[200] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_202_2 
+ bl[0] br[0] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_3 
+ bl[1] br[1] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_4 
+ bl[2] br[2] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_5 
+ bl[3] br[3] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_6 
+ bl[4] br[4] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_7 
+ bl[5] br[5] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_8 
+ bl[6] br[6] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_9 
+ bl[7] br[7] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_10 
+ bl[8] br[8] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_11 
+ bl[9] br[9] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_12 
+ bl[10] br[10] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_13 
+ bl[11] br[11] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_14 
+ bl[12] br[12] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_15 
+ bl[13] br[13] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_16 
+ bl[14] br[14] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_17 
+ bl[15] br[15] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_18 
+ bl[16] br[16] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_19 
+ bl[17] br[17] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_20 
+ bl[18] br[18] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_21 
+ bl[19] br[19] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_22 
+ bl[20] br[20] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_23 
+ bl[21] br[21] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_24 
+ bl[22] br[22] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_25 
+ bl[23] br[23] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_26 
+ bl[24] br[24] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_27 
+ bl[25] br[25] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_28 
+ bl[26] br[26] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_29 
+ bl[27] br[27] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_30 
+ bl[28] br[28] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_31 
+ bl[29] br[29] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_32 
+ bl[30] br[30] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_33 
+ bl[31] br[31] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_34 
+ bl[32] br[32] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_35 
+ bl[33] br[33] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_36 
+ bl[34] br[34] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_37 
+ bl[35] br[35] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_38 
+ bl[36] br[36] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_39 
+ bl[37] br[37] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_40 
+ bl[38] br[38] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_41 
+ bl[39] br[39] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_42 
+ bl[40] br[40] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_43 
+ bl[41] br[41] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_44 
+ bl[42] br[42] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_45 
+ bl[43] br[43] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_46 
+ bl[44] br[44] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_47 
+ bl[45] br[45] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_48 
+ bl[46] br[46] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_49 
+ bl[47] br[47] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_50 
+ bl[48] br[48] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_51 
+ bl[49] br[49] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_52 
+ bl[50] br[50] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_53 
+ bl[51] br[51] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_54 
+ bl[52] br[52] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_55 
+ bl[53] br[53] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_56 
+ bl[54] br[54] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_57 
+ bl[55] br[55] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_58 
+ bl[56] br[56] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_59 
+ bl[57] br[57] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_60 
+ bl[58] br[58] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_61 
+ bl[59] br[59] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_62 
+ bl[60] br[60] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_63 
+ bl[61] br[61] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_64 
+ bl[62] br[62] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_65 
+ bl[63] br[63] vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_66 
+ vdd vdd vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_202_67 
+ vdd vdd vdd vss wl[200] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_0 
+ vdd vdd vss vdd vpb vnb wl[201] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_203_1 
+ rbl rbr vss vdd vpb vnb wl[201] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_203_2 
+ bl[0] br[0] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_3 
+ bl[1] br[1] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_4 
+ bl[2] br[2] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_5 
+ bl[3] br[3] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_6 
+ bl[4] br[4] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_7 
+ bl[5] br[5] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_8 
+ bl[6] br[6] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_9 
+ bl[7] br[7] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_10 
+ bl[8] br[8] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_11 
+ bl[9] br[9] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_12 
+ bl[10] br[10] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_13 
+ bl[11] br[11] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_14 
+ bl[12] br[12] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_15 
+ bl[13] br[13] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_16 
+ bl[14] br[14] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_17 
+ bl[15] br[15] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_18 
+ bl[16] br[16] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_19 
+ bl[17] br[17] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_20 
+ bl[18] br[18] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_21 
+ bl[19] br[19] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_22 
+ bl[20] br[20] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_23 
+ bl[21] br[21] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_24 
+ bl[22] br[22] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_25 
+ bl[23] br[23] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_26 
+ bl[24] br[24] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_27 
+ bl[25] br[25] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_28 
+ bl[26] br[26] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_29 
+ bl[27] br[27] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_30 
+ bl[28] br[28] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_31 
+ bl[29] br[29] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_32 
+ bl[30] br[30] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_33 
+ bl[31] br[31] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_34 
+ bl[32] br[32] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_35 
+ bl[33] br[33] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_36 
+ bl[34] br[34] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_37 
+ bl[35] br[35] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_38 
+ bl[36] br[36] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_39 
+ bl[37] br[37] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_40 
+ bl[38] br[38] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_41 
+ bl[39] br[39] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_42 
+ bl[40] br[40] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_43 
+ bl[41] br[41] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_44 
+ bl[42] br[42] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_45 
+ bl[43] br[43] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_46 
+ bl[44] br[44] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_47 
+ bl[45] br[45] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_48 
+ bl[46] br[46] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_49 
+ bl[47] br[47] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_50 
+ bl[48] br[48] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_51 
+ bl[49] br[49] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_52 
+ bl[50] br[50] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_53 
+ bl[51] br[51] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_54 
+ bl[52] br[52] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_55 
+ bl[53] br[53] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_56 
+ bl[54] br[54] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_57 
+ bl[55] br[55] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_58 
+ bl[56] br[56] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_59 
+ bl[57] br[57] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_60 
+ bl[58] br[58] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_61 
+ bl[59] br[59] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_62 
+ bl[60] br[60] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_63 
+ bl[61] br[61] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_64 
+ bl[62] br[62] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_65 
+ bl[63] br[63] vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_66 
+ vdd vdd vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_203_67 
+ vdd vdd vdd vss wl[201] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_0 
+ vdd vdd vss vdd vpb vnb wl[202] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_204_1 
+ rbl rbr vss vdd vpb vnb wl[202] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_204_2 
+ bl[0] br[0] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_3 
+ bl[1] br[1] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_4 
+ bl[2] br[2] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_5 
+ bl[3] br[3] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_6 
+ bl[4] br[4] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_7 
+ bl[5] br[5] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_8 
+ bl[6] br[6] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_9 
+ bl[7] br[7] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_10 
+ bl[8] br[8] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_11 
+ bl[9] br[9] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_12 
+ bl[10] br[10] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_13 
+ bl[11] br[11] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_14 
+ bl[12] br[12] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_15 
+ bl[13] br[13] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_16 
+ bl[14] br[14] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_17 
+ bl[15] br[15] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_18 
+ bl[16] br[16] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_19 
+ bl[17] br[17] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_20 
+ bl[18] br[18] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_21 
+ bl[19] br[19] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_22 
+ bl[20] br[20] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_23 
+ bl[21] br[21] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_24 
+ bl[22] br[22] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_25 
+ bl[23] br[23] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_26 
+ bl[24] br[24] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_27 
+ bl[25] br[25] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_28 
+ bl[26] br[26] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_29 
+ bl[27] br[27] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_30 
+ bl[28] br[28] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_31 
+ bl[29] br[29] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_32 
+ bl[30] br[30] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_33 
+ bl[31] br[31] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_34 
+ bl[32] br[32] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_35 
+ bl[33] br[33] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_36 
+ bl[34] br[34] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_37 
+ bl[35] br[35] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_38 
+ bl[36] br[36] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_39 
+ bl[37] br[37] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_40 
+ bl[38] br[38] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_41 
+ bl[39] br[39] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_42 
+ bl[40] br[40] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_43 
+ bl[41] br[41] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_44 
+ bl[42] br[42] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_45 
+ bl[43] br[43] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_46 
+ bl[44] br[44] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_47 
+ bl[45] br[45] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_48 
+ bl[46] br[46] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_49 
+ bl[47] br[47] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_50 
+ bl[48] br[48] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_51 
+ bl[49] br[49] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_52 
+ bl[50] br[50] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_53 
+ bl[51] br[51] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_54 
+ bl[52] br[52] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_55 
+ bl[53] br[53] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_56 
+ bl[54] br[54] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_57 
+ bl[55] br[55] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_58 
+ bl[56] br[56] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_59 
+ bl[57] br[57] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_60 
+ bl[58] br[58] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_61 
+ bl[59] br[59] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_62 
+ bl[60] br[60] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_63 
+ bl[61] br[61] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_64 
+ bl[62] br[62] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_65 
+ bl[63] br[63] vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_66 
+ vdd vdd vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_204_67 
+ vdd vdd vdd vss wl[202] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_0 
+ vdd vdd vss vdd vpb vnb wl[203] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_205_1 
+ rbl rbr vss vdd vpb vnb wl[203] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_205_2 
+ bl[0] br[0] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_3 
+ bl[1] br[1] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_4 
+ bl[2] br[2] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_5 
+ bl[3] br[3] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_6 
+ bl[4] br[4] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_7 
+ bl[5] br[5] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_8 
+ bl[6] br[6] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_9 
+ bl[7] br[7] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_10 
+ bl[8] br[8] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_11 
+ bl[9] br[9] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_12 
+ bl[10] br[10] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_13 
+ bl[11] br[11] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_14 
+ bl[12] br[12] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_15 
+ bl[13] br[13] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_16 
+ bl[14] br[14] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_17 
+ bl[15] br[15] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_18 
+ bl[16] br[16] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_19 
+ bl[17] br[17] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_20 
+ bl[18] br[18] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_21 
+ bl[19] br[19] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_22 
+ bl[20] br[20] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_23 
+ bl[21] br[21] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_24 
+ bl[22] br[22] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_25 
+ bl[23] br[23] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_26 
+ bl[24] br[24] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_27 
+ bl[25] br[25] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_28 
+ bl[26] br[26] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_29 
+ bl[27] br[27] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_30 
+ bl[28] br[28] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_31 
+ bl[29] br[29] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_32 
+ bl[30] br[30] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_33 
+ bl[31] br[31] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_34 
+ bl[32] br[32] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_35 
+ bl[33] br[33] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_36 
+ bl[34] br[34] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_37 
+ bl[35] br[35] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_38 
+ bl[36] br[36] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_39 
+ bl[37] br[37] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_40 
+ bl[38] br[38] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_41 
+ bl[39] br[39] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_42 
+ bl[40] br[40] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_43 
+ bl[41] br[41] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_44 
+ bl[42] br[42] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_45 
+ bl[43] br[43] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_46 
+ bl[44] br[44] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_47 
+ bl[45] br[45] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_48 
+ bl[46] br[46] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_49 
+ bl[47] br[47] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_50 
+ bl[48] br[48] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_51 
+ bl[49] br[49] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_52 
+ bl[50] br[50] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_53 
+ bl[51] br[51] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_54 
+ bl[52] br[52] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_55 
+ bl[53] br[53] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_56 
+ bl[54] br[54] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_57 
+ bl[55] br[55] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_58 
+ bl[56] br[56] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_59 
+ bl[57] br[57] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_60 
+ bl[58] br[58] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_61 
+ bl[59] br[59] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_62 
+ bl[60] br[60] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_63 
+ bl[61] br[61] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_64 
+ bl[62] br[62] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_65 
+ bl[63] br[63] vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_66 
+ vdd vdd vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_205_67 
+ vdd vdd vdd vss wl[203] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_0 
+ vdd vdd vss vdd vpb vnb wl[204] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_206_1 
+ rbl rbr vss vdd vpb vnb wl[204] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_206_2 
+ bl[0] br[0] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_3 
+ bl[1] br[1] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_4 
+ bl[2] br[2] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_5 
+ bl[3] br[3] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_6 
+ bl[4] br[4] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_7 
+ bl[5] br[5] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_8 
+ bl[6] br[6] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_9 
+ bl[7] br[7] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_10 
+ bl[8] br[8] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_11 
+ bl[9] br[9] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_12 
+ bl[10] br[10] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_13 
+ bl[11] br[11] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_14 
+ bl[12] br[12] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_15 
+ bl[13] br[13] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_16 
+ bl[14] br[14] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_17 
+ bl[15] br[15] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_18 
+ bl[16] br[16] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_19 
+ bl[17] br[17] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_20 
+ bl[18] br[18] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_21 
+ bl[19] br[19] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_22 
+ bl[20] br[20] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_23 
+ bl[21] br[21] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_24 
+ bl[22] br[22] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_25 
+ bl[23] br[23] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_26 
+ bl[24] br[24] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_27 
+ bl[25] br[25] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_28 
+ bl[26] br[26] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_29 
+ bl[27] br[27] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_30 
+ bl[28] br[28] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_31 
+ bl[29] br[29] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_32 
+ bl[30] br[30] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_33 
+ bl[31] br[31] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_34 
+ bl[32] br[32] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_35 
+ bl[33] br[33] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_36 
+ bl[34] br[34] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_37 
+ bl[35] br[35] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_38 
+ bl[36] br[36] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_39 
+ bl[37] br[37] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_40 
+ bl[38] br[38] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_41 
+ bl[39] br[39] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_42 
+ bl[40] br[40] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_43 
+ bl[41] br[41] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_44 
+ bl[42] br[42] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_45 
+ bl[43] br[43] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_46 
+ bl[44] br[44] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_47 
+ bl[45] br[45] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_48 
+ bl[46] br[46] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_49 
+ bl[47] br[47] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_50 
+ bl[48] br[48] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_51 
+ bl[49] br[49] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_52 
+ bl[50] br[50] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_53 
+ bl[51] br[51] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_54 
+ bl[52] br[52] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_55 
+ bl[53] br[53] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_56 
+ bl[54] br[54] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_57 
+ bl[55] br[55] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_58 
+ bl[56] br[56] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_59 
+ bl[57] br[57] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_60 
+ bl[58] br[58] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_61 
+ bl[59] br[59] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_62 
+ bl[60] br[60] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_63 
+ bl[61] br[61] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_64 
+ bl[62] br[62] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_65 
+ bl[63] br[63] vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_66 
+ vdd vdd vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_206_67 
+ vdd vdd vdd vss wl[204] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_0 
+ vdd vdd vss vdd vpb vnb wl[205] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_207_1 
+ rbl rbr vss vdd vpb vnb wl[205] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_207_2 
+ bl[0] br[0] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_3 
+ bl[1] br[1] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_4 
+ bl[2] br[2] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_5 
+ bl[3] br[3] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_6 
+ bl[4] br[4] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_7 
+ bl[5] br[5] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_8 
+ bl[6] br[6] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_9 
+ bl[7] br[7] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_10 
+ bl[8] br[8] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_11 
+ bl[9] br[9] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_12 
+ bl[10] br[10] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_13 
+ bl[11] br[11] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_14 
+ bl[12] br[12] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_15 
+ bl[13] br[13] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_16 
+ bl[14] br[14] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_17 
+ bl[15] br[15] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_18 
+ bl[16] br[16] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_19 
+ bl[17] br[17] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_20 
+ bl[18] br[18] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_21 
+ bl[19] br[19] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_22 
+ bl[20] br[20] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_23 
+ bl[21] br[21] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_24 
+ bl[22] br[22] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_25 
+ bl[23] br[23] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_26 
+ bl[24] br[24] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_27 
+ bl[25] br[25] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_28 
+ bl[26] br[26] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_29 
+ bl[27] br[27] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_30 
+ bl[28] br[28] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_31 
+ bl[29] br[29] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_32 
+ bl[30] br[30] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_33 
+ bl[31] br[31] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_34 
+ bl[32] br[32] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_35 
+ bl[33] br[33] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_36 
+ bl[34] br[34] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_37 
+ bl[35] br[35] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_38 
+ bl[36] br[36] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_39 
+ bl[37] br[37] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_40 
+ bl[38] br[38] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_41 
+ bl[39] br[39] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_42 
+ bl[40] br[40] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_43 
+ bl[41] br[41] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_44 
+ bl[42] br[42] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_45 
+ bl[43] br[43] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_46 
+ bl[44] br[44] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_47 
+ bl[45] br[45] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_48 
+ bl[46] br[46] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_49 
+ bl[47] br[47] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_50 
+ bl[48] br[48] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_51 
+ bl[49] br[49] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_52 
+ bl[50] br[50] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_53 
+ bl[51] br[51] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_54 
+ bl[52] br[52] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_55 
+ bl[53] br[53] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_56 
+ bl[54] br[54] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_57 
+ bl[55] br[55] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_58 
+ bl[56] br[56] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_59 
+ bl[57] br[57] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_60 
+ bl[58] br[58] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_61 
+ bl[59] br[59] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_62 
+ bl[60] br[60] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_63 
+ bl[61] br[61] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_64 
+ bl[62] br[62] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_65 
+ bl[63] br[63] vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_66 
+ vdd vdd vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_207_67 
+ vdd vdd vdd vss wl[205] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_0 
+ vdd vdd vss vdd vpb vnb wl[206] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_208_1 
+ rbl rbr vss vdd vpb vnb wl[206] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_208_2 
+ bl[0] br[0] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_3 
+ bl[1] br[1] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_4 
+ bl[2] br[2] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_5 
+ bl[3] br[3] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_6 
+ bl[4] br[4] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_7 
+ bl[5] br[5] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_8 
+ bl[6] br[6] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_9 
+ bl[7] br[7] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_10 
+ bl[8] br[8] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_11 
+ bl[9] br[9] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_12 
+ bl[10] br[10] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_13 
+ bl[11] br[11] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_14 
+ bl[12] br[12] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_15 
+ bl[13] br[13] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_16 
+ bl[14] br[14] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_17 
+ bl[15] br[15] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_18 
+ bl[16] br[16] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_19 
+ bl[17] br[17] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_20 
+ bl[18] br[18] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_21 
+ bl[19] br[19] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_22 
+ bl[20] br[20] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_23 
+ bl[21] br[21] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_24 
+ bl[22] br[22] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_25 
+ bl[23] br[23] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_26 
+ bl[24] br[24] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_27 
+ bl[25] br[25] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_28 
+ bl[26] br[26] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_29 
+ bl[27] br[27] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_30 
+ bl[28] br[28] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_31 
+ bl[29] br[29] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_32 
+ bl[30] br[30] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_33 
+ bl[31] br[31] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_34 
+ bl[32] br[32] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_35 
+ bl[33] br[33] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_36 
+ bl[34] br[34] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_37 
+ bl[35] br[35] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_38 
+ bl[36] br[36] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_39 
+ bl[37] br[37] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_40 
+ bl[38] br[38] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_41 
+ bl[39] br[39] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_42 
+ bl[40] br[40] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_43 
+ bl[41] br[41] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_44 
+ bl[42] br[42] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_45 
+ bl[43] br[43] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_46 
+ bl[44] br[44] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_47 
+ bl[45] br[45] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_48 
+ bl[46] br[46] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_49 
+ bl[47] br[47] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_50 
+ bl[48] br[48] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_51 
+ bl[49] br[49] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_52 
+ bl[50] br[50] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_53 
+ bl[51] br[51] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_54 
+ bl[52] br[52] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_55 
+ bl[53] br[53] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_56 
+ bl[54] br[54] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_57 
+ bl[55] br[55] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_58 
+ bl[56] br[56] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_59 
+ bl[57] br[57] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_60 
+ bl[58] br[58] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_61 
+ bl[59] br[59] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_62 
+ bl[60] br[60] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_63 
+ bl[61] br[61] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_64 
+ bl[62] br[62] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_65 
+ bl[63] br[63] vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_66 
+ vdd vdd vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_208_67 
+ vdd vdd vdd vss wl[206] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_0 
+ vdd vdd vss vdd vpb vnb wl[207] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_209_1 
+ rbl rbr vss vdd vpb vnb wl[207] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_209_2 
+ bl[0] br[0] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_3 
+ bl[1] br[1] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_4 
+ bl[2] br[2] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_5 
+ bl[3] br[3] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_6 
+ bl[4] br[4] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_7 
+ bl[5] br[5] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_8 
+ bl[6] br[6] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_9 
+ bl[7] br[7] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_10 
+ bl[8] br[8] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_11 
+ bl[9] br[9] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_12 
+ bl[10] br[10] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_13 
+ bl[11] br[11] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_14 
+ bl[12] br[12] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_15 
+ bl[13] br[13] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_16 
+ bl[14] br[14] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_17 
+ bl[15] br[15] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_18 
+ bl[16] br[16] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_19 
+ bl[17] br[17] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_20 
+ bl[18] br[18] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_21 
+ bl[19] br[19] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_22 
+ bl[20] br[20] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_23 
+ bl[21] br[21] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_24 
+ bl[22] br[22] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_25 
+ bl[23] br[23] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_26 
+ bl[24] br[24] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_27 
+ bl[25] br[25] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_28 
+ bl[26] br[26] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_29 
+ bl[27] br[27] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_30 
+ bl[28] br[28] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_31 
+ bl[29] br[29] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_32 
+ bl[30] br[30] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_33 
+ bl[31] br[31] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_34 
+ bl[32] br[32] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_35 
+ bl[33] br[33] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_36 
+ bl[34] br[34] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_37 
+ bl[35] br[35] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_38 
+ bl[36] br[36] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_39 
+ bl[37] br[37] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_40 
+ bl[38] br[38] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_41 
+ bl[39] br[39] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_42 
+ bl[40] br[40] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_43 
+ bl[41] br[41] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_44 
+ bl[42] br[42] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_45 
+ bl[43] br[43] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_46 
+ bl[44] br[44] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_47 
+ bl[45] br[45] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_48 
+ bl[46] br[46] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_49 
+ bl[47] br[47] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_50 
+ bl[48] br[48] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_51 
+ bl[49] br[49] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_52 
+ bl[50] br[50] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_53 
+ bl[51] br[51] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_54 
+ bl[52] br[52] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_55 
+ bl[53] br[53] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_56 
+ bl[54] br[54] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_57 
+ bl[55] br[55] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_58 
+ bl[56] br[56] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_59 
+ bl[57] br[57] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_60 
+ bl[58] br[58] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_61 
+ bl[59] br[59] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_62 
+ bl[60] br[60] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_63 
+ bl[61] br[61] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_64 
+ bl[62] br[62] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_65 
+ bl[63] br[63] vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_66 
+ vdd vdd vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_209_67 
+ vdd vdd vdd vss wl[207] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_0 
+ vdd vdd vss vdd vpb vnb wl[208] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_210_1 
+ rbl rbr vss vdd vpb vnb wl[208] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_210_2 
+ bl[0] br[0] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_3 
+ bl[1] br[1] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_4 
+ bl[2] br[2] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_5 
+ bl[3] br[3] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_6 
+ bl[4] br[4] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_7 
+ bl[5] br[5] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_8 
+ bl[6] br[6] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_9 
+ bl[7] br[7] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_10 
+ bl[8] br[8] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_11 
+ bl[9] br[9] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_12 
+ bl[10] br[10] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_13 
+ bl[11] br[11] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_14 
+ bl[12] br[12] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_15 
+ bl[13] br[13] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_16 
+ bl[14] br[14] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_17 
+ bl[15] br[15] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_18 
+ bl[16] br[16] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_19 
+ bl[17] br[17] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_20 
+ bl[18] br[18] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_21 
+ bl[19] br[19] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_22 
+ bl[20] br[20] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_23 
+ bl[21] br[21] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_24 
+ bl[22] br[22] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_25 
+ bl[23] br[23] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_26 
+ bl[24] br[24] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_27 
+ bl[25] br[25] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_28 
+ bl[26] br[26] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_29 
+ bl[27] br[27] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_30 
+ bl[28] br[28] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_31 
+ bl[29] br[29] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_32 
+ bl[30] br[30] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_33 
+ bl[31] br[31] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_34 
+ bl[32] br[32] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_35 
+ bl[33] br[33] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_36 
+ bl[34] br[34] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_37 
+ bl[35] br[35] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_38 
+ bl[36] br[36] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_39 
+ bl[37] br[37] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_40 
+ bl[38] br[38] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_41 
+ bl[39] br[39] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_42 
+ bl[40] br[40] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_43 
+ bl[41] br[41] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_44 
+ bl[42] br[42] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_45 
+ bl[43] br[43] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_46 
+ bl[44] br[44] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_47 
+ bl[45] br[45] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_48 
+ bl[46] br[46] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_49 
+ bl[47] br[47] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_50 
+ bl[48] br[48] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_51 
+ bl[49] br[49] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_52 
+ bl[50] br[50] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_53 
+ bl[51] br[51] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_54 
+ bl[52] br[52] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_55 
+ bl[53] br[53] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_56 
+ bl[54] br[54] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_57 
+ bl[55] br[55] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_58 
+ bl[56] br[56] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_59 
+ bl[57] br[57] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_60 
+ bl[58] br[58] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_61 
+ bl[59] br[59] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_62 
+ bl[60] br[60] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_63 
+ bl[61] br[61] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_64 
+ bl[62] br[62] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_65 
+ bl[63] br[63] vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_66 
+ vdd vdd vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_210_67 
+ vdd vdd vdd vss wl[208] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_0 
+ vdd vdd vss vdd vpb vnb wl[209] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_211_1 
+ rbl rbr vss vdd vpb vnb wl[209] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_211_2 
+ bl[0] br[0] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_3 
+ bl[1] br[1] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_4 
+ bl[2] br[2] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_5 
+ bl[3] br[3] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_6 
+ bl[4] br[4] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_7 
+ bl[5] br[5] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_8 
+ bl[6] br[6] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_9 
+ bl[7] br[7] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_10 
+ bl[8] br[8] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_11 
+ bl[9] br[9] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_12 
+ bl[10] br[10] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_13 
+ bl[11] br[11] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_14 
+ bl[12] br[12] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_15 
+ bl[13] br[13] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_16 
+ bl[14] br[14] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_17 
+ bl[15] br[15] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_18 
+ bl[16] br[16] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_19 
+ bl[17] br[17] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_20 
+ bl[18] br[18] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_21 
+ bl[19] br[19] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_22 
+ bl[20] br[20] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_23 
+ bl[21] br[21] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_24 
+ bl[22] br[22] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_25 
+ bl[23] br[23] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_26 
+ bl[24] br[24] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_27 
+ bl[25] br[25] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_28 
+ bl[26] br[26] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_29 
+ bl[27] br[27] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_30 
+ bl[28] br[28] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_31 
+ bl[29] br[29] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_32 
+ bl[30] br[30] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_33 
+ bl[31] br[31] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_34 
+ bl[32] br[32] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_35 
+ bl[33] br[33] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_36 
+ bl[34] br[34] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_37 
+ bl[35] br[35] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_38 
+ bl[36] br[36] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_39 
+ bl[37] br[37] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_40 
+ bl[38] br[38] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_41 
+ bl[39] br[39] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_42 
+ bl[40] br[40] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_43 
+ bl[41] br[41] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_44 
+ bl[42] br[42] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_45 
+ bl[43] br[43] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_46 
+ bl[44] br[44] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_47 
+ bl[45] br[45] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_48 
+ bl[46] br[46] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_49 
+ bl[47] br[47] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_50 
+ bl[48] br[48] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_51 
+ bl[49] br[49] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_52 
+ bl[50] br[50] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_53 
+ bl[51] br[51] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_54 
+ bl[52] br[52] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_55 
+ bl[53] br[53] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_56 
+ bl[54] br[54] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_57 
+ bl[55] br[55] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_58 
+ bl[56] br[56] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_59 
+ bl[57] br[57] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_60 
+ bl[58] br[58] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_61 
+ bl[59] br[59] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_62 
+ bl[60] br[60] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_63 
+ bl[61] br[61] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_64 
+ bl[62] br[62] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_65 
+ bl[63] br[63] vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_66 
+ vdd vdd vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_211_67 
+ vdd vdd vdd vss wl[209] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_0 
+ vdd vdd vss vdd vpb vnb wl[210] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_212_1 
+ rbl rbr vss vdd vpb vnb wl[210] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_212_2 
+ bl[0] br[0] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_3 
+ bl[1] br[1] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_4 
+ bl[2] br[2] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_5 
+ bl[3] br[3] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_6 
+ bl[4] br[4] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_7 
+ bl[5] br[5] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_8 
+ bl[6] br[6] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_9 
+ bl[7] br[7] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_10 
+ bl[8] br[8] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_11 
+ bl[9] br[9] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_12 
+ bl[10] br[10] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_13 
+ bl[11] br[11] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_14 
+ bl[12] br[12] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_15 
+ bl[13] br[13] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_16 
+ bl[14] br[14] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_17 
+ bl[15] br[15] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_18 
+ bl[16] br[16] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_19 
+ bl[17] br[17] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_20 
+ bl[18] br[18] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_21 
+ bl[19] br[19] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_22 
+ bl[20] br[20] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_23 
+ bl[21] br[21] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_24 
+ bl[22] br[22] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_25 
+ bl[23] br[23] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_26 
+ bl[24] br[24] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_27 
+ bl[25] br[25] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_28 
+ bl[26] br[26] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_29 
+ bl[27] br[27] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_30 
+ bl[28] br[28] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_31 
+ bl[29] br[29] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_32 
+ bl[30] br[30] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_33 
+ bl[31] br[31] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_34 
+ bl[32] br[32] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_35 
+ bl[33] br[33] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_36 
+ bl[34] br[34] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_37 
+ bl[35] br[35] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_38 
+ bl[36] br[36] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_39 
+ bl[37] br[37] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_40 
+ bl[38] br[38] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_41 
+ bl[39] br[39] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_42 
+ bl[40] br[40] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_43 
+ bl[41] br[41] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_44 
+ bl[42] br[42] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_45 
+ bl[43] br[43] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_46 
+ bl[44] br[44] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_47 
+ bl[45] br[45] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_48 
+ bl[46] br[46] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_49 
+ bl[47] br[47] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_50 
+ bl[48] br[48] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_51 
+ bl[49] br[49] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_52 
+ bl[50] br[50] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_53 
+ bl[51] br[51] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_54 
+ bl[52] br[52] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_55 
+ bl[53] br[53] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_56 
+ bl[54] br[54] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_57 
+ bl[55] br[55] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_58 
+ bl[56] br[56] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_59 
+ bl[57] br[57] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_60 
+ bl[58] br[58] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_61 
+ bl[59] br[59] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_62 
+ bl[60] br[60] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_63 
+ bl[61] br[61] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_64 
+ bl[62] br[62] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_65 
+ bl[63] br[63] vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_66 
+ vdd vdd vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_212_67 
+ vdd vdd vdd vss wl[210] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_0 
+ vdd vdd vss vdd vpb vnb wl[211] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_213_1 
+ rbl rbr vss vdd vpb vnb wl[211] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_213_2 
+ bl[0] br[0] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_3 
+ bl[1] br[1] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_4 
+ bl[2] br[2] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_5 
+ bl[3] br[3] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_6 
+ bl[4] br[4] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_7 
+ bl[5] br[5] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_8 
+ bl[6] br[6] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_9 
+ bl[7] br[7] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_10 
+ bl[8] br[8] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_11 
+ bl[9] br[9] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_12 
+ bl[10] br[10] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_13 
+ bl[11] br[11] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_14 
+ bl[12] br[12] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_15 
+ bl[13] br[13] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_16 
+ bl[14] br[14] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_17 
+ bl[15] br[15] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_18 
+ bl[16] br[16] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_19 
+ bl[17] br[17] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_20 
+ bl[18] br[18] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_21 
+ bl[19] br[19] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_22 
+ bl[20] br[20] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_23 
+ bl[21] br[21] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_24 
+ bl[22] br[22] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_25 
+ bl[23] br[23] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_26 
+ bl[24] br[24] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_27 
+ bl[25] br[25] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_28 
+ bl[26] br[26] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_29 
+ bl[27] br[27] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_30 
+ bl[28] br[28] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_31 
+ bl[29] br[29] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_32 
+ bl[30] br[30] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_33 
+ bl[31] br[31] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_34 
+ bl[32] br[32] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_35 
+ bl[33] br[33] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_36 
+ bl[34] br[34] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_37 
+ bl[35] br[35] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_38 
+ bl[36] br[36] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_39 
+ bl[37] br[37] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_40 
+ bl[38] br[38] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_41 
+ bl[39] br[39] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_42 
+ bl[40] br[40] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_43 
+ bl[41] br[41] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_44 
+ bl[42] br[42] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_45 
+ bl[43] br[43] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_46 
+ bl[44] br[44] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_47 
+ bl[45] br[45] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_48 
+ bl[46] br[46] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_49 
+ bl[47] br[47] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_50 
+ bl[48] br[48] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_51 
+ bl[49] br[49] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_52 
+ bl[50] br[50] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_53 
+ bl[51] br[51] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_54 
+ bl[52] br[52] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_55 
+ bl[53] br[53] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_56 
+ bl[54] br[54] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_57 
+ bl[55] br[55] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_58 
+ bl[56] br[56] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_59 
+ bl[57] br[57] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_60 
+ bl[58] br[58] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_61 
+ bl[59] br[59] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_62 
+ bl[60] br[60] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_63 
+ bl[61] br[61] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_64 
+ bl[62] br[62] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_65 
+ bl[63] br[63] vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_66 
+ vdd vdd vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_213_67 
+ vdd vdd vdd vss wl[211] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_0 
+ vdd vdd vss vdd vpb vnb wl[212] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_214_1 
+ rbl rbr vss vdd vpb vnb wl[212] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_214_2 
+ bl[0] br[0] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_3 
+ bl[1] br[1] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_4 
+ bl[2] br[2] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_5 
+ bl[3] br[3] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_6 
+ bl[4] br[4] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_7 
+ bl[5] br[5] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_8 
+ bl[6] br[6] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_9 
+ bl[7] br[7] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_10 
+ bl[8] br[8] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_11 
+ bl[9] br[9] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_12 
+ bl[10] br[10] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_13 
+ bl[11] br[11] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_14 
+ bl[12] br[12] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_15 
+ bl[13] br[13] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_16 
+ bl[14] br[14] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_17 
+ bl[15] br[15] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_18 
+ bl[16] br[16] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_19 
+ bl[17] br[17] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_20 
+ bl[18] br[18] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_21 
+ bl[19] br[19] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_22 
+ bl[20] br[20] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_23 
+ bl[21] br[21] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_24 
+ bl[22] br[22] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_25 
+ bl[23] br[23] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_26 
+ bl[24] br[24] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_27 
+ bl[25] br[25] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_28 
+ bl[26] br[26] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_29 
+ bl[27] br[27] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_30 
+ bl[28] br[28] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_31 
+ bl[29] br[29] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_32 
+ bl[30] br[30] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_33 
+ bl[31] br[31] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_34 
+ bl[32] br[32] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_35 
+ bl[33] br[33] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_36 
+ bl[34] br[34] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_37 
+ bl[35] br[35] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_38 
+ bl[36] br[36] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_39 
+ bl[37] br[37] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_40 
+ bl[38] br[38] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_41 
+ bl[39] br[39] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_42 
+ bl[40] br[40] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_43 
+ bl[41] br[41] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_44 
+ bl[42] br[42] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_45 
+ bl[43] br[43] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_46 
+ bl[44] br[44] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_47 
+ bl[45] br[45] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_48 
+ bl[46] br[46] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_49 
+ bl[47] br[47] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_50 
+ bl[48] br[48] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_51 
+ bl[49] br[49] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_52 
+ bl[50] br[50] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_53 
+ bl[51] br[51] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_54 
+ bl[52] br[52] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_55 
+ bl[53] br[53] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_56 
+ bl[54] br[54] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_57 
+ bl[55] br[55] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_58 
+ bl[56] br[56] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_59 
+ bl[57] br[57] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_60 
+ bl[58] br[58] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_61 
+ bl[59] br[59] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_62 
+ bl[60] br[60] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_63 
+ bl[61] br[61] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_64 
+ bl[62] br[62] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_65 
+ bl[63] br[63] vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_66 
+ vdd vdd vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_214_67 
+ vdd vdd vdd vss wl[212] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_0 
+ vdd vdd vss vdd vpb vnb wl[213] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_215_1 
+ rbl rbr vss vdd vpb vnb wl[213] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_215_2 
+ bl[0] br[0] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_3 
+ bl[1] br[1] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_4 
+ bl[2] br[2] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_5 
+ bl[3] br[3] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_6 
+ bl[4] br[4] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_7 
+ bl[5] br[5] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_8 
+ bl[6] br[6] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_9 
+ bl[7] br[7] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_10 
+ bl[8] br[8] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_11 
+ bl[9] br[9] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_12 
+ bl[10] br[10] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_13 
+ bl[11] br[11] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_14 
+ bl[12] br[12] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_15 
+ bl[13] br[13] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_16 
+ bl[14] br[14] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_17 
+ bl[15] br[15] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_18 
+ bl[16] br[16] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_19 
+ bl[17] br[17] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_20 
+ bl[18] br[18] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_21 
+ bl[19] br[19] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_22 
+ bl[20] br[20] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_23 
+ bl[21] br[21] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_24 
+ bl[22] br[22] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_25 
+ bl[23] br[23] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_26 
+ bl[24] br[24] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_27 
+ bl[25] br[25] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_28 
+ bl[26] br[26] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_29 
+ bl[27] br[27] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_30 
+ bl[28] br[28] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_31 
+ bl[29] br[29] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_32 
+ bl[30] br[30] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_33 
+ bl[31] br[31] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_34 
+ bl[32] br[32] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_35 
+ bl[33] br[33] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_36 
+ bl[34] br[34] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_37 
+ bl[35] br[35] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_38 
+ bl[36] br[36] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_39 
+ bl[37] br[37] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_40 
+ bl[38] br[38] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_41 
+ bl[39] br[39] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_42 
+ bl[40] br[40] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_43 
+ bl[41] br[41] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_44 
+ bl[42] br[42] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_45 
+ bl[43] br[43] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_46 
+ bl[44] br[44] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_47 
+ bl[45] br[45] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_48 
+ bl[46] br[46] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_49 
+ bl[47] br[47] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_50 
+ bl[48] br[48] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_51 
+ bl[49] br[49] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_52 
+ bl[50] br[50] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_53 
+ bl[51] br[51] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_54 
+ bl[52] br[52] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_55 
+ bl[53] br[53] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_56 
+ bl[54] br[54] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_57 
+ bl[55] br[55] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_58 
+ bl[56] br[56] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_59 
+ bl[57] br[57] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_60 
+ bl[58] br[58] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_61 
+ bl[59] br[59] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_62 
+ bl[60] br[60] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_63 
+ bl[61] br[61] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_64 
+ bl[62] br[62] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_65 
+ bl[63] br[63] vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_66 
+ vdd vdd vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_215_67 
+ vdd vdd vdd vss wl[213] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_0 
+ vdd vdd vss vdd vpb vnb wl[214] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_216_1 
+ rbl rbr vss vdd vpb vnb wl[214] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_216_2 
+ bl[0] br[0] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_3 
+ bl[1] br[1] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_4 
+ bl[2] br[2] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_5 
+ bl[3] br[3] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_6 
+ bl[4] br[4] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_7 
+ bl[5] br[5] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_8 
+ bl[6] br[6] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_9 
+ bl[7] br[7] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_10 
+ bl[8] br[8] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_11 
+ bl[9] br[9] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_12 
+ bl[10] br[10] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_13 
+ bl[11] br[11] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_14 
+ bl[12] br[12] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_15 
+ bl[13] br[13] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_16 
+ bl[14] br[14] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_17 
+ bl[15] br[15] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_18 
+ bl[16] br[16] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_19 
+ bl[17] br[17] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_20 
+ bl[18] br[18] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_21 
+ bl[19] br[19] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_22 
+ bl[20] br[20] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_23 
+ bl[21] br[21] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_24 
+ bl[22] br[22] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_25 
+ bl[23] br[23] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_26 
+ bl[24] br[24] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_27 
+ bl[25] br[25] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_28 
+ bl[26] br[26] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_29 
+ bl[27] br[27] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_30 
+ bl[28] br[28] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_31 
+ bl[29] br[29] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_32 
+ bl[30] br[30] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_33 
+ bl[31] br[31] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_34 
+ bl[32] br[32] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_35 
+ bl[33] br[33] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_36 
+ bl[34] br[34] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_37 
+ bl[35] br[35] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_38 
+ bl[36] br[36] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_39 
+ bl[37] br[37] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_40 
+ bl[38] br[38] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_41 
+ bl[39] br[39] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_42 
+ bl[40] br[40] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_43 
+ bl[41] br[41] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_44 
+ bl[42] br[42] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_45 
+ bl[43] br[43] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_46 
+ bl[44] br[44] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_47 
+ bl[45] br[45] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_48 
+ bl[46] br[46] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_49 
+ bl[47] br[47] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_50 
+ bl[48] br[48] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_51 
+ bl[49] br[49] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_52 
+ bl[50] br[50] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_53 
+ bl[51] br[51] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_54 
+ bl[52] br[52] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_55 
+ bl[53] br[53] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_56 
+ bl[54] br[54] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_57 
+ bl[55] br[55] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_58 
+ bl[56] br[56] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_59 
+ bl[57] br[57] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_60 
+ bl[58] br[58] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_61 
+ bl[59] br[59] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_62 
+ bl[60] br[60] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_63 
+ bl[61] br[61] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_64 
+ bl[62] br[62] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_65 
+ bl[63] br[63] vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_66 
+ vdd vdd vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_216_67 
+ vdd vdd vdd vss wl[214] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_0 
+ vdd vdd vss vdd vpb vnb wl[215] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_217_1 
+ rbl rbr vss vdd vpb vnb wl[215] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_217_2 
+ bl[0] br[0] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_3 
+ bl[1] br[1] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_4 
+ bl[2] br[2] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_5 
+ bl[3] br[3] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_6 
+ bl[4] br[4] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_7 
+ bl[5] br[5] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_8 
+ bl[6] br[6] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_9 
+ bl[7] br[7] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_10 
+ bl[8] br[8] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_11 
+ bl[9] br[9] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_12 
+ bl[10] br[10] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_13 
+ bl[11] br[11] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_14 
+ bl[12] br[12] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_15 
+ bl[13] br[13] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_16 
+ bl[14] br[14] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_17 
+ bl[15] br[15] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_18 
+ bl[16] br[16] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_19 
+ bl[17] br[17] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_20 
+ bl[18] br[18] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_21 
+ bl[19] br[19] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_22 
+ bl[20] br[20] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_23 
+ bl[21] br[21] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_24 
+ bl[22] br[22] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_25 
+ bl[23] br[23] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_26 
+ bl[24] br[24] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_27 
+ bl[25] br[25] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_28 
+ bl[26] br[26] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_29 
+ bl[27] br[27] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_30 
+ bl[28] br[28] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_31 
+ bl[29] br[29] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_32 
+ bl[30] br[30] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_33 
+ bl[31] br[31] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_34 
+ bl[32] br[32] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_35 
+ bl[33] br[33] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_36 
+ bl[34] br[34] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_37 
+ bl[35] br[35] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_38 
+ bl[36] br[36] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_39 
+ bl[37] br[37] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_40 
+ bl[38] br[38] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_41 
+ bl[39] br[39] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_42 
+ bl[40] br[40] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_43 
+ bl[41] br[41] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_44 
+ bl[42] br[42] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_45 
+ bl[43] br[43] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_46 
+ bl[44] br[44] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_47 
+ bl[45] br[45] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_48 
+ bl[46] br[46] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_49 
+ bl[47] br[47] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_50 
+ bl[48] br[48] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_51 
+ bl[49] br[49] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_52 
+ bl[50] br[50] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_53 
+ bl[51] br[51] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_54 
+ bl[52] br[52] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_55 
+ bl[53] br[53] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_56 
+ bl[54] br[54] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_57 
+ bl[55] br[55] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_58 
+ bl[56] br[56] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_59 
+ bl[57] br[57] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_60 
+ bl[58] br[58] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_61 
+ bl[59] br[59] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_62 
+ bl[60] br[60] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_63 
+ bl[61] br[61] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_64 
+ bl[62] br[62] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_65 
+ bl[63] br[63] vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_66 
+ vdd vdd vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_217_67 
+ vdd vdd vdd vss wl[215] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_0 
+ vdd vdd vss vdd vpb vnb wl[216] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_218_1 
+ rbl rbr vss vdd vpb vnb wl[216] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_218_2 
+ bl[0] br[0] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_3 
+ bl[1] br[1] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_4 
+ bl[2] br[2] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_5 
+ bl[3] br[3] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_6 
+ bl[4] br[4] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_7 
+ bl[5] br[5] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_8 
+ bl[6] br[6] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_9 
+ bl[7] br[7] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_10 
+ bl[8] br[8] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_11 
+ bl[9] br[9] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_12 
+ bl[10] br[10] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_13 
+ bl[11] br[11] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_14 
+ bl[12] br[12] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_15 
+ bl[13] br[13] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_16 
+ bl[14] br[14] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_17 
+ bl[15] br[15] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_18 
+ bl[16] br[16] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_19 
+ bl[17] br[17] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_20 
+ bl[18] br[18] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_21 
+ bl[19] br[19] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_22 
+ bl[20] br[20] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_23 
+ bl[21] br[21] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_24 
+ bl[22] br[22] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_25 
+ bl[23] br[23] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_26 
+ bl[24] br[24] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_27 
+ bl[25] br[25] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_28 
+ bl[26] br[26] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_29 
+ bl[27] br[27] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_30 
+ bl[28] br[28] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_31 
+ bl[29] br[29] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_32 
+ bl[30] br[30] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_33 
+ bl[31] br[31] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_34 
+ bl[32] br[32] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_35 
+ bl[33] br[33] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_36 
+ bl[34] br[34] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_37 
+ bl[35] br[35] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_38 
+ bl[36] br[36] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_39 
+ bl[37] br[37] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_40 
+ bl[38] br[38] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_41 
+ bl[39] br[39] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_42 
+ bl[40] br[40] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_43 
+ bl[41] br[41] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_44 
+ bl[42] br[42] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_45 
+ bl[43] br[43] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_46 
+ bl[44] br[44] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_47 
+ bl[45] br[45] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_48 
+ bl[46] br[46] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_49 
+ bl[47] br[47] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_50 
+ bl[48] br[48] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_51 
+ bl[49] br[49] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_52 
+ bl[50] br[50] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_53 
+ bl[51] br[51] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_54 
+ bl[52] br[52] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_55 
+ bl[53] br[53] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_56 
+ bl[54] br[54] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_57 
+ bl[55] br[55] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_58 
+ bl[56] br[56] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_59 
+ bl[57] br[57] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_60 
+ bl[58] br[58] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_61 
+ bl[59] br[59] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_62 
+ bl[60] br[60] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_63 
+ bl[61] br[61] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_64 
+ bl[62] br[62] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_65 
+ bl[63] br[63] vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_66 
+ vdd vdd vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_218_67 
+ vdd vdd vdd vss wl[216] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_0 
+ vdd vdd vss vdd vpb vnb wl[217] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_219_1 
+ rbl rbr vss vdd vpb vnb wl[217] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_219_2 
+ bl[0] br[0] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_3 
+ bl[1] br[1] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_4 
+ bl[2] br[2] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_5 
+ bl[3] br[3] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_6 
+ bl[4] br[4] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_7 
+ bl[5] br[5] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_8 
+ bl[6] br[6] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_9 
+ bl[7] br[7] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_10 
+ bl[8] br[8] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_11 
+ bl[9] br[9] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_12 
+ bl[10] br[10] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_13 
+ bl[11] br[11] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_14 
+ bl[12] br[12] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_15 
+ bl[13] br[13] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_16 
+ bl[14] br[14] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_17 
+ bl[15] br[15] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_18 
+ bl[16] br[16] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_19 
+ bl[17] br[17] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_20 
+ bl[18] br[18] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_21 
+ bl[19] br[19] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_22 
+ bl[20] br[20] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_23 
+ bl[21] br[21] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_24 
+ bl[22] br[22] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_25 
+ bl[23] br[23] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_26 
+ bl[24] br[24] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_27 
+ bl[25] br[25] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_28 
+ bl[26] br[26] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_29 
+ bl[27] br[27] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_30 
+ bl[28] br[28] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_31 
+ bl[29] br[29] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_32 
+ bl[30] br[30] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_33 
+ bl[31] br[31] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_34 
+ bl[32] br[32] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_35 
+ bl[33] br[33] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_36 
+ bl[34] br[34] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_37 
+ bl[35] br[35] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_38 
+ bl[36] br[36] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_39 
+ bl[37] br[37] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_40 
+ bl[38] br[38] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_41 
+ bl[39] br[39] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_42 
+ bl[40] br[40] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_43 
+ bl[41] br[41] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_44 
+ bl[42] br[42] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_45 
+ bl[43] br[43] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_46 
+ bl[44] br[44] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_47 
+ bl[45] br[45] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_48 
+ bl[46] br[46] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_49 
+ bl[47] br[47] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_50 
+ bl[48] br[48] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_51 
+ bl[49] br[49] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_52 
+ bl[50] br[50] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_53 
+ bl[51] br[51] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_54 
+ bl[52] br[52] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_55 
+ bl[53] br[53] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_56 
+ bl[54] br[54] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_57 
+ bl[55] br[55] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_58 
+ bl[56] br[56] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_59 
+ bl[57] br[57] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_60 
+ bl[58] br[58] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_61 
+ bl[59] br[59] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_62 
+ bl[60] br[60] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_63 
+ bl[61] br[61] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_64 
+ bl[62] br[62] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_65 
+ bl[63] br[63] vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_66 
+ vdd vdd vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_219_67 
+ vdd vdd vdd vss wl[217] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_0 
+ vdd vdd vss vdd vpb vnb wl[218] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_220_1 
+ rbl rbr vss vdd vpb vnb wl[218] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_220_2 
+ bl[0] br[0] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_3 
+ bl[1] br[1] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_4 
+ bl[2] br[2] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_5 
+ bl[3] br[3] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_6 
+ bl[4] br[4] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_7 
+ bl[5] br[5] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_8 
+ bl[6] br[6] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_9 
+ bl[7] br[7] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_10 
+ bl[8] br[8] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_11 
+ bl[9] br[9] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_12 
+ bl[10] br[10] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_13 
+ bl[11] br[11] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_14 
+ bl[12] br[12] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_15 
+ bl[13] br[13] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_16 
+ bl[14] br[14] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_17 
+ bl[15] br[15] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_18 
+ bl[16] br[16] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_19 
+ bl[17] br[17] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_20 
+ bl[18] br[18] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_21 
+ bl[19] br[19] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_22 
+ bl[20] br[20] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_23 
+ bl[21] br[21] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_24 
+ bl[22] br[22] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_25 
+ bl[23] br[23] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_26 
+ bl[24] br[24] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_27 
+ bl[25] br[25] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_28 
+ bl[26] br[26] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_29 
+ bl[27] br[27] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_30 
+ bl[28] br[28] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_31 
+ bl[29] br[29] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_32 
+ bl[30] br[30] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_33 
+ bl[31] br[31] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_34 
+ bl[32] br[32] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_35 
+ bl[33] br[33] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_36 
+ bl[34] br[34] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_37 
+ bl[35] br[35] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_38 
+ bl[36] br[36] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_39 
+ bl[37] br[37] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_40 
+ bl[38] br[38] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_41 
+ bl[39] br[39] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_42 
+ bl[40] br[40] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_43 
+ bl[41] br[41] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_44 
+ bl[42] br[42] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_45 
+ bl[43] br[43] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_46 
+ bl[44] br[44] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_47 
+ bl[45] br[45] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_48 
+ bl[46] br[46] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_49 
+ bl[47] br[47] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_50 
+ bl[48] br[48] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_51 
+ bl[49] br[49] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_52 
+ bl[50] br[50] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_53 
+ bl[51] br[51] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_54 
+ bl[52] br[52] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_55 
+ bl[53] br[53] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_56 
+ bl[54] br[54] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_57 
+ bl[55] br[55] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_58 
+ bl[56] br[56] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_59 
+ bl[57] br[57] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_60 
+ bl[58] br[58] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_61 
+ bl[59] br[59] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_62 
+ bl[60] br[60] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_63 
+ bl[61] br[61] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_64 
+ bl[62] br[62] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_65 
+ bl[63] br[63] vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_66 
+ vdd vdd vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_220_67 
+ vdd vdd vdd vss wl[218] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_0 
+ vdd vdd vss vdd vpb vnb wl[219] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_221_1 
+ rbl rbr vss vdd vpb vnb wl[219] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_221_2 
+ bl[0] br[0] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_3 
+ bl[1] br[1] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_4 
+ bl[2] br[2] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_5 
+ bl[3] br[3] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_6 
+ bl[4] br[4] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_7 
+ bl[5] br[5] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_8 
+ bl[6] br[6] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_9 
+ bl[7] br[7] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_10 
+ bl[8] br[8] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_11 
+ bl[9] br[9] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_12 
+ bl[10] br[10] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_13 
+ bl[11] br[11] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_14 
+ bl[12] br[12] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_15 
+ bl[13] br[13] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_16 
+ bl[14] br[14] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_17 
+ bl[15] br[15] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_18 
+ bl[16] br[16] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_19 
+ bl[17] br[17] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_20 
+ bl[18] br[18] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_21 
+ bl[19] br[19] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_22 
+ bl[20] br[20] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_23 
+ bl[21] br[21] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_24 
+ bl[22] br[22] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_25 
+ bl[23] br[23] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_26 
+ bl[24] br[24] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_27 
+ bl[25] br[25] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_28 
+ bl[26] br[26] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_29 
+ bl[27] br[27] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_30 
+ bl[28] br[28] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_31 
+ bl[29] br[29] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_32 
+ bl[30] br[30] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_33 
+ bl[31] br[31] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_34 
+ bl[32] br[32] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_35 
+ bl[33] br[33] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_36 
+ bl[34] br[34] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_37 
+ bl[35] br[35] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_38 
+ bl[36] br[36] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_39 
+ bl[37] br[37] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_40 
+ bl[38] br[38] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_41 
+ bl[39] br[39] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_42 
+ bl[40] br[40] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_43 
+ bl[41] br[41] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_44 
+ bl[42] br[42] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_45 
+ bl[43] br[43] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_46 
+ bl[44] br[44] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_47 
+ bl[45] br[45] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_48 
+ bl[46] br[46] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_49 
+ bl[47] br[47] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_50 
+ bl[48] br[48] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_51 
+ bl[49] br[49] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_52 
+ bl[50] br[50] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_53 
+ bl[51] br[51] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_54 
+ bl[52] br[52] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_55 
+ bl[53] br[53] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_56 
+ bl[54] br[54] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_57 
+ bl[55] br[55] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_58 
+ bl[56] br[56] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_59 
+ bl[57] br[57] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_60 
+ bl[58] br[58] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_61 
+ bl[59] br[59] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_62 
+ bl[60] br[60] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_63 
+ bl[61] br[61] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_64 
+ bl[62] br[62] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_65 
+ bl[63] br[63] vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_66 
+ vdd vdd vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_221_67 
+ vdd vdd vdd vss wl[219] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_0 
+ vdd vdd vss vdd vpb vnb wl[220] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_222_1 
+ rbl rbr vss vdd vpb vnb wl[220] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_222_2 
+ bl[0] br[0] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_3 
+ bl[1] br[1] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_4 
+ bl[2] br[2] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_5 
+ bl[3] br[3] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_6 
+ bl[4] br[4] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_7 
+ bl[5] br[5] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_8 
+ bl[6] br[6] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_9 
+ bl[7] br[7] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_10 
+ bl[8] br[8] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_11 
+ bl[9] br[9] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_12 
+ bl[10] br[10] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_13 
+ bl[11] br[11] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_14 
+ bl[12] br[12] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_15 
+ bl[13] br[13] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_16 
+ bl[14] br[14] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_17 
+ bl[15] br[15] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_18 
+ bl[16] br[16] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_19 
+ bl[17] br[17] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_20 
+ bl[18] br[18] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_21 
+ bl[19] br[19] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_22 
+ bl[20] br[20] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_23 
+ bl[21] br[21] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_24 
+ bl[22] br[22] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_25 
+ bl[23] br[23] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_26 
+ bl[24] br[24] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_27 
+ bl[25] br[25] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_28 
+ bl[26] br[26] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_29 
+ bl[27] br[27] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_30 
+ bl[28] br[28] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_31 
+ bl[29] br[29] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_32 
+ bl[30] br[30] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_33 
+ bl[31] br[31] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_34 
+ bl[32] br[32] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_35 
+ bl[33] br[33] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_36 
+ bl[34] br[34] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_37 
+ bl[35] br[35] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_38 
+ bl[36] br[36] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_39 
+ bl[37] br[37] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_40 
+ bl[38] br[38] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_41 
+ bl[39] br[39] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_42 
+ bl[40] br[40] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_43 
+ bl[41] br[41] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_44 
+ bl[42] br[42] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_45 
+ bl[43] br[43] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_46 
+ bl[44] br[44] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_47 
+ bl[45] br[45] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_48 
+ bl[46] br[46] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_49 
+ bl[47] br[47] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_50 
+ bl[48] br[48] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_51 
+ bl[49] br[49] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_52 
+ bl[50] br[50] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_53 
+ bl[51] br[51] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_54 
+ bl[52] br[52] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_55 
+ bl[53] br[53] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_56 
+ bl[54] br[54] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_57 
+ bl[55] br[55] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_58 
+ bl[56] br[56] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_59 
+ bl[57] br[57] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_60 
+ bl[58] br[58] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_61 
+ bl[59] br[59] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_62 
+ bl[60] br[60] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_63 
+ bl[61] br[61] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_64 
+ bl[62] br[62] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_65 
+ bl[63] br[63] vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_66 
+ vdd vdd vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_222_67 
+ vdd vdd vdd vss wl[220] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_0 
+ vdd vdd vss vdd vpb vnb wl[221] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_223_1 
+ rbl rbr vss vdd vpb vnb wl[221] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_223_2 
+ bl[0] br[0] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_3 
+ bl[1] br[1] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_4 
+ bl[2] br[2] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_5 
+ bl[3] br[3] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_6 
+ bl[4] br[4] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_7 
+ bl[5] br[5] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_8 
+ bl[6] br[6] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_9 
+ bl[7] br[7] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_10 
+ bl[8] br[8] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_11 
+ bl[9] br[9] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_12 
+ bl[10] br[10] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_13 
+ bl[11] br[11] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_14 
+ bl[12] br[12] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_15 
+ bl[13] br[13] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_16 
+ bl[14] br[14] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_17 
+ bl[15] br[15] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_18 
+ bl[16] br[16] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_19 
+ bl[17] br[17] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_20 
+ bl[18] br[18] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_21 
+ bl[19] br[19] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_22 
+ bl[20] br[20] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_23 
+ bl[21] br[21] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_24 
+ bl[22] br[22] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_25 
+ bl[23] br[23] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_26 
+ bl[24] br[24] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_27 
+ bl[25] br[25] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_28 
+ bl[26] br[26] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_29 
+ bl[27] br[27] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_30 
+ bl[28] br[28] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_31 
+ bl[29] br[29] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_32 
+ bl[30] br[30] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_33 
+ bl[31] br[31] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_34 
+ bl[32] br[32] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_35 
+ bl[33] br[33] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_36 
+ bl[34] br[34] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_37 
+ bl[35] br[35] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_38 
+ bl[36] br[36] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_39 
+ bl[37] br[37] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_40 
+ bl[38] br[38] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_41 
+ bl[39] br[39] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_42 
+ bl[40] br[40] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_43 
+ bl[41] br[41] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_44 
+ bl[42] br[42] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_45 
+ bl[43] br[43] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_46 
+ bl[44] br[44] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_47 
+ bl[45] br[45] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_48 
+ bl[46] br[46] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_49 
+ bl[47] br[47] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_50 
+ bl[48] br[48] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_51 
+ bl[49] br[49] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_52 
+ bl[50] br[50] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_53 
+ bl[51] br[51] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_54 
+ bl[52] br[52] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_55 
+ bl[53] br[53] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_56 
+ bl[54] br[54] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_57 
+ bl[55] br[55] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_58 
+ bl[56] br[56] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_59 
+ bl[57] br[57] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_60 
+ bl[58] br[58] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_61 
+ bl[59] br[59] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_62 
+ bl[60] br[60] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_63 
+ bl[61] br[61] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_64 
+ bl[62] br[62] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_65 
+ bl[63] br[63] vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_66 
+ vdd vdd vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_223_67 
+ vdd vdd vdd vss wl[221] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_0 
+ vdd vdd vss vdd vpb vnb wl[222] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_224_1 
+ rbl rbr vss vdd vpb vnb wl[222] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_224_2 
+ bl[0] br[0] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_3 
+ bl[1] br[1] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_4 
+ bl[2] br[2] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_5 
+ bl[3] br[3] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_6 
+ bl[4] br[4] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_7 
+ bl[5] br[5] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_8 
+ bl[6] br[6] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_9 
+ bl[7] br[7] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_10 
+ bl[8] br[8] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_11 
+ bl[9] br[9] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_12 
+ bl[10] br[10] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_13 
+ bl[11] br[11] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_14 
+ bl[12] br[12] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_15 
+ bl[13] br[13] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_16 
+ bl[14] br[14] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_17 
+ bl[15] br[15] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_18 
+ bl[16] br[16] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_19 
+ bl[17] br[17] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_20 
+ bl[18] br[18] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_21 
+ bl[19] br[19] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_22 
+ bl[20] br[20] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_23 
+ bl[21] br[21] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_24 
+ bl[22] br[22] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_25 
+ bl[23] br[23] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_26 
+ bl[24] br[24] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_27 
+ bl[25] br[25] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_28 
+ bl[26] br[26] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_29 
+ bl[27] br[27] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_30 
+ bl[28] br[28] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_31 
+ bl[29] br[29] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_32 
+ bl[30] br[30] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_33 
+ bl[31] br[31] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_34 
+ bl[32] br[32] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_35 
+ bl[33] br[33] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_36 
+ bl[34] br[34] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_37 
+ bl[35] br[35] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_38 
+ bl[36] br[36] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_39 
+ bl[37] br[37] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_40 
+ bl[38] br[38] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_41 
+ bl[39] br[39] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_42 
+ bl[40] br[40] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_43 
+ bl[41] br[41] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_44 
+ bl[42] br[42] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_45 
+ bl[43] br[43] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_46 
+ bl[44] br[44] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_47 
+ bl[45] br[45] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_48 
+ bl[46] br[46] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_49 
+ bl[47] br[47] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_50 
+ bl[48] br[48] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_51 
+ bl[49] br[49] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_52 
+ bl[50] br[50] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_53 
+ bl[51] br[51] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_54 
+ bl[52] br[52] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_55 
+ bl[53] br[53] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_56 
+ bl[54] br[54] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_57 
+ bl[55] br[55] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_58 
+ bl[56] br[56] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_59 
+ bl[57] br[57] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_60 
+ bl[58] br[58] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_61 
+ bl[59] br[59] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_62 
+ bl[60] br[60] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_63 
+ bl[61] br[61] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_64 
+ bl[62] br[62] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_65 
+ bl[63] br[63] vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_66 
+ vdd vdd vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_224_67 
+ vdd vdd vdd vss wl[222] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_0 
+ vdd vdd vss vdd vpb vnb wl[223] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_225_1 
+ rbl rbr vss vdd vpb vnb wl[223] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_225_2 
+ bl[0] br[0] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_3 
+ bl[1] br[1] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_4 
+ bl[2] br[2] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_5 
+ bl[3] br[3] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_6 
+ bl[4] br[4] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_7 
+ bl[5] br[5] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_8 
+ bl[6] br[6] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_9 
+ bl[7] br[7] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_10 
+ bl[8] br[8] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_11 
+ bl[9] br[9] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_12 
+ bl[10] br[10] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_13 
+ bl[11] br[11] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_14 
+ bl[12] br[12] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_15 
+ bl[13] br[13] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_16 
+ bl[14] br[14] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_17 
+ bl[15] br[15] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_18 
+ bl[16] br[16] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_19 
+ bl[17] br[17] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_20 
+ bl[18] br[18] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_21 
+ bl[19] br[19] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_22 
+ bl[20] br[20] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_23 
+ bl[21] br[21] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_24 
+ bl[22] br[22] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_25 
+ bl[23] br[23] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_26 
+ bl[24] br[24] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_27 
+ bl[25] br[25] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_28 
+ bl[26] br[26] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_29 
+ bl[27] br[27] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_30 
+ bl[28] br[28] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_31 
+ bl[29] br[29] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_32 
+ bl[30] br[30] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_33 
+ bl[31] br[31] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_34 
+ bl[32] br[32] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_35 
+ bl[33] br[33] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_36 
+ bl[34] br[34] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_37 
+ bl[35] br[35] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_38 
+ bl[36] br[36] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_39 
+ bl[37] br[37] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_40 
+ bl[38] br[38] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_41 
+ bl[39] br[39] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_42 
+ bl[40] br[40] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_43 
+ bl[41] br[41] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_44 
+ bl[42] br[42] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_45 
+ bl[43] br[43] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_46 
+ bl[44] br[44] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_47 
+ bl[45] br[45] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_48 
+ bl[46] br[46] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_49 
+ bl[47] br[47] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_50 
+ bl[48] br[48] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_51 
+ bl[49] br[49] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_52 
+ bl[50] br[50] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_53 
+ bl[51] br[51] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_54 
+ bl[52] br[52] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_55 
+ bl[53] br[53] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_56 
+ bl[54] br[54] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_57 
+ bl[55] br[55] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_58 
+ bl[56] br[56] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_59 
+ bl[57] br[57] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_60 
+ bl[58] br[58] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_61 
+ bl[59] br[59] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_62 
+ bl[60] br[60] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_63 
+ bl[61] br[61] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_64 
+ bl[62] br[62] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_65 
+ bl[63] br[63] vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_66 
+ vdd vdd vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_225_67 
+ vdd vdd vdd vss wl[223] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_0 
+ vdd vdd vss vdd vpb vnb wl[224] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_226_1 
+ rbl rbr vss vdd vpb vnb wl[224] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_226_2 
+ bl[0] br[0] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_3 
+ bl[1] br[1] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_4 
+ bl[2] br[2] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_5 
+ bl[3] br[3] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_6 
+ bl[4] br[4] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_7 
+ bl[5] br[5] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_8 
+ bl[6] br[6] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_9 
+ bl[7] br[7] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_10 
+ bl[8] br[8] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_11 
+ bl[9] br[9] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_12 
+ bl[10] br[10] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_13 
+ bl[11] br[11] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_14 
+ bl[12] br[12] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_15 
+ bl[13] br[13] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_16 
+ bl[14] br[14] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_17 
+ bl[15] br[15] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_18 
+ bl[16] br[16] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_19 
+ bl[17] br[17] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_20 
+ bl[18] br[18] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_21 
+ bl[19] br[19] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_22 
+ bl[20] br[20] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_23 
+ bl[21] br[21] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_24 
+ bl[22] br[22] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_25 
+ bl[23] br[23] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_26 
+ bl[24] br[24] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_27 
+ bl[25] br[25] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_28 
+ bl[26] br[26] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_29 
+ bl[27] br[27] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_30 
+ bl[28] br[28] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_31 
+ bl[29] br[29] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_32 
+ bl[30] br[30] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_33 
+ bl[31] br[31] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_34 
+ bl[32] br[32] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_35 
+ bl[33] br[33] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_36 
+ bl[34] br[34] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_37 
+ bl[35] br[35] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_38 
+ bl[36] br[36] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_39 
+ bl[37] br[37] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_40 
+ bl[38] br[38] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_41 
+ bl[39] br[39] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_42 
+ bl[40] br[40] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_43 
+ bl[41] br[41] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_44 
+ bl[42] br[42] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_45 
+ bl[43] br[43] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_46 
+ bl[44] br[44] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_47 
+ bl[45] br[45] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_48 
+ bl[46] br[46] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_49 
+ bl[47] br[47] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_50 
+ bl[48] br[48] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_51 
+ bl[49] br[49] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_52 
+ bl[50] br[50] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_53 
+ bl[51] br[51] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_54 
+ bl[52] br[52] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_55 
+ bl[53] br[53] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_56 
+ bl[54] br[54] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_57 
+ bl[55] br[55] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_58 
+ bl[56] br[56] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_59 
+ bl[57] br[57] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_60 
+ bl[58] br[58] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_61 
+ bl[59] br[59] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_62 
+ bl[60] br[60] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_63 
+ bl[61] br[61] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_64 
+ bl[62] br[62] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_65 
+ bl[63] br[63] vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_66 
+ vdd vdd vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_226_67 
+ vdd vdd vdd vss wl[224] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_0 
+ vdd vdd vss vdd vpb vnb wl[225] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_227_1 
+ rbl rbr vss vdd vpb vnb wl[225] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_227_2 
+ bl[0] br[0] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_3 
+ bl[1] br[1] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_4 
+ bl[2] br[2] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_5 
+ bl[3] br[3] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_6 
+ bl[4] br[4] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_7 
+ bl[5] br[5] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_8 
+ bl[6] br[6] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_9 
+ bl[7] br[7] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_10 
+ bl[8] br[8] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_11 
+ bl[9] br[9] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_12 
+ bl[10] br[10] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_13 
+ bl[11] br[11] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_14 
+ bl[12] br[12] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_15 
+ bl[13] br[13] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_16 
+ bl[14] br[14] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_17 
+ bl[15] br[15] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_18 
+ bl[16] br[16] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_19 
+ bl[17] br[17] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_20 
+ bl[18] br[18] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_21 
+ bl[19] br[19] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_22 
+ bl[20] br[20] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_23 
+ bl[21] br[21] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_24 
+ bl[22] br[22] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_25 
+ bl[23] br[23] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_26 
+ bl[24] br[24] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_27 
+ bl[25] br[25] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_28 
+ bl[26] br[26] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_29 
+ bl[27] br[27] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_30 
+ bl[28] br[28] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_31 
+ bl[29] br[29] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_32 
+ bl[30] br[30] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_33 
+ bl[31] br[31] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_34 
+ bl[32] br[32] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_35 
+ bl[33] br[33] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_36 
+ bl[34] br[34] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_37 
+ bl[35] br[35] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_38 
+ bl[36] br[36] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_39 
+ bl[37] br[37] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_40 
+ bl[38] br[38] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_41 
+ bl[39] br[39] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_42 
+ bl[40] br[40] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_43 
+ bl[41] br[41] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_44 
+ bl[42] br[42] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_45 
+ bl[43] br[43] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_46 
+ bl[44] br[44] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_47 
+ bl[45] br[45] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_48 
+ bl[46] br[46] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_49 
+ bl[47] br[47] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_50 
+ bl[48] br[48] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_51 
+ bl[49] br[49] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_52 
+ bl[50] br[50] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_53 
+ bl[51] br[51] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_54 
+ bl[52] br[52] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_55 
+ bl[53] br[53] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_56 
+ bl[54] br[54] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_57 
+ bl[55] br[55] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_58 
+ bl[56] br[56] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_59 
+ bl[57] br[57] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_60 
+ bl[58] br[58] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_61 
+ bl[59] br[59] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_62 
+ bl[60] br[60] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_63 
+ bl[61] br[61] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_64 
+ bl[62] br[62] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_65 
+ bl[63] br[63] vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_66 
+ vdd vdd vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_227_67 
+ vdd vdd vdd vss wl[225] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_0 
+ vdd vdd vss vdd vpb vnb wl[226] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_228_1 
+ rbl rbr vss vdd vpb vnb wl[226] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_228_2 
+ bl[0] br[0] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_3 
+ bl[1] br[1] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_4 
+ bl[2] br[2] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_5 
+ bl[3] br[3] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_6 
+ bl[4] br[4] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_7 
+ bl[5] br[5] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_8 
+ bl[6] br[6] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_9 
+ bl[7] br[7] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_10 
+ bl[8] br[8] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_11 
+ bl[9] br[9] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_12 
+ bl[10] br[10] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_13 
+ bl[11] br[11] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_14 
+ bl[12] br[12] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_15 
+ bl[13] br[13] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_16 
+ bl[14] br[14] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_17 
+ bl[15] br[15] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_18 
+ bl[16] br[16] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_19 
+ bl[17] br[17] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_20 
+ bl[18] br[18] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_21 
+ bl[19] br[19] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_22 
+ bl[20] br[20] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_23 
+ bl[21] br[21] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_24 
+ bl[22] br[22] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_25 
+ bl[23] br[23] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_26 
+ bl[24] br[24] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_27 
+ bl[25] br[25] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_28 
+ bl[26] br[26] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_29 
+ bl[27] br[27] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_30 
+ bl[28] br[28] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_31 
+ bl[29] br[29] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_32 
+ bl[30] br[30] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_33 
+ bl[31] br[31] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_34 
+ bl[32] br[32] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_35 
+ bl[33] br[33] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_36 
+ bl[34] br[34] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_37 
+ bl[35] br[35] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_38 
+ bl[36] br[36] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_39 
+ bl[37] br[37] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_40 
+ bl[38] br[38] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_41 
+ bl[39] br[39] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_42 
+ bl[40] br[40] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_43 
+ bl[41] br[41] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_44 
+ bl[42] br[42] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_45 
+ bl[43] br[43] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_46 
+ bl[44] br[44] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_47 
+ bl[45] br[45] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_48 
+ bl[46] br[46] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_49 
+ bl[47] br[47] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_50 
+ bl[48] br[48] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_51 
+ bl[49] br[49] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_52 
+ bl[50] br[50] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_53 
+ bl[51] br[51] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_54 
+ bl[52] br[52] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_55 
+ bl[53] br[53] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_56 
+ bl[54] br[54] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_57 
+ bl[55] br[55] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_58 
+ bl[56] br[56] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_59 
+ bl[57] br[57] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_60 
+ bl[58] br[58] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_61 
+ bl[59] br[59] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_62 
+ bl[60] br[60] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_63 
+ bl[61] br[61] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_64 
+ bl[62] br[62] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_65 
+ bl[63] br[63] vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_66 
+ vdd vdd vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_228_67 
+ vdd vdd vdd vss wl[226] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_0 
+ vdd vdd vss vdd vpb vnb wl[227] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_229_1 
+ rbl rbr vss vdd vpb vnb wl[227] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_229_2 
+ bl[0] br[0] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_3 
+ bl[1] br[1] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_4 
+ bl[2] br[2] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_5 
+ bl[3] br[3] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_6 
+ bl[4] br[4] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_7 
+ bl[5] br[5] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_8 
+ bl[6] br[6] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_9 
+ bl[7] br[7] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_10 
+ bl[8] br[8] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_11 
+ bl[9] br[9] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_12 
+ bl[10] br[10] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_13 
+ bl[11] br[11] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_14 
+ bl[12] br[12] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_15 
+ bl[13] br[13] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_16 
+ bl[14] br[14] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_17 
+ bl[15] br[15] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_18 
+ bl[16] br[16] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_19 
+ bl[17] br[17] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_20 
+ bl[18] br[18] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_21 
+ bl[19] br[19] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_22 
+ bl[20] br[20] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_23 
+ bl[21] br[21] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_24 
+ bl[22] br[22] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_25 
+ bl[23] br[23] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_26 
+ bl[24] br[24] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_27 
+ bl[25] br[25] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_28 
+ bl[26] br[26] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_29 
+ bl[27] br[27] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_30 
+ bl[28] br[28] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_31 
+ bl[29] br[29] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_32 
+ bl[30] br[30] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_33 
+ bl[31] br[31] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_34 
+ bl[32] br[32] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_35 
+ bl[33] br[33] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_36 
+ bl[34] br[34] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_37 
+ bl[35] br[35] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_38 
+ bl[36] br[36] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_39 
+ bl[37] br[37] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_40 
+ bl[38] br[38] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_41 
+ bl[39] br[39] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_42 
+ bl[40] br[40] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_43 
+ bl[41] br[41] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_44 
+ bl[42] br[42] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_45 
+ bl[43] br[43] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_46 
+ bl[44] br[44] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_47 
+ bl[45] br[45] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_48 
+ bl[46] br[46] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_49 
+ bl[47] br[47] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_50 
+ bl[48] br[48] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_51 
+ bl[49] br[49] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_52 
+ bl[50] br[50] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_53 
+ bl[51] br[51] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_54 
+ bl[52] br[52] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_55 
+ bl[53] br[53] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_56 
+ bl[54] br[54] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_57 
+ bl[55] br[55] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_58 
+ bl[56] br[56] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_59 
+ bl[57] br[57] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_60 
+ bl[58] br[58] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_61 
+ bl[59] br[59] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_62 
+ bl[60] br[60] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_63 
+ bl[61] br[61] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_64 
+ bl[62] br[62] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_65 
+ bl[63] br[63] vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_66 
+ vdd vdd vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_229_67 
+ vdd vdd vdd vss wl[227] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_0 
+ vdd vdd vss vdd vpb vnb wl[228] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_230_1 
+ rbl rbr vss vdd vpb vnb wl[228] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_230_2 
+ bl[0] br[0] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_3 
+ bl[1] br[1] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_4 
+ bl[2] br[2] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_5 
+ bl[3] br[3] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_6 
+ bl[4] br[4] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_7 
+ bl[5] br[5] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_8 
+ bl[6] br[6] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_9 
+ bl[7] br[7] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_10 
+ bl[8] br[8] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_11 
+ bl[9] br[9] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_12 
+ bl[10] br[10] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_13 
+ bl[11] br[11] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_14 
+ bl[12] br[12] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_15 
+ bl[13] br[13] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_16 
+ bl[14] br[14] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_17 
+ bl[15] br[15] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_18 
+ bl[16] br[16] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_19 
+ bl[17] br[17] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_20 
+ bl[18] br[18] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_21 
+ bl[19] br[19] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_22 
+ bl[20] br[20] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_23 
+ bl[21] br[21] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_24 
+ bl[22] br[22] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_25 
+ bl[23] br[23] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_26 
+ bl[24] br[24] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_27 
+ bl[25] br[25] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_28 
+ bl[26] br[26] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_29 
+ bl[27] br[27] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_30 
+ bl[28] br[28] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_31 
+ bl[29] br[29] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_32 
+ bl[30] br[30] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_33 
+ bl[31] br[31] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_34 
+ bl[32] br[32] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_35 
+ bl[33] br[33] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_36 
+ bl[34] br[34] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_37 
+ bl[35] br[35] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_38 
+ bl[36] br[36] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_39 
+ bl[37] br[37] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_40 
+ bl[38] br[38] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_41 
+ bl[39] br[39] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_42 
+ bl[40] br[40] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_43 
+ bl[41] br[41] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_44 
+ bl[42] br[42] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_45 
+ bl[43] br[43] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_46 
+ bl[44] br[44] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_47 
+ bl[45] br[45] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_48 
+ bl[46] br[46] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_49 
+ bl[47] br[47] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_50 
+ bl[48] br[48] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_51 
+ bl[49] br[49] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_52 
+ bl[50] br[50] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_53 
+ bl[51] br[51] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_54 
+ bl[52] br[52] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_55 
+ bl[53] br[53] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_56 
+ bl[54] br[54] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_57 
+ bl[55] br[55] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_58 
+ bl[56] br[56] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_59 
+ bl[57] br[57] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_60 
+ bl[58] br[58] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_61 
+ bl[59] br[59] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_62 
+ bl[60] br[60] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_63 
+ bl[61] br[61] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_64 
+ bl[62] br[62] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_65 
+ bl[63] br[63] vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_66 
+ vdd vdd vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_230_67 
+ vdd vdd vdd vss wl[228] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_0 
+ vdd vdd vss vdd vpb vnb wl[229] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_231_1 
+ rbl rbr vss vdd vpb vnb wl[229] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_231_2 
+ bl[0] br[0] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_3 
+ bl[1] br[1] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_4 
+ bl[2] br[2] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_5 
+ bl[3] br[3] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_6 
+ bl[4] br[4] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_7 
+ bl[5] br[5] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_8 
+ bl[6] br[6] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_9 
+ bl[7] br[7] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_10 
+ bl[8] br[8] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_11 
+ bl[9] br[9] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_12 
+ bl[10] br[10] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_13 
+ bl[11] br[11] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_14 
+ bl[12] br[12] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_15 
+ bl[13] br[13] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_16 
+ bl[14] br[14] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_17 
+ bl[15] br[15] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_18 
+ bl[16] br[16] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_19 
+ bl[17] br[17] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_20 
+ bl[18] br[18] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_21 
+ bl[19] br[19] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_22 
+ bl[20] br[20] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_23 
+ bl[21] br[21] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_24 
+ bl[22] br[22] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_25 
+ bl[23] br[23] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_26 
+ bl[24] br[24] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_27 
+ bl[25] br[25] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_28 
+ bl[26] br[26] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_29 
+ bl[27] br[27] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_30 
+ bl[28] br[28] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_31 
+ bl[29] br[29] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_32 
+ bl[30] br[30] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_33 
+ bl[31] br[31] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_34 
+ bl[32] br[32] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_35 
+ bl[33] br[33] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_36 
+ bl[34] br[34] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_37 
+ bl[35] br[35] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_38 
+ bl[36] br[36] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_39 
+ bl[37] br[37] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_40 
+ bl[38] br[38] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_41 
+ bl[39] br[39] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_42 
+ bl[40] br[40] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_43 
+ bl[41] br[41] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_44 
+ bl[42] br[42] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_45 
+ bl[43] br[43] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_46 
+ bl[44] br[44] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_47 
+ bl[45] br[45] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_48 
+ bl[46] br[46] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_49 
+ bl[47] br[47] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_50 
+ bl[48] br[48] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_51 
+ bl[49] br[49] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_52 
+ bl[50] br[50] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_53 
+ bl[51] br[51] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_54 
+ bl[52] br[52] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_55 
+ bl[53] br[53] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_56 
+ bl[54] br[54] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_57 
+ bl[55] br[55] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_58 
+ bl[56] br[56] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_59 
+ bl[57] br[57] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_60 
+ bl[58] br[58] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_61 
+ bl[59] br[59] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_62 
+ bl[60] br[60] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_63 
+ bl[61] br[61] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_64 
+ bl[62] br[62] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_65 
+ bl[63] br[63] vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_66 
+ vdd vdd vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_231_67 
+ vdd vdd vdd vss wl[229] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_0 
+ vdd vdd vss vdd vpb vnb wl[230] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_232_1 
+ rbl rbr vss vdd vpb vnb wl[230] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_232_2 
+ bl[0] br[0] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_3 
+ bl[1] br[1] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_4 
+ bl[2] br[2] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_5 
+ bl[3] br[3] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_6 
+ bl[4] br[4] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_7 
+ bl[5] br[5] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_8 
+ bl[6] br[6] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_9 
+ bl[7] br[7] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_10 
+ bl[8] br[8] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_11 
+ bl[9] br[9] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_12 
+ bl[10] br[10] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_13 
+ bl[11] br[11] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_14 
+ bl[12] br[12] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_15 
+ bl[13] br[13] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_16 
+ bl[14] br[14] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_17 
+ bl[15] br[15] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_18 
+ bl[16] br[16] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_19 
+ bl[17] br[17] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_20 
+ bl[18] br[18] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_21 
+ bl[19] br[19] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_22 
+ bl[20] br[20] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_23 
+ bl[21] br[21] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_24 
+ bl[22] br[22] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_25 
+ bl[23] br[23] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_26 
+ bl[24] br[24] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_27 
+ bl[25] br[25] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_28 
+ bl[26] br[26] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_29 
+ bl[27] br[27] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_30 
+ bl[28] br[28] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_31 
+ bl[29] br[29] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_32 
+ bl[30] br[30] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_33 
+ bl[31] br[31] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_34 
+ bl[32] br[32] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_35 
+ bl[33] br[33] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_36 
+ bl[34] br[34] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_37 
+ bl[35] br[35] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_38 
+ bl[36] br[36] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_39 
+ bl[37] br[37] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_40 
+ bl[38] br[38] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_41 
+ bl[39] br[39] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_42 
+ bl[40] br[40] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_43 
+ bl[41] br[41] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_44 
+ bl[42] br[42] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_45 
+ bl[43] br[43] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_46 
+ bl[44] br[44] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_47 
+ bl[45] br[45] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_48 
+ bl[46] br[46] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_49 
+ bl[47] br[47] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_50 
+ bl[48] br[48] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_51 
+ bl[49] br[49] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_52 
+ bl[50] br[50] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_53 
+ bl[51] br[51] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_54 
+ bl[52] br[52] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_55 
+ bl[53] br[53] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_56 
+ bl[54] br[54] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_57 
+ bl[55] br[55] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_58 
+ bl[56] br[56] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_59 
+ bl[57] br[57] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_60 
+ bl[58] br[58] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_61 
+ bl[59] br[59] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_62 
+ bl[60] br[60] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_63 
+ bl[61] br[61] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_64 
+ bl[62] br[62] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_65 
+ bl[63] br[63] vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_66 
+ vdd vdd vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_232_67 
+ vdd vdd vdd vss wl[230] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_0 
+ vdd vdd vss vdd vpb vnb wl[231] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_233_1 
+ rbl rbr vss vdd vpb vnb wl[231] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_233_2 
+ bl[0] br[0] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_3 
+ bl[1] br[1] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_4 
+ bl[2] br[2] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_5 
+ bl[3] br[3] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_6 
+ bl[4] br[4] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_7 
+ bl[5] br[5] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_8 
+ bl[6] br[6] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_9 
+ bl[7] br[7] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_10 
+ bl[8] br[8] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_11 
+ bl[9] br[9] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_12 
+ bl[10] br[10] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_13 
+ bl[11] br[11] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_14 
+ bl[12] br[12] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_15 
+ bl[13] br[13] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_16 
+ bl[14] br[14] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_17 
+ bl[15] br[15] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_18 
+ bl[16] br[16] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_19 
+ bl[17] br[17] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_20 
+ bl[18] br[18] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_21 
+ bl[19] br[19] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_22 
+ bl[20] br[20] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_23 
+ bl[21] br[21] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_24 
+ bl[22] br[22] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_25 
+ bl[23] br[23] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_26 
+ bl[24] br[24] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_27 
+ bl[25] br[25] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_28 
+ bl[26] br[26] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_29 
+ bl[27] br[27] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_30 
+ bl[28] br[28] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_31 
+ bl[29] br[29] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_32 
+ bl[30] br[30] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_33 
+ bl[31] br[31] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_34 
+ bl[32] br[32] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_35 
+ bl[33] br[33] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_36 
+ bl[34] br[34] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_37 
+ bl[35] br[35] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_38 
+ bl[36] br[36] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_39 
+ bl[37] br[37] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_40 
+ bl[38] br[38] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_41 
+ bl[39] br[39] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_42 
+ bl[40] br[40] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_43 
+ bl[41] br[41] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_44 
+ bl[42] br[42] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_45 
+ bl[43] br[43] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_46 
+ bl[44] br[44] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_47 
+ bl[45] br[45] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_48 
+ bl[46] br[46] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_49 
+ bl[47] br[47] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_50 
+ bl[48] br[48] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_51 
+ bl[49] br[49] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_52 
+ bl[50] br[50] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_53 
+ bl[51] br[51] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_54 
+ bl[52] br[52] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_55 
+ bl[53] br[53] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_56 
+ bl[54] br[54] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_57 
+ bl[55] br[55] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_58 
+ bl[56] br[56] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_59 
+ bl[57] br[57] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_60 
+ bl[58] br[58] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_61 
+ bl[59] br[59] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_62 
+ bl[60] br[60] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_63 
+ bl[61] br[61] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_64 
+ bl[62] br[62] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_65 
+ bl[63] br[63] vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_66 
+ vdd vdd vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_233_67 
+ vdd vdd vdd vss wl[231] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_0 
+ vdd vdd vss vdd vpb vnb wl[232] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_234_1 
+ rbl rbr vss vdd vpb vnb wl[232] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_234_2 
+ bl[0] br[0] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_3 
+ bl[1] br[1] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_4 
+ bl[2] br[2] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_5 
+ bl[3] br[3] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_6 
+ bl[4] br[4] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_7 
+ bl[5] br[5] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_8 
+ bl[6] br[6] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_9 
+ bl[7] br[7] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_10 
+ bl[8] br[8] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_11 
+ bl[9] br[9] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_12 
+ bl[10] br[10] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_13 
+ bl[11] br[11] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_14 
+ bl[12] br[12] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_15 
+ bl[13] br[13] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_16 
+ bl[14] br[14] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_17 
+ bl[15] br[15] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_18 
+ bl[16] br[16] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_19 
+ bl[17] br[17] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_20 
+ bl[18] br[18] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_21 
+ bl[19] br[19] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_22 
+ bl[20] br[20] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_23 
+ bl[21] br[21] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_24 
+ bl[22] br[22] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_25 
+ bl[23] br[23] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_26 
+ bl[24] br[24] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_27 
+ bl[25] br[25] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_28 
+ bl[26] br[26] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_29 
+ bl[27] br[27] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_30 
+ bl[28] br[28] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_31 
+ bl[29] br[29] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_32 
+ bl[30] br[30] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_33 
+ bl[31] br[31] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_34 
+ bl[32] br[32] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_35 
+ bl[33] br[33] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_36 
+ bl[34] br[34] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_37 
+ bl[35] br[35] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_38 
+ bl[36] br[36] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_39 
+ bl[37] br[37] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_40 
+ bl[38] br[38] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_41 
+ bl[39] br[39] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_42 
+ bl[40] br[40] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_43 
+ bl[41] br[41] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_44 
+ bl[42] br[42] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_45 
+ bl[43] br[43] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_46 
+ bl[44] br[44] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_47 
+ bl[45] br[45] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_48 
+ bl[46] br[46] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_49 
+ bl[47] br[47] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_50 
+ bl[48] br[48] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_51 
+ bl[49] br[49] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_52 
+ bl[50] br[50] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_53 
+ bl[51] br[51] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_54 
+ bl[52] br[52] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_55 
+ bl[53] br[53] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_56 
+ bl[54] br[54] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_57 
+ bl[55] br[55] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_58 
+ bl[56] br[56] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_59 
+ bl[57] br[57] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_60 
+ bl[58] br[58] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_61 
+ bl[59] br[59] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_62 
+ bl[60] br[60] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_63 
+ bl[61] br[61] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_64 
+ bl[62] br[62] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_65 
+ bl[63] br[63] vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_66 
+ vdd vdd vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_234_67 
+ vdd vdd vdd vss wl[232] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_0 
+ vdd vdd vss vdd vpb vnb wl[233] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_235_1 
+ rbl rbr vss vdd vpb vnb wl[233] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_235_2 
+ bl[0] br[0] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_3 
+ bl[1] br[1] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_4 
+ bl[2] br[2] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_5 
+ bl[3] br[3] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_6 
+ bl[4] br[4] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_7 
+ bl[5] br[5] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_8 
+ bl[6] br[6] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_9 
+ bl[7] br[7] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_10 
+ bl[8] br[8] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_11 
+ bl[9] br[9] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_12 
+ bl[10] br[10] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_13 
+ bl[11] br[11] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_14 
+ bl[12] br[12] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_15 
+ bl[13] br[13] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_16 
+ bl[14] br[14] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_17 
+ bl[15] br[15] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_18 
+ bl[16] br[16] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_19 
+ bl[17] br[17] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_20 
+ bl[18] br[18] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_21 
+ bl[19] br[19] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_22 
+ bl[20] br[20] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_23 
+ bl[21] br[21] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_24 
+ bl[22] br[22] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_25 
+ bl[23] br[23] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_26 
+ bl[24] br[24] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_27 
+ bl[25] br[25] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_28 
+ bl[26] br[26] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_29 
+ bl[27] br[27] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_30 
+ bl[28] br[28] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_31 
+ bl[29] br[29] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_32 
+ bl[30] br[30] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_33 
+ bl[31] br[31] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_34 
+ bl[32] br[32] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_35 
+ bl[33] br[33] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_36 
+ bl[34] br[34] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_37 
+ bl[35] br[35] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_38 
+ bl[36] br[36] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_39 
+ bl[37] br[37] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_40 
+ bl[38] br[38] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_41 
+ bl[39] br[39] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_42 
+ bl[40] br[40] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_43 
+ bl[41] br[41] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_44 
+ bl[42] br[42] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_45 
+ bl[43] br[43] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_46 
+ bl[44] br[44] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_47 
+ bl[45] br[45] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_48 
+ bl[46] br[46] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_49 
+ bl[47] br[47] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_50 
+ bl[48] br[48] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_51 
+ bl[49] br[49] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_52 
+ bl[50] br[50] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_53 
+ bl[51] br[51] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_54 
+ bl[52] br[52] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_55 
+ bl[53] br[53] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_56 
+ bl[54] br[54] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_57 
+ bl[55] br[55] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_58 
+ bl[56] br[56] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_59 
+ bl[57] br[57] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_60 
+ bl[58] br[58] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_61 
+ bl[59] br[59] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_62 
+ bl[60] br[60] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_63 
+ bl[61] br[61] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_64 
+ bl[62] br[62] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_65 
+ bl[63] br[63] vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_66 
+ vdd vdd vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_235_67 
+ vdd vdd vdd vss wl[233] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_0 
+ vdd vdd vss vdd vpb vnb wl[234] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_236_1 
+ rbl rbr vss vdd vpb vnb wl[234] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_236_2 
+ bl[0] br[0] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_3 
+ bl[1] br[1] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_4 
+ bl[2] br[2] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_5 
+ bl[3] br[3] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_6 
+ bl[4] br[4] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_7 
+ bl[5] br[5] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_8 
+ bl[6] br[6] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_9 
+ bl[7] br[7] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_10 
+ bl[8] br[8] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_11 
+ bl[9] br[9] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_12 
+ bl[10] br[10] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_13 
+ bl[11] br[11] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_14 
+ bl[12] br[12] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_15 
+ bl[13] br[13] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_16 
+ bl[14] br[14] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_17 
+ bl[15] br[15] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_18 
+ bl[16] br[16] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_19 
+ bl[17] br[17] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_20 
+ bl[18] br[18] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_21 
+ bl[19] br[19] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_22 
+ bl[20] br[20] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_23 
+ bl[21] br[21] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_24 
+ bl[22] br[22] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_25 
+ bl[23] br[23] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_26 
+ bl[24] br[24] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_27 
+ bl[25] br[25] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_28 
+ bl[26] br[26] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_29 
+ bl[27] br[27] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_30 
+ bl[28] br[28] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_31 
+ bl[29] br[29] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_32 
+ bl[30] br[30] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_33 
+ bl[31] br[31] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_34 
+ bl[32] br[32] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_35 
+ bl[33] br[33] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_36 
+ bl[34] br[34] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_37 
+ bl[35] br[35] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_38 
+ bl[36] br[36] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_39 
+ bl[37] br[37] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_40 
+ bl[38] br[38] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_41 
+ bl[39] br[39] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_42 
+ bl[40] br[40] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_43 
+ bl[41] br[41] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_44 
+ bl[42] br[42] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_45 
+ bl[43] br[43] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_46 
+ bl[44] br[44] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_47 
+ bl[45] br[45] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_48 
+ bl[46] br[46] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_49 
+ bl[47] br[47] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_50 
+ bl[48] br[48] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_51 
+ bl[49] br[49] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_52 
+ bl[50] br[50] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_53 
+ bl[51] br[51] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_54 
+ bl[52] br[52] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_55 
+ bl[53] br[53] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_56 
+ bl[54] br[54] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_57 
+ bl[55] br[55] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_58 
+ bl[56] br[56] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_59 
+ bl[57] br[57] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_60 
+ bl[58] br[58] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_61 
+ bl[59] br[59] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_62 
+ bl[60] br[60] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_63 
+ bl[61] br[61] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_64 
+ bl[62] br[62] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_65 
+ bl[63] br[63] vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_66 
+ vdd vdd vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_236_67 
+ vdd vdd vdd vss wl[234] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_0 
+ vdd vdd vss vdd vpb vnb wl[235] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_237_1 
+ rbl rbr vss vdd vpb vnb wl[235] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_237_2 
+ bl[0] br[0] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_3 
+ bl[1] br[1] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_4 
+ bl[2] br[2] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_5 
+ bl[3] br[3] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_6 
+ bl[4] br[4] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_7 
+ bl[5] br[5] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_8 
+ bl[6] br[6] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_9 
+ bl[7] br[7] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_10 
+ bl[8] br[8] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_11 
+ bl[9] br[9] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_12 
+ bl[10] br[10] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_13 
+ bl[11] br[11] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_14 
+ bl[12] br[12] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_15 
+ bl[13] br[13] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_16 
+ bl[14] br[14] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_17 
+ bl[15] br[15] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_18 
+ bl[16] br[16] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_19 
+ bl[17] br[17] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_20 
+ bl[18] br[18] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_21 
+ bl[19] br[19] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_22 
+ bl[20] br[20] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_23 
+ bl[21] br[21] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_24 
+ bl[22] br[22] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_25 
+ bl[23] br[23] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_26 
+ bl[24] br[24] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_27 
+ bl[25] br[25] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_28 
+ bl[26] br[26] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_29 
+ bl[27] br[27] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_30 
+ bl[28] br[28] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_31 
+ bl[29] br[29] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_32 
+ bl[30] br[30] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_33 
+ bl[31] br[31] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_34 
+ bl[32] br[32] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_35 
+ bl[33] br[33] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_36 
+ bl[34] br[34] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_37 
+ bl[35] br[35] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_38 
+ bl[36] br[36] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_39 
+ bl[37] br[37] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_40 
+ bl[38] br[38] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_41 
+ bl[39] br[39] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_42 
+ bl[40] br[40] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_43 
+ bl[41] br[41] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_44 
+ bl[42] br[42] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_45 
+ bl[43] br[43] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_46 
+ bl[44] br[44] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_47 
+ bl[45] br[45] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_48 
+ bl[46] br[46] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_49 
+ bl[47] br[47] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_50 
+ bl[48] br[48] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_51 
+ bl[49] br[49] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_52 
+ bl[50] br[50] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_53 
+ bl[51] br[51] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_54 
+ bl[52] br[52] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_55 
+ bl[53] br[53] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_56 
+ bl[54] br[54] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_57 
+ bl[55] br[55] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_58 
+ bl[56] br[56] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_59 
+ bl[57] br[57] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_60 
+ bl[58] br[58] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_61 
+ bl[59] br[59] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_62 
+ bl[60] br[60] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_63 
+ bl[61] br[61] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_64 
+ bl[62] br[62] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_65 
+ bl[63] br[63] vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_66 
+ vdd vdd vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_237_67 
+ vdd vdd vdd vss wl[235] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_0 
+ vdd vdd vss vdd vpb vnb wl[236] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_238_1 
+ rbl rbr vss vdd vpb vnb wl[236] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_238_2 
+ bl[0] br[0] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_3 
+ bl[1] br[1] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_4 
+ bl[2] br[2] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_5 
+ bl[3] br[3] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_6 
+ bl[4] br[4] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_7 
+ bl[5] br[5] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_8 
+ bl[6] br[6] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_9 
+ bl[7] br[7] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_10 
+ bl[8] br[8] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_11 
+ bl[9] br[9] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_12 
+ bl[10] br[10] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_13 
+ bl[11] br[11] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_14 
+ bl[12] br[12] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_15 
+ bl[13] br[13] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_16 
+ bl[14] br[14] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_17 
+ bl[15] br[15] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_18 
+ bl[16] br[16] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_19 
+ bl[17] br[17] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_20 
+ bl[18] br[18] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_21 
+ bl[19] br[19] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_22 
+ bl[20] br[20] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_23 
+ bl[21] br[21] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_24 
+ bl[22] br[22] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_25 
+ bl[23] br[23] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_26 
+ bl[24] br[24] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_27 
+ bl[25] br[25] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_28 
+ bl[26] br[26] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_29 
+ bl[27] br[27] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_30 
+ bl[28] br[28] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_31 
+ bl[29] br[29] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_32 
+ bl[30] br[30] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_33 
+ bl[31] br[31] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_34 
+ bl[32] br[32] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_35 
+ bl[33] br[33] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_36 
+ bl[34] br[34] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_37 
+ bl[35] br[35] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_38 
+ bl[36] br[36] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_39 
+ bl[37] br[37] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_40 
+ bl[38] br[38] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_41 
+ bl[39] br[39] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_42 
+ bl[40] br[40] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_43 
+ bl[41] br[41] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_44 
+ bl[42] br[42] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_45 
+ bl[43] br[43] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_46 
+ bl[44] br[44] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_47 
+ bl[45] br[45] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_48 
+ bl[46] br[46] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_49 
+ bl[47] br[47] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_50 
+ bl[48] br[48] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_51 
+ bl[49] br[49] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_52 
+ bl[50] br[50] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_53 
+ bl[51] br[51] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_54 
+ bl[52] br[52] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_55 
+ bl[53] br[53] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_56 
+ bl[54] br[54] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_57 
+ bl[55] br[55] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_58 
+ bl[56] br[56] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_59 
+ bl[57] br[57] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_60 
+ bl[58] br[58] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_61 
+ bl[59] br[59] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_62 
+ bl[60] br[60] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_63 
+ bl[61] br[61] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_64 
+ bl[62] br[62] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_65 
+ bl[63] br[63] vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_66 
+ vdd vdd vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_238_67 
+ vdd vdd vdd vss wl[236] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_0 
+ vdd vdd vss vdd vpb vnb wl[237] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_239_1 
+ rbl rbr vss vdd vpb vnb wl[237] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_239_2 
+ bl[0] br[0] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_3 
+ bl[1] br[1] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_4 
+ bl[2] br[2] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_5 
+ bl[3] br[3] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_6 
+ bl[4] br[4] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_7 
+ bl[5] br[5] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_8 
+ bl[6] br[6] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_9 
+ bl[7] br[7] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_10 
+ bl[8] br[8] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_11 
+ bl[9] br[9] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_12 
+ bl[10] br[10] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_13 
+ bl[11] br[11] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_14 
+ bl[12] br[12] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_15 
+ bl[13] br[13] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_16 
+ bl[14] br[14] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_17 
+ bl[15] br[15] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_18 
+ bl[16] br[16] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_19 
+ bl[17] br[17] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_20 
+ bl[18] br[18] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_21 
+ bl[19] br[19] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_22 
+ bl[20] br[20] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_23 
+ bl[21] br[21] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_24 
+ bl[22] br[22] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_25 
+ bl[23] br[23] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_26 
+ bl[24] br[24] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_27 
+ bl[25] br[25] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_28 
+ bl[26] br[26] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_29 
+ bl[27] br[27] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_30 
+ bl[28] br[28] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_31 
+ bl[29] br[29] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_32 
+ bl[30] br[30] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_33 
+ bl[31] br[31] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_34 
+ bl[32] br[32] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_35 
+ bl[33] br[33] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_36 
+ bl[34] br[34] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_37 
+ bl[35] br[35] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_38 
+ bl[36] br[36] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_39 
+ bl[37] br[37] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_40 
+ bl[38] br[38] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_41 
+ bl[39] br[39] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_42 
+ bl[40] br[40] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_43 
+ bl[41] br[41] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_44 
+ bl[42] br[42] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_45 
+ bl[43] br[43] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_46 
+ bl[44] br[44] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_47 
+ bl[45] br[45] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_48 
+ bl[46] br[46] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_49 
+ bl[47] br[47] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_50 
+ bl[48] br[48] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_51 
+ bl[49] br[49] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_52 
+ bl[50] br[50] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_53 
+ bl[51] br[51] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_54 
+ bl[52] br[52] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_55 
+ bl[53] br[53] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_56 
+ bl[54] br[54] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_57 
+ bl[55] br[55] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_58 
+ bl[56] br[56] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_59 
+ bl[57] br[57] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_60 
+ bl[58] br[58] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_61 
+ bl[59] br[59] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_62 
+ bl[60] br[60] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_63 
+ bl[61] br[61] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_64 
+ bl[62] br[62] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_65 
+ bl[63] br[63] vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_66 
+ vdd vdd vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_239_67 
+ vdd vdd vdd vss wl[237] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_0 
+ vdd vdd vss vdd vpb vnb wl[238] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_240_1 
+ rbl rbr vss vdd vpb vnb wl[238] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_240_2 
+ bl[0] br[0] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_3 
+ bl[1] br[1] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_4 
+ bl[2] br[2] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_5 
+ bl[3] br[3] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_6 
+ bl[4] br[4] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_7 
+ bl[5] br[5] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_8 
+ bl[6] br[6] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_9 
+ bl[7] br[7] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_10 
+ bl[8] br[8] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_11 
+ bl[9] br[9] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_12 
+ bl[10] br[10] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_13 
+ bl[11] br[11] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_14 
+ bl[12] br[12] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_15 
+ bl[13] br[13] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_16 
+ bl[14] br[14] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_17 
+ bl[15] br[15] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_18 
+ bl[16] br[16] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_19 
+ bl[17] br[17] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_20 
+ bl[18] br[18] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_21 
+ bl[19] br[19] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_22 
+ bl[20] br[20] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_23 
+ bl[21] br[21] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_24 
+ bl[22] br[22] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_25 
+ bl[23] br[23] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_26 
+ bl[24] br[24] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_27 
+ bl[25] br[25] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_28 
+ bl[26] br[26] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_29 
+ bl[27] br[27] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_30 
+ bl[28] br[28] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_31 
+ bl[29] br[29] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_32 
+ bl[30] br[30] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_33 
+ bl[31] br[31] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_34 
+ bl[32] br[32] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_35 
+ bl[33] br[33] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_36 
+ bl[34] br[34] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_37 
+ bl[35] br[35] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_38 
+ bl[36] br[36] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_39 
+ bl[37] br[37] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_40 
+ bl[38] br[38] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_41 
+ bl[39] br[39] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_42 
+ bl[40] br[40] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_43 
+ bl[41] br[41] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_44 
+ bl[42] br[42] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_45 
+ bl[43] br[43] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_46 
+ bl[44] br[44] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_47 
+ bl[45] br[45] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_48 
+ bl[46] br[46] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_49 
+ bl[47] br[47] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_50 
+ bl[48] br[48] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_51 
+ bl[49] br[49] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_52 
+ bl[50] br[50] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_53 
+ bl[51] br[51] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_54 
+ bl[52] br[52] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_55 
+ bl[53] br[53] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_56 
+ bl[54] br[54] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_57 
+ bl[55] br[55] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_58 
+ bl[56] br[56] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_59 
+ bl[57] br[57] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_60 
+ bl[58] br[58] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_61 
+ bl[59] br[59] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_62 
+ bl[60] br[60] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_63 
+ bl[61] br[61] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_64 
+ bl[62] br[62] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_65 
+ bl[63] br[63] vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_66 
+ vdd vdd vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_240_67 
+ vdd vdd vdd vss wl[238] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_0 
+ vdd vdd vss vdd vpb vnb wl[239] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_241_1 
+ rbl rbr vss vdd vpb vnb wl[239] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_241_2 
+ bl[0] br[0] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_3 
+ bl[1] br[1] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_4 
+ bl[2] br[2] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_5 
+ bl[3] br[3] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_6 
+ bl[4] br[4] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_7 
+ bl[5] br[5] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_8 
+ bl[6] br[6] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_9 
+ bl[7] br[7] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_10 
+ bl[8] br[8] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_11 
+ bl[9] br[9] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_12 
+ bl[10] br[10] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_13 
+ bl[11] br[11] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_14 
+ bl[12] br[12] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_15 
+ bl[13] br[13] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_16 
+ bl[14] br[14] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_17 
+ bl[15] br[15] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_18 
+ bl[16] br[16] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_19 
+ bl[17] br[17] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_20 
+ bl[18] br[18] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_21 
+ bl[19] br[19] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_22 
+ bl[20] br[20] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_23 
+ bl[21] br[21] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_24 
+ bl[22] br[22] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_25 
+ bl[23] br[23] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_26 
+ bl[24] br[24] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_27 
+ bl[25] br[25] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_28 
+ bl[26] br[26] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_29 
+ bl[27] br[27] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_30 
+ bl[28] br[28] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_31 
+ bl[29] br[29] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_32 
+ bl[30] br[30] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_33 
+ bl[31] br[31] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_34 
+ bl[32] br[32] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_35 
+ bl[33] br[33] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_36 
+ bl[34] br[34] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_37 
+ bl[35] br[35] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_38 
+ bl[36] br[36] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_39 
+ bl[37] br[37] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_40 
+ bl[38] br[38] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_41 
+ bl[39] br[39] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_42 
+ bl[40] br[40] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_43 
+ bl[41] br[41] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_44 
+ bl[42] br[42] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_45 
+ bl[43] br[43] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_46 
+ bl[44] br[44] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_47 
+ bl[45] br[45] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_48 
+ bl[46] br[46] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_49 
+ bl[47] br[47] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_50 
+ bl[48] br[48] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_51 
+ bl[49] br[49] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_52 
+ bl[50] br[50] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_53 
+ bl[51] br[51] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_54 
+ bl[52] br[52] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_55 
+ bl[53] br[53] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_56 
+ bl[54] br[54] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_57 
+ bl[55] br[55] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_58 
+ bl[56] br[56] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_59 
+ bl[57] br[57] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_60 
+ bl[58] br[58] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_61 
+ bl[59] br[59] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_62 
+ bl[60] br[60] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_63 
+ bl[61] br[61] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_64 
+ bl[62] br[62] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_65 
+ bl[63] br[63] vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_66 
+ vdd vdd vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_241_67 
+ vdd vdd vdd vss wl[239] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_0 
+ vdd vdd vss vdd vpb vnb wl[240] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_242_1 
+ rbl rbr vss vdd vpb vnb wl[240] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_242_2 
+ bl[0] br[0] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_3 
+ bl[1] br[1] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_4 
+ bl[2] br[2] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_5 
+ bl[3] br[3] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_6 
+ bl[4] br[4] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_7 
+ bl[5] br[5] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_8 
+ bl[6] br[6] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_9 
+ bl[7] br[7] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_10 
+ bl[8] br[8] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_11 
+ bl[9] br[9] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_12 
+ bl[10] br[10] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_13 
+ bl[11] br[11] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_14 
+ bl[12] br[12] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_15 
+ bl[13] br[13] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_16 
+ bl[14] br[14] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_17 
+ bl[15] br[15] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_18 
+ bl[16] br[16] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_19 
+ bl[17] br[17] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_20 
+ bl[18] br[18] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_21 
+ bl[19] br[19] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_22 
+ bl[20] br[20] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_23 
+ bl[21] br[21] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_24 
+ bl[22] br[22] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_25 
+ bl[23] br[23] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_26 
+ bl[24] br[24] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_27 
+ bl[25] br[25] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_28 
+ bl[26] br[26] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_29 
+ bl[27] br[27] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_30 
+ bl[28] br[28] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_31 
+ bl[29] br[29] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_32 
+ bl[30] br[30] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_33 
+ bl[31] br[31] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_34 
+ bl[32] br[32] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_35 
+ bl[33] br[33] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_36 
+ bl[34] br[34] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_37 
+ bl[35] br[35] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_38 
+ bl[36] br[36] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_39 
+ bl[37] br[37] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_40 
+ bl[38] br[38] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_41 
+ bl[39] br[39] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_42 
+ bl[40] br[40] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_43 
+ bl[41] br[41] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_44 
+ bl[42] br[42] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_45 
+ bl[43] br[43] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_46 
+ bl[44] br[44] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_47 
+ bl[45] br[45] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_48 
+ bl[46] br[46] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_49 
+ bl[47] br[47] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_50 
+ bl[48] br[48] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_51 
+ bl[49] br[49] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_52 
+ bl[50] br[50] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_53 
+ bl[51] br[51] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_54 
+ bl[52] br[52] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_55 
+ bl[53] br[53] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_56 
+ bl[54] br[54] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_57 
+ bl[55] br[55] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_58 
+ bl[56] br[56] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_59 
+ bl[57] br[57] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_60 
+ bl[58] br[58] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_61 
+ bl[59] br[59] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_62 
+ bl[60] br[60] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_63 
+ bl[61] br[61] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_64 
+ bl[62] br[62] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_65 
+ bl[63] br[63] vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_66 
+ vdd vdd vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_242_67 
+ vdd vdd vdd vss wl[240] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_0 
+ vdd vdd vss vdd vpb vnb wl[241] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_243_1 
+ rbl rbr vss vdd vpb vnb wl[241] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_243_2 
+ bl[0] br[0] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_3 
+ bl[1] br[1] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_4 
+ bl[2] br[2] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_5 
+ bl[3] br[3] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_6 
+ bl[4] br[4] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_7 
+ bl[5] br[5] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_8 
+ bl[6] br[6] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_9 
+ bl[7] br[7] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_10 
+ bl[8] br[8] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_11 
+ bl[9] br[9] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_12 
+ bl[10] br[10] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_13 
+ bl[11] br[11] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_14 
+ bl[12] br[12] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_15 
+ bl[13] br[13] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_16 
+ bl[14] br[14] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_17 
+ bl[15] br[15] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_18 
+ bl[16] br[16] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_19 
+ bl[17] br[17] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_20 
+ bl[18] br[18] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_21 
+ bl[19] br[19] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_22 
+ bl[20] br[20] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_23 
+ bl[21] br[21] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_24 
+ bl[22] br[22] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_25 
+ bl[23] br[23] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_26 
+ bl[24] br[24] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_27 
+ bl[25] br[25] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_28 
+ bl[26] br[26] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_29 
+ bl[27] br[27] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_30 
+ bl[28] br[28] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_31 
+ bl[29] br[29] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_32 
+ bl[30] br[30] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_33 
+ bl[31] br[31] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_34 
+ bl[32] br[32] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_35 
+ bl[33] br[33] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_36 
+ bl[34] br[34] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_37 
+ bl[35] br[35] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_38 
+ bl[36] br[36] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_39 
+ bl[37] br[37] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_40 
+ bl[38] br[38] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_41 
+ bl[39] br[39] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_42 
+ bl[40] br[40] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_43 
+ bl[41] br[41] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_44 
+ bl[42] br[42] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_45 
+ bl[43] br[43] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_46 
+ bl[44] br[44] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_47 
+ bl[45] br[45] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_48 
+ bl[46] br[46] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_49 
+ bl[47] br[47] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_50 
+ bl[48] br[48] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_51 
+ bl[49] br[49] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_52 
+ bl[50] br[50] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_53 
+ bl[51] br[51] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_54 
+ bl[52] br[52] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_55 
+ bl[53] br[53] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_56 
+ bl[54] br[54] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_57 
+ bl[55] br[55] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_58 
+ bl[56] br[56] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_59 
+ bl[57] br[57] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_60 
+ bl[58] br[58] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_61 
+ bl[59] br[59] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_62 
+ bl[60] br[60] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_63 
+ bl[61] br[61] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_64 
+ bl[62] br[62] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_65 
+ bl[63] br[63] vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_66 
+ vdd vdd vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_243_67 
+ vdd vdd vdd vss wl[241] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_0 
+ vdd vdd vss vdd vpb vnb wl[242] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_244_1 
+ rbl rbr vss vdd vpb vnb wl[242] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_244_2 
+ bl[0] br[0] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_3 
+ bl[1] br[1] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_4 
+ bl[2] br[2] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_5 
+ bl[3] br[3] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_6 
+ bl[4] br[4] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_7 
+ bl[5] br[5] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_8 
+ bl[6] br[6] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_9 
+ bl[7] br[7] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_10 
+ bl[8] br[8] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_11 
+ bl[9] br[9] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_12 
+ bl[10] br[10] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_13 
+ bl[11] br[11] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_14 
+ bl[12] br[12] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_15 
+ bl[13] br[13] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_16 
+ bl[14] br[14] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_17 
+ bl[15] br[15] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_18 
+ bl[16] br[16] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_19 
+ bl[17] br[17] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_20 
+ bl[18] br[18] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_21 
+ bl[19] br[19] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_22 
+ bl[20] br[20] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_23 
+ bl[21] br[21] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_24 
+ bl[22] br[22] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_25 
+ bl[23] br[23] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_26 
+ bl[24] br[24] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_27 
+ bl[25] br[25] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_28 
+ bl[26] br[26] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_29 
+ bl[27] br[27] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_30 
+ bl[28] br[28] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_31 
+ bl[29] br[29] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_32 
+ bl[30] br[30] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_33 
+ bl[31] br[31] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_34 
+ bl[32] br[32] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_35 
+ bl[33] br[33] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_36 
+ bl[34] br[34] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_37 
+ bl[35] br[35] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_38 
+ bl[36] br[36] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_39 
+ bl[37] br[37] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_40 
+ bl[38] br[38] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_41 
+ bl[39] br[39] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_42 
+ bl[40] br[40] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_43 
+ bl[41] br[41] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_44 
+ bl[42] br[42] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_45 
+ bl[43] br[43] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_46 
+ bl[44] br[44] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_47 
+ bl[45] br[45] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_48 
+ bl[46] br[46] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_49 
+ bl[47] br[47] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_50 
+ bl[48] br[48] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_51 
+ bl[49] br[49] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_52 
+ bl[50] br[50] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_53 
+ bl[51] br[51] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_54 
+ bl[52] br[52] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_55 
+ bl[53] br[53] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_56 
+ bl[54] br[54] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_57 
+ bl[55] br[55] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_58 
+ bl[56] br[56] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_59 
+ bl[57] br[57] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_60 
+ bl[58] br[58] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_61 
+ bl[59] br[59] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_62 
+ bl[60] br[60] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_63 
+ bl[61] br[61] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_64 
+ bl[62] br[62] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_65 
+ bl[63] br[63] vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_66 
+ vdd vdd vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_244_67 
+ vdd vdd vdd vss wl[242] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_0 
+ vdd vdd vss vdd vpb vnb wl[243] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_245_1 
+ rbl rbr vss vdd vpb vnb wl[243] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_245_2 
+ bl[0] br[0] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_3 
+ bl[1] br[1] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_4 
+ bl[2] br[2] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_5 
+ bl[3] br[3] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_6 
+ bl[4] br[4] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_7 
+ bl[5] br[5] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_8 
+ bl[6] br[6] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_9 
+ bl[7] br[7] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_10 
+ bl[8] br[8] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_11 
+ bl[9] br[9] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_12 
+ bl[10] br[10] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_13 
+ bl[11] br[11] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_14 
+ bl[12] br[12] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_15 
+ bl[13] br[13] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_16 
+ bl[14] br[14] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_17 
+ bl[15] br[15] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_18 
+ bl[16] br[16] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_19 
+ bl[17] br[17] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_20 
+ bl[18] br[18] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_21 
+ bl[19] br[19] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_22 
+ bl[20] br[20] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_23 
+ bl[21] br[21] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_24 
+ bl[22] br[22] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_25 
+ bl[23] br[23] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_26 
+ bl[24] br[24] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_27 
+ bl[25] br[25] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_28 
+ bl[26] br[26] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_29 
+ bl[27] br[27] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_30 
+ bl[28] br[28] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_31 
+ bl[29] br[29] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_32 
+ bl[30] br[30] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_33 
+ bl[31] br[31] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_34 
+ bl[32] br[32] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_35 
+ bl[33] br[33] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_36 
+ bl[34] br[34] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_37 
+ bl[35] br[35] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_38 
+ bl[36] br[36] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_39 
+ bl[37] br[37] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_40 
+ bl[38] br[38] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_41 
+ bl[39] br[39] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_42 
+ bl[40] br[40] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_43 
+ bl[41] br[41] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_44 
+ bl[42] br[42] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_45 
+ bl[43] br[43] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_46 
+ bl[44] br[44] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_47 
+ bl[45] br[45] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_48 
+ bl[46] br[46] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_49 
+ bl[47] br[47] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_50 
+ bl[48] br[48] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_51 
+ bl[49] br[49] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_52 
+ bl[50] br[50] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_53 
+ bl[51] br[51] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_54 
+ bl[52] br[52] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_55 
+ bl[53] br[53] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_56 
+ bl[54] br[54] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_57 
+ bl[55] br[55] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_58 
+ bl[56] br[56] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_59 
+ bl[57] br[57] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_60 
+ bl[58] br[58] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_61 
+ bl[59] br[59] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_62 
+ bl[60] br[60] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_63 
+ bl[61] br[61] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_64 
+ bl[62] br[62] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_65 
+ bl[63] br[63] vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_66 
+ vdd vdd vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_245_67 
+ vdd vdd vdd vss wl[243] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_0 
+ vdd vdd vss vdd vpb vnb wl[244] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_246_1 
+ rbl rbr vss vdd vpb vnb wl[244] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_246_2 
+ bl[0] br[0] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_3 
+ bl[1] br[1] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_4 
+ bl[2] br[2] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_5 
+ bl[3] br[3] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_6 
+ bl[4] br[4] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_7 
+ bl[5] br[5] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_8 
+ bl[6] br[6] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_9 
+ bl[7] br[7] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_10 
+ bl[8] br[8] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_11 
+ bl[9] br[9] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_12 
+ bl[10] br[10] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_13 
+ bl[11] br[11] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_14 
+ bl[12] br[12] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_15 
+ bl[13] br[13] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_16 
+ bl[14] br[14] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_17 
+ bl[15] br[15] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_18 
+ bl[16] br[16] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_19 
+ bl[17] br[17] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_20 
+ bl[18] br[18] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_21 
+ bl[19] br[19] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_22 
+ bl[20] br[20] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_23 
+ bl[21] br[21] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_24 
+ bl[22] br[22] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_25 
+ bl[23] br[23] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_26 
+ bl[24] br[24] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_27 
+ bl[25] br[25] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_28 
+ bl[26] br[26] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_29 
+ bl[27] br[27] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_30 
+ bl[28] br[28] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_31 
+ bl[29] br[29] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_32 
+ bl[30] br[30] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_33 
+ bl[31] br[31] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_34 
+ bl[32] br[32] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_35 
+ bl[33] br[33] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_36 
+ bl[34] br[34] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_37 
+ bl[35] br[35] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_38 
+ bl[36] br[36] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_39 
+ bl[37] br[37] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_40 
+ bl[38] br[38] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_41 
+ bl[39] br[39] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_42 
+ bl[40] br[40] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_43 
+ bl[41] br[41] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_44 
+ bl[42] br[42] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_45 
+ bl[43] br[43] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_46 
+ bl[44] br[44] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_47 
+ bl[45] br[45] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_48 
+ bl[46] br[46] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_49 
+ bl[47] br[47] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_50 
+ bl[48] br[48] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_51 
+ bl[49] br[49] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_52 
+ bl[50] br[50] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_53 
+ bl[51] br[51] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_54 
+ bl[52] br[52] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_55 
+ bl[53] br[53] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_56 
+ bl[54] br[54] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_57 
+ bl[55] br[55] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_58 
+ bl[56] br[56] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_59 
+ bl[57] br[57] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_60 
+ bl[58] br[58] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_61 
+ bl[59] br[59] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_62 
+ bl[60] br[60] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_63 
+ bl[61] br[61] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_64 
+ bl[62] br[62] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_65 
+ bl[63] br[63] vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_66 
+ vdd vdd vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_246_67 
+ vdd vdd vdd vss wl[244] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_0 
+ vdd vdd vss vdd vpb vnb wl[245] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_247_1 
+ rbl rbr vss vdd vpb vnb wl[245] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_247_2 
+ bl[0] br[0] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_3 
+ bl[1] br[1] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_4 
+ bl[2] br[2] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_5 
+ bl[3] br[3] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_6 
+ bl[4] br[4] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_7 
+ bl[5] br[5] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_8 
+ bl[6] br[6] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_9 
+ bl[7] br[7] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_10 
+ bl[8] br[8] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_11 
+ bl[9] br[9] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_12 
+ bl[10] br[10] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_13 
+ bl[11] br[11] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_14 
+ bl[12] br[12] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_15 
+ bl[13] br[13] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_16 
+ bl[14] br[14] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_17 
+ bl[15] br[15] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_18 
+ bl[16] br[16] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_19 
+ bl[17] br[17] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_20 
+ bl[18] br[18] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_21 
+ bl[19] br[19] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_22 
+ bl[20] br[20] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_23 
+ bl[21] br[21] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_24 
+ bl[22] br[22] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_25 
+ bl[23] br[23] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_26 
+ bl[24] br[24] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_27 
+ bl[25] br[25] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_28 
+ bl[26] br[26] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_29 
+ bl[27] br[27] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_30 
+ bl[28] br[28] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_31 
+ bl[29] br[29] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_32 
+ bl[30] br[30] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_33 
+ bl[31] br[31] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_34 
+ bl[32] br[32] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_35 
+ bl[33] br[33] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_36 
+ bl[34] br[34] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_37 
+ bl[35] br[35] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_38 
+ bl[36] br[36] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_39 
+ bl[37] br[37] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_40 
+ bl[38] br[38] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_41 
+ bl[39] br[39] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_42 
+ bl[40] br[40] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_43 
+ bl[41] br[41] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_44 
+ bl[42] br[42] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_45 
+ bl[43] br[43] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_46 
+ bl[44] br[44] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_47 
+ bl[45] br[45] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_48 
+ bl[46] br[46] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_49 
+ bl[47] br[47] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_50 
+ bl[48] br[48] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_51 
+ bl[49] br[49] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_52 
+ bl[50] br[50] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_53 
+ bl[51] br[51] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_54 
+ bl[52] br[52] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_55 
+ bl[53] br[53] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_56 
+ bl[54] br[54] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_57 
+ bl[55] br[55] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_58 
+ bl[56] br[56] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_59 
+ bl[57] br[57] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_60 
+ bl[58] br[58] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_61 
+ bl[59] br[59] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_62 
+ bl[60] br[60] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_63 
+ bl[61] br[61] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_64 
+ bl[62] br[62] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_65 
+ bl[63] br[63] vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_66 
+ vdd vdd vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_247_67 
+ vdd vdd vdd vss wl[245] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_0 
+ vdd vdd vss vdd vpb vnb wl[246] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_248_1 
+ rbl rbr vss vdd vpb vnb wl[246] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_248_2 
+ bl[0] br[0] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_3 
+ bl[1] br[1] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_4 
+ bl[2] br[2] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_5 
+ bl[3] br[3] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_6 
+ bl[4] br[4] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_7 
+ bl[5] br[5] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_8 
+ bl[6] br[6] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_9 
+ bl[7] br[7] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_10 
+ bl[8] br[8] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_11 
+ bl[9] br[9] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_12 
+ bl[10] br[10] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_13 
+ bl[11] br[11] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_14 
+ bl[12] br[12] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_15 
+ bl[13] br[13] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_16 
+ bl[14] br[14] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_17 
+ bl[15] br[15] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_18 
+ bl[16] br[16] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_19 
+ bl[17] br[17] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_20 
+ bl[18] br[18] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_21 
+ bl[19] br[19] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_22 
+ bl[20] br[20] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_23 
+ bl[21] br[21] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_24 
+ bl[22] br[22] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_25 
+ bl[23] br[23] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_26 
+ bl[24] br[24] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_27 
+ bl[25] br[25] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_28 
+ bl[26] br[26] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_29 
+ bl[27] br[27] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_30 
+ bl[28] br[28] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_31 
+ bl[29] br[29] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_32 
+ bl[30] br[30] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_33 
+ bl[31] br[31] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_34 
+ bl[32] br[32] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_35 
+ bl[33] br[33] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_36 
+ bl[34] br[34] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_37 
+ bl[35] br[35] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_38 
+ bl[36] br[36] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_39 
+ bl[37] br[37] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_40 
+ bl[38] br[38] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_41 
+ bl[39] br[39] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_42 
+ bl[40] br[40] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_43 
+ bl[41] br[41] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_44 
+ bl[42] br[42] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_45 
+ bl[43] br[43] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_46 
+ bl[44] br[44] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_47 
+ bl[45] br[45] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_48 
+ bl[46] br[46] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_49 
+ bl[47] br[47] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_50 
+ bl[48] br[48] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_51 
+ bl[49] br[49] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_52 
+ bl[50] br[50] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_53 
+ bl[51] br[51] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_54 
+ bl[52] br[52] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_55 
+ bl[53] br[53] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_56 
+ bl[54] br[54] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_57 
+ bl[55] br[55] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_58 
+ bl[56] br[56] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_59 
+ bl[57] br[57] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_60 
+ bl[58] br[58] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_61 
+ bl[59] br[59] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_62 
+ bl[60] br[60] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_63 
+ bl[61] br[61] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_64 
+ bl[62] br[62] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_65 
+ bl[63] br[63] vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_66 
+ vdd vdd vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_248_67 
+ vdd vdd vdd vss wl[246] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_0 
+ vdd vdd vss vdd vpb vnb wl[247] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_249_1 
+ rbl rbr vss vdd vpb vnb wl[247] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_249_2 
+ bl[0] br[0] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_3 
+ bl[1] br[1] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_4 
+ bl[2] br[2] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_5 
+ bl[3] br[3] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_6 
+ bl[4] br[4] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_7 
+ bl[5] br[5] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_8 
+ bl[6] br[6] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_9 
+ bl[7] br[7] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_10 
+ bl[8] br[8] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_11 
+ bl[9] br[9] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_12 
+ bl[10] br[10] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_13 
+ bl[11] br[11] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_14 
+ bl[12] br[12] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_15 
+ bl[13] br[13] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_16 
+ bl[14] br[14] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_17 
+ bl[15] br[15] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_18 
+ bl[16] br[16] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_19 
+ bl[17] br[17] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_20 
+ bl[18] br[18] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_21 
+ bl[19] br[19] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_22 
+ bl[20] br[20] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_23 
+ bl[21] br[21] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_24 
+ bl[22] br[22] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_25 
+ bl[23] br[23] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_26 
+ bl[24] br[24] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_27 
+ bl[25] br[25] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_28 
+ bl[26] br[26] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_29 
+ bl[27] br[27] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_30 
+ bl[28] br[28] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_31 
+ bl[29] br[29] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_32 
+ bl[30] br[30] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_33 
+ bl[31] br[31] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_34 
+ bl[32] br[32] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_35 
+ bl[33] br[33] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_36 
+ bl[34] br[34] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_37 
+ bl[35] br[35] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_38 
+ bl[36] br[36] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_39 
+ bl[37] br[37] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_40 
+ bl[38] br[38] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_41 
+ bl[39] br[39] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_42 
+ bl[40] br[40] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_43 
+ bl[41] br[41] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_44 
+ bl[42] br[42] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_45 
+ bl[43] br[43] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_46 
+ bl[44] br[44] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_47 
+ bl[45] br[45] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_48 
+ bl[46] br[46] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_49 
+ bl[47] br[47] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_50 
+ bl[48] br[48] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_51 
+ bl[49] br[49] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_52 
+ bl[50] br[50] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_53 
+ bl[51] br[51] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_54 
+ bl[52] br[52] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_55 
+ bl[53] br[53] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_56 
+ bl[54] br[54] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_57 
+ bl[55] br[55] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_58 
+ bl[56] br[56] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_59 
+ bl[57] br[57] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_60 
+ bl[58] br[58] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_61 
+ bl[59] br[59] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_62 
+ bl[60] br[60] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_63 
+ bl[61] br[61] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_64 
+ bl[62] br[62] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_65 
+ bl[63] br[63] vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_66 
+ vdd vdd vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_249_67 
+ vdd vdd vdd vss wl[247] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_0 
+ vdd vdd vss vdd vpb vnb wl[248] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_250_1 
+ rbl rbr vss vdd vpb vnb wl[248] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_250_2 
+ bl[0] br[0] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_3 
+ bl[1] br[1] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_4 
+ bl[2] br[2] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_5 
+ bl[3] br[3] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_6 
+ bl[4] br[4] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_7 
+ bl[5] br[5] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_8 
+ bl[6] br[6] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_9 
+ bl[7] br[7] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_10 
+ bl[8] br[8] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_11 
+ bl[9] br[9] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_12 
+ bl[10] br[10] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_13 
+ bl[11] br[11] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_14 
+ bl[12] br[12] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_15 
+ bl[13] br[13] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_16 
+ bl[14] br[14] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_17 
+ bl[15] br[15] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_18 
+ bl[16] br[16] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_19 
+ bl[17] br[17] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_20 
+ bl[18] br[18] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_21 
+ bl[19] br[19] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_22 
+ bl[20] br[20] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_23 
+ bl[21] br[21] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_24 
+ bl[22] br[22] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_25 
+ bl[23] br[23] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_26 
+ bl[24] br[24] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_27 
+ bl[25] br[25] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_28 
+ bl[26] br[26] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_29 
+ bl[27] br[27] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_30 
+ bl[28] br[28] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_31 
+ bl[29] br[29] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_32 
+ bl[30] br[30] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_33 
+ bl[31] br[31] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_34 
+ bl[32] br[32] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_35 
+ bl[33] br[33] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_36 
+ bl[34] br[34] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_37 
+ bl[35] br[35] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_38 
+ bl[36] br[36] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_39 
+ bl[37] br[37] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_40 
+ bl[38] br[38] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_41 
+ bl[39] br[39] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_42 
+ bl[40] br[40] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_43 
+ bl[41] br[41] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_44 
+ bl[42] br[42] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_45 
+ bl[43] br[43] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_46 
+ bl[44] br[44] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_47 
+ bl[45] br[45] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_48 
+ bl[46] br[46] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_49 
+ bl[47] br[47] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_50 
+ bl[48] br[48] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_51 
+ bl[49] br[49] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_52 
+ bl[50] br[50] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_53 
+ bl[51] br[51] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_54 
+ bl[52] br[52] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_55 
+ bl[53] br[53] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_56 
+ bl[54] br[54] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_57 
+ bl[55] br[55] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_58 
+ bl[56] br[56] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_59 
+ bl[57] br[57] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_60 
+ bl[58] br[58] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_61 
+ bl[59] br[59] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_62 
+ bl[60] br[60] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_63 
+ bl[61] br[61] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_64 
+ bl[62] br[62] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_65 
+ bl[63] br[63] vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_66 
+ vdd vdd vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_250_67 
+ vdd vdd vdd vss wl[248] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_0 
+ vdd vdd vss vdd vpb vnb wl[249] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_251_1 
+ rbl rbr vss vdd vpb vnb wl[249] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_251_2 
+ bl[0] br[0] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_3 
+ bl[1] br[1] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_4 
+ bl[2] br[2] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_5 
+ bl[3] br[3] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_6 
+ bl[4] br[4] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_7 
+ bl[5] br[5] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_8 
+ bl[6] br[6] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_9 
+ bl[7] br[7] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_10 
+ bl[8] br[8] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_11 
+ bl[9] br[9] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_12 
+ bl[10] br[10] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_13 
+ bl[11] br[11] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_14 
+ bl[12] br[12] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_15 
+ bl[13] br[13] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_16 
+ bl[14] br[14] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_17 
+ bl[15] br[15] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_18 
+ bl[16] br[16] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_19 
+ bl[17] br[17] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_20 
+ bl[18] br[18] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_21 
+ bl[19] br[19] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_22 
+ bl[20] br[20] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_23 
+ bl[21] br[21] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_24 
+ bl[22] br[22] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_25 
+ bl[23] br[23] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_26 
+ bl[24] br[24] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_27 
+ bl[25] br[25] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_28 
+ bl[26] br[26] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_29 
+ bl[27] br[27] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_30 
+ bl[28] br[28] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_31 
+ bl[29] br[29] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_32 
+ bl[30] br[30] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_33 
+ bl[31] br[31] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_34 
+ bl[32] br[32] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_35 
+ bl[33] br[33] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_36 
+ bl[34] br[34] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_37 
+ bl[35] br[35] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_38 
+ bl[36] br[36] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_39 
+ bl[37] br[37] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_40 
+ bl[38] br[38] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_41 
+ bl[39] br[39] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_42 
+ bl[40] br[40] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_43 
+ bl[41] br[41] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_44 
+ bl[42] br[42] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_45 
+ bl[43] br[43] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_46 
+ bl[44] br[44] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_47 
+ bl[45] br[45] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_48 
+ bl[46] br[46] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_49 
+ bl[47] br[47] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_50 
+ bl[48] br[48] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_51 
+ bl[49] br[49] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_52 
+ bl[50] br[50] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_53 
+ bl[51] br[51] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_54 
+ bl[52] br[52] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_55 
+ bl[53] br[53] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_56 
+ bl[54] br[54] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_57 
+ bl[55] br[55] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_58 
+ bl[56] br[56] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_59 
+ bl[57] br[57] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_60 
+ bl[58] br[58] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_61 
+ bl[59] br[59] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_62 
+ bl[60] br[60] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_63 
+ bl[61] br[61] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_64 
+ bl[62] br[62] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_65 
+ bl[63] br[63] vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_66 
+ vdd vdd vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_251_67 
+ vdd vdd vdd vss wl[249] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_0 
+ vdd vdd vss vdd vpb vnb wl[250] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_252_1 
+ rbl rbr vss vdd vpb vnb wl[250] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_252_2 
+ bl[0] br[0] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_3 
+ bl[1] br[1] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_4 
+ bl[2] br[2] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_5 
+ bl[3] br[3] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_6 
+ bl[4] br[4] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_7 
+ bl[5] br[5] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_8 
+ bl[6] br[6] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_9 
+ bl[7] br[7] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_10 
+ bl[8] br[8] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_11 
+ bl[9] br[9] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_12 
+ bl[10] br[10] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_13 
+ bl[11] br[11] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_14 
+ bl[12] br[12] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_15 
+ bl[13] br[13] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_16 
+ bl[14] br[14] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_17 
+ bl[15] br[15] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_18 
+ bl[16] br[16] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_19 
+ bl[17] br[17] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_20 
+ bl[18] br[18] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_21 
+ bl[19] br[19] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_22 
+ bl[20] br[20] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_23 
+ bl[21] br[21] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_24 
+ bl[22] br[22] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_25 
+ bl[23] br[23] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_26 
+ bl[24] br[24] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_27 
+ bl[25] br[25] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_28 
+ bl[26] br[26] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_29 
+ bl[27] br[27] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_30 
+ bl[28] br[28] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_31 
+ bl[29] br[29] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_32 
+ bl[30] br[30] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_33 
+ bl[31] br[31] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_34 
+ bl[32] br[32] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_35 
+ bl[33] br[33] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_36 
+ bl[34] br[34] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_37 
+ bl[35] br[35] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_38 
+ bl[36] br[36] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_39 
+ bl[37] br[37] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_40 
+ bl[38] br[38] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_41 
+ bl[39] br[39] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_42 
+ bl[40] br[40] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_43 
+ bl[41] br[41] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_44 
+ bl[42] br[42] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_45 
+ bl[43] br[43] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_46 
+ bl[44] br[44] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_47 
+ bl[45] br[45] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_48 
+ bl[46] br[46] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_49 
+ bl[47] br[47] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_50 
+ bl[48] br[48] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_51 
+ bl[49] br[49] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_52 
+ bl[50] br[50] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_53 
+ bl[51] br[51] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_54 
+ bl[52] br[52] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_55 
+ bl[53] br[53] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_56 
+ bl[54] br[54] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_57 
+ bl[55] br[55] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_58 
+ bl[56] br[56] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_59 
+ bl[57] br[57] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_60 
+ bl[58] br[58] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_61 
+ bl[59] br[59] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_62 
+ bl[60] br[60] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_63 
+ bl[61] br[61] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_64 
+ bl[62] br[62] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_65 
+ bl[63] br[63] vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_66 
+ vdd vdd vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_252_67 
+ vdd vdd vdd vss wl[250] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_0 
+ vdd vdd vss vdd vpb vnb wl[251] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_253_1 
+ rbl rbr vss vdd vpb vnb wl[251] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_253_2 
+ bl[0] br[0] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_3 
+ bl[1] br[1] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_4 
+ bl[2] br[2] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_5 
+ bl[3] br[3] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_6 
+ bl[4] br[4] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_7 
+ bl[5] br[5] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_8 
+ bl[6] br[6] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_9 
+ bl[7] br[7] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_10 
+ bl[8] br[8] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_11 
+ bl[9] br[9] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_12 
+ bl[10] br[10] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_13 
+ bl[11] br[11] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_14 
+ bl[12] br[12] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_15 
+ bl[13] br[13] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_16 
+ bl[14] br[14] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_17 
+ bl[15] br[15] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_18 
+ bl[16] br[16] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_19 
+ bl[17] br[17] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_20 
+ bl[18] br[18] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_21 
+ bl[19] br[19] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_22 
+ bl[20] br[20] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_23 
+ bl[21] br[21] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_24 
+ bl[22] br[22] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_25 
+ bl[23] br[23] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_26 
+ bl[24] br[24] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_27 
+ bl[25] br[25] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_28 
+ bl[26] br[26] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_29 
+ bl[27] br[27] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_30 
+ bl[28] br[28] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_31 
+ bl[29] br[29] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_32 
+ bl[30] br[30] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_33 
+ bl[31] br[31] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_34 
+ bl[32] br[32] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_35 
+ bl[33] br[33] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_36 
+ bl[34] br[34] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_37 
+ bl[35] br[35] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_38 
+ bl[36] br[36] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_39 
+ bl[37] br[37] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_40 
+ bl[38] br[38] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_41 
+ bl[39] br[39] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_42 
+ bl[40] br[40] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_43 
+ bl[41] br[41] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_44 
+ bl[42] br[42] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_45 
+ bl[43] br[43] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_46 
+ bl[44] br[44] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_47 
+ bl[45] br[45] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_48 
+ bl[46] br[46] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_49 
+ bl[47] br[47] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_50 
+ bl[48] br[48] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_51 
+ bl[49] br[49] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_52 
+ bl[50] br[50] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_53 
+ bl[51] br[51] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_54 
+ bl[52] br[52] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_55 
+ bl[53] br[53] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_56 
+ bl[54] br[54] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_57 
+ bl[55] br[55] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_58 
+ bl[56] br[56] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_59 
+ bl[57] br[57] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_60 
+ bl[58] br[58] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_61 
+ bl[59] br[59] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_62 
+ bl[60] br[60] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_63 
+ bl[61] br[61] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_64 
+ bl[62] br[62] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_65 
+ bl[63] br[63] vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_66 
+ vdd vdd vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_253_67 
+ vdd vdd vdd vss wl[251] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_0 
+ vdd vdd vss vdd vpb vnb wl[252] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_254_1 
+ rbl rbr vss vdd vpb vnb wl[252] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_254_2 
+ bl[0] br[0] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_3 
+ bl[1] br[1] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_4 
+ bl[2] br[2] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_5 
+ bl[3] br[3] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_6 
+ bl[4] br[4] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_7 
+ bl[5] br[5] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_8 
+ bl[6] br[6] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_9 
+ bl[7] br[7] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_10 
+ bl[8] br[8] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_11 
+ bl[9] br[9] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_12 
+ bl[10] br[10] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_13 
+ bl[11] br[11] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_14 
+ bl[12] br[12] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_15 
+ bl[13] br[13] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_16 
+ bl[14] br[14] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_17 
+ bl[15] br[15] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_18 
+ bl[16] br[16] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_19 
+ bl[17] br[17] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_20 
+ bl[18] br[18] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_21 
+ bl[19] br[19] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_22 
+ bl[20] br[20] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_23 
+ bl[21] br[21] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_24 
+ bl[22] br[22] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_25 
+ bl[23] br[23] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_26 
+ bl[24] br[24] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_27 
+ bl[25] br[25] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_28 
+ bl[26] br[26] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_29 
+ bl[27] br[27] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_30 
+ bl[28] br[28] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_31 
+ bl[29] br[29] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_32 
+ bl[30] br[30] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_33 
+ bl[31] br[31] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_34 
+ bl[32] br[32] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_35 
+ bl[33] br[33] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_36 
+ bl[34] br[34] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_37 
+ bl[35] br[35] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_38 
+ bl[36] br[36] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_39 
+ bl[37] br[37] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_40 
+ bl[38] br[38] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_41 
+ bl[39] br[39] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_42 
+ bl[40] br[40] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_43 
+ bl[41] br[41] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_44 
+ bl[42] br[42] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_45 
+ bl[43] br[43] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_46 
+ bl[44] br[44] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_47 
+ bl[45] br[45] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_48 
+ bl[46] br[46] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_49 
+ bl[47] br[47] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_50 
+ bl[48] br[48] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_51 
+ bl[49] br[49] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_52 
+ bl[50] br[50] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_53 
+ bl[51] br[51] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_54 
+ bl[52] br[52] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_55 
+ bl[53] br[53] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_56 
+ bl[54] br[54] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_57 
+ bl[55] br[55] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_58 
+ bl[56] br[56] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_59 
+ bl[57] br[57] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_60 
+ bl[58] br[58] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_61 
+ bl[59] br[59] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_62 
+ bl[60] br[60] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_63 
+ bl[61] br[61] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_64 
+ bl[62] br[62] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_65 
+ bl[63] br[63] vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_66 
+ vdd vdd vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_254_67 
+ vdd vdd vdd vss wl[252] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_0 
+ vdd vdd vss vdd vpb vnb wl[253] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_255_1 
+ rbl rbr vss vdd vpb vnb wl[253] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_255_2 
+ bl[0] br[0] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_3 
+ bl[1] br[1] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_4 
+ bl[2] br[2] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_5 
+ bl[3] br[3] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_6 
+ bl[4] br[4] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_7 
+ bl[5] br[5] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_8 
+ bl[6] br[6] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_9 
+ bl[7] br[7] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_10 
+ bl[8] br[8] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_11 
+ bl[9] br[9] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_12 
+ bl[10] br[10] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_13 
+ bl[11] br[11] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_14 
+ bl[12] br[12] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_15 
+ bl[13] br[13] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_16 
+ bl[14] br[14] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_17 
+ bl[15] br[15] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_18 
+ bl[16] br[16] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_19 
+ bl[17] br[17] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_20 
+ bl[18] br[18] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_21 
+ bl[19] br[19] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_22 
+ bl[20] br[20] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_23 
+ bl[21] br[21] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_24 
+ bl[22] br[22] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_25 
+ bl[23] br[23] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_26 
+ bl[24] br[24] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_27 
+ bl[25] br[25] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_28 
+ bl[26] br[26] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_29 
+ bl[27] br[27] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_30 
+ bl[28] br[28] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_31 
+ bl[29] br[29] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_32 
+ bl[30] br[30] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_33 
+ bl[31] br[31] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_34 
+ bl[32] br[32] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_35 
+ bl[33] br[33] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_36 
+ bl[34] br[34] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_37 
+ bl[35] br[35] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_38 
+ bl[36] br[36] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_39 
+ bl[37] br[37] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_40 
+ bl[38] br[38] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_41 
+ bl[39] br[39] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_42 
+ bl[40] br[40] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_43 
+ bl[41] br[41] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_44 
+ bl[42] br[42] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_45 
+ bl[43] br[43] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_46 
+ bl[44] br[44] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_47 
+ bl[45] br[45] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_48 
+ bl[46] br[46] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_49 
+ bl[47] br[47] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_50 
+ bl[48] br[48] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_51 
+ bl[49] br[49] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_52 
+ bl[50] br[50] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_53 
+ bl[51] br[51] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_54 
+ bl[52] br[52] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_55 
+ bl[53] br[53] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_56 
+ bl[54] br[54] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_57 
+ bl[55] br[55] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_58 
+ bl[56] br[56] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_59 
+ bl[57] br[57] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_60 
+ bl[58] br[58] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_61 
+ bl[59] br[59] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_62 
+ bl[60] br[60] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_63 
+ bl[61] br[61] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_64 
+ bl[62] br[62] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_65 
+ bl[63] br[63] vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_66 
+ vdd vdd vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_255_67 
+ vdd vdd vdd vss wl[253] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_0 
+ vdd vdd vss vdd vpb vnb wl[254] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_256_1 
+ rbl rbr vss vdd vpb vnb wl[254] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_256_2 
+ bl[0] br[0] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_3 
+ bl[1] br[1] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_4 
+ bl[2] br[2] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_5 
+ bl[3] br[3] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_6 
+ bl[4] br[4] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_7 
+ bl[5] br[5] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_8 
+ bl[6] br[6] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_9 
+ bl[7] br[7] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_10 
+ bl[8] br[8] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_11 
+ bl[9] br[9] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_12 
+ bl[10] br[10] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_13 
+ bl[11] br[11] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_14 
+ bl[12] br[12] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_15 
+ bl[13] br[13] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_16 
+ bl[14] br[14] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_17 
+ bl[15] br[15] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_18 
+ bl[16] br[16] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_19 
+ bl[17] br[17] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_20 
+ bl[18] br[18] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_21 
+ bl[19] br[19] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_22 
+ bl[20] br[20] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_23 
+ bl[21] br[21] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_24 
+ bl[22] br[22] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_25 
+ bl[23] br[23] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_26 
+ bl[24] br[24] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_27 
+ bl[25] br[25] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_28 
+ bl[26] br[26] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_29 
+ bl[27] br[27] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_30 
+ bl[28] br[28] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_31 
+ bl[29] br[29] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_32 
+ bl[30] br[30] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_33 
+ bl[31] br[31] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_34 
+ bl[32] br[32] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_35 
+ bl[33] br[33] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_36 
+ bl[34] br[34] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_37 
+ bl[35] br[35] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_38 
+ bl[36] br[36] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_39 
+ bl[37] br[37] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_40 
+ bl[38] br[38] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_41 
+ bl[39] br[39] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_42 
+ bl[40] br[40] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_43 
+ bl[41] br[41] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_44 
+ bl[42] br[42] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_45 
+ bl[43] br[43] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_46 
+ bl[44] br[44] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_47 
+ bl[45] br[45] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_48 
+ bl[46] br[46] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_49 
+ bl[47] br[47] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_50 
+ bl[48] br[48] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_51 
+ bl[49] br[49] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_52 
+ bl[50] br[50] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_53 
+ bl[51] br[51] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_54 
+ bl[52] br[52] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_55 
+ bl[53] br[53] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_56 
+ bl[54] br[54] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_57 
+ bl[55] br[55] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_58 
+ bl[56] br[56] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_59 
+ bl[57] br[57] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_60 
+ bl[58] br[58] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_61 
+ bl[59] br[59] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_62 
+ bl[60] br[60] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_63 
+ bl[61] br[61] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_64 
+ bl[62] br[62] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_65 
+ bl[63] br[63] vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_66 
+ vdd vdd vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_256_67 
+ vdd vdd vdd vss wl[254] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_0 
+ vdd vdd vss vdd vpb vnb wl[255] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_257_1 
+ rbl rbr vss vdd vpb vnb wl[255] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_257_2 
+ bl[0] br[0] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_3 
+ bl[1] br[1] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_4 
+ bl[2] br[2] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_5 
+ bl[3] br[3] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_6 
+ bl[4] br[4] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_7 
+ bl[5] br[5] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_8 
+ bl[6] br[6] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_9 
+ bl[7] br[7] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_10 
+ bl[8] br[8] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_11 
+ bl[9] br[9] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_12 
+ bl[10] br[10] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_13 
+ bl[11] br[11] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_14 
+ bl[12] br[12] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_15 
+ bl[13] br[13] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_16 
+ bl[14] br[14] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_17 
+ bl[15] br[15] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_18 
+ bl[16] br[16] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_19 
+ bl[17] br[17] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_20 
+ bl[18] br[18] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_21 
+ bl[19] br[19] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_22 
+ bl[20] br[20] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_23 
+ bl[21] br[21] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_24 
+ bl[22] br[22] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_25 
+ bl[23] br[23] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_26 
+ bl[24] br[24] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_27 
+ bl[25] br[25] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_28 
+ bl[26] br[26] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_29 
+ bl[27] br[27] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_30 
+ bl[28] br[28] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_31 
+ bl[29] br[29] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_32 
+ bl[30] br[30] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_33 
+ bl[31] br[31] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_34 
+ bl[32] br[32] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_35 
+ bl[33] br[33] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_36 
+ bl[34] br[34] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_37 
+ bl[35] br[35] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_38 
+ bl[36] br[36] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_39 
+ bl[37] br[37] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_40 
+ bl[38] br[38] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_41 
+ bl[39] br[39] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_42 
+ bl[40] br[40] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_43 
+ bl[41] br[41] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_44 
+ bl[42] br[42] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_45 
+ bl[43] br[43] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_46 
+ bl[44] br[44] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_47 
+ bl[45] br[45] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_48 
+ bl[46] br[46] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_49 
+ bl[47] br[47] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_50 
+ bl[48] br[48] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_51 
+ bl[49] br[49] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_52 
+ bl[50] br[50] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_53 
+ bl[51] br[51] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_54 
+ bl[52] br[52] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_55 
+ bl[53] br[53] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_56 
+ bl[54] br[54] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_57 
+ bl[55] br[55] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_58 
+ bl[56] br[56] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_59 
+ bl[57] br[57] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_60 
+ bl[58] br[58] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_61 
+ bl[59] br[59] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_62 
+ bl[60] br[60] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_63 
+ bl[61] br[61] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_64 
+ bl[62] br[62] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_65 
+ bl[63] br[63] vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_66 
+ vdd vdd vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_257_67 
+ vdd vdd vdd vss wl[255] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_0 
+ vdd vdd vss vdd vpb vnb wl[256] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_258_1 
+ rbl rbr vss vdd vpb vnb wl[256] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_258_2 
+ bl[0] br[0] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_3 
+ bl[1] br[1] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_4 
+ bl[2] br[2] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_5 
+ bl[3] br[3] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_6 
+ bl[4] br[4] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_7 
+ bl[5] br[5] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_8 
+ bl[6] br[6] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_9 
+ bl[7] br[7] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_10 
+ bl[8] br[8] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_11 
+ bl[9] br[9] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_12 
+ bl[10] br[10] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_13 
+ bl[11] br[11] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_14 
+ bl[12] br[12] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_15 
+ bl[13] br[13] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_16 
+ bl[14] br[14] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_17 
+ bl[15] br[15] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_18 
+ bl[16] br[16] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_19 
+ bl[17] br[17] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_20 
+ bl[18] br[18] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_21 
+ bl[19] br[19] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_22 
+ bl[20] br[20] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_23 
+ bl[21] br[21] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_24 
+ bl[22] br[22] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_25 
+ bl[23] br[23] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_26 
+ bl[24] br[24] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_27 
+ bl[25] br[25] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_28 
+ bl[26] br[26] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_29 
+ bl[27] br[27] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_30 
+ bl[28] br[28] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_31 
+ bl[29] br[29] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_32 
+ bl[30] br[30] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_33 
+ bl[31] br[31] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_34 
+ bl[32] br[32] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_35 
+ bl[33] br[33] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_36 
+ bl[34] br[34] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_37 
+ bl[35] br[35] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_38 
+ bl[36] br[36] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_39 
+ bl[37] br[37] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_40 
+ bl[38] br[38] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_41 
+ bl[39] br[39] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_42 
+ bl[40] br[40] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_43 
+ bl[41] br[41] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_44 
+ bl[42] br[42] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_45 
+ bl[43] br[43] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_46 
+ bl[44] br[44] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_47 
+ bl[45] br[45] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_48 
+ bl[46] br[46] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_49 
+ bl[47] br[47] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_50 
+ bl[48] br[48] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_51 
+ bl[49] br[49] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_52 
+ bl[50] br[50] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_53 
+ bl[51] br[51] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_54 
+ bl[52] br[52] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_55 
+ bl[53] br[53] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_56 
+ bl[54] br[54] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_57 
+ bl[55] br[55] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_58 
+ bl[56] br[56] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_59 
+ bl[57] br[57] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_60 
+ bl[58] br[58] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_61 
+ bl[59] br[59] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_62 
+ bl[60] br[60] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_63 
+ bl[61] br[61] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_64 
+ bl[62] br[62] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_65 
+ bl[63] br[63] vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_66 
+ vdd vdd vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_258_67 
+ vdd vdd vdd vss wl[256] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_0 
+ vdd vdd vss vdd vpb vnb wl[257] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_259_1 
+ rbl rbr vss vdd vpb vnb wl[257] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_259_2 
+ bl[0] br[0] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_3 
+ bl[1] br[1] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_4 
+ bl[2] br[2] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_5 
+ bl[3] br[3] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_6 
+ bl[4] br[4] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_7 
+ bl[5] br[5] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_8 
+ bl[6] br[6] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_9 
+ bl[7] br[7] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_10 
+ bl[8] br[8] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_11 
+ bl[9] br[9] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_12 
+ bl[10] br[10] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_13 
+ bl[11] br[11] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_14 
+ bl[12] br[12] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_15 
+ bl[13] br[13] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_16 
+ bl[14] br[14] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_17 
+ bl[15] br[15] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_18 
+ bl[16] br[16] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_19 
+ bl[17] br[17] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_20 
+ bl[18] br[18] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_21 
+ bl[19] br[19] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_22 
+ bl[20] br[20] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_23 
+ bl[21] br[21] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_24 
+ bl[22] br[22] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_25 
+ bl[23] br[23] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_26 
+ bl[24] br[24] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_27 
+ bl[25] br[25] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_28 
+ bl[26] br[26] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_29 
+ bl[27] br[27] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_30 
+ bl[28] br[28] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_31 
+ bl[29] br[29] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_32 
+ bl[30] br[30] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_33 
+ bl[31] br[31] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_34 
+ bl[32] br[32] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_35 
+ bl[33] br[33] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_36 
+ bl[34] br[34] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_37 
+ bl[35] br[35] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_38 
+ bl[36] br[36] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_39 
+ bl[37] br[37] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_40 
+ bl[38] br[38] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_41 
+ bl[39] br[39] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_42 
+ bl[40] br[40] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_43 
+ bl[41] br[41] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_44 
+ bl[42] br[42] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_45 
+ bl[43] br[43] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_46 
+ bl[44] br[44] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_47 
+ bl[45] br[45] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_48 
+ bl[46] br[46] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_49 
+ bl[47] br[47] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_50 
+ bl[48] br[48] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_51 
+ bl[49] br[49] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_52 
+ bl[50] br[50] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_53 
+ bl[51] br[51] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_54 
+ bl[52] br[52] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_55 
+ bl[53] br[53] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_56 
+ bl[54] br[54] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_57 
+ bl[55] br[55] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_58 
+ bl[56] br[56] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_59 
+ bl[57] br[57] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_60 
+ bl[58] br[58] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_61 
+ bl[59] br[59] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_62 
+ bl[60] br[60] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_63 
+ bl[61] br[61] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_64 
+ bl[62] br[62] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_65 
+ bl[63] br[63] vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_66 
+ vdd vdd vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_259_67 
+ vdd vdd vdd vss wl[257] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_0 
+ vdd vdd vss vdd vpb vnb wl[258] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_260_1 
+ rbl rbr vss vdd vpb vnb wl[258] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_260_2 
+ bl[0] br[0] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_3 
+ bl[1] br[1] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_4 
+ bl[2] br[2] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_5 
+ bl[3] br[3] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_6 
+ bl[4] br[4] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_7 
+ bl[5] br[5] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_8 
+ bl[6] br[6] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_9 
+ bl[7] br[7] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_10 
+ bl[8] br[8] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_11 
+ bl[9] br[9] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_12 
+ bl[10] br[10] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_13 
+ bl[11] br[11] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_14 
+ bl[12] br[12] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_15 
+ bl[13] br[13] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_16 
+ bl[14] br[14] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_17 
+ bl[15] br[15] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_18 
+ bl[16] br[16] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_19 
+ bl[17] br[17] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_20 
+ bl[18] br[18] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_21 
+ bl[19] br[19] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_22 
+ bl[20] br[20] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_23 
+ bl[21] br[21] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_24 
+ bl[22] br[22] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_25 
+ bl[23] br[23] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_26 
+ bl[24] br[24] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_27 
+ bl[25] br[25] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_28 
+ bl[26] br[26] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_29 
+ bl[27] br[27] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_30 
+ bl[28] br[28] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_31 
+ bl[29] br[29] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_32 
+ bl[30] br[30] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_33 
+ bl[31] br[31] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_34 
+ bl[32] br[32] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_35 
+ bl[33] br[33] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_36 
+ bl[34] br[34] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_37 
+ bl[35] br[35] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_38 
+ bl[36] br[36] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_39 
+ bl[37] br[37] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_40 
+ bl[38] br[38] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_41 
+ bl[39] br[39] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_42 
+ bl[40] br[40] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_43 
+ bl[41] br[41] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_44 
+ bl[42] br[42] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_45 
+ bl[43] br[43] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_46 
+ bl[44] br[44] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_47 
+ bl[45] br[45] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_48 
+ bl[46] br[46] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_49 
+ bl[47] br[47] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_50 
+ bl[48] br[48] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_51 
+ bl[49] br[49] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_52 
+ bl[50] br[50] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_53 
+ bl[51] br[51] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_54 
+ bl[52] br[52] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_55 
+ bl[53] br[53] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_56 
+ bl[54] br[54] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_57 
+ bl[55] br[55] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_58 
+ bl[56] br[56] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_59 
+ bl[57] br[57] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_60 
+ bl[58] br[58] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_61 
+ bl[59] br[59] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_62 
+ bl[60] br[60] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_63 
+ bl[61] br[61] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_64 
+ bl[62] br[62] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_65 
+ bl[63] br[63] vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_66 
+ vdd vdd vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_260_67 
+ vdd vdd vdd vss wl[258] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_0 
+ vdd vdd vss vdd vpb vnb wl[259] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_261_1 
+ rbl rbr vss vdd vpb vnb wl[259] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_261_2 
+ bl[0] br[0] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_3 
+ bl[1] br[1] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_4 
+ bl[2] br[2] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_5 
+ bl[3] br[3] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_6 
+ bl[4] br[4] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_7 
+ bl[5] br[5] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_8 
+ bl[6] br[6] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_9 
+ bl[7] br[7] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_10 
+ bl[8] br[8] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_11 
+ bl[9] br[9] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_12 
+ bl[10] br[10] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_13 
+ bl[11] br[11] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_14 
+ bl[12] br[12] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_15 
+ bl[13] br[13] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_16 
+ bl[14] br[14] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_17 
+ bl[15] br[15] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_18 
+ bl[16] br[16] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_19 
+ bl[17] br[17] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_20 
+ bl[18] br[18] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_21 
+ bl[19] br[19] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_22 
+ bl[20] br[20] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_23 
+ bl[21] br[21] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_24 
+ bl[22] br[22] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_25 
+ bl[23] br[23] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_26 
+ bl[24] br[24] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_27 
+ bl[25] br[25] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_28 
+ bl[26] br[26] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_29 
+ bl[27] br[27] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_30 
+ bl[28] br[28] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_31 
+ bl[29] br[29] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_32 
+ bl[30] br[30] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_33 
+ bl[31] br[31] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_34 
+ bl[32] br[32] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_35 
+ bl[33] br[33] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_36 
+ bl[34] br[34] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_37 
+ bl[35] br[35] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_38 
+ bl[36] br[36] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_39 
+ bl[37] br[37] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_40 
+ bl[38] br[38] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_41 
+ bl[39] br[39] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_42 
+ bl[40] br[40] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_43 
+ bl[41] br[41] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_44 
+ bl[42] br[42] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_45 
+ bl[43] br[43] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_46 
+ bl[44] br[44] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_47 
+ bl[45] br[45] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_48 
+ bl[46] br[46] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_49 
+ bl[47] br[47] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_50 
+ bl[48] br[48] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_51 
+ bl[49] br[49] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_52 
+ bl[50] br[50] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_53 
+ bl[51] br[51] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_54 
+ bl[52] br[52] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_55 
+ bl[53] br[53] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_56 
+ bl[54] br[54] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_57 
+ bl[55] br[55] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_58 
+ bl[56] br[56] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_59 
+ bl[57] br[57] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_60 
+ bl[58] br[58] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_61 
+ bl[59] br[59] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_62 
+ bl[60] br[60] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_63 
+ bl[61] br[61] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_64 
+ bl[62] br[62] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_65 
+ bl[63] br[63] vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_66 
+ vdd vdd vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_261_67 
+ vdd vdd vdd vss wl[259] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_0 
+ vdd vdd vss vdd vpb vnb wl[260] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_262_1 
+ rbl rbr vss vdd vpb vnb wl[260] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_262_2 
+ bl[0] br[0] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_3 
+ bl[1] br[1] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_4 
+ bl[2] br[2] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_5 
+ bl[3] br[3] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_6 
+ bl[4] br[4] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_7 
+ bl[5] br[5] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_8 
+ bl[6] br[6] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_9 
+ bl[7] br[7] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_10 
+ bl[8] br[8] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_11 
+ bl[9] br[9] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_12 
+ bl[10] br[10] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_13 
+ bl[11] br[11] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_14 
+ bl[12] br[12] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_15 
+ bl[13] br[13] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_16 
+ bl[14] br[14] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_17 
+ bl[15] br[15] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_18 
+ bl[16] br[16] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_19 
+ bl[17] br[17] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_20 
+ bl[18] br[18] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_21 
+ bl[19] br[19] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_22 
+ bl[20] br[20] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_23 
+ bl[21] br[21] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_24 
+ bl[22] br[22] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_25 
+ bl[23] br[23] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_26 
+ bl[24] br[24] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_27 
+ bl[25] br[25] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_28 
+ bl[26] br[26] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_29 
+ bl[27] br[27] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_30 
+ bl[28] br[28] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_31 
+ bl[29] br[29] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_32 
+ bl[30] br[30] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_33 
+ bl[31] br[31] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_34 
+ bl[32] br[32] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_35 
+ bl[33] br[33] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_36 
+ bl[34] br[34] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_37 
+ bl[35] br[35] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_38 
+ bl[36] br[36] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_39 
+ bl[37] br[37] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_40 
+ bl[38] br[38] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_41 
+ bl[39] br[39] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_42 
+ bl[40] br[40] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_43 
+ bl[41] br[41] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_44 
+ bl[42] br[42] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_45 
+ bl[43] br[43] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_46 
+ bl[44] br[44] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_47 
+ bl[45] br[45] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_48 
+ bl[46] br[46] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_49 
+ bl[47] br[47] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_50 
+ bl[48] br[48] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_51 
+ bl[49] br[49] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_52 
+ bl[50] br[50] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_53 
+ bl[51] br[51] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_54 
+ bl[52] br[52] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_55 
+ bl[53] br[53] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_56 
+ bl[54] br[54] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_57 
+ bl[55] br[55] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_58 
+ bl[56] br[56] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_59 
+ bl[57] br[57] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_60 
+ bl[58] br[58] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_61 
+ bl[59] br[59] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_62 
+ bl[60] br[60] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_63 
+ bl[61] br[61] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_64 
+ bl[62] br[62] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_65 
+ bl[63] br[63] vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_66 
+ vdd vdd vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_262_67 
+ vdd vdd vdd vss wl[260] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_0 
+ vdd vdd vss vdd vpb vnb wl[261] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_263_1 
+ rbl rbr vss vdd vpb vnb wl[261] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_263_2 
+ bl[0] br[0] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_3 
+ bl[1] br[1] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_4 
+ bl[2] br[2] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_5 
+ bl[3] br[3] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_6 
+ bl[4] br[4] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_7 
+ bl[5] br[5] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_8 
+ bl[6] br[6] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_9 
+ bl[7] br[7] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_10 
+ bl[8] br[8] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_11 
+ bl[9] br[9] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_12 
+ bl[10] br[10] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_13 
+ bl[11] br[11] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_14 
+ bl[12] br[12] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_15 
+ bl[13] br[13] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_16 
+ bl[14] br[14] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_17 
+ bl[15] br[15] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_18 
+ bl[16] br[16] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_19 
+ bl[17] br[17] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_20 
+ bl[18] br[18] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_21 
+ bl[19] br[19] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_22 
+ bl[20] br[20] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_23 
+ bl[21] br[21] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_24 
+ bl[22] br[22] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_25 
+ bl[23] br[23] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_26 
+ bl[24] br[24] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_27 
+ bl[25] br[25] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_28 
+ bl[26] br[26] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_29 
+ bl[27] br[27] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_30 
+ bl[28] br[28] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_31 
+ bl[29] br[29] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_32 
+ bl[30] br[30] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_33 
+ bl[31] br[31] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_34 
+ bl[32] br[32] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_35 
+ bl[33] br[33] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_36 
+ bl[34] br[34] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_37 
+ bl[35] br[35] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_38 
+ bl[36] br[36] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_39 
+ bl[37] br[37] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_40 
+ bl[38] br[38] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_41 
+ bl[39] br[39] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_42 
+ bl[40] br[40] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_43 
+ bl[41] br[41] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_44 
+ bl[42] br[42] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_45 
+ bl[43] br[43] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_46 
+ bl[44] br[44] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_47 
+ bl[45] br[45] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_48 
+ bl[46] br[46] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_49 
+ bl[47] br[47] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_50 
+ bl[48] br[48] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_51 
+ bl[49] br[49] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_52 
+ bl[50] br[50] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_53 
+ bl[51] br[51] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_54 
+ bl[52] br[52] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_55 
+ bl[53] br[53] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_56 
+ bl[54] br[54] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_57 
+ bl[55] br[55] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_58 
+ bl[56] br[56] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_59 
+ bl[57] br[57] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_60 
+ bl[58] br[58] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_61 
+ bl[59] br[59] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_62 
+ bl[60] br[60] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_63 
+ bl[61] br[61] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_64 
+ bl[62] br[62] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_65 
+ bl[63] br[63] vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_66 
+ vdd vdd vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_263_67 
+ vdd vdd vdd vss wl[261] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_0 
+ vdd vdd vss vdd vpb vnb wl[262] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_264_1 
+ rbl rbr vss vdd vpb vnb wl[262] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_264_2 
+ bl[0] br[0] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_3 
+ bl[1] br[1] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_4 
+ bl[2] br[2] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_5 
+ bl[3] br[3] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_6 
+ bl[4] br[4] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_7 
+ bl[5] br[5] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_8 
+ bl[6] br[6] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_9 
+ bl[7] br[7] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_10 
+ bl[8] br[8] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_11 
+ bl[9] br[9] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_12 
+ bl[10] br[10] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_13 
+ bl[11] br[11] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_14 
+ bl[12] br[12] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_15 
+ bl[13] br[13] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_16 
+ bl[14] br[14] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_17 
+ bl[15] br[15] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_18 
+ bl[16] br[16] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_19 
+ bl[17] br[17] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_20 
+ bl[18] br[18] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_21 
+ bl[19] br[19] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_22 
+ bl[20] br[20] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_23 
+ bl[21] br[21] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_24 
+ bl[22] br[22] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_25 
+ bl[23] br[23] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_26 
+ bl[24] br[24] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_27 
+ bl[25] br[25] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_28 
+ bl[26] br[26] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_29 
+ bl[27] br[27] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_30 
+ bl[28] br[28] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_31 
+ bl[29] br[29] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_32 
+ bl[30] br[30] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_33 
+ bl[31] br[31] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_34 
+ bl[32] br[32] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_35 
+ bl[33] br[33] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_36 
+ bl[34] br[34] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_37 
+ bl[35] br[35] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_38 
+ bl[36] br[36] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_39 
+ bl[37] br[37] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_40 
+ bl[38] br[38] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_41 
+ bl[39] br[39] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_42 
+ bl[40] br[40] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_43 
+ bl[41] br[41] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_44 
+ bl[42] br[42] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_45 
+ bl[43] br[43] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_46 
+ bl[44] br[44] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_47 
+ bl[45] br[45] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_48 
+ bl[46] br[46] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_49 
+ bl[47] br[47] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_50 
+ bl[48] br[48] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_51 
+ bl[49] br[49] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_52 
+ bl[50] br[50] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_53 
+ bl[51] br[51] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_54 
+ bl[52] br[52] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_55 
+ bl[53] br[53] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_56 
+ bl[54] br[54] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_57 
+ bl[55] br[55] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_58 
+ bl[56] br[56] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_59 
+ bl[57] br[57] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_60 
+ bl[58] br[58] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_61 
+ bl[59] br[59] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_62 
+ bl[60] br[60] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_63 
+ bl[61] br[61] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_64 
+ bl[62] br[62] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_65 
+ bl[63] br[63] vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_66 
+ vdd vdd vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_264_67 
+ vdd vdd vdd vss wl[262] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_0 
+ vdd vdd vss vdd vpb vnb wl[263] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_265_1 
+ rbl rbr vss vdd vpb vnb wl[263] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_265_2 
+ bl[0] br[0] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_3 
+ bl[1] br[1] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_4 
+ bl[2] br[2] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_5 
+ bl[3] br[3] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_6 
+ bl[4] br[4] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_7 
+ bl[5] br[5] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_8 
+ bl[6] br[6] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_9 
+ bl[7] br[7] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_10 
+ bl[8] br[8] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_11 
+ bl[9] br[9] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_12 
+ bl[10] br[10] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_13 
+ bl[11] br[11] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_14 
+ bl[12] br[12] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_15 
+ bl[13] br[13] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_16 
+ bl[14] br[14] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_17 
+ bl[15] br[15] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_18 
+ bl[16] br[16] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_19 
+ bl[17] br[17] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_20 
+ bl[18] br[18] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_21 
+ bl[19] br[19] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_22 
+ bl[20] br[20] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_23 
+ bl[21] br[21] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_24 
+ bl[22] br[22] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_25 
+ bl[23] br[23] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_26 
+ bl[24] br[24] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_27 
+ bl[25] br[25] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_28 
+ bl[26] br[26] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_29 
+ bl[27] br[27] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_30 
+ bl[28] br[28] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_31 
+ bl[29] br[29] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_32 
+ bl[30] br[30] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_33 
+ bl[31] br[31] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_34 
+ bl[32] br[32] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_35 
+ bl[33] br[33] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_36 
+ bl[34] br[34] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_37 
+ bl[35] br[35] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_38 
+ bl[36] br[36] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_39 
+ bl[37] br[37] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_40 
+ bl[38] br[38] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_41 
+ bl[39] br[39] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_42 
+ bl[40] br[40] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_43 
+ bl[41] br[41] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_44 
+ bl[42] br[42] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_45 
+ bl[43] br[43] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_46 
+ bl[44] br[44] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_47 
+ bl[45] br[45] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_48 
+ bl[46] br[46] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_49 
+ bl[47] br[47] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_50 
+ bl[48] br[48] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_51 
+ bl[49] br[49] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_52 
+ bl[50] br[50] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_53 
+ bl[51] br[51] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_54 
+ bl[52] br[52] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_55 
+ bl[53] br[53] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_56 
+ bl[54] br[54] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_57 
+ bl[55] br[55] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_58 
+ bl[56] br[56] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_59 
+ bl[57] br[57] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_60 
+ bl[58] br[58] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_61 
+ bl[59] br[59] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_62 
+ bl[60] br[60] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_63 
+ bl[61] br[61] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_64 
+ bl[62] br[62] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_65 
+ bl[63] br[63] vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_66 
+ vdd vdd vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_265_67 
+ vdd vdd vdd vss wl[263] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_0 
+ vdd vdd vss vdd vpb vnb wl[264] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_266_1 
+ rbl rbr vss vdd vpb vnb wl[264] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_266_2 
+ bl[0] br[0] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_3 
+ bl[1] br[1] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_4 
+ bl[2] br[2] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_5 
+ bl[3] br[3] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_6 
+ bl[4] br[4] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_7 
+ bl[5] br[5] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_8 
+ bl[6] br[6] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_9 
+ bl[7] br[7] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_10 
+ bl[8] br[8] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_11 
+ bl[9] br[9] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_12 
+ bl[10] br[10] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_13 
+ bl[11] br[11] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_14 
+ bl[12] br[12] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_15 
+ bl[13] br[13] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_16 
+ bl[14] br[14] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_17 
+ bl[15] br[15] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_18 
+ bl[16] br[16] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_19 
+ bl[17] br[17] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_20 
+ bl[18] br[18] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_21 
+ bl[19] br[19] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_22 
+ bl[20] br[20] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_23 
+ bl[21] br[21] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_24 
+ bl[22] br[22] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_25 
+ bl[23] br[23] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_26 
+ bl[24] br[24] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_27 
+ bl[25] br[25] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_28 
+ bl[26] br[26] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_29 
+ bl[27] br[27] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_30 
+ bl[28] br[28] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_31 
+ bl[29] br[29] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_32 
+ bl[30] br[30] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_33 
+ bl[31] br[31] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_34 
+ bl[32] br[32] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_35 
+ bl[33] br[33] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_36 
+ bl[34] br[34] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_37 
+ bl[35] br[35] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_38 
+ bl[36] br[36] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_39 
+ bl[37] br[37] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_40 
+ bl[38] br[38] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_41 
+ bl[39] br[39] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_42 
+ bl[40] br[40] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_43 
+ bl[41] br[41] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_44 
+ bl[42] br[42] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_45 
+ bl[43] br[43] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_46 
+ bl[44] br[44] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_47 
+ bl[45] br[45] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_48 
+ bl[46] br[46] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_49 
+ bl[47] br[47] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_50 
+ bl[48] br[48] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_51 
+ bl[49] br[49] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_52 
+ bl[50] br[50] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_53 
+ bl[51] br[51] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_54 
+ bl[52] br[52] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_55 
+ bl[53] br[53] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_56 
+ bl[54] br[54] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_57 
+ bl[55] br[55] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_58 
+ bl[56] br[56] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_59 
+ bl[57] br[57] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_60 
+ bl[58] br[58] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_61 
+ bl[59] br[59] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_62 
+ bl[60] br[60] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_63 
+ bl[61] br[61] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_64 
+ bl[62] br[62] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_65 
+ bl[63] br[63] vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_66 
+ vdd vdd vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_266_67 
+ vdd vdd vdd vss wl[264] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_0 
+ vdd vdd vss vdd vpb vnb wl[265] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_267_1 
+ rbl rbr vss vdd vpb vnb wl[265] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_267_2 
+ bl[0] br[0] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_3 
+ bl[1] br[1] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_4 
+ bl[2] br[2] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_5 
+ bl[3] br[3] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_6 
+ bl[4] br[4] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_7 
+ bl[5] br[5] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_8 
+ bl[6] br[6] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_9 
+ bl[7] br[7] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_10 
+ bl[8] br[8] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_11 
+ bl[9] br[9] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_12 
+ bl[10] br[10] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_13 
+ bl[11] br[11] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_14 
+ bl[12] br[12] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_15 
+ bl[13] br[13] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_16 
+ bl[14] br[14] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_17 
+ bl[15] br[15] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_18 
+ bl[16] br[16] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_19 
+ bl[17] br[17] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_20 
+ bl[18] br[18] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_21 
+ bl[19] br[19] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_22 
+ bl[20] br[20] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_23 
+ bl[21] br[21] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_24 
+ bl[22] br[22] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_25 
+ bl[23] br[23] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_26 
+ bl[24] br[24] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_27 
+ bl[25] br[25] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_28 
+ bl[26] br[26] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_29 
+ bl[27] br[27] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_30 
+ bl[28] br[28] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_31 
+ bl[29] br[29] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_32 
+ bl[30] br[30] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_33 
+ bl[31] br[31] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_34 
+ bl[32] br[32] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_35 
+ bl[33] br[33] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_36 
+ bl[34] br[34] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_37 
+ bl[35] br[35] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_38 
+ bl[36] br[36] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_39 
+ bl[37] br[37] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_40 
+ bl[38] br[38] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_41 
+ bl[39] br[39] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_42 
+ bl[40] br[40] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_43 
+ bl[41] br[41] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_44 
+ bl[42] br[42] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_45 
+ bl[43] br[43] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_46 
+ bl[44] br[44] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_47 
+ bl[45] br[45] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_48 
+ bl[46] br[46] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_49 
+ bl[47] br[47] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_50 
+ bl[48] br[48] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_51 
+ bl[49] br[49] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_52 
+ bl[50] br[50] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_53 
+ bl[51] br[51] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_54 
+ bl[52] br[52] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_55 
+ bl[53] br[53] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_56 
+ bl[54] br[54] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_57 
+ bl[55] br[55] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_58 
+ bl[56] br[56] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_59 
+ bl[57] br[57] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_60 
+ bl[58] br[58] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_61 
+ bl[59] br[59] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_62 
+ bl[60] br[60] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_63 
+ bl[61] br[61] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_64 
+ bl[62] br[62] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_65 
+ bl[63] br[63] vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_66 
+ vdd vdd vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_267_67 
+ vdd vdd vdd vss wl[265] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_0 
+ vdd vdd vss vdd vpb vnb wl[266] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_268_1 
+ rbl rbr vss vdd vpb vnb wl[266] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_268_2 
+ bl[0] br[0] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_3 
+ bl[1] br[1] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_4 
+ bl[2] br[2] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_5 
+ bl[3] br[3] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_6 
+ bl[4] br[4] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_7 
+ bl[5] br[5] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_8 
+ bl[6] br[6] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_9 
+ bl[7] br[7] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_10 
+ bl[8] br[8] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_11 
+ bl[9] br[9] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_12 
+ bl[10] br[10] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_13 
+ bl[11] br[11] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_14 
+ bl[12] br[12] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_15 
+ bl[13] br[13] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_16 
+ bl[14] br[14] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_17 
+ bl[15] br[15] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_18 
+ bl[16] br[16] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_19 
+ bl[17] br[17] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_20 
+ bl[18] br[18] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_21 
+ bl[19] br[19] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_22 
+ bl[20] br[20] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_23 
+ bl[21] br[21] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_24 
+ bl[22] br[22] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_25 
+ bl[23] br[23] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_26 
+ bl[24] br[24] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_27 
+ bl[25] br[25] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_28 
+ bl[26] br[26] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_29 
+ bl[27] br[27] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_30 
+ bl[28] br[28] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_31 
+ bl[29] br[29] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_32 
+ bl[30] br[30] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_33 
+ bl[31] br[31] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_34 
+ bl[32] br[32] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_35 
+ bl[33] br[33] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_36 
+ bl[34] br[34] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_37 
+ bl[35] br[35] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_38 
+ bl[36] br[36] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_39 
+ bl[37] br[37] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_40 
+ bl[38] br[38] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_41 
+ bl[39] br[39] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_42 
+ bl[40] br[40] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_43 
+ bl[41] br[41] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_44 
+ bl[42] br[42] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_45 
+ bl[43] br[43] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_46 
+ bl[44] br[44] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_47 
+ bl[45] br[45] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_48 
+ bl[46] br[46] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_49 
+ bl[47] br[47] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_50 
+ bl[48] br[48] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_51 
+ bl[49] br[49] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_52 
+ bl[50] br[50] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_53 
+ bl[51] br[51] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_54 
+ bl[52] br[52] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_55 
+ bl[53] br[53] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_56 
+ bl[54] br[54] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_57 
+ bl[55] br[55] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_58 
+ bl[56] br[56] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_59 
+ bl[57] br[57] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_60 
+ bl[58] br[58] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_61 
+ bl[59] br[59] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_62 
+ bl[60] br[60] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_63 
+ bl[61] br[61] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_64 
+ bl[62] br[62] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_65 
+ bl[63] br[63] vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_66 
+ vdd vdd vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_268_67 
+ vdd vdd vdd vss wl[266] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_0 
+ vdd vdd vss vdd vpb vnb wl[267] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_269_1 
+ rbl rbr vss vdd vpb vnb wl[267] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_269_2 
+ bl[0] br[0] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_3 
+ bl[1] br[1] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_4 
+ bl[2] br[2] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_5 
+ bl[3] br[3] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_6 
+ bl[4] br[4] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_7 
+ bl[5] br[5] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_8 
+ bl[6] br[6] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_9 
+ bl[7] br[7] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_10 
+ bl[8] br[8] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_11 
+ bl[9] br[9] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_12 
+ bl[10] br[10] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_13 
+ bl[11] br[11] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_14 
+ bl[12] br[12] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_15 
+ bl[13] br[13] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_16 
+ bl[14] br[14] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_17 
+ bl[15] br[15] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_18 
+ bl[16] br[16] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_19 
+ bl[17] br[17] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_20 
+ bl[18] br[18] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_21 
+ bl[19] br[19] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_22 
+ bl[20] br[20] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_23 
+ bl[21] br[21] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_24 
+ bl[22] br[22] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_25 
+ bl[23] br[23] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_26 
+ bl[24] br[24] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_27 
+ bl[25] br[25] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_28 
+ bl[26] br[26] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_29 
+ bl[27] br[27] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_30 
+ bl[28] br[28] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_31 
+ bl[29] br[29] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_32 
+ bl[30] br[30] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_33 
+ bl[31] br[31] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_34 
+ bl[32] br[32] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_35 
+ bl[33] br[33] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_36 
+ bl[34] br[34] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_37 
+ bl[35] br[35] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_38 
+ bl[36] br[36] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_39 
+ bl[37] br[37] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_40 
+ bl[38] br[38] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_41 
+ bl[39] br[39] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_42 
+ bl[40] br[40] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_43 
+ bl[41] br[41] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_44 
+ bl[42] br[42] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_45 
+ bl[43] br[43] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_46 
+ bl[44] br[44] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_47 
+ bl[45] br[45] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_48 
+ bl[46] br[46] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_49 
+ bl[47] br[47] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_50 
+ bl[48] br[48] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_51 
+ bl[49] br[49] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_52 
+ bl[50] br[50] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_53 
+ bl[51] br[51] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_54 
+ bl[52] br[52] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_55 
+ bl[53] br[53] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_56 
+ bl[54] br[54] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_57 
+ bl[55] br[55] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_58 
+ bl[56] br[56] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_59 
+ bl[57] br[57] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_60 
+ bl[58] br[58] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_61 
+ bl[59] br[59] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_62 
+ bl[60] br[60] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_63 
+ bl[61] br[61] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_64 
+ bl[62] br[62] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_65 
+ bl[63] br[63] vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_66 
+ vdd vdd vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_269_67 
+ vdd vdd vdd vss wl[267] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_0 
+ vdd vdd vss vdd vpb vnb wl[268] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_270_1 
+ rbl rbr vss vdd vpb vnb wl[268] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_270_2 
+ bl[0] br[0] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_3 
+ bl[1] br[1] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_4 
+ bl[2] br[2] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_5 
+ bl[3] br[3] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_6 
+ bl[4] br[4] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_7 
+ bl[5] br[5] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_8 
+ bl[6] br[6] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_9 
+ bl[7] br[7] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_10 
+ bl[8] br[8] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_11 
+ bl[9] br[9] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_12 
+ bl[10] br[10] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_13 
+ bl[11] br[11] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_14 
+ bl[12] br[12] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_15 
+ bl[13] br[13] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_16 
+ bl[14] br[14] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_17 
+ bl[15] br[15] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_18 
+ bl[16] br[16] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_19 
+ bl[17] br[17] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_20 
+ bl[18] br[18] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_21 
+ bl[19] br[19] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_22 
+ bl[20] br[20] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_23 
+ bl[21] br[21] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_24 
+ bl[22] br[22] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_25 
+ bl[23] br[23] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_26 
+ bl[24] br[24] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_27 
+ bl[25] br[25] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_28 
+ bl[26] br[26] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_29 
+ bl[27] br[27] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_30 
+ bl[28] br[28] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_31 
+ bl[29] br[29] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_32 
+ bl[30] br[30] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_33 
+ bl[31] br[31] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_34 
+ bl[32] br[32] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_35 
+ bl[33] br[33] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_36 
+ bl[34] br[34] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_37 
+ bl[35] br[35] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_38 
+ bl[36] br[36] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_39 
+ bl[37] br[37] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_40 
+ bl[38] br[38] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_41 
+ bl[39] br[39] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_42 
+ bl[40] br[40] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_43 
+ bl[41] br[41] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_44 
+ bl[42] br[42] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_45 
+ bl[43] br[43] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_46 
+ bl[44] br[44] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_47 
+ bl[45] br[45] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_48 
+ bl[46] br[46] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_49 
+ bl[47] br[47] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_50 
+ bl[48] br[48] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_51 
+ bl[49] br[49] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_52 
+ bl[50] br[50] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_53 
+ bl[51] br[51] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_54 
+ bl[52] br[52] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_55 
+ bl[53] br[53] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_56 
+ bl[54] br[54] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_57 
+ bl[55] br[55] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_58 
+ bl[56] br[56] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_59 
+ bl[57] br[57] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_60 
+ bl[58] br[58] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_61 
+ bl[59] br[59] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_62 
+ bl[60] br[60] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_63 
+ bl[61] br[61] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_64 
+ bl[62] br[62] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_65 
+ bl[63] br[63] vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_66 
+ vdd vdd vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_270_67 
+ vdd vdd vdd vss wl[268] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_0 
+ vdd vdd vss vdd vpb vnb wl[269] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_271_1 
+ rbl rbr vss vdd vpb vnb wl[269] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_271_2 
+ bl[0] br[0] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_3 
+ bl[1] br[1] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_4 
+ bl[2] br[2] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_5 
+ bl[3] br[3] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_6 
+ bl[4] br[4] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_7 
+ bl[5] br[5] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_8 
+ bl[6] br[6] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_9 
+ bl[7] br[7] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_10 
+ bl[8] br[8] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_11 
+ bl[9] br[9] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_12 
+ bl[10] br[10] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_13 
+ bl[11] br[11] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_14 
+ bl[12] br[12] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_15 
+ bl[13] br[13] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_16 
+ bl[14] br[14] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_17 
+ bl[15] br[15] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_18 
+ bl[16] br[16] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_19 
+ bl[17] br[17] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_20 
+ bl[18] br[18] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_21 
+ bl[19] br[19] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_22 
+ bl[20] br[20] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_23 
+ bl[21] br[21] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_24 
+ bl[22] br[22] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_25 
+ bl[23] br[23] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_26 
+ bl[24] br[24] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_27 
+ bl[25] br[25] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_28 
+ bl[26] br[26] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_29 
+ bl[27] br[27] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_30 
+ bl[28] br[28] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_31 
+ bl[29] br[29] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_32 
+ bl[30] br[30] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_33 
+ bl[31] br[31] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_34 
+ bl[32] br[32] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_35 
+ bl[33] br[33] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_36 
+ bl[34] br[34] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_37 
+ bl[35] br[35] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_38 
+ bl[36] br[36] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_39 
+ bl[37] br[37] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_40 
+ bl[38] br[38] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_41 
+ bl[39] br[39] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_42 
+ bl[40] br[40] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_43 
+ bl[41] br[41] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_44 
+ bl[42] br[42] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_45 
+ bl[43] br[43] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_46 
+ bl[44] br[44] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_47 
+ bl[45] br[45] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_48 
+ bl[46] br[46] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_49 
+ bl[47] br[47] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_50 
+ bl[48] br[48] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_51 
+ bl[49] br[49] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_52 
+ bl[50] br[50] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_53 
+ bl[51] br[51] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_54 
+ bl[52] br[52] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_55 
+ bl[53] br[53] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_56 
+ bl[54] br[54] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_57 
+ bl[55] br[55] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_58 
+ bl[56] br[56] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_59 
+ bl[57] br[57] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_60 
+ bl[58] br[58] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_61 
+ bl[59] br[59] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_62 
+ bl[60] br[60] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_63 
+ bl[61] br[61] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_64 
+ bl[62] br[62] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_65 
+ bl[63] br[63] vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_66 
+ vdd vdd vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_271_67 
+ vdd vdd vdd vss wl[269] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_0 
+ vdd vdd vss vdd vpb vnb wl[270] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_272_1 
+ rbl rbr vss vdd vpb vnb wl[270] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_272_2 
+ bl[0] br[0] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_3 
+ bl[1] br[1] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_4 
+ bl[2] br[2] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_5 
+ bl[3] br[3] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_6 
+ bl[4] br[4] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_7 
+ bl[5] br[5] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_8 
+ bl[6] br[6] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_9 
+ bl[7] br[7] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_10 
+ bl[8] br[8] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_11 
+ bl[9] br[9] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_12 
+ bl[10] br[10] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_13 
+ bl[11] br[11] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_14 
+ bl[12] br[12] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_15 
+ bl[13] br[13] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_16 
+ bl[14] br[14] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_17 
+ bl[15] br[15] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_18 
+ bl[16] br[16] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_19 
+ bl[17] br[17] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_20 
+ bl[18] br[18] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_21 
+ bl[19] br[19] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_22 
+ bl[20] br[20] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_23 
+ bl[21] br[21] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_24 
+ bl[22] br[22] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_25 
+ bl[23] br[23] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_26 
+ bl[24] br[24] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_27 
+ bl[25] br[25] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_28 
+ bl[26] br[26] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_29 
+ bl[27] br[27] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_30 
+ bl[28] br[28] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_31 
+ bl[29] br[29] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_32 
+ bl[30] br[30] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_33 
+ bl[31] br[31] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_34 
+ bl[32] br[32] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_35 
+ bl[33] br[33] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_36 
+ bl[34] br[34] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_37 
+ bl[35] br[35] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_38 
+ bl[36] br[36] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_39 
+ bl[37] br[37] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_40 
+ bl[38] br[38] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_41 
+ bl[39] br[39] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_42 
+ bl[40] br[40] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_43 
+ bl[41] br[41] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_44 
+ bl[42] br[42] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_45 
+ bl[43] br[43] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_46 
+ bl[44] br[44] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_47 
+ bl[45] br[45] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_48 
+ bl[46] br[46] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_49 
+ bl[47] br[47] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_50 
+ bl[48] br[48] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_51 
+ bl[49] br[49] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_52 
+ bl[50] br[50] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_53 
+ bl[51] br[51] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_54 
+ bl[52] br[52] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_55 
+ bl[53] br[53] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_56 
+ bl[54] br[54] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_57 
+ bl[55] br[55] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_58 
+ bl[56] br[56] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_59 
+ bl[57] br[57] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_60 
+ bl[58] br[58] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_61 
+ bl[59] br[59] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_62 
+ bl[60] br[60] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_63 
+ bl[61] br[61] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_64 
+ bl[62] br[62] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_65 
+ bl[63] br[63] vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_66 
+ vdd vdd vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_272_67 
+ vdd vdd vdd vss wl[270] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_0 
+ vdd vdd vss vdd vpb vnb wl[271] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_273_1 
+ rbl rbr vss vdd vpb vnb wl[271] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_273_2 
+ bl[0] br[0] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_3 
+ bl[1] br[1] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_4 
+ bl[2] br[2] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_5 
+ bl[3] br[3] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_6 
+ bl[4] br[4] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_7 
+ bl[5] br[5] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_8 
+ bl[6] br[6] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_9 
+ bl[7] br[7] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_10 
+ bl[8] br[8] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_11 
+ bl[9] br[9] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_12 
+ bl[10] br[10] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_13 
+ bl[11] br[11] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_14 
+ bl[12] br[12] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_15 
+ bl[13] br[13] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_16 
+ bl[14] br[14] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_17 
+ bl[15] br[15] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_18 
+ bl[16] br[16] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_19 
+ bl[17] br[17] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_20 
+ bl[18] br[18] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_21 
+ bl[19] br[19] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_22 
+ bl[20] br[20] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_23 
+ bl[21] br[21] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_24 
+ bl[22] br[22] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_25 
+ bl[23] br[23] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_26 
+ bl[24] br[24] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_27 
+ bl[25] br[25] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_28 
+ bl[26] br[26] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_29 
+ bl[27] br[27] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_30 
+ bl[28] br[28] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_31 
+ bl[29] br[29] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_32 
+ bl[30] br[30] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_33 
+ bl[31] br[31] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_34 
+ bl[32] br[32] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_35 
+ bl[33] br[33] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_36 
+ bl[34] br[34] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_37 
+ bl[35] br[35] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_38 
+ bl[36] br[36] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_39 
+ bl[37] br[37] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_40 
+ bl[38] br[38] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_41 
+ bl[39] br[39] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_42 
+ bl[40] br[40] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_43 
+ bl[41] br[41] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_44 
+ bl[42] br[42] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_45 
+ bl[43] br[43] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_46 
+ bl[44] br[44] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_47 
+ bl[45] br[45] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_48 
+ bl[46] br[46] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_49 
+ bl[47] br[47] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_50 
+ bl[48] br[48] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_51 
+ bl[49] br[49] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_52 
+ bl[50] br[50] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_53 
+ bl[51] br[51] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_54 
+ bl[52] br[52] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_55 
+ bl[53] br[53] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_56 
+ bl[54] br[54] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_57 
+ bl[55] br[55] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_58 
+ bl[56] br[56] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_59 
+ bl[57] br[57] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_60 
+ bl[58] br[58] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_61 
+ bl[59] br[59] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_62 
+ bl[60] br[60] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_63 
+ bl[61] br[61] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_64 
+ bl[62] br[62] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_65 
+ bl[63] br[63] vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_66 
+ vdd vdd vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_273_67 
+ vdd vdd vdd vss wl[271] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_0 
+ vdd vdd vss vdd vpb vnb wl[272] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_274_1 
+ rbl rbr vss vdd vpb vnb wl[272] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_274_2 
+ bl[0] br[0] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_3 
+ bl[1] br[1] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_4 
+ bl[2] br[2] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_5 
+ bl[3] br[3] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_6 
+ bl[4] br[4] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_7 
+ bl[5] br[5] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_8 
+ bl[6] br[6] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_9 
+ bl[7] br[7] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_10 
+ bl[8] br[8] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_11 
+ bl[9] br[9] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_12 
+ bl[10] br[10] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_13 
+ bl[11] br[11] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_14 
+ bl[12] br[12] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_15 
+ bl[13] br[13] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_16 
+ bl[14] br[14] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_17 
+ bl[15] br[15] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_18 
+ bl[16] br[16] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_19 
+ bl[17] br[17] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_20 
+ bl[18] br[18] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_21 
+ bl[19] br[19] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_22 
+ bl[20] br[20] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_23 
+ bl[21] br[21] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_24 
+ bl[22] br[22] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_25 
+ bl[23] br[23] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_26 
+ bl[24] br[24] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_27 
+ bl[25] br[25] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_28 
+ bl[26] br[26] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_29 
+ bl[27] br[27] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_30 
+ bl[28] br[28] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_31 
+ bl[29] br[29] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_32 
+ bl[30] br[30] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_33 
+ bl[31] br[31] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_34 
+ bl[32] br[32] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_35 
+ bl[33] br[33] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_36 
+ bl[34] br[34] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_37 
+ bl[35] br[35] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_38 
+ bl[36] br[36] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_39 
+ bl[37] br[37] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_40 
+ bl[38] br[38] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_41 
+ bl[39] br[39] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_42 
+ bl[40] br[40] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_43 
+ bl[41] br[41] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_44 
+ bl[42] br[42] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_45 
+ bl[43] br[43] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_46 
+ bl[44] br[44] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_47 
+ bl[45] br[45] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_48 
+ bl[46] br[46] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_49 
+ bl[47] br[47] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_50 
+ bl[48] br[48] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_51 
+ bl[49] br[49] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_52 
+ bl[50] br[50] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_53 
+ bl[51] br[51] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_54 
+ bl[52] br[52] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_55 
+ bl[53] br[53] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_56 
+ bl[54] br[54] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_57 
+ bl[55] br[55] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_58 
+ bl[56] br[56] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_59 
+ bl[57] br[57] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_60 
+ bl[58] br[58] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_61 
+ bl[59] br[59] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_62 
+ bl[60] br[60] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_63 
+ bl[61] br[61] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_64 
+ bl[62] br[62] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_65 
+ bl[63] br[63] vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_66 
+ vdd vdd vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_274_67 
+ vdd vdd vdd vss wl[272] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_0 
+ vdd vdd vss vdd vpb vnb wl[273] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_275_1 
+ rbl rbr vss vdd vpb vnb wl[273] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_275_2 
+ bl[0] br[0] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_3 
+ bl[1] br[1] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_4 
+ bl[2] br[2] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_5 
+ bl[3] br[3] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_6 
+ bl[4] br[4] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_7 
+ bl[5] br[5] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_8 
+ bl[6] br[6] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_9 
+ bl[7] br[7] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_10 
+ bl[8] br[8] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_11 
+ bl[9] br[9] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_12 
+ bl[10] br[10] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_13 
+ bl[11] br[11] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_14 
+ bl[12] br[12] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_15 
+ bl[13] br[13] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_16 
+ bl[14] br[14] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_17 
+ bl[15] br[15] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_18 
+ bl[16] br[16] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_19 
+ bl[17] br[17] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_20 
+ bl[18] br[18] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_21 
+ bl[19] br[19] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_22 
+ bl[20] br[20] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_23 
+ bl[21] br[21] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_24 
+ bl[22] br[22] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_25 
+ bl[23] br[23] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_26 
+ bl[24] br[24] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_27 
+ bl[25] br[25] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_28 
+ bl[26] br[26] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_29 
+ bl[27] br[27] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_30 
+ bl[28] br[28] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_31 
+ bl[29] br[29] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_32 
+ bl[30] br[30] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_33 
+ bl[31] br[31] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_34 
+ bl[32] br[32] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_35 
+ bl[33] br[33] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_36 
+ bl[34] br[34] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_37 
+ bl[35] br[35] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_38 
+ bl[36] br[36] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_39 
+ bl[37] br[37] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_40 
+ bl[38] br[38] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_41 
+ bl[39] br[39] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_42 
+ bl[40] br[40] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_43 
+ bl[41] br[41] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_44 
+ bl[42] br[42] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_45 
+ bl[43] br[43] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_46 
+ bl[44] br[44] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_47 
+ bl[45] br[45] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_48 
+ bl[46] br[46] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_49 
+ bl[47] br[47] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_50 
+ bl[48] br[48] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_51 
+ bl[49] br[49] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_52 
+ bl[50] br[50] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_53 
+ bl[51] br[51] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_54 
+ bl[52] br[52] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_55 
+ bl[53] br[53] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_56 
+ bl[54] br[54] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_57 
+ bl[55] br[55] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_58 
+ bl[56] br[56] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_59 
+ bl[57] br[57] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_60 
+ bl[58] br[58] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_61 
+ bl[59] br[59] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_62 
+ bl[60] br[60] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_63 
+ bl[61] br[61] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_64 
+ bl[62] br[62] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_65 
+ bl[63] br[63] vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_66 
+ vdd vdd vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_275_67 
+ vdd vdd vdd vss wl[273] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_0 
+ vdd vdd vss vdd vpb vnb wl[274] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_276_1 
+ rbl rbr vss vdd vpb vnb wl[274] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_276_2 
+ bl[0] br[0] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_3 
+ bl[1] br[1] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_4 
+ bl[2] br[2] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_5 
+ bl[3] br[3] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_6 
+ bl[4] br[4] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_7 
+ bl[5] br[5] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_8 
+ bl[6] br[6] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_9 
+ bl[7] br[7] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_10 
+ bl[8] br[8] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_11 
+ bl[9] br[9] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_12 
+ bl[10] br[10] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_13 
+ bl[11] br[11] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_14 
+ bl[12] br[12] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_15 
+ bl[13] br[13] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_16 
+ bl[14] br[14] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_17 
+ bl[15] br[15] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_18 
+ bl[16] br[16] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_19 
+ bl[17] br[17] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_20 
+ bl[18] br[18] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_21 
+ bl[19] br[19] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_22 
+ bl[20] br[20] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_23 
+ bl[21] br[21] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_24 
+ bl[22] br[22] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_25 
+ bl[23] br[23] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_26 
+ bl[24] br[24] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_27 
+ bl[25] br[25] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_28 
+ bl[26] br[26] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_29 
+ bl[27] br[27] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_30 
+ bl[28] br[28] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_31 
+ bl[29] br[29] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_32 
+ bl[30] br[30] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_33 
+ bl[31] br[31] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_34 
+ bl[32] br[32] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_35 
+ bl[33] br[33] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_36 
+ bl[34] br[34] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_37 
+ bl[35] br[35] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_38 
+ bl[36] br[36] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_39 
+ bl[37] br[37] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_40 
+ bl[38] br[38] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_41 
+ bl[39] br[39] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_42 
+ bl[40] br[40] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_43 
+ bl[41] br[41] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_44 
+ bl[42] br[42] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_45 
+ bl[43] br[43] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_46 
+ bl[44] br[44] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_47 
+ bl[45] br[45] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_48 
+ bl[46] br[46] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_49 
+ bl[47] br[47] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_50 
+ bl[48] br[48] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_51 
+ bl[49] br[49] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_52 
+ bl[50] br[50] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_53 
+ bl[51] br[51] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_54 
+ bl[52] br[52] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_55 
+ bl[53] br[53] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_56 
+ bl[54] br[54] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_57 
+ bl[55] br[55] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_58 
+ bl[56] br[56] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_59 
+ bl[57] br[57] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_60 
+ bl[58] br[58] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_61 
+ bl[59] br[59] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_62 
+ bl[60] br[60] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_63 
+ bl[61] br[61] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_64 
+ bl[62] br[62] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_65 
+ bl[63] br[63] vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_66 
+ vdd vdd vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_276_67 
+ vdd vdd vdd vss wl[274] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_0 
+ vdd vdd vss vdd vpb vnb wl[275] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_277_1 
+ rbl rbr vss vdd vpb vnb wl[275] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_277_2 
+ bl[0] br[0] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_3 
+ bl[1] br[1] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_4 
+ bl[2] br[2] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_5 
+ bl[3] br[3] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_6 
+ bl[4] br[4] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_7 
+ bl[5] br[5] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_8 
+ bl[6] br[6] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_9 
+ bl[7] br[7] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_10 
+ bl[8] br[8] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_11 
+ bl[9] br[9] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_12 
+ bl[10] br[10] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_13 
+ bl[11] br[11] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_14 
+ bl[12] br[12] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_15 
+ bl[13] br[13] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_16 
+ bl[14] br[14] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_17 
+ bl[15] br[15] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_18 
+ bl[16] br[16] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_19 
+ bl[17] br[17] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_20 
+ bl[18] br[18] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_21 
+ bl[19] br[19] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_22 
+ bl[20] br[20] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_23 
+ bl[21] br[21] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_24 
+ bl[22] br[22] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_25 
+ bl[23] br[23] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_26 
+ bl[24] br[24] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_27 
+ bl[25] br[25] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_28 
+ bl[26] br[26] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_29 
+ bl[27] br[27] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_30 
+ bl[28] br[28] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_31 
+ bl[29] br[29] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_32 
+ bl[30] br[30] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_33 
+ bl[31] br[31] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_34 
+ bl[32] br[32] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_35 
+ bl[33] br[33] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_36 
+ bl[34] br[34] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_37 
+ bl[35] br[35] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_38 
+ bl[36] br[36] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_39 
+ bl[37] br[37] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_40 
+ bl[38] br[38] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_41 
+ bl[39] br[39] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_42 
+ bl[40] br[40] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_43 
+ bl[41] br[41] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_44 
+ bl[42] br[42] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_45 
+ bl[43] br[43] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_46 
+ bl[44] br[44] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_47 
+ bl[45] br[45] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_48 
+ bl[46] br[46] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_49 
+ bl[47] br[47] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_50 
+ bl[48] br[48] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_51 
+ bl[49] br[49] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_52 
+ bl[50] br[50] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_53 
+ bl[51] br[51] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_54 
+ bl[52] br[52] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_55 
+ bl[53] br[53] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_56 
+ bl[54] br[54] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_57 
+ bl[55] br[55] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_58 
+ bl[56] br[56] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_59 
+ bl[57] br[57] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_60 
+ bl[58] br[58] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_61 
+ bl[59] br[59] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_62 
+ bl[60] br[60] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_63 
+ bl[61] br[61] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_64 
+ bl[62] br[62] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_65 
+ bl[63] br[63] vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_66 
+ vdd vdd vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_277_67 
+ vdd vdd vdd vss wl[275] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_0 
+ vdd vdd vss vdd vpb vnb wl[276] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_278_1 
+ rbl rbr vss vdd vpb vnb wl[276] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_278_2 
+ bl[0] br[0] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_3 
+ bl[1] br[1] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_4 
+ bl[2] br[2] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_5 
+ bl[3] br[3] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_6 
+ bl[4] br[4] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_7 
+ bl[5] br[5] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_8 
+ bl[6] br[6] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_9 
+ bl[7] br[7] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_10 
+ bl[8] br[8] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_11 
+ bl[9] br[9] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_12 
+ bl[10] br[10] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_13 
+ bl[11] br[11] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_14 
+ bl[12] br[12] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_15 
+ bl[13] br[13] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_16 
+ bl[14] br[14] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_17 
+ bl[15] br[15] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_18 
+ bl[16] br[16] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_19 
+ bl[17] br[17] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_20 
+ bl[18] br[18] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_21 
+ bl[19] br[19] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_22 
+ bl[20] br[20] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_23 
+ bl[21] br[21] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_24 
+ bl[22] br[22] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_25 
+ bl[23] br[23] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_26 
+ bl[24] br[24] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_27 
+ bl[25] br[25] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_28 
+ bl[26] br[26] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_29 
+ bl[27] br[27] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_30 
+ bl[28] br[28] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_31 
+ bl[29] br[29] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_32 
+ bl[30] br[30] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_33 
+ bl[31] br[31] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_34 
+ bl[32] br[32] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_35 
+ bl[33] br[33] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_36 
+ bl[34] br[34] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_37 
+ bl[35] br[35] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_38 
+ bl[36] br[36] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_39 
+ bl[37] br[37] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_40 
+ bl[38] br[38] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_41 
+ bl[39] br[39] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_42 
+ bl[40] br[40] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_43 
+ bl[41] br[41] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_44 
+ bl[42] br[42] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_45 
+ bl[43] br[43] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_46 
+ bl[44] br[44] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_47 
+ bl[45] br[45] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_48 
+ bl[46] br[46] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_49 
+ bl[47] br[47] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_50 
+ bl[48] br[48] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_51 
+ bl[49] br[49] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_52 
+ bl[50] br[50] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_53 
+ bl[51] br[51] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_54 
+ bl[52] br[52] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_55 
+ bl[53] br[53] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_56 
+ bl[54] br[54] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_57 
+ bl[55] br[55] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_58 
+ bl[56] br[56] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_59 
+ bl[57] br[57] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_60 
+ bl[58] br[58] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_61 
+ bl[59] br[59] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_62 
+ bl[60] br[60] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_63 
+ bl[61] br[61] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_64 
+ bl[62] br[62] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_65 
+ bl[63] br[63] vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_66 
+ vdd vdd vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_278_67 
+ vdd vdd vdd vss wl[276] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_0 
+ vdd vdd vss vdd vpb vnb wl[277] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_279_1 
+ rbl rbr vss vdd vpb vnb wl[277] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_279_2 
+ bl[0] br[0] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_3 
+ bl[1] br[1] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_4 
+ bl[2] br[2] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_5 
+ bl[3] br[3] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_6 
+ bl[4] br[4] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_7 
+ bl[5] br[5] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_8 
+ bl[6] br[6] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_9 
+ bl[7] br[7] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_10 
+ bl[8] br[8] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_11 
+ bl[9] br[9] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_12 
+ bl[10] br[10] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_13 
+ bl[11] br[11] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_14 
+ bl[12] br[12] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_15 
+ bl[13] br[13] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_16 
+ bl[14] br[14] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_17 
+ bl[15] br[15] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_18 
+ bl[16] br[16] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_19 
+ bl[17] br[17] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_20 
+ bl[18] br[18] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_21 
+ bl[19] br[19] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_22 
+ bl[20] br[20] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_23 
+ bl[21] br[21] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_24 
+ bl[22] br[22] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_25 
+ bl[23] br[23] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_26 
+ bl[24] br[24] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_27 
+ bl[25] br[25] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_28 
+ bl[26] br[26] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_29 
+ bl[27] br[27] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_30 
+ bl[28] br[28] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_31 
+ bl[29] br[29] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_32 
+ bl[30] br[30] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_33 
+ bl[31] br[31] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_34 
+ bl[32] br[32] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_35 
+ bl[33] br[33] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_36 
+ bl[34] br[34] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_37 
+ bl[35] br[35] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_38 
+ bl[36] br[36] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_39 
+ bl[37] br[37] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_40 
+ bl[38] br[38] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_41 
+ bl[39] br[39] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_42 
+ bl[40] br[40] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_43 
+ bl[41] br[41] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_44 
+ bl[42] br[42] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_45 
+ bl[43] br[43] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_46 
+ bl[44] br[44] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_47 
+ bl[45] br[45] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_48 
+ bl[46] br[46] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_49 
+ bl[47] br[47] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_50 
+ bl[48] br[48] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_51 
+ bl[49] br[49] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_52 
+ bl[50] br[50] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_53 
+ bl[51] br[51] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_54 
+ bl[52] br[52] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_55 
+ bl[53] br[53] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_56 
+ bl[54] br[54] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_57 
+ bl[55] br[55] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_58 
+ bl[56] br[56] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_59 
+ bl[57] br[57] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_60 
+ bl[58] br[58] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_61 
+ bl[59] br[59] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_62 
+ bl[60] br[60] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_63 
+ bl[61] br[61] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_64 
+ bl[62] br[62] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_65 
+ bl[63] br[63] vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_66 
+ vdd vdd vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_279_67 
+ vdd vdd vdd vss wl[277] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_0 
+ vdd vdd vss vdd vpb vnb wl[278] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_280_1 
+ rbl rbr vss vdd vpb vnb wl[278] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_280_2 
+ bl[0] br[0] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_3 
+ bl[1] br[1] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_4 
+ bl[2] br[2] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_5 
+ bl[3] br[3] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_6 
+ bl[4] br[4] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_7 
+ bl[5] br[5] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_8 
+ bl[6] br[6] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_9 
+ bl[7] br[7] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_10 
+ bl[8] br[8] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_11 
+ bl[9] br[9] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_12 
+ bl[10] br[10] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_13 
+ bl[11] br[11] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_14 
+ bl[12] br[12] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_15 
+ bl[13] br[13] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_16 
+ bl[14] br[14] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_17 
+ bl[15] br[15] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_18 
+ bl[16] br[16] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_19 
+ bl[17] br[17] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_20 
+ bl[18] br[18] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_21 
+ bl[19] br[19] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_22 
+ bl[20] br[20] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_23 
+ bl[21] br[21] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_24 
+ bl[22] br[22] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_25 
+ bl[23] br[23] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_26 
+ bl[24] br[24] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_27 
+ bl[25] br[25] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_28 
+ bl[26] br[26] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_29 
+ bl[27] br[27] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_30 
+ bl[28] br[28] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_31 
+ bl[29] br[29] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_32 
+ bl[30] br[30] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_33 
+ bl[31] br[31] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_34 
+ bl[32] br[32] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_35 
+ bl[33] br[33] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_36 
+ bl[34] br[34] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_37 
+ bl[35] br[35] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_38 
+ bl[36] br[36] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_39 
+ bl[37] br[37] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_40 
+ bl[38] br[38] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_41 
+ bl[39] br[39] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_42 
+ bl[40] br[40] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_43 
+ bl[41] br[41] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_44 
+ bl[42] br[42] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_45 
+ bl[43] br[43] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_46 
+ bl[44] br[44] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_47 
+ bl[45] br[45] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_48 
+ bl[46] br[46] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_49 
+ bl[47] br[47] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_50 
+ bl[48] br[48] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_51 
+ bl[49] br[49] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_52 
+ bl[50] br[50] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_53 
+ bl[51] br[51] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_54 
+ bl[52] br[52] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_55 
+ bl[53] br[53] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_56 
+ bl[54] br[54] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_57 
+ bl[55] br[55] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_58 
+ bl[56] br[56] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_59 
+ bl[57] br[57] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_60 
+ bl[58] br[58] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_61 
+ bl[59] br[59] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_62 
+ bl[60] br[60] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_63 
+ bl[61] br[61] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_64 
+ bl[62] br[62] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_65 
+ bl[63] br[63] vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_66 
+ vdd vdd vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_280_67 
+ vdd vdd vdd vss wl[278] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_0 
+ vdd vdd vss vdd vpb vnb wl[279] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_281_1 
+ rbl rbr vss vdd vpb vnb wl[279] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_281_2 
+ bl[0] br[0] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_3 
+ bl[1] br[1] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_4 
+ bl[2] br[2] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_5 
+ bl[3] br[3] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_6 
+ bl[4] br[4] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_7 
+ bl[5] br[5] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_8 
+ bl[6] br[6] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_9 
+ bl[7] br[7] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_10 
+ bl[8] br[8] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_11 
+ bl[9] br[9] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_12 
+ bl[10] br[10] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_13 
+ bl[11] br[11] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_14 
+ bl[12] br[12] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_15 
+ bl[13] br[13] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_16 
+ bl[14] br[14] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_17 
+ bl[15] br[15] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_18 
+ bl[16] br[16] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_19 
+ bl[17] br[17] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_20 
+ bl[18] br[18] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_21 
+ bl[19] br[19] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_22 
+ bl[20] br[20] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_23 
+ bl[21] br[21] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_24 
+ bl[22] br[22] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_25 
+ bl[23] br[23] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_26 
+ bl[24] br[24] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_27 
+ bl[25] br[25] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_28 
+ bl[26] br[26] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_29 
+ bl[27] br[27] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_30 
+ bl[28] br[28] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_31 
+ bl[29] br[29] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_32 
+ bl[30] br[30] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_33 
+ bl[31] br[31] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_34 
+ bl[32] br[32] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_35 
+ bl[33] br[33] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_36 
+ bl[34] br[34] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_37 
+ bl[35] br[35] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_38 
+ bl[36] br[36] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_39 
+ bl[37] br[37] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_40 
+ bl[38] br[38] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_41 
+ bl[39] br[39] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_42 
+ bl[40] br[40] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_43 
+ bl[41] br[41] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_44 
+ bl[42] br[42] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_45 
+ bl[43] br[43] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_46 
+ bl[44] br[44] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_47 
+ bl[45] br[45] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_48 
+ bl[46] br[46] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_49 
+ bl[47] br[47] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_50 
+ bl[48] br[48] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_51 
+ bl[49] br[49] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_52 
+ bl[50] br[50] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_53 
+ bl[51] br[51] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_54 
+ bl[52] br[52] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_55 
+ bl[53] br[53] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_56 
+ bl[54] br[54] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_57 
+ bl[55] br[55] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_58 
+ bl[56] br[56] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_59 
+ bl[57] br[57] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_60 
+ bl[58] br[58] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_61 
+ bl[59] br[59] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_62 
+ bl[60] br[60] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_63 
+ bl[61] br[61] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_64 
+ bl[62] br[62] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_65 
+ bl[63] br[63] vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_66 
+ vdd vdd vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_281_67 
+ vdd vdd vdd vss wl[279] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_0 
+ vdd vdd vss vdd vpb vnb wl[280] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_282_1 
+ rbl rbr vss vdd vpb vnb wl[280] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_282_2 
+ bl[0] br[0] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_3 
+ bl[1] br[1] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_4 
+ bl[2] br[2] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_5 
+ bl[3] br[3] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_6 
+ bl[4] br[4] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_7 
+ bl[5] br[5] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_8 
+ bl[6] br[6] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_9 
+ bl[7] br[7] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_10 
+ bl[8] br[8] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_11 
+ bl[9] br[9] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_12 
+ bl[10] br[10] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_13 
+ bl[11] br[11] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_14 
+ bl[12] br[12] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_15 
+ bl[13] br[13] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_16 
+ bl[14] br[14] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_17 
+ bl[15] br[15] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_18 
+ bl[16] br[16] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_19 
+ bl[17] br[17] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_20 
+ bl[18] br[18] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_21 
+ bl[19] br[19] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_22 
+ bl[20] br[20] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_23 
+ bl[21] br[21] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_24 
+ bl[22] br[22] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_25 
+ bl[23] br[23] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_26 
+ bl[24] br[24] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_27 
+ bl[25] br[25] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_28 
+ bl[26] br[26] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_29 
+ bl[27] br[27] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_30 
+ bl[28] br[28] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_31 
+ bl[29] br[29] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_32 
+ bl[30] br[30] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_33 
+ bl[31] br[31] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_34 
+ bl[32] br[32] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_35 
+ bl[33] br[33] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_36 
+ bl[34] br[34] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_37 
+ bl[35] br[35] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_38 
+ bl[36] br[36] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_39 
+ bl[37] br[37] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_40 
+ bl[38] br[38] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_41 
+ bl[39] br[39] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_42 
+ bl[40] br[40] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_43 
+ bl[41] br[41] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_44 
+ bl[42] br[42] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_45 
+ bl[43] br[43] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_46 
+ bl[44] br[44] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_47 
+ bl[45] br[45] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_48 
+ bl[46] br[46] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_49 
+ bl[47] br[47] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_50 
+ bl[48] br[48] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_51 
+ bl[49] br[49] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_52 
+ bl[50] br[50] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_53 
+ bl[51] br[51] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_54 
+ bl[52] br[52] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_55 
+ bl[53] br[53] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_56 
+ bl[54] br[54] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_57 
+ bl[55] br[55] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_58 
+ bl[56] br[56] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_59 
+ bl[57] br[57] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_60 
+ bl[58] br[58] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_61 
+ bl[59] br[59] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_62 
+ bl[60] br[60] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_63 
+ bl[61] br[61] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_64 
+ bl[62] br[62] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_65 
+ bl[63] br[63] vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_66 
+ vdd vdd vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_282_67 
+ vdd vdd vdd vss wl[280] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_0 
+ vdd vdd vss vdd vpb vnb wl[281] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_283_1 
+ rbl rbr vss vdd vpb vnb wl[281] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_283_2 
+ bl[0] br[0] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_3 
+ bl[1] br[1] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_4 
+ bl[2] br[2] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_5 
+ bl[3] br[3] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_6 
+ bl[4] br[4] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_7 
+ bl[5] br[5] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_8 
+ bl[6] br[6] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_9 
+ bl[7] br[7] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_10 
+ bl[8] br[8] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_11 
+ bl[9] br[9] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_12 
+ bl[10] br[10] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_13 
+ bl[11] br[11] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_14 
+ bl[12] br[12] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_15 
+ bl[13] br[13] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_16 
+ bl[14] br[14] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_17 
+ bl[15] br[15] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_18 
+ bl[16] br[16] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_19 
+ bl[17] br[17] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_20 
+ bl[18] br[18] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_21 
+ bl[19] br[19] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_22 
+ bl[20] br[20] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_23 
+ bl[21] br[21] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_24 
+ bl[22] br[22] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_25 
+ bl[23] br[23] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_26 
+ bl[24] br[24] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_27 
+ bl[25] br[25] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_28 
+ bl[26] br[26] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_29 
+ bl[27] br[27] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_30 
+ bl[28] br[28] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_31 
+ bl[29] br[29] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_32 
+ bl[30] br[30] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_33 
+ bl[31] br[31] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_34 
+ bl[32] br[32] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_35 
+ bl[33] br[33] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_36 
+ bl[34] br[34] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_37 
+ bl[35] br[35] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_38 
+ bl[36] br[36] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_39 
+ bl[37] br[37] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_40 
+ bl[38] br[38] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_41 
+ bl[39] br[39] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_42 
+ bl[40] br[40] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_43 
+ bl[41] br[41] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_44 
+ bl[42] br[42] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_45 
+ bl[43] br[43] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_46 
+ bl[44] br[44] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_47 
+ bl[45] br[45] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_48 
+ bl[46] br[46] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_49 
+ bl[47] br[47] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_50 
+ bl[48] br[48] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_51 
+ bl[49] br[49] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_52 
+ bl[50] br[50] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_53 
+ bl[51] br[51] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_54 
+ bl[52] br[52] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_55 
+ bl[53] br[53] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_56 
+ bl[54] br[54] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_57 
+ bl[55] br[55] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_58 
+ bl[56] br[56] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_59 
+ bl[57] br[57] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_60 
+ bl[58] br[58] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_61 
+ bl[59] br[59] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_62 
+ bl[60] br[60] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_63 
+ bl[61] br[61] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_64 
+ bl[62] br[62] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_65 
+ bl[63] br[63] vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_66 
+ vdd vdd vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_283_67 
+ vdd vdd vdd vss wl[281] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_0 
+ vdd vdd vss vdd vpb vnb wl[282] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_284_1 
+ rbl rbr vss vdd vpb vnb wl[282] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_284_2 
+ bl[0] br[0] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_3 
+ bl[1] br[1] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_4 
+ bl[2] br[2] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_5 
+ bl[3] br[3] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_6 
+ bl[4] br[4] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_7 
+ bl[5] br[5] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_8 
+ bl[6] br[6] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_9 
+ bl[7] br[7] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_10 
+ bl[8] br[8] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_11 
+ bl[9] br[9] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_12 
+ bl[10] br[10] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_13 
+ bl[11] br[11] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_14 
+ bl[12] br[12] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_15 
+ bl[13] br[13] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_16 
+ bl[14] br[14] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_17 
+ bl[15] br[15] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_18 
+ bl[16] br[16] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_19 
+ bl[17] br[17] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_20 
+ bl[18] br[18] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_21 
+ bl[19] br[19] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_22 
+ bl[20] br[20] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_23 
+ bl[21] br[21] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_24 
+ bl[22] br[22] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_25 
+ bl[23] br[23] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_26 
+ bl[24] br[24] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_27 
+ bl[25] br[25] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_28 
+ bl[26] br[26] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_29 
+ bl[27] br[27] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_30 
+ bl[28] br[28] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_31 
+ bl[29] br[29] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_32 
+ bl[30] br[30] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_33 
+ bl[31] br[31] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_34 
+ bl[32] br[32] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_35 
+ bl[33] br[33] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_36 
+ bl[34] br[34] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_37 
+ bl[35] br[35] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_38 
+ bl[36] br[36] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_39 
+ bl[37] br[37] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_40 
+ bl[38] br[38] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_41 
+ bl[39] br[39] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_42 
+ bl[40] br[40] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_43 
+ bl[41] br[41] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_44 
+ bl[42] br[42] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_45 
+ bl[43] br[43] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_46 
+ bl[44] br[44] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_47 
+ bl[45] br[45] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_48 
+ bl[46] br[46] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_49 
+ bl[47] br[47] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_50 
+ bl[48] br[48] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_51 
+ bl[49] br[49] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_52 
+ bl[50] br[50] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_53 
+ bl[51] br[51] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_54 
+ bl[52] br[52] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_55 
+ bl[53] br[53] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_56 
+ bl[54] br[54] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_57 
+ bl[55] br[55] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_58 
+ bl[56] br[56] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_59 
+ bl[57] br[57] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_60 
+ bl[58] br[58] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_61 
+ bl[59] br[59] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_62 
+ bl[60] br[60] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_63 
+ bl[61] br[61] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_64 
+ bl[62] br[62] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_65 
+ bl[63] br[63] vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_66 
+ vdd vdd vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_284_67 
+ vdd vdd vdd vss wl[282] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_0 
+ vdd vdd vss vdd vpb vnb wl[283] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_285_1 
+ rbl rbr vss vdd vpb vnb wl[283] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_285_2 
+ bl[0] br[0] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_3 
+ bl[1] br[1] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_4 
+ bl[2] br[2] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_5 
+ bl[3] br[3] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_6 
+ bl[4] br[4] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_7 
+ bl[5] br[5] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_8 
+ bl[6] br[6] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_9 
+ bl[7] br[7] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_10 
+ bl[8] br[8] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_11 
+ bl[9] br[9] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_12 
+ bl[10] br[10] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_13 
+ bl[11] br[11] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_14 
+ bl[12] br[12] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_15 
+ bl[13] br[13] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_16 
+ bl[14] br[14] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_17 
+ bl[15] br[15] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_18 
+ bl[16] br[16] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_19 
+ bl[17] br[17] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_20 
+ bl[18] br[18] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_21 
+ bl[19] br[19] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_22 
+ bl[20] br[20] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_23 
+ bl[21] br[21] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_24 
+ bl[22] br[22] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_25 
+ bl[23] br[23] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_26 
+ bl[24] br[24] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_27 
+ bl[25] br[25] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_28 
+ bl[26] br[26] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_29 
+ bl[27] br[27] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_30 
+ bl[28] br[28] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_31 
+ bl[29] br[29] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_32 
+ bl[30] br[30] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_33 
+ bl[31] br[31] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_34 
+ bl[32] br[32] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_35 
+ bl[33] br[33] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_36 
+ bl[34] br[34] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_37 
+ bl[35] br[35] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_38 
+ bl[36] br[36] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_39 
+ bl[37] br[37] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_40 
+ bl[38] br[38] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_41 
+ bl[39] br[39] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_42 
+ bl[40] br[40] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_43 
+ bl[41] br[41] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_44 
+ bl[42] br[42] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_45 
+ bl[43] br[43] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_46 
+ bl[44] br[44] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_47 
+ bl[45] br[45] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_48 
+ bl[46] br[46] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_49 
+ bl[47] br[47] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_50 
+ bl[48] br[48] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_51 
+ bl[49] br[49] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_52 
+ bl[50] br[50] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_53 
+ bl[51] br[51] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_54 
+ bl[52] br[52] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_55 
+ bl[53] br[53] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_56 
+ bl[54] br[54] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_57 
+ bl[55] br[55] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_58 
+ bl[56] br[56] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_59 
+ bl[57] br[57] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_60 
+ bl[58] br[58] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_61 
+ bl[59] br[59] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_62 
+ bl[60] br[60] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_63 
+ bl[61] br[61] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_64 
+ bl[62] br[62] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_65 
+ bl[63] br[63] vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_66 
+ vdd vdd vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_285_67 
+ vdd vdd vdd vss wl[283] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_0 
+ vdd vdd vss vdd vpb vnb wl[284] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_286_1 
+ rbl rbr vss vdd vpb vnb wl[284] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_286_2 
+ bl[0] br[0] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_3 
+ bl[1] br[1] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_4 
+ bl[2] br[2] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_5 
+ bl[3] br[3] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_6 
+ bl[4] br[4] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_7 
+ bl[5] br[5] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_8 
+ bl[6] br[6] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_9 
+ bl[7] br[7] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_10 
+ bl[8] br[8] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_11 
+ bl[9] br[9] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_12 
+ bl[10] br[10] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_13 
+ bl[11] br[11] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_14 
+ bl[12] br[12] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_15 
+ bl[13] br[13] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_16 
+ bl[14] br[14] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_17 
+ bl[15] br[15] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_18 
+ bl[16] br[16] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_19 
+ bl[17] br[17] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_20 
+ bl[18] br[18] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_21 
+ bl[19] br[19] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_22 
+ bl[20] br[20] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_23 
+ bl[21] br[21] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_24 
+ bl[22] br[22] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_25 
+ bl[23] br[23] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_26 
+ bl[24] br[24] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_27 
+ bl[25] br[25] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_28 
+ bl[26] br[26] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_29 
+ bl[27] br[27] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_30 
+ bl[28] br[28] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_31 
+ bl[29] br[29] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_32 
+ bl[30] br[30] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_33 
+ bl[31] br[31] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_34 
+ bl[32] br[32] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_35 
+ bl[33] br[33] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_36 
+ bl[34] br[34] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_37 
+ bl[35] br[35] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_38 
+ bl[36] br[36] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_39 
+ bl[37] br[37] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_40 
+ bl[38] br[38] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_41 
+ bl[39] br[39] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_42 
+ bl[40] br[40] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_43 
+ bl[41] br[41] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_44 
+ bl[42] br[42] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_45 
+ bl[43] br[43] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_46 
+ bl[44] br[44] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_47 
+ bl[45] br[45] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_48 
+ bl[46] br[46] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_49 
+ bl[47] br[47] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_50 
+ bl[48] br[48] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_51 
+ bl[49] br[49] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_52 
+ bl[50] br[50] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_53 
+ bl[51] br[51] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_54 
+ bl[52] br[52] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_55 
+ bl[53] br[53] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_56 
+ bl[54] br[54] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_57 
+ bl[55] br[55] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_58 
+ bl[56] br[56] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_59 
+ bl[57] br[57] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_60 
+ bl[58] br[58] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_61 
+ bl[59] br[59] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_62 
+ bl[60] br[60] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_63 
+ bl[61] br[61] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_64 
+ bl[62] br[62] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_65 
+ bl[63] br[63] vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_66 
+ vdd vdd vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_286_67 
+ vdd vdd vdd vss wl[284] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_0 
+ vdd vdd vss vdd vpb vnb wl[285] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_287_1 
+ rbl rbr vss vdd vpb vnb wl[285] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_287_2 
+ bl[0] br[0] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_3 
+ bl[1] br[1] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_4 
+ bl[2] br[2] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_5 
+ bl[3] br[3] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_6 
+ bl[4] br[4] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_7 
+ bl[5] br[5] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_8 
+ bl[6] br[6] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_9 
+ bl[7] br[7] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_10 
+ bl[8] br[8] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_11 
+ bl[9] br[9] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_12 
+ bl[10] br[10] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_13 
+ bl[11] br[11] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_14 
+ bl[12] br[12] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_15 
+ bl[13] br[13] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_16 
+ bl[14] br[14] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_17 
+ bl[15] br[15] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_18 
+ bl[16] br[16] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_19 
+ bl[17] br[17] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_20 
+ bl[18] br[18] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_21 
+ bl[19] br[19] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_22 
+ bl[20] br[20] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_23 
+ bl[21] br[21] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_24 
+ bl[22] br[22] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_25 
+ bl[23] br[23] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_26 
+ bl[24] br[24] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_27 
+ bl[25] br[25] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_28 
+ bl[26] br[26] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_29 
+ bl[27] br[27] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_30 
+ bl[28] br[28] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_31 
+ bl[29] br[29] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_32 
+ bl[30] br[30] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_33 
+ bl[31] br[31] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_34 
+ bl[32] br[32] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_35 
+ bl[33] br[33] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_36 
+ bl[34] br[34] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_37 
+ bl[35] br[35] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_38 
+ bl[36] br[36] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_39 
+ bl[37] br[37] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_40 
+ bl[38] br[38] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_41 
+ bl[39] br[39] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_42 
+ bl[40] br[40] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_43 
+ bl[41] br[41] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_44 
+ bl[42] br[42] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_45 
+ bl[43] br[43] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_46 
+ bl[44] br[44] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_47 
+ bl[45] br[45] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_48 
+ bl[46] br[46] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_49 
+ bl[47] br[47] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_50 
+ bl[48] br[48] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_51 
+ bl[49] br[49] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_52 
+ bl[50] br[50] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_53 
+ bl[51] br[51] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_54 
+ bl[52] br[52] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_55 
+ bl[53] br[53] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_56 
+ bl[54] br[54] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_57 
+ bl[55] br[55] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_58 
+ bl[56] br[56] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_59 
+ bl[57] br[57] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_60 
+ bl[58] br[58] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_61 
+ bl[59] br[59] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_62 
+ bl[60] br[60] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_63 
+ bl[61] br[61] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_64 
+ bl[62] br[62] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_65 
+ bl[63] br[63] vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_66 
+ vdd vdd vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_287_67 
+ vdd vdd vdd vss wl[285] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_0 
+ vdd vdd vss vdd vpb vnb wl[286] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_288_1 
+ rbl rbr vss vdd vpb vnb wl[286] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_288_2 
+ bl[0] br[0] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_3 
+ bl[1] br[1] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_4 
+ bl[2] br[2] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_5 
+ bl[3] br[3] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_6 
+ bl[4] br[4] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_7 
+ bl[5] br[5] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_8 
+ bl[6] br[6] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_9 
+ bl[7] br[7] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_10 
+ bl[8] br[8] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_11 
+ bl[9] br[9] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_12 
+ bl[10] br[10] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_13 
+ bl[11] br[11] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_14 
+ bl[12] br[12] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_15 
+ bl[13] br[13] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_16 
+ bl[14] br[14] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_17 
+ bl[15] br[15] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_18 
+ bl[16] br[16] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_19 
+ bl[17] br[17] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_20 
+ bl[18] br[18] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_21 
+ bl[19] br[19] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_22 
+ bl[20] br[20] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_23 
+ bl[21] br[21] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_24 
+ bl[22] br[22] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_25 
+ bl[23] br[23] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_26 
+ bl[24] br[24] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_27 
+ bl[25] br[25] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_28 
+ bl[26] br[26] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_29 
+ bl[27] br[27] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_30 
+ bl[28] br[28] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_31 
+ bl[29] br[29] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_32 
+ bl[30] br[30] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_33 
+ bl[31] br[31] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_34 
+ bl[32] br[32] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_35 
+ bl[33] br[33] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_36 
+ bl[34] br[34] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_37 
+ bl[35] br[35] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_38 
+ bl[36] br[36] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_39 
+ bl[37] br[37] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_40 
+ bl[38] br[38] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_41 
+ bl[39] br[39] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_42 
+ bl[40] br[40] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_43 
+ bl[41] br[41] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_44 
+ bl[42] br[42] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_45 
+ bl[43] br[43] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_46 
+ bl[44] br[44] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_47 
+ bl[45] br[45] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_48 
+ bl[46] br[46] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_49 
+ bl[47] br[47] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_50 
+ bl[48] br[48] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_51 
+ bl[49] br[49] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_52 
+ bl[50] br[50] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_53 
+ bl[51] br[51] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_54 
+ bl[52] br[52] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_55 
+ bl[53] br[53] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_56 
+ bl[54] br[54] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_57 
+ bl[55] br[55] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_58 
+ bl[56] br[56] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_59 
+ bl[57] br[57] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_60 
+ bl[58] br[58] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_61 
+ bl[59] br[59] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_62 
+ bl[60] br[60] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_63 
+ bl[61] br[61] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_64 
+ bl[62] br[62] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_65 
+ bl[63] br[63] vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_66 
+ vdd vdd vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_288_67 
+ vdd vdd vdd vss wl[286] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_0 
+ vdd vdd vss vdd vpb vnb wl[287] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_289_1 
+ rbl rbr vss vdd vpb vnb wl[287] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_289_2 
+ bl[0] br[0] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_3 
+ bl[1] br[1] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_4 
+ bl[2] br[2] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_5 
+ bl[3] br[3] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_6 
+ bl[4] br[4] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_7 
+ bl[5] br[5] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_8 
+ bl[6] br[6] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_9 
+ bl[7] br[7] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_10 
+ bl[8] br[8] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_11 
+ bl[9] br[9] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_12 
+ bl[10] br[10] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_13 
+ bl[11] br[11] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_14 
+ bl[12] br[12] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_15 
+ bl[13] br[13] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_16 
+ bl[14] br[14] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_17 
+ bl[15] br[15] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_18 
+ bl[16] br[16] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_19 
+ bl[17] br[17] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_20 
+ bl[18] br[18] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_21 
+ bl[19] br[19] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_22 
+ bl[20] br[20] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_23 
+ bl[21] br[21] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_24 
+ bl[22] br[22] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_25 
+ bl[23] br[23] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_26 
+ bl[24] br[24] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_27 
+ bl[25] br[25] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_28 
+ bl[26] br[26] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_29 
+ bl[27] br[27] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_30 
+ bl[28] br[28] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_31 
+ bl[29] br[29] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_32 
+ bl[30] br[30] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_33 
+ bl[31] br[31] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_34 
+ bl[32] br[32] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_35 
+ bl[33] br[33] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_36 
+ bl[34] br[34] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_37 
+ bl[35] br[35] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_38 
+ bl[36] br[36] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_39 
+ bl[37] br[37] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_40 
+ bl[38] br[38] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_41 
+ bl[39] br[39] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_42 
+ bl[40] br[40] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_43 
+ bl[41] br[41] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_44 
+ bl[42] br[42] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_45 
+ bl[43] br[43] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_46 
+ bl[44] br[44] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_47 
+ bl[45] br[45] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_48 
+ bl[46] br[46] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_49 
+ bl[47] br[47] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_50 
+ bl[48] br[48] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_51 
+ bl[49] br[49] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_52 
+ bl[50] br[50] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_53 
+ bl[51] br[51] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_54 
+ bl[52] br[52] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_55 
+ bl[53] br[53] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_56 
+ bl[54] br[54] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_57 
+ bl[55] br[55] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_58 
+ bl[56] br[56] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_59 
+ bl[57] br[57] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_60 
+ bl[58] br[58] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_61 
+ bl[59] br[59] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_62 
+ bl[60] br[60] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_63 
+ bl[61] br[61] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_64 
+ bl[62] br[62] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_65 
+ bl[63] br[63] vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_66 
+ vdd vdd vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_289_67 
+ vdd vdd vdd vss wl[287] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_0 
+ vdd vdd vss vdd vpb vnb wl[288] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_290_1 
+ rbl rbr vss vdd vpb vnb wl[288] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_290_2 
+ bl[0] br[0] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_3 
+ bl[1] br[1] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_4 
+ bl[2] br[2] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_5 
+ bl[3] br[3] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_6 
+ bl[4] br[4] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_7 
+ bl[5] br[5] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_8 
+ bl[6] br[6] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_9 
+ bl[7] br[7] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_10 
+ bl[8] br[8] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_11 
+ bl[9] br[9] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_12 
+ bl[10] br[10] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_13 
+ bl[11] br[11] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_14 
+ bl[12] br[12] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_15 
+ bl[13] br[13] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_16 
+ bl[14] br[14] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_17 
+ bl[15] br[15] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_18 
+ bl[16] br[16] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_19 
+ bl[17] br[17] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_20 
+ bl[18] br[18] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_21 
+ bl[19] br[19] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_22 
+ bl[20] br[20] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_23 
+ bl[21] br[21] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_24 
+ bl[22] br[22] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_25 
+ bl[23] br[23] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_26 
+ bl[24] br[24] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_27 
+ bl[25] br[25] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_28 
+ bl[26] br[26] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_29 
+ bl[27] br[27] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_30 
+ bl[28] br[28] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_31 
+ bl[29] br[29] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_32 
+ bl[30] br[30] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_33 
+ bl[31] br[31] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_34 
+ bl[32] br[32] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_35 
+ bl[33] br[33] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_36 
+ bl[34] br[34] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_37 
+ bl[35] br[35] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_38 
+ bl[36] br[36] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_39 
+ bl[37] br[37] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_40 
+ bl[38] br[38] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_41 
+ bl[39] br[39] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_42 
+ bl[40] br[40] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_43 
+ bl[41] br[41] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_44 
+ bl[42] br[42] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_45 
+ bl[43] br[43] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_46 
+ bl[44] br[44] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_47 
+ bl[45] br[45] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_48 
+ bl[46] br[46] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_49 
+ bl[47] br[47] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_50 
+ bl[48] br[48] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_51 
+ bl[49] br[49] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_52 
+ bl[50] br[50] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_53 
+ bl[51] br[51] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_54 
+ bl[52] br[52] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_55 
+ bl[53] br[53] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_56 
+ bl[54] br[54] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_57 
+ bl[55] br[55] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_58 
+ bl[56] br[56] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_59 
+ bl[57] br[57] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_60 
+ bl[58] br[58] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_61 
+ bl[59] br[59] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_62 
+ bl[60] br[60] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_63 
+ bl[61] br[61] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_64 
+ bl[62] br[62] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_65 
+ bl[63] br[63] vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_66 
+ vdd vdd vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_290_67 
+ vdd vdd vdd vss wl[288] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_0 
+ vdd vdd vss vdd vpb vnb wl[289] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_291_1 
+ rbl rbr vss vdd vpb vnb wl[289] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_291_2 
+ bl[0] br[0] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_3 
+ bl[1] br[1] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_4 
+ bl[2] br[2] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_5 
+ bl[3] br[3] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_6 
+ bl[4] br[4] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_7 
+ bl[5] br[5] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_8 
+ bl[6] br[6] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_9 
+ bl[7] br[7] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_10 
+ bl[8] br[8] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_11 
+ bl[9] br[9] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_12 
+ bl[10] br[10] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_13 
+ bl[11] br[11] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_14 
+ bl[12] br[12] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_15 
+ bl[13] br[13] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_16 
+ bl[14] br[14] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_17 
+ bl[15] br[15] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_18 
+ bl[16] br[16] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_19 
+ bl[17] br[17] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_20 
+ bl[18] br[18] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_21 
+ bl[19] br[19] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_22 
+ bl[20] br[20] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_23 
+ bl[21] br[21] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_24 
+ bl[22] br[22] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_25 
+ bl[23] br[23] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_26 
+ bl[24] br[24] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_27 
+ bl[25] br[25] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_28 
+ bl[26] br[26] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_29 
+ bl[27] br[27] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_30 
+ bl[28] br[28] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_31 
+ bl[29] br[29] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_32 
+ bl[30] br[30] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_33 
+ bl[31] br[31] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_34 
+ bl[32] br[32] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_35 
+ bl[33] br[33] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_36 
+ bl[34] br[34] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_37 
+ bl[35] br[35] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_38 
+ bl[36] br[36] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_39 
+ bl[37] br[37] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_40 
+ bl[38] br[38] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_41 
+ bl[39] br[39] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_42 
+ bl[40] br[40] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_43 
+ bl[41] br[41] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_44 
+ bl[42] br[42] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_45 
+ bl[43] br[43] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_46 
+ bl[44] br[44] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_47 
+ bl[45] br[45] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_48 
+ bl[46] br[46] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_49 
+ bl[47] br[47] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_50 
+ bl[48] br[48] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_51 
+ bl[49] br[49] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_52 
+ bl[50] br[50] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_53 
+ bl[51] br[51] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_54 
+ bl[52] br[52] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_55 
+ bl[53] br[53] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_56 
+ bl[54] br[54] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_57 
+ bl[55] br[55] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_58 
+ bl[56] br[56] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_59 
+ bl[57] br[57] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_60 
+ bl[58] br[58] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_61 
+ bl[59] br[59] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_62 
+ bl[60] br[60] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_63 
+ bl[61] br[61] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_64 
+ bl[62] br[62] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_65 
+ bl[63] br[63] vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_66 
+ vdd vdd vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_291_67 
+ vdd vdd vdd vss wl[289] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_0 
+ vdd vdd vss vdd vpb vnb wl[290] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_292_1 
+ rbl rbr vss vdd vpb vnb wl[290] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_292_2 
+ bl[0] br[0] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_3 
+ bl[1] br[1] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_4 
+ bl[2] br[2] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_5 
+ bl[3] br[3] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_6 
+ bl[4] br[4] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_7 
+ bl[5] br[5] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_8 
+ bl[6] br[6] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_9 
+ bl[7] br[7] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_10 
+ bl[8] br[8] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_11 
+ bl[9] br[9] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_12 
+ bl[10] br[10] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_13 
+ bl[11] br[11] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_14 
+ bl[12] br[12] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_15 
+ bl[13] br[13] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_16 
+ bl[14] br[14] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_17 
+ bl[15] br[15] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_18 
+ bl[16] br[16] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_19 
+ bl[17] br[17] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_20 
+ bl[18] br[18] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_21 
+ bl[19] br[19] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_22 
+ bl[20] br[20] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_23 
+ bl[21] br[21] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_24 
+ bl[22] br[22] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_25 
+ bl[23] br[23] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_26 
+ bl[24] br[24] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_27 
+ bl[25] br[25] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_28 
+ bl[26] br[26] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_29 
+ bl[27] br[27] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_30 
+ bl[28] br[28] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_31 
+ bl[29] br[29] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_32 
+ bl[30] br[30] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_33 
+ bl[31] br[31] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_34 
+ bl[32] br[32] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_35 
+ bl[33] br[33] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_36 
+ bl[34] br[34] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_37 
+ bl[35] br[35] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_38 
+ bl[36] br[36] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_39 
+ bl[37] br[37] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_40 
+ bl[38] br[38] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_41 
+ bl[39] br[39] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_42 
+ bl[40] br[40] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_43 
+ bl[41] br[41] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_44 
+ bl[42] br[42] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_45 
+ bl[43] br[43] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_46 
+ bl[44] br[44] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_47 
+ bl[45] br[45] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_48 
+ bl[46] br[46] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_49 
+ bl[47] br[47] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_50 
+ bl[48] br[48] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_51 
+ bl[49] br[49] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_52 
+ bl[50] br[50] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_53 
+ bl[51] br[51] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_54 
+ bl[52] br[52] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_55 
+ bl[53] br[53] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_56 
+ bl[54] br[54] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_57 
+ bl[55] br[55] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_58 
+ bl[56] br[56] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_59 
+ bl[57] br[57] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_60 
+ bl[58] br[58] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_61 
+ bl[59] br[59] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_62 
+ bl[60] br[60] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_63 
+ bl[61] br[61] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_64 
+ bl[62] br[62] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_65 
+ bl[63] br[63] vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_66 
+ vdd vdd vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_292_67 
+ vdd vdd vdd vss wl[290] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_0 
+ vdd vdd vss vdd vpb vnb wl[291] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_293_1 
+ rbl rbr vss vdd vpb vnb wl[291] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_293_2 
+ bl[0] br[0] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_3 
+ bl[1] br[1] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_4 
+ bl[2] br[2] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_5 
+ bl[3] br[3] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_6 
+ bl[4] br[4] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_7 
+ bl[5] br[5] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_8 
+ bl[6] br[6] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_9 
+ bl[7] br[7] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_10 
+ bl[8] br[8] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_11 
+ bl[9] br[9] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_12 
+ bl[10] br[10] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_13 
+ bl[11] br[11] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_14 
+ bl[12] br[12] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_15 
+ bl[13] br[13] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_16 
+ bl[14] br[14] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_17 
+ bl[15] br[15] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_18 
+ bl[16] br[16] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_19 
+ bl[17] br[17] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_20 
+ bl[18] br[18] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_21 
+ bl[19] br[19] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_22 
+ bl[20] br[20] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_23 
+ bl[21] br[21] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_24 
+ bl[22] br[22] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_25 
+ bl[23] br[23] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_26 
+ bl[24] br[24] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_27 
+ bl[25] br[25] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_28 
+ bl[26] br[26] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_29 
+ bl[27] br[27] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_30 
+ bl[28] br[28] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_31 
+ bl[29] br[29] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_32 
+ bl[30] br[30] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_33 
+ bl[31] br[31] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_34 
+ bl[32] br[32] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_35 
+ bl[33] br[33] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_36 
+ bl[34] br[34] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_37 
+ bl[35] br[35] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_38 
+ bl[36] br[36] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_39 
+ bl[37] br[37] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_40 
+ bl[38] br[38] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_41 
+ bl[39] br[39] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_42 
+ bl[40] br[40] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_43 
+ bl[41] br[41] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_44 
+ bl[42] br[42] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_45 
+ bl[43] br[43] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_46 
+ bl[44] br[44] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_47 
+ bl[45] br[45] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_48 
+ bl[46] br[46] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_49 
+ bl[47] br[47] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_50 
+ bl[48] br[48] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_51 
+ bl[49] br[49] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_52 
+ bl[50] br[50] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_53 
+ bl[51] br[51] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_54 
+ bl[52] br[52] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_55 
+ bl[53] br[53] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_56 
+ bl[54] br[54] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_57 
+ bl[55] br[55] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_58 
+ bl[56] br[56] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_59 
+ bl[57] br[57] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_60 
+ bl[58] br[58] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_61 
+ bl[59] br[59] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_62 
+ bl[60] br[60] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_63 
+ bl[61] br[61] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_64 
+ bl[62] br[62] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_65 
+ bl[63] br[63] vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_66 
+ vdd vdd vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_293_67 
+ vdd vdd vdd vss wl[291] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_0 
+ vdd vdd vss vdd vpb vnb wl[292] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_294_1 
+ rbl rbr vss vdd vpb vnb wl[292] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_294_2 
+ bl[0] br[0] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_3 
+ bl[1] br[1] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_4 
+ bl[2] br[2] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_5 
+ bl[3] br[3] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_6 
+ bl[4] br[4] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_7 
+ bl[5] br[5] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_8 
+ bl[6] br[6] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_9 
+ bl[7] br[7] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_10 
+ bl[8] br[8] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_11 
+ bl[9] br[9] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_12 
+ bl[10] br[10] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_13 
+ bl[11] br[11] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_14 
+ bl[12] br[12] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_15 
+ bl[13] br[13] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_16 
+ bl[14] br[14] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_17 
+ bl[15] br[15] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_18 
+ bl[16] br[16] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_19 
+ bl[17] br[17] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_20 
+ bl[18] br[18] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_21 
+ bl[19] br[19] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_22 
+ bl[20] br[20] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_23 
+ bl[21] br[21] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_24 
+ bl[22] br[22] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_25 
+ bl[23] br[23] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_26 
+ bl[24] br[24] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_27 
+ bl[25] br[25] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_28 
+ bl[26] br[26] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_29 
+ bl[27] br[27] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_30 
+ bl[28] br[28] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_31 
+ bl[29] br[29] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_32 
+ bl[30] br[30] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_33 
+ bl[31] br[31] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_34 
+ bl[32] br[32] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_35 
+ bl[33] br[33] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_36 
+ bl[34] br[34] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_37 
+ bl[35] br[35] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_38 
+ bl[36] br[36] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_39 
+ bl[37] br[37] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_40 
+ bl[38] br[38] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_41 
+ bl[39] br[39] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_42 
+ bl[40] br[40] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_43 
+ bl[41] br[41] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_44 
+ bl[42] br[42] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_45 
+ bl[43] br[43] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_46 
+ bl[44] br[44] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_47 
+ bl[45] br[45] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_48 
+ bl[46] br[46] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_49 
+ bl[47] br[47] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_50 
+ bl[48] br[48] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_51 
+ bl[49] br[49] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_52 
+ bl[50] br[50] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_53 
+ bl[51] br[51] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_54 
+ bl[52] br[52] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_55 
+ bl[53] br[53] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_56 
+ bl[54] br[54] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_57 
+ bl[55] br[55] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_58 
+ bl[56] br[56] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_59 
+ bl[57] br[57] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_60 
+ bl[58] br[58] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_61 
+ bl[59] br[59] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_62 
+ bl[60] br[60] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_63 
+ bl[61] br[61] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_64 
+ bl[62] br[62] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_65 
+ bl[63] br[63] vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_66 
+ vdd vdd vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_294_67 
+ vdd vdd vdd vss wl[292] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_0 
+ vdd vdd vss vdd vpb vnb wl[293] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_295_1 
+ rbl rbr vss vdd vpb vnb wl[293] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_295_2 
+ bl[0] br[0] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_3 
+ bl[1] br[1] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_4 
+ bl[2] br[2] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_5 
+ bl[3] br[3] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_6 
+ bl[4] br[4] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_7 
+ bl[5] br[5] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_8 
+ bl[6] br[6] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_9 
+ bl[7] br[7] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_10 
+ bl[8] br[8] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_11 
+ bl[9] br[9] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_12 
+ bl[10] br[10] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_13 
+ bl[11] br[11] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_14 
+ bl[12] br[12] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_15 
+ bl[13] br[13] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_16 
+ bl[14] br[14] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_17 
+ bl[15] br[15] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_18 
+ bl[16] br[16] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_19 
+ bl[17] br[17] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_20 
+ bl[18] br[18] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_21 
+ bl[19] br[19] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_22 
+ bl[20] br[20] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_23 
+ bl[21] br[21] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_24 
+ bl[22] br[22] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_25 
+ bl[23] br[23] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_26 
+ bl[24] br[24] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_27 
+ bl[25] br[25] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_28 
+ bl[26] br[26] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_29 
+ bl[27] br[27] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_30 
+ bl[28] br[28] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_31 
+ bl[29] br[29] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_32 
+ bl[30] br[30] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_33 
+ bl[31] br[31] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_34 
+ bl[32] br[32] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_35 
+ bl[33] br[33] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_36 
+ bl[34] br[34] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_37 
+ bl[35] br[35] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_38 
+ bl[36] br[36] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_39 
+ bl[37] br[37] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_40 
+ bl[38] br[38] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_41 
+ bl[39] br[39] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_42 
+ bl[40] br[40] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_43 
+ bl[41] br[41] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_44 
+ bl[42] br[42] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_45 
+ bl[43] br[43] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_46 
+ bl[44] br[44] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_47 
+ bl[45] br[45] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_48 
+ bl[46] br[46] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_49 
+ bl[47] br[47] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_50 
+ bl[48] br[48] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_51 
+ bl[49] br[49] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_52 
+ bl[50] br[50] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_53 
+ bl[51] br[51] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_54 
+ bl[52] br[52] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_55 
+ bl[53] br[53] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_56 
+ bl[54] br[54] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_57 
+ bl[55] br[55] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_58 
+ bl[56] br[56] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_59 
+ bl[57] br[57] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_60 
+ bl[58] br[58] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_61 
+ bl[59] br[59] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_62 
+ bl[60] br[60] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_63 
+ bl[61] br[61] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_64 
+ bl[62] br[62] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_65 
+ bl[63] br[63] vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_66 
+ vdd vdd vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_295_67 
+ vdd vdd vdd vss wl[293] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_0 
+ vdd vdd vss vdd vpb vnb wl[294] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_296_1 
+ rbl rbr vss vdd vpb vnb wl[294] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_296_2 
+ bl[0] br[0] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_3 
+ bl[1] br[1] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_4 
+ bl[2] br[2] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_5 
+ bl[3] br[3] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_6 
+ bl[4] br[4] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_7 
+ bl[5] br[5] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_8 
+ bl[6] br[6] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_9 
+ bl[7] br[7] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_10 
+ bl[8] br[8] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_11 
+ bl[9] br[9] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_12 
+ bl[10] br[10] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_13 
+ bl[11] br[11] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_14 
+ bl[12] br[12] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_15 
+ bl[13] br[13] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_16 
+ bl[14] br[14] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_17 
+ bl[15] br[15] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_18 
+ bl[16] br[16] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_19 
+ bl[17] br[17] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_20 
+ bl[18] br[18] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_21 
+ bl[19] br[19] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_22 
+ bl[20] br[20] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_23 
+ bl[21] br[21] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_24 
+ bl[22] br[22] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_25 
+ bl[23] br[23] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_26 
+ bl[24] br[24] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_27 
+ bl[25] br[25] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_28 
+ bl[26] br[26] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_29 
+ bl[27] br[27] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_30 
+ bl[28] br[28] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_31 
+ bl[29] br[29] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_32 
+ bl[30] br[30] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_33 
+ bl[31] br[31] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_34 
+ bl[32] br[32] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_35 
+ bl[33] br[33] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_36 
+ bl[34] br[34] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_37 
+ bl[35] br[35] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_38 
+ bl[36] br[36] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_39 
+ bl[37] br[37] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_40 
+ bl[38] br[38] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_41 
+ bl[39] br[39] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_42 
+ bl[40] br[40] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_43 
+ bl[41] br[41] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_44 
+ bl[42] br[42] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_45 
+ bl[43] br[43] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_46 
+ bl[44] br[44] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_47 
+ bl[45] br[45] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_48 
+ bl[46] br[46] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_49 
+ bl[47] br[47] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_50 
+ bl[48] br[48] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_51 
+ bl[49] br[49] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_52 
+ bl[50] br[50] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_53 
+ bl[51] br[51] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_54 
+ bl[52] br[52] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_55 
+ bl[53] br[53] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_56 
+ bl[54] br[54] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_57 
+ bl[55] br[55] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_58 
+ bl[56] br[56] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_59 
+ bl[57] br[57] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_60 
+ bl[58] br[58] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_61 
+ bl[59] br[59] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_62 
+ bl[60] br[60] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_63 
+ bl[61] br[61] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_64 
+ bl[62] br[62] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_65 
+ bl[63] br[63] vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_66 
+ vdd vdd vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_296_67 
+ vdd vdd vdd vss wl[294] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_0 
+ vdd vdd vss vdd vpb vnb wl[295] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_297_1 
+ rbl rbr vss vdd vpb vnb wl[295] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_297_2 
+ bl[0] br[0] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_3 
+ bl[1] br[1] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_4 
+ bl[2] br[2] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_5 
+ bl[3] br[3] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_6 
+ bl[4] br[4] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_7 
+ bl[5] br[5] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_8 
+ bl[6] br[6] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_9 
+ bl[7] br[7] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_10 
+ bl[8] br[8] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_11 
+ bl[9] br[9] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_12 
+ bl[10] br[10] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_13 
+ bl[11] br[11] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_14 
+ bl[12] br[12] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_15 
+ bl[13] br[13] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_16 
+ bl[14] br[14] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_17 
+ bl[15] br[15] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_18 
+ bl[16] br[16] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_19 
+ bl[17] br[17] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_20 
+ bl[18] br[18] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_21 
+ bl[19] br[19] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_22 
+ bl[20] br[20] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_23 
+ bl[21] br[21] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_24 
+ bl[22] br[22] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_25 
+ bl[23] br[23] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_26 
+ bl[24] br[24] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_27 
+ bl[25] br[25] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_28 
+ bl[26] br[26] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_29 
+ bl[27] br[27] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_30 
+ bl[28] br[28] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_31 
+ bl[29] br[29] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_32 
+ bl[30] br[30] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_33 
+ bl[31] br[31] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_34 
+ bl[32] br[32] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_35 
+ bl[33] br[33] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_36 
+ bl[34] br[34] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_37 
+ bl[35] br[35] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_38 
+ bl[36] br[36] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_39 
+ bl[37] br[37] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_40 
+ bl[38] br[38] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_41 
+ bl[39] br[39] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_42 
+ bl[40] br[40] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_43 
+ bl[41] br[41] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_44 
+ bl[42] br[42] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_45 
+ bl[43] br[43] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_46 
+ bl[44] br[44] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_47 
+ bl[45] br[45] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_48 
+ bl[46] br[46] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_49 
+ bl[47] br[47] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_50 
+ bl[48] br[48] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_51 
+ bl[49] br[49] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_52 
+ bl[50] br[50] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_53 
+ bl[51] br[51] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_54 
+ bl[52] br[52] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_55 
+ bl[53] br[53] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_56 
+ bl[54] br[54] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_57 
+ bl[55] br[55] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_58 
+ bl[56] br[56] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_59 
+ bl[57] br[57] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_60 
+ bl[58] br[58] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_61 
+ bl[59] br[59] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_62 
+ bl[60] br[60] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_63 
+ bl[61] br[61] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_64 
+ bl[62] br[62] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_65 
+ bl[63] br[63] vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_66 
+ vdd vdd vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_297_67 
+ vdd vdd vdd vss wl[295] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_0 
+ vdd vdd vss vdd vpb vnb wl[296] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_298_1 
+ rbl rbr vss vdd vpb vnb wl[296] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_298_2 
+ bl[0] br[0] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_3 
+ bl[1] br[1] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_4 
+ bl[2] br[2] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_5 
+ bl[3] br[3] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_6 
+ bl[4] br[4] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_7 
+ bl[5] br[5] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_8 
+ bl[6] br[6] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_9 
+ bl[7] br[7] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_10 
+ bl[8] br[8] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_11 
+ bl[9] br[9] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_12 
+ bl[10] br[10] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_13 
+ bl[11] br[11] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_14 
+ bl[12] br[12] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_15 
+ bl[13] br[13] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_16 
+ bl[14] br[14] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_17 
+ bl[15] br[15] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_18 
+ bl[16] br[16] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_19 
+ bl[17] br[17] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_20 
+ bl[18] br[18] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_21 
+ bl[19] br[19] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_22 
+ bl[20] br[20] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_23 
+ bl[21] br[21] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_24 
+ bl[22] br[22] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_25 
+ bl[23] br[23] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_26 
+ bl[24] br[24] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_27 
+ bl[25] br[25] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_28 
+ bl[26] br[26] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_29 
+ bl[27] br[27] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_30 
+ bl[28] br[28] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_31 
+ bl[29] br[29] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_32 
+ bl[30] br[30] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_33 
+ bl[31] br[31] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_34 
+ bl[32] br[32] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_35 
+ bl[33] br[33] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_36 
+ bl[34] br[34] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_37 
+ bl[35] br[35] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_38 
+ bl[36] br[36] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_39 
+ bl[37] br[37] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_40 
+ bl[38] br[38] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_41 
+ bl[39] br[39] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_42 
+ bl[40] br[40] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_43 
+ bl[41] br[41] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_44 
+ bl[42] br[42] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_45 
+ bl[43] br[43] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_46 
+ bl[44] br[44] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_47 
+ bl[45] br[45] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_48 
+ bl[46] br[46] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_49 
+ bl[47] br[47] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_50 
+ bl[48] br[48] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_51 
+ bl[49] br[49] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_52 
+ bl[50] br[50] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_53 
+ bl[51] br[51] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_54 
+ bl[52] br[52] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_55 
+ bl[53] br[53] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_56 
+ bl[54] br[54] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_57 
+ bl[55] br[55] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_58 
+ bl[56] br[56] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_59 
+ bl[57] br[57] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_60 
+ bl[58] br[58] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_61 
+ bl[59] br[59] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_62 
+ bl[60] br[60] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_63 
+ bl[61] br[61] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_64 
+ bl[62] br[62] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_65 
+ bl[63] br[63] vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_66 
+ vdd vdd vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_298_67 
+ vdd vdd vdd vss wl[296] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_0 
+ vdd vdd vss vdd vpb vnb wl[297] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_299_1 
+ rbl rbr vss vdd vpb vnb wl[297] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_299_2 
+ bl[0] br[0] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_3 
+ bl[1] br[1] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_4 
+ bl[2] br[2] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_5 
+ bl[3] br[3] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_6 
+ bl[4] br[4] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_7 
+ bl[5] br[5] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_8 
+ bl[6] br[6] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_9 
+ bl[7] br[7] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_10 
+ bl[8] br[8] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_11 
+ bl[9] br[9] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_12 
+ bl[10] br[10] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_13 
+ bl[11] br[11] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_14 
+ bl[12] br[12] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_15 
+ bl[13] br[13] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_16 
+ bl[14] br[14] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_17 
+ bl[15] br[15] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_18 
+ bl[16] br[16] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_19 
+ bl[17] br[17] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_20 
+ bl[18] br[18] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_21 
+ bl[19] br[19] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_22 
+ bl[20] br[20] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_23 
+ bl[21] br[21] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_24 
+ bl[22] br[22] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_25 
+ bl[23] br[23] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_26 
+ bl[24] br[24] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_27 
+ bl[25] br[25] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_28 
+ bl[26] br[26] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_29 
+ bl[27] br[27] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_30 
+ bl[28] br[28] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_31 
+ bl[29] br[29] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_32 
+ bl[30] br[30] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_33 
+ bl[31] br[31] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_34 
+ bl[32] br[32] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_35 
+ bl[33] br[33] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_36 
+ bl[34] br[34] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_37 
+ bl[35] br[35] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_38 
+ bl[36] br[36] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_39 
+ bl[37] br[37] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_40 
+ bl[38] br[38] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_41 
+ bl[39] br[39] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_42 
+ bl[40] br[40] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_43 
+ bl[41] br[41] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_44 
+ bl[42] br[42] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_45 
+ bl[43] br[43] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_46 
+ bl[44] br[44] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_47 
+ bl[45] br[45] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_48 
+ bl[46] br[46] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_49 
+ bl[47] br[47] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_50 
+ bl[48] br[48] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_51 
+ bl[49] br[49] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_52 
+ bl[50] br[50] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_53 
+ bl[51] br[51] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_54 
+ bl[52] br[52] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_55 
+ bl[53] br[53] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_56 
+ bl[54] br[54] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_57 
+ bl[55] br[55] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_58 
+ bl[56] br[56] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_59 
+ bl[57] br[57] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_60 
+ bl[58] br[58] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_61 
+ bl[59] br[59] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_62 
+ bl[60] br[60] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_63 
+ bl[61] br[61] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_64 
+ bl[62] br[62] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_65 
+ bl[63] br[63] vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_66 
+ vdd vdd vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_299_67 
+ vdd vdd vdd vss wl[297] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_0 
+ vdd vdd vss vdd vpb vnb wl[298] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_300_1 
+ rbl rbr vss vdd vpb vnb wl[298] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_300_2 
+ bl[0] br[0] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_3 
+ bl[1] br[1] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_4 
+ bl[2] br[2] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_5 
+ bl[3] br[3] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_6 
+ bl[4] br[4] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_7 
+ bl[5] br[5] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_8 
+ bl[6] br[6] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_9 
+ bl[7] br[7] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_10 
+ bl[8] br[8] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_11 
+ bl[9] br[9] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_12 
+ bl[10] br[10] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_13 
+ bl[11] br[11] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_14 
+ bl[12] br[12] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_15 
+ bl[13] br[13] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_16 
+ bl[14] br[14] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_17 
+ bl[15] br[15] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_18 
+ bl[16] br[16] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_19 
+ bl[17] br[17] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_20 
+ bl[18] br[18] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_21 
+ bl[19] br[19] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_22 
+ bl[20] br[20] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_23 
+ bl[21] br[21] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_24 
+ bl[22] br[22] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_25 
+ bl[23] br[23] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_26 
+ bl[24] br[24] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_27 
+ bl[25] br[25] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_28 
+ bl[26] br[26] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_29 
+ bl[27] br[27] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_30 
+ bl[28] br[28] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_31 
+ bl[29] br[29] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_32 
+ bl[30] br[30] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_33 
+ bl[31] br[31] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_34 
+ bl[32] br[32] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_35 
+ bl[33] br[33] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_36 
+ bl[34] br[34] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_37 
+ bl[35] br[35] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_38 
+ bl[36] br[36] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_39 
+ bl[37] br[37] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_40 
+ bl[38] br[38] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_41 
+ bl[39] br[39] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_42 
+ bl[40] br[40] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_43 
+ bl[41] br[41] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_44 
+ bl[42] br[42] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_45 
+ bl[43] br[43] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_46 
+ bl[44] br[44] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_47 
+ bl[45] br[45] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_48 
+ bl[46] br[46] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_49 
+ bl[47] br[47] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_50 
+ bl[48] br[48] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_51 
+ bl[49] br[49] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_52 
+ bl[50] br[50] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_53 
+ bl[51] br[51] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_54 
+ bl[52] br[52] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_55 
+ bl[53] br[53] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_56 
+ bl[54] br[54] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_57 
+ bl[55] br[55] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_58 
+ bl[56] br[56] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_59 
+ bl[57] br[57] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_60 
+ bl[58] br[58] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_61 
+ bl[59] br[59] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_62 
+ bl[60] br[60] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_63 
+ bl[61] br[61] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_64 
+ bl[62] br[62] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_65 
+ bl[63] br[63] vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_66 
+ vdd vdd vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_300_67 
+ vdd vdd vdd vss wl[298] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_0 
+ vdd vdd vss vdd vpb vnb wl[299] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_301_1 
+ rbl rbr vss vdd vpb vnb wl[299] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_301_2 
+ bl[0] br[0] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_3 
+ bl[1] br[1] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_4 
+ bl[2] br[2] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_5 
+ bl[3] br[3] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_6 
+ bl[4] br[4] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_7 
+ bl[5] br[5] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_8 
+ bl[6] br[6] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_9 
+ bl[7] br[7] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_10 
+ bl[8] br[8] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_11 
+ bl[9] br[9] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_12 
+ bl[10] br[10] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_13 
+ bl[11] br[11] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_14 
+ bl[12] br[12] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_15 
+ bl[13] br[13] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_16 
+ bl[14] br[14] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_17 
+ bl[15] br[15] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_18 
+ bl[16] br[16] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_19 
+ bl[17] br[17] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_20 
+ bl[18] br[18] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_21 
+ bl[19] br[19] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_22 
+ bl[20] br[20] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_23 
+ bl[21] br[21] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_24 
+ bl[22] br[22] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_25 
+ bl[23] br[23] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_26 
+ bl[24] br[24] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_27 
+ bl[25] br[25] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_28 
+ bl[26] br[26] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_29 
+ bl[27] br[27] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_30 
+ bl[28] br[28] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_31 
+ bl[29] br[29] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_32 
+ bl[30] br[30] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_33 
+ bl[31] br[31] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_34 
+ bl[32] br[32] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_35 
+ bl[33] br[33] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_36 
+ bl[34] br[34] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_37 
+ bl[35] br[35] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_38 
+ bl[36] br[36] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_39 
+ bl[37] br[37] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_40 
+ bl[38] br[38] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_41 
+ bl[39] br[39] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_42 
+ bl[40] br[40] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_43 
+ bl[41] br[41] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_44 
+ bl[42] br[42] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_45 
+ bl[43] br[43] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_46 
+ bl[44] br[44] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_47 
+ bl[45] br[45] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_48 
+ bl[46] br[46] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_49 
+ bl[47] br[47] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_50 
+ bl[48] br[48] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_51 
+ bl[49] br[49] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_52 
+ bl[50] br[50] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_53 
+ bl[51] br[51] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_54 
+ bl[52] br[52] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_55 
+ bl[53] br[53] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_56 
+ bl[54] br[54] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_57 
+ bl[55] br[55] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_58 
+ bl[56] br[56] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_59 
+ bl[57] br[57] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_60 
+ bl[58] br[58] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_61 
+ bl[59] br[59] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_62 
+ bl[60] br[60] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_63 
+ bl[61] br[61] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_64 
+ bl[62] br[62] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_65 
+ bl[63] br[63] vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_66 
+ vdd vdd vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_301_67 
+ vdd vdd vdd vss wl[299] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_0 
+ vdd vdd vss vdd vpb vnb wl[300] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_302_1 
+ rbl rbr vss vdd vpb vnb wl[300] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_302_2 
+ bl[0] br[0] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_3 
+ bl[1] br[1] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_4 
+ bl[2] br[2] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_5 
+ bl[3] br[3] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_6 
+ bl[4] br[4] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_7 
+ bl[5] br[5] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_8 
+ bl[6] br[6] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_9 
+ bl[7] br[7] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_10 
+ bl[8] br[8] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_11 
+ bl[9] br[9] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_12 
+ bl[10] br[10] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_13 
+ bl[11] br[11] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_14 
+ bl[12] br[12] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_15 
+ bl[13] br[13] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_16 
+ bl[14] br[14] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_17 
+ bl[15] br[15] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_18 
+ bl[16] br[16] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_19 
+ bl[17] br[17] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_20 
+ bl[18] br[18] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_21 
+ bl[19] br[19] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_22 
+ bl[20] br[20] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_23 
+ bl[21] br[21] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_24 
+ bl[22] br[22] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_25 
+ bl[23] br[23] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_26 
+ bl[24] br[24] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_27 
+ bl[25] br[25] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_28 
+ bl[26] br[26] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_29 
+ bl[27] br[27] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_30 
+ bl[28] br[28] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_31 
+ bl[29] br[29] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_32 
+ bl[30] br[30] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_33 
+ bl[31] br[31] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_34 
+ bl[32] br[32] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_35 
+ bl[33] br[33] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_36 
+ bl[34] br[34] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_37 
+ bl[35] br[35] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_38 
+ bl[36] br[36] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_39 
+ bl[37] br[37] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_40 
+ bl[38] br[38] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_41 
+ bl[39] br[39] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_42 
+ bl[40] br[40] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_43 
+ bl[41] br[41] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_44 
+ bl[42] br[42] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_45 
+ bl[43] br[43] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_46 
+ bl[44] br[44] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_47 
+ bl[45] br[45] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_48 
+ bl[46] br[46] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_49 
+ bl[47] br[47] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_50 
+ bl[48] br[48] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_51 
+ bl[49] br[49] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_52 
+ bl[50] br[50] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_53 
+ bl[51] br[51] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_54 
+ bl[52] br[52] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_55 
+ bl[53] br[53] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_56 
+ bl[54] br[54] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_57 
+ bl[55] br[55] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_58 
+ bl[56] br[56] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_59 
+ bl[57] br[57] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_60 
+ bl[58] br[58] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_61 
+ bl[59] br[59] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_62 
+ bl[60] br[60] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_63 
+ bl[61] br[61] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_64 
+ bl[62] br[62] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_65 
+ bl[63] br[63] vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_66 
+ vdd vdd vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_302_67 
+ vdd vdd vdd vss wl[300] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_0 
+ vdd vdd vss vdd vpb vnb wl[301] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_303_1 
+ rbl rbr vss vdd vpb vnb wl[301] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_303_2 
+ bl[0] br[0] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_3 
+ bl[1] br[1] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_4 
+ bl[2] br[2] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_5 
+ bl[3] br[3] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_6 
+ bl[4] br[4] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_7 
+ bl[5] br[5] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_8 
+ bl[6] br[6] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_9 
+ bl[7] br[7] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_10 
+ bl[8] br[8] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_11 
+ bl[9] br[9] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_12 
+ bl[10] br[10] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_13 
+ bl[11] br[11] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_14 
+ bl[12] br[12] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_15 
+ bl[13] br[13] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_16 
+ bl[14] br[14] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_17 
+ bl[15] br[15] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_18 
+ bl[16] br[16] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_19 
+ bl[17] br[17] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_20 
+ bl[18] br[18] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_21 
+ bl[19] br[19] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_22 
+ bl[20] br[20] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_23 
+ bl[21] br[21] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_24 
+ bl[22] br[22] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_25 
+ bl[23] br[23] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_26 
+ bl[24] br[24] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_27 
+ bl[25] br[25] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_28 
+ bl[26] br[26] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_29 
+ bl[27] br[27] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_30 
+ bl[28] br[28] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_31 
+ bl[29] br[29] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_32 
+ bl[30] br[30] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_33 
+ bl[31] br[31] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_34 
+ bl[32] br[32] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_35 
+ bl[33] br[33] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_36 
+ bl[34] br[34] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_37 
+ bl[35] br[35] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_38 
+ bl[36] br[36] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_39 
+ bl[37] br[37] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_40 
+ bl[38] br[38] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_41 
+ bl[39] br[39] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_42 
+ bl[40] br[40] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_43 
+ bl[41] br[41] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_44 
+ bl[42] br[42] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_45 
+ bl[43] br[43] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_46 
+ bl[44] br[44] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_47 
+ bl[45] br[45] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_48 
+ bl[46] br[46] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_49 
+ bl[47] br[47] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_50 
+ bl[48] br[48] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_51 
+ bl[49] br[49] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_52 
+ bl[50] br[50] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_53 
+ bl[51] br[51] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_54 
+ bl[52] br[52] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_55 
+ bl[53] br[53] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_56 
+ bl[54] br[54] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_57 
+ bl[55] br[55] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_58 
+ bl[56] br[56] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_59 
+ bl[57] br[57] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_60 
+ bl[58] br[58] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_61 
+ bl[59] br[59] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_62 
+ bl[60] br[60] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_63 
+ bl[61] br[61] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_64 
+ bl[62] br[62] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_65 
+ bl[63] br[63] vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_66 
+ vdd vdd vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_303_67 
+ vdd vdd vdd vss wl[301] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_0 
+ vdd vdd vss vdd vpb vnb wl[302] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_304_1 
+ rbl rbr vss vdd vpb vnb wl[302] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_304_2 
+ bl[0] br[0] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_3 
+ bl[1] br[1] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_4 
+ bl[2] br[2] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_5 
+ bl[3] br[3] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_6 
+ bl[4] br[4] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_7 
+ bl[5] br[5] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_8 
+ bl[6] br[6] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_9 
+ bl[7] br[7] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_10 
+ bl[8] br[8] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_11 
+ bl[9] br[9] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_12 
+ bl[10] br[10] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_13 
+ bl[11] br[11] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_14 
+ bl[12] br[12] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_15 
+ bl[13] br[13] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_16 
+ bl[14] br[14] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_17 
+ bl[15] br[15] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_18 
+ bl[16] br[16] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_19 
+ bl[17] br[17] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_20 
+ bl[18] br[18] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_21 
+ bl[19] br[19] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_22 
+ bl[20] br[20] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_23 
+ bl[21] br[21] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_24 
+ bl[22] br[22] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_25 
+ bl[23] br[23] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_26 
+ bl[24] br[24] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_27 
+ bl[25] br[25] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_28 
+ bl[26] br[26] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_29 
+ bl[27] br[27] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_30 
+ bl[28] br[28] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_31 
+ bl[29] br[29] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_32 
+ bl[30] br[30] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_33 
+ bl[31] br[31] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_34 
+ bl[32] br[32] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_35 
+ bl[33] br[33] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_36 
+ bl[34] br[34] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_37 
+ bl[35] br[35] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_38 
+ bl[36] br[36] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_39 
+ bl[37] br[37] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_40 
+ bl[38] br[38] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_41 
+ bl[39] br[39] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_42 
+ bl[40] br[40] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_43 
+ bl[41] br[41] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_44 
+ bl[42] br[42] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_45 
+ bl[43] br[43] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_46 
+ bl[44] br[44] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_47 
+ bl[45] br[45] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_48 
+ bl[46] br[46] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_49 
+ bl[47] br[47] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_50 
+ bl[48] br[48] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_51 
+ bl[49] br[49] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_52 
+ bl[50] br[50] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_53 
+ bl[51] br[51] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_54 
+ bl[52] br[52] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_55 
+ bl[53] br[53] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_56 
+ bl[54] br[54] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_57 
+ bl[55] br[55] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_58 
+ bl[56] br[56] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_59 
+ bl[57] br[57] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_60 
+ bl[58] br[58] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_61 
+ bl[59] br[59] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_62 
+ bl[60] br[60] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_63 
+ bl[61] br[61] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_64 
+ bl[62] br[62] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_65 
+ bl[63] br[63] vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_66 
+ vdd vdd vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_304_67 
+ vdd vdd vdd vss wl[302] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_0 
+ vdd vdd vss vdd vpb vnb wl[303] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_305_1 
+ rbl rbr vss vdd vpb vnb wl[303] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_305_2 
+ bl[0] br[0] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_3 
+ bl[1] br[1] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_4 
+ bl[2] br[2] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_5 
+ bl[3] br[3] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_6 
+ bl[4] br[4] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_7 
+ bl[5] br[5] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_8 
+ bl[6] br[6] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_9 
+ bl[7] br[7] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_10 
+ bl[8] br[8] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_11 
+ bl[9] br[9] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_12 
+ bl[10] br[10] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_13 
+ bl[11] br[11] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_14 
+ bl[12] br[12] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_15 
+ bl[13] br[13] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_16 
+ bl[14] br[14] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_17 
+ bl[15] br[15] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_18 
+ bl[16] br[16] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_19 
+ bl[17] br[17] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_20 
+ bl[18] br[18] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_21 
+ bl[19] br[19] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_22 
+ bl[20] br[20] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_23 
+ bl[21] br[21] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_24 
+ bl[22] br[22] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_25 
+ bl[23] br[23] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_26 
+ bl[24] br[24] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_27 
+ bl[25] br[25] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_28 
+ bl[26] br[26] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_29 
+ bl[27] br[27] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_30 
+ bl[28] br[28] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_31 
+ bl[29] br[29] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_32 
+ bl[30] br[30] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_33 
+ bl[31] br[31] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_34 
+ bl[32] br[32] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_35 
+ bl[33] br[33] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_36 
+ bl[34] br[34] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_37 
+ bl[35] br[35] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_38 
+ bl[36] br[36] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_39 
+ bl[37] br[37] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_40 
+ bl[38] br[38] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_41 
+ bl[39] br[39] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_42 
+ bl[40] br[40] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_43 
+ bl[41] br[41] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_44 
+ bl[42] br[42] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_45 
+ bl[43] br[43] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_46 
+ bl[44] br[44] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_47 
+ bl[45] br[45] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_48 
+ bl[46] br[46] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_49 
+ bl[47] br[47] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_50 
+ bl[48] br[48] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_51 
+ bl[49] br[49] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_52 
+ bl[50] br[50] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_53 
+ bl[51] br[51] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_54 
+ bl[52] br[52] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_55 
+ bl[53] br[53] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_56 
+ bl[54] br[54] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_57 
+ bl[55] br[55] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_58 
+ bl[56] br[56] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_59 
+ bl[57] br[57] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_60 
+ bl[58] br[58] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_61 
+ bl[59] br[59] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_62 
+ bl[60] br[60] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_63 
+ bl[61] br[61] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_64 
+ bl[62] br[62] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_65 
+ bl[63] br[63] vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_66 
+ vdd vdd vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_305_67 
+ vdd vdd vdd vss wl[303] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_0 
+ vdd vdd vss vdd vpb vnb wl[304] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_306_1 
+ rbl rbr vss vdd vpb vnb wl[304] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_306_2 
+ bl[0] br[0] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_3 
+ bl[1] br[1] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_4 
+ bl[2] br[2] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_5 
+ bl[3] br[3] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_6 
+ bl[4] br[4] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_7 
+ bl[5] br[5] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_8 
+ bl[6] br[6] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_9 
+ bl[7] br[7] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_10 
+ bl[8] br[8] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_11 
+ bl[9] br[9] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_12 
+ bl[10] br[10] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_13 
+ bl[11] br[11] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_14 
+ bl[12] br[12] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_15 
+ bl[13] br[13] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_16 
+ bl[14] br[14] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_17 
+ bl[15] br[15] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_18 
+ bl[16] br[16] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_19 
+ bl[17] br[17] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_20 
+ bl[18] br[18] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_21 
+ bl[19] br[19] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_22 
+ bl[20] br[20] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_23 
+ bl[21] br[21] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_24 
+ bl[22] br[22] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_25 
+ bl[23] br[23] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_26 
+ bl[24] br[24] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_27 
+ bl[25] br[25] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_28 
+ bl[26] br[26] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_29 
+ bl[27] br[27] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_30 
+ bl[28] br[28] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_31 
+ bl[29] br[29] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_32 
+ bl[30] br[30] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_33 
+ bl[31] br[31] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_34 
+ bl[32] br[32] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_35 
+ bl[33] br[33] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_36 
+ bl[34] br[34] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_37 
+ bl[35] br[35] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_38 
+ bl[36] br[36] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_39 
+ bl[37] br[37] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_40 
+ bl[38] br[38] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_41 
+ bl[39] br[39] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_42 
+ bl[40] br[40] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_43 
+ bl[41] br[41] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_44 
+ bl[42] br[42] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_45 
+ bl[43] br[43] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_46 
+ bl[44] br[44] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_47 
+ bl[45] br[45] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_48 
+ bl[46] br[46] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_49 
+ bl[47] br[47] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_50 
+ bl[48] br[48] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_51 
+ bl[49] br[49] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_52 
+ bl[50] br[50] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_53 
+ bl[51] br[51] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_54 
+ bl[52] br[52] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_55 
+ bl[53] br[53] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_56 
+ bl[54] br[54] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_57 
+ bl[55] br[55] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_58 
+ bl[56] br[56] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_59 
+ bl[57] br[57] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_60 
+ bl[58] br[58] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_61 
+ bl[59] br[59] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_62 
+ bl[60] br[60] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_63 
+ bl[61] br[61] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_64 
+ bl[62] br[62] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_65 
+ bl[63] br[63] vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_66 
+ vdd vdd vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_306_67 
+ vdd vdd vdd vss wl[304] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_0 
+ vdd vdd vss vdd vpb vnb wl[305] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_307_1 
+ rbl rbr vss vdd vpb vnb wl[305] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_307_2 
+ bl[0] br[0] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_3 
+ bl[1] br[1] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_4 
+ bl[2] br[2] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_5 
+ bl[3] br[3] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_6 
+ bl[4] br[4] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_7 
+ bl[5] br[5] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_8 
+ bl[6] br[6] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_9 
+ bl[7] br[7] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_10 
+ bl[8] br[8] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_11 
+ bl[9] br[9] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_12 
+ bl[10] br[10] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_13 
+ bl[11] br[11] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_14 
+ bl[12] br[12] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_15 
+ bl[13] br[13] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_16 
+ bl[14] br[14] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_17 
+ bl[15] br[15] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_18 
+ bl[16] br[16] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_19 
+ bl[17] br[17] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_20 
+ bl[18] br[18] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_21 
+ bl[19] br[19] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_22 
+ bl[20] br[20] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_23 
+ bl[21] br[21] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_24 
+ bl[22] br[22] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_25 
+ bl[23] br[23] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_26 
+ bl[24] br[24] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_27 
+ bl[25] br[25] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_28 
+ bl[26] br[26] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_29 
+ bl[27] br[27] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_30 
+ bl[28] br[28] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_31 
+ bl[29] br[29] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_32 
+ bl[30] br[30] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_33 
+ bl[31] br[31] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_34 
+ bl[32] br[32] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_35 
+ bl[33] br[33] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_36 
+ bl[34] br[34] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_37 
+ bl[35] br[35] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_38 
+ bl[36] br[36] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_39 
+ bl[37] br[37] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_40 
+ bl[38] br[38] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_41 
+ bl[39] br[39] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_42 
+ bl[40] br[40] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_43 
+ bl[41] br[41] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_44 
+ bl[42] br[42] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_45 
+ bl[43] br[43] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_46 
+ bl[44] br[44] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_47 
+ bl[45] br[45] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_48 
+ bl[46] br[46] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_49 
+ bl[47] br[47] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_50 
+ bl[48] br[48] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_51 
+ bl[49] br[49] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_52 
+ bl[50] br[50] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_53 
+ bl[51] br[51] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_54 
+ bl[52] br[52] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_55 
+ bl[53] br[53] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_56 
+ bl[54] br[54] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_57 
+ bl[55] br[55] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_58 
+ bl[56] br[56] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_59 
+ bl[57] br[57] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_60 
+ bl[58] br[58] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_61 
+ bl[59] br[59] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_62 
+ bl[60] br[60] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_63 
+ bl[61] br[61] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_64 
+ bl[62] br[62] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_65 
+ bl[63] br[63] vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_66 
+ vdd vdd vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_307_67 
+ vdd vdd vdd vss wl[305] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_0 
+ vdd vdd vss vdd vpb vnb wl[306] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_308_1 
+ rbl rbr vss vdd vpb vnb wl[306] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_308_2 
+ bl[0] br[0] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_3 
+ bl[1] br[1] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_4 
+ bl[2] br[2] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_5 
+ bl[3] br[3] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_6 
+ bl[4] br[4] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_7 
+ bl[5] br[5] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_8 
+ bl[6] br[6] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_9 
+ bl[7] br[7] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_10 
+ bl[8] br[8] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_11 
+ bl[9] br[9] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_12 
+ bl[10] br[10] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_13 
+ bl[11] br[11] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_14 
+ bl[12] br[12] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_15 
+ bl[13] br[13] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_16 
+ bl[14] br[14] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_17 
+ bl[15] br[15] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_18 
+ bl[16] br[16] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_19 
+ bl[17] br[17] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_20 
+ bl[18] br[18] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_21 
+ bl[19] br[19] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_22 
+ bl[20] br[20] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_23 
+ bl[21] br[21] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_24 
+ bl[22] br[22] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_25 
+ bl[23] br[23] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_26 
+ bl[24] br[24] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_27 
+ bl[25] br[25] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_28 
+ bl[26] br[26] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_29 
+ bl[27] br[27] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_30 
+ bl[28] br[28] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_31 
+ bl[29] br[29] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_32 
+ bl[30] br[30] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_33 
+ bl[31] br[31] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_34 
+ bl[32] br[32] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_35 
+ bl[33] br[33] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_36 
+ bl[34] br[34] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_37 
+ bl[35] br[35] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_38 
+ bl[36] br[36] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_39 
+ bl[37] br[37] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_40 
+ bl[38] br[38] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_41 
+ bl[39] br[39] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_42 
+ bl[40] br[40] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_43 
+ bl[41] br[41] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_44 
+ bl[42] br[42] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_45 
+ bl[43] br[43] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_46 
+ bl[44] br[44] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_47 
+ bl[45] br[45] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_48 
+ bl[46] br[46] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_49 
+ bl[47] br[47] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_50 
+ bl[48] br[48] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_51 
+ bl[49] br[49] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_52 
+ bl[50] br[50] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_53 
+ bl[51] br[51] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_54 
+ bl[52] br[52] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_55 
+ bl[53] br[53] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_56 
+ bl[54] br[54] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_57 
+ bl[55] br[55] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_58 
+ bl[56] br[56] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_59 
+ bl[57] br[57] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_60 
+ bl[58] br[58] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_61 
+ bl[59] br[59] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_62 
+ bl[60] br[60] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_63 
+ bl[61] br[61] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_64 
+ bl[62] br[62] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_65 
+ bl[63] br[63] vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_66 
+ vdd vdd vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_308_67 
+ vdd vdd vdd vss wl[306] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_0 
+ vdd vdd vss vdd vpb vnb wl[307] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_309_1 
+ rbl rbr vss vdd vpb vnb wl[307] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_309_2 
+ bl[0] br[0] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_3 
+ bl[1] br[1] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_4 
+ bl[2] br[2] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_5 
+ bl[3] br[3] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_6 
+ bl[4] br[4] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_7 
+ bl[5] br[5] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_8 
+ bl[6] br[6] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_9 
+ bl[7] br[7] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_10 
+ bl[8] br[8] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_11 
+ bl[9] br[9] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_12 
+ bl[10] br[10] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_13 
+ bl[11] br[11] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_14 
+ bl[12] br[12] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_15 
+ bl[13] br[13] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_16 
+ bl[14] br[14] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_17 
+ bl[15] br[15] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_18 
+ bl[16] br[16] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_19 
+ bl[17] br[17] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_20 
+ bl[18] br[18] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_21 
+ bl[19] br[19] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_22 
+ bl[20] br[20] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_23 
+ bl[21] br[21] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_24 
+ bl[22] br[22] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_25 
+ bl[23] br[23] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_26 
+ bl[24] br[24] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_27 
+ bl[25] br[25] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_28 
+ bl[26] br[26] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_29 
+ bl[27] br[27] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_30 
+ bl[28] br[28] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_31 
+ bl[29] br[29] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_32 
+ bl[30] br[30] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_33 
+ bl[31] br[31] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_34 
+ bl[32] br[32] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_35 
+ bl[33] br[33] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_36 
+ bl[34] br[34] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_37 
+ bl[35] br[35] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_38 
+ bl[36] br[36] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_39 
+ bl[37] br[37] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_40 
+ bl[38] br[38] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_41 
+ bl[39] br[39] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_42 
+ bl[40] br[40] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_43 
+ bl[41] br[41] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_44 
+ bl[42] br[42] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_45 
+ bl[43] br[43] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_46 
+ bl[44] br[44] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_47 
+ bl[45] br[45] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_48 
+ bl[46] br[46] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_49 
+ bl[47] br[47] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_50 
+ bl[48] br[48] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_51 
+ bl[49] br[49] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_52 
+ bl[50] br[50] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_53 
+ bl[51] br[51] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_54 
+ bl[52] br[52] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_55 
+ bl[53] br[53] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_56 
+ bl[54] br[54] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_57 
+ bl[55] br[55] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_58 
+ bl[56] br[56] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_59 
+ bl[57] br[57] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_60 
+ bl[58] br[58] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_61 
+ bl[59] br[59] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_62 
+ bl[60] br[60] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_63 
+ bl[61] br[61] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_64 
+ bl[62] br[62] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_65 
+ bl[63] br[63] vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_66 
+ vdd vdd vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_309_67 
+ vdd vdd vdd vss wl[307] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_0 
+ vdd vdd vss vdd vpb vnb wl[308] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_310_1 
+ rbl rbr vss vdd vpb vnb wl[308] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_310_2 
+ bl[0] br[0] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_3 
+ bl[1] br[1] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_4 
+ bl[2] br[2] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_5 
+ bl[3] br[3] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_6 
+ bl[4] br[4] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_7 
+ bl[5] br[5] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_8 
+ bl[6] br[6] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_9 
+ bl[7] br[7] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_10 
+ bl[8] br[8] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_11 
+ bl[9] br[9] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_12 
+ bl[10] br[10] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_13 
+ bl[11] br[11] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_14 
+ bl[12] br[12] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_15 
+ bl[13] br[13] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_16 
+ bl[14] br[14] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_17 
+ bl[15] br[15] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_18 
+ bl[16] br[16] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_19 
+ bl[17] br[17] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_20 
+ bl[18] br[18] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_21 
+ bl[19] br[19] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_22 
+ bl[20] br[20] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_23 
+ bl[21] br[21] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_24 
+ bl[22] br[22] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_25 
+ bl[23] br[23] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_26 
+ bl[24] br[24] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_27 
+ bl[25] br[25] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_28 
+ bl[26] br[26] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_29 
+ bl[27] br[27] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_30 
+ bl[28] br[28] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_31 
+ bl[29] br[29] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_32 
+ bl[30] br[30] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_33 
+ bl[31] br[31] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_34 
+ bl[32] br[32] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_35 
+ bl[33] br[33] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_36 
+ bl[34] br[34] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_37 
+ bl[35] br[35] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_38 
+ bl[36] br[36] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_39 
+ bl[37] br[37] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_40 
+ bl[38] br[38] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_41 
+ bl[39] br[39] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_42 
+ bl[40] br[40] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_43 
+ bl[41] br[41] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_44 
+ bl[42] br[42] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_45 
+ bl[43] br[43] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_46 
+ bl[44] br[44] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_47 
+ bl[45] br[45] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_48 
+ bl[46] br[46] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_49 
+ bl[47] br[47] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_50 
+ bl[48] br[48] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_51 
+ bl[49] br[49] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_52 
+ bl[50] br[50] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_53 
+ bl[51] br[51] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_54 
+ bl[52] br[52] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_55 
+ bl[53] br[53] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_56 
+ bl[54] br[54] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_57 
+ bl[55] br[55] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_58 
+ bl[56] br[56] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_59 
+ bl[57] br[57] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_60 
+ bl[58] br[58] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_61 
+ bl[59] br[59] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_62 
+ bl[60] br[60] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_63 
+ bl[61] br[61] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_64 
+ bl[62] br[62] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_65 
+ bl[63] br[63] vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_66 
+ vdd vdd vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_310_67 
+ vdd vdd vdd vss wl[308] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_0 
+ vdd vdd vss vdd vpb vnb wl[309] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_311_1 
+ rbl rbr vss vdd vpb vnb wl[309] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_311_2 
+ bl[0] br[0] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_3 
+ bl[1] br[1] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_4 
+ bl[2] br[2] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_5 
+ bl[3] br[3] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_6 
+ bl[4] br[4] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_7 
+ bl[5] br[5] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_8 
+ bl[6] br[6] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_9 
+ bl[7] br[7] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_10 
+ bl[8] br[8] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_11 
+ bl[9] br[9] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_12 
+ bl[10] br[10] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_13 
+ bl[11] br[11] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_14 
+ bl[12] br[12] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_15 
+ bl[13] br[13] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_16 
+ bl[14] br[14] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_17 
+ bl[15] br[15] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_18 
+ bl[16] br[16] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_19 
+ bl[17] br[17] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_20 
+ bl[18] br[18] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_21 
+ bl[19] br[19] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_22 
+ bl[20] br[20] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_23 
+ bl[21] br[21] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_24 
+ bl[22] br[22] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_25 
+ bl[23] br[23] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_26 
+ bl[24] br[24] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_27 
+ bl[25] br[25] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_28 
+ bl[26] br[26] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_29 
+ bl[27] br[27] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_30 
+ bl[28] br[28] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_31 
+ bl[29] br[29] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_32 
+ bl[30] br[30] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_33 
+ bl[31] br[31] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_34 
+ bl[32] br[32] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_35 
+ bl[33] br[33] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_36 
+ bl[34] br[34] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_37 
+ bl[35] br[35] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_38 
+ bl[36] br[36] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_39 
+ bl[37] br[37] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_40 
+ bl[38] br[38] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_41 
+ bl[39] br[39] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_42 
+ bl[40] br[40] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_43 
+ bl[41] br[41] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_44 
+ bl[42] br[42] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_45 
+ bl[43] br[43] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_46 
+ bl[44] br[44] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_47 
+ bl[45] br[45] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_48 
+ bl[46] br[46] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_49 
+ bl[47] br[47] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_50 
+ bl[48] br[48] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_51 
+ bl[49] br[49] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_52 
+ bl[50] br[50] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_53 
+ bl[51] br[51] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_54 
+ bl[52] br[52] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_55 
+ bl[53] br[53] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_56 
+ bl[54] br[54] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_57 
+ bl[55] br[55] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_58 
+ bl[56] br[56] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_59 
+ bl[57] br[57] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_60 
+ bl[58] br[58] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_61 
+ bl[59] br[59] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_62 
+ bl[60] br[60] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_63 
+ bl[61] br[61] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_64 
+ bl[62] br[62] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_65 
+ bl[63] br[63] vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_66 
+ vdd vdd vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_311_67 
+ vdd vdd vdd vss wl[309] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_0 
+ vdd vdd vss vdd vpb vnb wl[310] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_312_1 
+ rbl rbr vss vdd vpb vnb wl[310] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_312_2 
+ bl[0] br[0] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_3 
+ bl[1] br[1] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_4 
+ bl[2] br[2] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_5 
+ bl[3] br[3] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_6 
+ bl[4] br[4] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_7 
+ bl[5] br[5] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_8 
+ bl[6] br[6] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_9 
+ bl[7] br[7] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_10 
+ bl[8] br[8] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_11 
+ bl[9] br[9] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_12 
+ bl[10] br[10] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_13 
+ bl[11] br[11] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_14 
+ bl[12] br[12] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_15 
+ bl[13] br[13] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_16 
+ bl[14] br[14] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_17 
+ bl[15] br[15] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_18 
+ bl[16] br[16] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_19 
+ bl[17] br[17] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_20 
+ bl[18] br[18] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_21 
+ bl[19] br[19] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_22 
+ bl[20] br[20] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_23 
+ bl[21] br[21] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_24 
+ bl[22] br[22] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_25 
+ bl[23] br[23] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_26 
+ bl[24] br[24] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_27 
+ bl[25] br[25] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_28 
+ bl[26] br[26] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_29 
+ bl[27] br[27] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_30 
+ bl[28] br[28] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_31 
+ bl[29] br[29] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_32 
+ bl[30] br[30] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_33 
+ bl[31] br[31] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_34 
+ bl[32] br[32] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_35 
+ bl[33] br[33] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_36 
+ bl[34] br[34] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_37 
+ bl[35] br[35] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_38 
+ bl[36] br[36] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_39 
+ bl[37] br[37] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_40 
+ bl[38] br[38] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_41 
+ bl[39] br[39] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_42 
+ bl[40] br[40] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_43 
+ bl[41] br[41] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_44 
+ bl[42] br[42] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_45 
+ bl[43] br[43] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_46 
+ bl[44] br[44] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_47 
+ bl[45] br[45] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_48 
+ bl[46] br[46] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_49 
+ bl[47] br[47] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_50 
+ bl[48] br[48] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_51 
+ bl[49] br[49] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_52 
+ bl[50] br[50] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_53 
+ bl[51] br[51] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_54 
+ bl[52] br[52] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_55 
+ bl[53] br[53] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_56 
+ bl[54] br[54] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_57 
+ bl[55] br[55] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_58 
+ bl[56] br[56] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_59 
+ bl[57] br[57] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_60 
+ bl[58] br[58] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_61 
+ bl[59] br[59] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_62 
+ bl[60] br[60] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_63 
+ bl[61] br[61] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_64 
+ bl[62] br[62] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_65 
+ bl[63] br[63] vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_66 
+ vdd vdd vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_312_67 
+ vdd vdd vdd vss wl[310] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_0 
+ vdd vdd vss vdd vpb vnb wl[311] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_313_1 
+ rbl rbr vss vdd vpb vnb wl[311] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_313_2 
+ bl[0] br[0] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_3 
+ bl[1] br[1] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_4 
+ bl[2] br[2] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_5 
+ bl[3] br[3] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_6 
+ bl[4] br[4] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_7 
+ bl[5] br[5] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_8 
+ bl[6] br[6] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_9 
+ bl[7] br[7] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_10 
+ bl[8] br[8] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_11 
+ bl[9] br[9] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_12 
+ bl[10] br[10] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_13 
+ bl[11] br[11] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_14 
+ bl[12] br[12] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_15 
+ bl[13] br[13] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_16 
+ bl[14] br[14] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_17 
+ bl[15] br[15] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_18 
+ bl[16] br[16] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_19 
+ bl[17] br[17] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_20 
+ bl[18] br[18] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_21 
+ bl[19] br[19] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_22 
+ bl[20] br[20] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_23 
+ bl[21] br[21] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_24 
+ bl[22] br[22] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_25 
+ bl[23] br[23] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_26 
+ bl[24] br[24] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_27 
+ bl[25] br[25] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_28 
+ bl[26] br[26] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_29 
+ bl[27] br[27] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_30 
+ bl[28] br[28] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_31 
+ bl[29] br[29] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_32 
+ bl[30] br[30] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_33 
+ bl[31] br[31] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_34 
+ bl[32] br[32] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_35 
+ bl[33] br[33] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_36 
+ bl[34] br[34] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_37 
+ bl[35] br[35] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_38 
+ bl[36] br[36] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_39 
+ bl[37] br[37] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_40 
+ bl[38] br[38] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_41 
+ bl[39] br[39] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_42 
+ bl[40] br[40] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_43 
+ bl[41] br[41] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_44 
+ bl[42] br[42] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_45 
+ bl[43] br[43] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_46 
+ bl[44] br[44] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_47 
+ bl[45] br[45] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_48 
+ bl[46] br[46] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_49 
+ bl[47] br[47] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_50 
+ bl[48] br[48] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_51 
+ bl[49] br[49] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_52 
+ bl[50] br[50] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_53 
+ bl[51] br[51] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_54 
+ bl[52] br[52] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_55 
+ bl[53] br[53] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_56 
+ bl[54] br[54] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_57 
+ bl[55] br[55] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_58 
+ bl[56] br[56] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_59 
+ bl[57] br[57] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_60 
+ bl[58] br[58] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_61 
+ bl[59] br[59] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_62 
+ bl[60] br[60] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_63 
+ bl[61] br[61] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_64 
+ bl[62] br[62] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_65 
+ bl[63] br[63] vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_66 
+ vdd vdd vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_313_67 
+ vdd vdd vdd vss wl[311] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_0 
+ vdd vdd vss vdd vpb vnb wl[312] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_314_1 
+ rbl rbr vss vdd vpb vnb wl[312] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_314_2 
+ bl[0] br[0] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_3 
+ bl[1] br[1] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_4 
+ bl[2] br[2] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_5 
+ bl[3] br[3] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_6 
+ bl[4] br[4] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_7 
+ bl[5] br[5] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_8 
+ bl[6] br[6] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_9 
+ bl[7] br[7] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_10 
+ bl[8] br[8] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_11 
+ bl[9] br[9] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_12 
+ bl[10] br[10] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_13 
+ bl[11] br[11] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_14 
+ bl[12] br[12] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_15 
+ bl[13] br[13] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_16 
+ bl[14] br[14] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_17 
+ bl[15] br[15] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_18 
+ bl[16] br[16] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_19 
+ bl[17] br[17] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_20 
+ bl[18] br[18] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_21 
+ bl[19] br[19] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_22 
+ bl[20] br[20] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_23 
+ bl[21] br[21] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_24 
+ bl[22] br[22] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_25 
+ bl[23] br[23] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_26 
+ bl[24] br[24] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_27 
+ bl[25] br[25] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_28 
+ bl[26] br[26] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_29 
+ bl[27] br[27] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_30 
+ bl[28] br[28] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_31 
+ bl[29] br[29] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_32 
+ bl[30] br[30] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_33 
+ bl[31] br[31] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_34 
+ bl[32] br[32] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_35 
+ bl[33] br[33] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_36 
+ bl[34] br[34] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_37 
+ bl[35] br[35] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_38 
+ bl[36] br[36] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_39 
+ bl[37] br[37] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_40 
+ bl[38] br[38] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_41 
+ bl[39] br[39] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_42 
+ bl[40] br[40] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_43 
+ bl[41] br[41] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_44 
+ bl[42] br[42] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_45 
+ bl[43] br[43] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_46 
+ bl[44] br[44] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_47 
+ bl[45] br[45] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_48 
+ bl[46] br[46] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_49 
+ bl[47] br[47] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_50 
+ bl[48] br[48] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_51 
+ bl[49] br[49] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_52 
+ bl[50] br[50] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_53 
+ bl[51] br[51] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_54 
+ bl[52] br[52] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_55 
+ bl[53] br[53] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_56 
+ bl[54] br[54] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_57 
+ bl[55] br[55] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_58 
+ bl[56] br[56] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_59 
+ bl[57] br[57] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_60 
+ bl[58] br[58] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_61 
+ bl[59] br[59] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_62 
+ bl[60] br[60] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_63 
+ bl[61] br[61] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_64 
+ bl[62] br[62] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_65 
+ bl[63] br[63] vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_66 
+ vdd vdd vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_314_67 
+ vdd vdd vdd vss wl[312] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_0 
+ vdd vdd vss vdd vpb vnb wl[313] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_315_1 
+ rbl rbr vss vdd vpb vnb wl[313] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_315_2 
+ bl[0] br[0] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_3 
+ bl[1] br[1] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_4 
+ bl[2] br[2] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_5 
+ bl[3] br[3] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_6 
+ bl[4] br[4] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_7 
+ bl[5] br[5] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_8 
+ bl[6] br[6] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_9 
+ bl[7] br[7] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_10 
+ bl[8] br[8] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_11 
+ bl[9] br[9] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_12 
+ bl[10] br[10] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_13 
+ bl[11] br[11] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_14 
+ bl[12] br[12] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_15 
+ bl[13] br[13] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_16 
+ bl[14] br[14] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_17 
+ bl[15] br[15] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_18 
+ bl[16] br[16] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_19 
+ bl[17] br[17] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_20 
+ bl[18] br[18] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_21 
+ bl[19] br[19] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_22 
+ bl[20] br[20] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_23 
+ bl[21] br[21] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_24 
+ bl[22] br[22] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_25 
+ bl[23] br[23] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_26 
+ bl[24] br[24] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_27 
+ bl[25] br[25] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_28 
+ bl[26] br[26] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_29 
+ bl[27] br[27] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_30 
+ bl[28] br[28] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_31 
+ bl[29] br[29] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_32 
+ bl[30] br[30] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_33 
+ bl[31] br[31] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_34 
+ bl[32] br[32] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_35 
+ bl[33] br[33] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_36 
+ bl[34] br[34] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_37 
+ bl[35] br[35] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_38 
+ bl[36] br[36] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_39 
+ bl[37] br[37] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_40 
+ bl[38] br[38] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_41 
+ bl[39] br[39] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_42 
+ bl[40] br[40] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_43 
+ bl[41] br[41] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_44 
+ bl[42] br[42] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_45 
+ bl[43] br[43] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_46 
+ bl[44] br[44] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_47 
+ bl[45] br[45] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_48 
+ bl[46] br[46] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_49 
+ bl[47] br[47] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_50 
+ bl[48] br[48] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_51 
+ bl[49] br[49] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_52 
+ bl[50] br[50] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_53 
+ bl[51] br[51] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_54 
+ bl[52] br[52] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_55 
+ bl[53] br[53] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_56 
+ bl[54] br[54] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_57 
+ bl[55] br[55] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_58 
+ bl[56] br[56] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_59 
+ bl[57] br[57] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_60 
+ bl[58] br[58] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_61 
+ bl[59] br[59] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_62 
+ bl[60] br[60] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_63 
+ bl[61] br[61] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_64 
+ bl[62] br[62] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_65 
+ bl[63] br[63] vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_66 
+ vdd vdd vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_315_67 
+ vdd vdd vdd vss wl[313] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_0 
+ vdd vdd vss vdd vpb vnb wl[314] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_316_1 
+ rbl rbr vss vdd vpb vnb wl[314] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_316_2 
+ bl[0] br[0] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_3 
+ bl[1] br[1] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_4 
+ bl[2] br[2] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_5 
+ bl[3] br[3] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_6 
+ bl[4] br[4] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_7 
+ bl[5] br[5] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_8 
+ bl[6] br[6] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_9 
+ bl[7] br[7] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_10 
+ bl[8] br[8] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_11 
+ bl[9] br[9] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_12 
+ bl[10] br[10] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_13 
+ bl[11] br[11] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_14 
+ bl[12] br[12] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_15 
+ bl[13] br[13] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_16 
+ bl[14] br[14] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_17 
+ bl[15] br[15] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_18 
+ bl[16] br[16] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_19 
+ bl[17] br[17] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_20 
+ bl[18] br[18] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_21 
+ bl[19] br[19] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_22 
+ bl[20] br[20] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_23 
+ bl[21] br[21] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_24 
+ bl[22] br[22] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_25 
+ bl[23] br[23] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_26 
+ bl[24] br[24] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_27 
+ bl[25] br[25] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_28 
+ bl[26] br[26] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_29 
+ bl[27] br[27] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_30 
+ bl[28] br[28] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_31 
+ bl[29] br[29] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_32 
+ bl[30] br[30] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_33 
+ bl[31] br[31] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_34 
+ bl[32] br[32] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_35 
+ bl[33] br[33] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_36 
+ bl[34] br[34] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_37 
+ bl[35] br[35] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_38 
+ bl[36] br[36] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_39 
+ bl[37] br[37] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_40 
+ bl[38] br[38] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_41 
+ bl[39] br[39] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_42 
+ bl[40] br[40] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_43 
+ bl[41] br[41] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_44 
+ bl[42] br[42] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_45 
+ bl[43] br[43] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_46 
+ bl[44] br[44] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_47 
+ bl[45] br[45] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_48 
+ bl[46] br[46] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_49 
+ bl[47] br[47] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_50 
+ bl[48] br[48] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_51 
+ bl[49] br[49] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_52 
+ bl[50] br[50] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_53 
+ bl[51] br[51] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_54 
+ bl[52] br[52] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_55 
+ bl[53] br[53] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_56 
+ bl[54] br[54] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_57 
+ bl[55] br[55] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_58 
+ bl[56] br[56] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_59 
+ bl[57] br[57] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_60 
+ bl[58] br[58] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_61 
+ bl[59] br[59] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_62 
+ bl[60] br[60] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_63 
+ bl[61] br[61] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_64 
+ bl[62] br[62] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_65 
+ bl[63] br[63] vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_66 
+ vdd vdd vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_316_67 
+ vdd vdd vdd vss wl[314] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_0 
+ vdd vdd vss vdd vpb vnb wl[315] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_317_1 
+ rbl rbr vss vdd vpb vnb wl[315] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_317_2 
+ bl[0] br[0] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_3 
+ bl[1] br[1] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_4 
+ bl[2] br[2] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_5 
+ bl[3] br[3] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_6 
+ bl[4] br[4] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_7 
+ bl[5] br[5] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_8 
+ bl[6] br[6] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_9 
+ bl[7] br[7] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_10 
+ bl[8] br[8] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_11 
+ bl[9] br[9] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_12 
+ bl[10] br[10] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_13 
+ bl[11] br[11] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_14 
+ bl[12] br[12] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_15 
+ bl[13] br[13] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_16 
+ bl[14] br[14] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_17 
+ bl[15] br[15] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_18 
+ bl[16] br[16] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_19 
+ bl[17] br[17] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_20 
+ bl[18] br[18] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_21 
+ bl[19] br[19] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_22 
+ bl[20] br[20] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_23 
+ bl[21] br[21] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_24 
+ bl[22] br[22] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_25 
+ bl[23] br[23] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_26 
+ bl[24] br[24] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_27 
+ bl[25] br[25] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_28 
+ bl[26] br[26] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_29 
+ bl[27] br[27] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_30 
+ bl[28] br[28] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_31 
+ bl[29] br[29] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_32 
+ bl[30] br[30] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_33 
+ bl[31] br[31] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_34 
+ bl[32] br[32] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_35 
+ bl[33] br[33] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_36 
+ bl[34] br[34] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_37 
+ bl[35] br[35] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_38 
+ bl[36] br[36] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_39 
+ bl[37] br[37] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_40 
+ bl[38] br[38] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_41 
+ bl[39] br[39] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_42 
+ bl[40] br[40] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_43 
+ bl[41] br[41] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_44 
+ bl[42] br[42] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_45 
+ bl[43] br[43] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_46 
+ bl[44] br[44] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_47 
+ bl[45] br[45] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_48 
+ bl[46] br[46] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_49 
+ bl[47] br[47] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_50 
+ bl[48] br[48] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_51 
+ bl[49] br[49] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_52 
+ bl[50] br[50] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_53 
+ bl[51] br[51] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_54 
+ bl[52] br[52] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_55 
+ bl[53] br[53] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_56 
+ bl[54] br[54] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_57 
+ bl[55] br[55] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_58 
+ bl[56] br[56] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_59 
+ bl[57] br[57] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_60 
+ bl[58] br[58] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_61 
+ bl[59] br[59] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_62 
+ bl[60] br[60] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_63 
+ bl[61] br[61] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_64 
+ bl[62] br[62] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_65 
+ bl[63] br[63] vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_66 
+ vdd vdd vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_317_67 
+ vdd vdd vdd vss wl[315] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_0 
+ vdd vdd vss vdd vpb vnb wl[316] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_318_1 
+ rbl rbr vss vdd vpb vnb wl[316] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_318_2 
+ bl[0] br[0] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_3 
+ bl[1] br[1] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_4 
+ bl[2] br[2] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_5 
+ bl[3] br[3] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_6 
+ bl[4] br[4] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_7 
+ bl[5] br[5] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_8 
+ bl[6] br[6] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_9 
+ bl[7] br[7] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_10 
+ bl[8] br[8] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_11 
+ bl[9] br[9] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_12 
+ bl[10] br[10] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_13 
+ bl[11] br[11] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_14 
+ bl[12] br[12] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_15 
+ bl[13] br[13] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_16 
+ bl[14] br[14] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_17 
+ bl[15] br[15] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_18 
+ bl[16] br[16] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_19 
+ bl[17] br[17] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_20 
+ bl[18] br[18] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_21 
+ bl[19] br[19] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_22 
+ bl[20] br[20] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_23 
+ bl[21] br[21] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_24 
+ bl[22] br[22] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_25 
+ bl[23] br[23] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_26 
+ bl[24] br[24] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_27 
+ bl[25] br[25] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_28 
+ bl[26] br[26] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_29 
+ bl[27] br[27] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_30 
+ bl[28] br[28] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_31 
+ bl[29] br[29] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_32 
+ bl[30] br[30] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_33 
+ bl[31] br[31] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_34 
+ bl[32] br[32] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_35 
+ bl[33] br[33] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_36 
+ bl[34] br[34] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_37 
+ bl[35] br[35] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_38 
+ bl[36] br[36] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_39 
+ bl[37] br[37] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_40 
+ bl[38] br[38] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_41 
+ bl[39] br[39] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_42 
+ bl[40] br[40] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_43 
+ bl[41] br[41] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_44 
+ bl[42] br[42] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_45 
+ bl[43] br[43] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_46 
+ bl[44] br[44] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_47 
+ bl[45] br[45] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_48 
+ bl[46] br[46] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_49 
+ bl[47] br[47] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_50 
+ bl[48] br[48] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_51 
+ bl[49] br[49] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_52 
+ bl[50] br[50] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_53 
+ bl[51] br[51] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_54 
+ bl[52] br[52] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_55 
+ bl[53] br[53] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_56 
+ bl[54] br[54] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_57 
+ bl[55] br[55] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_58 
+ bl[56] br[56] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_59 
+ bl[57] br[57] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_60 
+ bl[58] br[58] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_61 
+ bl[59] br[59] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_62 
+ bl[60] br[60] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_63 
+ bl[61] br[61] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_64 
+ bl[62] br[62] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_65 
+ bl[63] br[63] vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_66 
+ vdd vdd vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_318_67 
+ vdd vdd vdd vss wl[316] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_0 
+ vdd vdd vss vdd vpb vnb wl[317] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_319_1 
+ rbl rbr vss vdd vpb vnb wl[317] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_319_2 
+ bl[0] br[0] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_3 
+ bl[1] br[1] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_4 
+ bl[2] br[2] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_5 
+ bl[3] br[3] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_6 
+ bl[4] br[4] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_7 
+ bl[5] br[5] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_8 
+ bl[6] br[6] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_9 
+ bl[7] br[7] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_10 
+ bl[8] br[8] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_11 
+ bl[9] br[9] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_12 
+ bl[10] br[10] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_13 
+ bl[11] br[11] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_14 
+ bl[12] br[12] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_15 
+ bl[13] br[13] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_16 
+ bl[14] br[14] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_17 
+ bl[15] br[15] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_18 
+ bl[16] br[16] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_19 
+ bl[17] br[17] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_20 
+ bl[18] br[18] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_21 
+ bl[19] br[19] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_22 
+ bl[20] br[20] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_23 
+ bl[21] br[21] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_24 
+ bl[22] br[22] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_25 
+ bl[23] br[23] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_26 
+ bl[24] br[24] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_27 
+ bl[25] br[25] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_28 
+ bl[26] br[26] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_29 
+ bl[27] br[27] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_30 
+ bl[28] br[28] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_31 
+ bl[29] br[29] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_32 
+ bl[30] br[30] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_33 
+ bl[31] br[31] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_34 
+ bl[32] br[32] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_35 
+ bl[33] br[33] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_36 
+ bl[34] br[34] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_37 
+ bl[35] br[35] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_38 
+ bl[36] br[36] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_39 
+ bl[37] br[37] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_40 
+ bl[38] br[38] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_41 
+ bl[39] br[39] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_42 
+ bl[40] br[40] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_43 
+ bl[41] br[41] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_44 
+ bl[42] br[42] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_45 
+ bl[43] br[43] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_46 
+ bl[44] br[44] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_47 
+ bl[45] br[45] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_48 
+ bl[46] br[46] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_49 
+ bl[47] br[47] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_50 
+ bl[48] br[48] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_51 
+ bl[49] br[49] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_52 
+ bl[50] br[50] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_53 
+ bl[51] br[51] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_54 
+ bl[52] br[52] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_55 
+ bl[53] br[53] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_56 
+ bl[54] br[54] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_57 
+ bl[55] br[55] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_58 
+ bl[56] br[56] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_59 
+ bl[57] br[57] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_60 
+ bl[58] br[58] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_61 
+ bl[59] br[59] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_62 
+ bl[60] br[60] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_63 
+ bl[61] br[61] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_64 
+ bl[62] br[62] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_65 
+ bl[63] br[63] vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_66 
+ vdd vdd vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_319_67 
+ vdd vdd vdd vss wl[317] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_0 
+ vdd vdd vss vdd vpb vnb wl[318] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_320_1 
+ rbl rbr vss vdd vpb vnb wl[318] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_320_2 
+ bl[0] br[0] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_3 
+ bl[1] br[1] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_4 
+ bl[2] br[2] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_5 
+ bl[3] br[3] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_6 
+ bl[4] br[4] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_7 
+ bl[5] br[5] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_8 
+ bl[6] br[6] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_9 
+ bl[7] br[7] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_10 
+ bl[8] br[8] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_11 
+ bl[9] br[9] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_12 
+ bl[10] br[10] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_13 
+ bl[11] br[11] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_14 
+ bl[12] br[12] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_15 
+ bl[13] br[13] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_16 
+ bl[14] br[14] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_17 
+ bl[15] br[15] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_18 
+ bl[16] br[16] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_19 
+ bl[17] br[17] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_20 
+ bl[18] br[18] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_21 
+ bl[19] br[19] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_22 
+ bl[20] br[20] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_23 
+ bl[21] br[21] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_24 
+ bl[22] br[22] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_25 
+ bl[23] br[23] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_26 
+ bl[24] br[24] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_27 
+ bl[25] br[25] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_28 
+ bl[26] br[26] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_29 
+ bl[27] br[27] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_30 
+ bl[28] br[28] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_31 
+ bl[29] br[29] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_32 
+ bl[30] br[30] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_33 
+ bl[31] br[31] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_34 
+ bl[32] br[32] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_35 
+ bl[33] br[33] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_36 
+ bl[34] br[34] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_37 
+ bl[35] br[35] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_38 
+ bl[36] br[36] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_39 
+ bl[37] br[37] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_40 
+ bl[38] br[38] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_41 
+ bl[39] br[39] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_42 
+ bl[40] br[40] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_43 
+ bl[41] br[41] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_44 
+ bl[42] br[42] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_45 
+ bl[43] br[43] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_46 
+ bl[44] br[44] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_47 
+ bl[45] br[45] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_48 
+ bl[46] br[46] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_49 
+ bl[47] br[47] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_50 
+ bl[48] br[48] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_51 
+ bl[49] br[49] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_52 
+ bl[50] br[50] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_53 
+ bl[51] br[51] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_54 
+ bl[52] br[52] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_55 
+ bl[53] br[53] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_56 
+ bl[54] br[54] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_57 
+ bl[55] br[55] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_58 
+ bl[56] br[56] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_59 
+ bl[57] br[57] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_60 
+ bl[58] br[58] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_61 
+ bl[59] br[59] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_62 
+ bl[60] br[60] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_63 
+ bl[61] br[61] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_64 
+ bl[62] br[62] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_65 
+ bl[63] br[63] vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_66 
+ vdd vdd vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_320_67 
+ vdd vdd vdd vss wl[318] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_0 
+ vdd vdd vss vdd vpb vnb wl[319] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_321_1 
+ rbl rbr vss vdd vpb vnb wl[319] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_321_2 
+ bl[0] br[0] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_3 
+ bl[1] br[1] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_4 
+ bl[2] br[2] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_5 
+ bl[3] br[3] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_6 
+ bl[4] br[4] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_7 
+ bl[5] br[5] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_8 
+ bl[6] br[6] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_9 
+ bl[7] br[7] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_10 
+ bl[8] br[8] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_11 
+ bl[9] br[9] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_12 
+ bl[10] br[10] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_13 
+ bl[11] br[11] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_14 
+ bl[12] br[12] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_15 
+ bl[13] br[13] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_16 
+ bl[14] br[14] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_17 
+ bl[15] br[15] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_18 
+ bl[16] br[16] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_19 
+ bl[17] br[17] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_20 
+ bl[18] br[18] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_21 
+ bl[19] br[19] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_22 
+ bl[20] br[20] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_23 
+ bl[21] br[21] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_24 
+ bl[22] br[22] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_25 
+ bl[23] br[23] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_26 
+ bl[24] br[24] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_27 
+ bl[25] br[25] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_28 
+ bl[26] br[26] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_29 
+ bl[27] br[27] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_30 
+ bl[28] br[28] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_31 
+ bl[29] br[29] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_32 
+ bl[30] br[30] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_33 
+ bl[31] br[31] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_34 
+ bl[32] br[32] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_35 
+ bl[33] br[33] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_36 
+ bl[34] br[34] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_37 
+ bl[35] br[35] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_38 
+ bl[36] br[36] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_39 
+ bl[37] br[37] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_40 
+ bl[38] br[38] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_41 
+ bl[39] br[39] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_42 
+ bl[40] br[40] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_43 
+ bl[41] br[41] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_44 
+ bl[42] br[42] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_45 
+ bl[43] br[43] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_46 
+ bl[44] br[44] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_47 
+ bl[45] br[45] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_48 
+ bl[46] br[46] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_49 
+ bl[47] br[47] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_50 
+ bl[48] br[48] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_51 
+ bl[49] br[49] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_52 
+ bl[50] br[50] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_53 
+ bl[51] br[51] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_54 
+ bl[52] br[52] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_55 
+ bl[53] br[53] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_56 
+ bl[54] br[54] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_57 
+ bl[55] br[55] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_58 
+ bl[56] br[56] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_59 
+ bl[57] br[57] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_60 
+ bl[58] br[58] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_61 
+ bl[59] br[59] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_62 
+ bl[60] br[60] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_63 
+ bl[61] br[61] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_64 
+ bl[62] br[62] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_65 
+ bl[63] br[63] vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_66 
+ vdd vdd vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_321_67 
+ vdd vdd vdd vss wl[319] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_0 
+ vdd vdd vss vdd vpb vnb wl[320] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_322_1 
+ rbl rbr vss vdd vpb vnb wl[320] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_322_2 
+ bl[0] br[0] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_3 
+ bl[1] br[1] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_4 
+ bl[2] br[2] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_5 
+ bl[3] br[3] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_6 
+ bl[4] br[4] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_7 
+ bl[5] br[5] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_8 
+ bl[6] br[6] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_9 
+ bl[7] br[7] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_10 
+ bl[8] br[8] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_11 
+ bl[9] br[9] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_12 
+ bl[10] br[10] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_13 
+ bl[11] br[11] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_14 
+ bl[12] br[12] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_15 
+ bl[13] br[13] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_16 
+ bl[14] br[14] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_17 
+ bl[15] br[15] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_18 
+ bl[16] br[16] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_19 
+ bl[17] br[17] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_20 
+ bl[18] br[18] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_21 
+ bl[19] br[19] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_22 
+ bl[20] br[20] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_23 
+ bl[21] br[21] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_24 
+ bl[22] br[22] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_25 
+ bl[23] br[23] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_26 
+ bl[24] br[24] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_27 
+ bl[25] br[25] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_28 
+ bl[26] br[26] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_29 
+ bl[27] br[27] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_30 
+ bl[28] br[28] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_31 
+ bl[29] br[29] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_32 
+ bl[30] br[30] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_33 
+ bl[31] br[31] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_34 
+ bl[32] br[32] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_35 
+ bl[33] br[33] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_36 
+ bl[34] br[34] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_37 
+ bl[35] br[35] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_38 
+ bl[36] br[36] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_39 
+ bl[37] br[37] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_40 
+ bl[38] br[38] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_41 
+ bl[39] br[39] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_42 
+ bl[40] br[40] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_43 
+ bl[41] br[41] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_44 
+ bl[42] br[42] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_45 
+ bl[43] br[43] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_46 
+ bl[44] br[44] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_47 
+ bl[45] br[45] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_48 
+ bl[46] br[46] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_49 
+ bl[47] br[47] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_50 
+ bl[48] br[48] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_51 
+ bl[49] br[49] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_52 
+ bl[50] br[50] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_53 
+ bl[51] br[51] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_54 
+ bl[52] br[52] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_55 
+ bl[53] br[53] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_56 
+ bl[54] br[54] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_57 
+ bl[55] br[55] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_58 
+ bl[56] br[56] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_59 
+ bl[57] br[57] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_60 
+ bl[58] br[58] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_61 
+ bl[59] br[59] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_62 
+ bl[60] br[60] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_63 
+ bl[61] br[61] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_64 
+ bl[62] br[62] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_65 
+ bl[63] br[63] vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_66 
+ vdd vdd vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_322_67 
+ vdd vdd vdd vss wl[320] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_0 
+ vdd vdd vss vdd vpb vnb wl[321] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_323_1 
+ rbl rbr vss vdd vpb vnb wl[321] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_323_2 
+ bl[0] br[0] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_3 
+ bl[1] br[1] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_4 
+ bl[2] br[2] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_5 
+ bl[3] br[3] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_6 
+ bl[4] br[4] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_7 
+ bl[5] br[5] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_8 
+ bl[6] br[6] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_9 
+ bl[7] br[7] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_10 
+ bl[8] br[8] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_11 
+ bl[9] br[9] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_12 
+ bl[10] br[10] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_13 
+ bl[11] br[11] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_14 
+ bl[12] br[12] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_15 
+ bl[13] br[13] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_16 
+ bl[14] br[14] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_17 
+ bl[15] br[15] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_18 
+ bl[16] br[16] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_19 
+ bl[17] br[17] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_20 
+ bl[18] br[18] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_21 
+ bl[19] br[19] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_22 
+ bl[20] br[20] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_23 
+ bl[21] br[21] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_24 
+ bl[22] br[22] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_25 
+ bl[23] br[23] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_26 
+ bl[24] br[24] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_27 
+ bl[25] br[25] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_28 
+ bl[26] br[26] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_29 
+ bl[27] br[27] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_30 
+ bl[28] br[28] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_31 
+ bl[29] br[29] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_32 
+ bl[30] br[30] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_33 
+ bl[31] br[31] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_34 
+ bl[32] br[32] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_35 
+ bl[33] br[33] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_36 
+ bl[34] br[34] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_37 
+ bl[35] br[35] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_38 
+ bl[36] br[36] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_39 
+ bl[37] br[37] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_40 
+ bl[38] br[38] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_41 
+ bl[39] br[39] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_42 
+ bl[40] br[40] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_43 
+ bl[41] br[41] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_44 
+ bl[42] br[42] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_45 
+ bl[43] br[43] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_46 
+ bl[44] br[44] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_47 
+ bl[45] br[45] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_48 
+ bl[46] br[46] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_49 
+ bl[47] br[47] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_50 
+ bl[48] br[48] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_51 
+ bl[49] br[49] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_52 
+ bl[50] br[50] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_53 
+ bl[51] br[51] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_54 
+ bl[52] br[52] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_55 
+ bl[53] br[53] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_56 
+ bl[54] br[54] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_57 
+ bl[55] br[55] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_58 
+ bl[56] br[56] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_59 
+ bl[57] br[57] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_60 
+ bl[58] br[58] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_61 
+ bl[59] br[59] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_62 
+ bl[60] br[60] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_63 
+ bl[61] br[61] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_64 
+ bl[62] br[62] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_65 
+ bl[63] br[63] vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_66 
+ vdd vdd vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_323_67 
+ vdd vdd vdd vss wl[321] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_0 
+ vdd vdd vss vdd vpb vnb wl[322] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_324_1 
+ rbl rbr vss vdd vpb vnb wl[322] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_324_2 
+ bl[0] br[0] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_3 
+ bl[1] br[1] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_4 
+ bl[2] br[2] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_5 
+ bl[3] br[3] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_6 
+ bl[4] br[4] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_7 
+ bl[5] br[5] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_8 
+ bl[6] br[6] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_9 
+ bl[7] br[7] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_10 
+ bl[8] br[8] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_11 
+ bl[9] br[9] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_12 
+ bl[10] br[10] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_13 
+ bl[11] br[11] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_14 
+ bl[12] br[12] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_15 
+ bl[13] br[13] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_16 
+ bl[14] br[14] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_17 
+ bl[15] br[15] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_18 
+ bl[16] br[16] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_19 
+ bl[17] br[17] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_20 
+ bl[18] br[18] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_21 
+ bl[19] br[19] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_22 
+ bl[20] br[20] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_23 
+ bl[21] br[21] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_24 
+ bl[22] br[22] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_25 
+ bl[23] br[23] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_26 
+ bl[24] br[24] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_27 
+ bl[25] br[25] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_28 
+ bl[26] br[26] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_29 
+ bl[27] br[27] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_30 
+ bl[28] br[28] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_31 
+ bl[29] br[29] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_32 
+ bl[30] br[30] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_33 
+ bl[31] br[31] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_34 
+ bl[32] br[32] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_35 
+ bl[33] br[33] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_36 
+ bl[34] br[34] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_37 
+ bl[35] br[35] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_38 
+ bl[36] br[36] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_39 
+ bl[37] br[37] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_40 
+ bl[38] br[38] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_41 
+ bl[39] br[39] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_42 
+ bl[40] br[40] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_43 
+ bl[41] br[41] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_44 
+ bl[42] br[42] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_45 
+ bl[43] br[43] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_46 
+ bl[44] br[44] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_47 
+ bl[45] br[45] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_48 
+ bl[46] br[46] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_49 
+ bl[47] br[47] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_50 
+ bl[48] br[48] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_51 
+ bl[49] br[49] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_52 
+ bl[50] br[50] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_53 
+ bl[51] br[51] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_54 
+ bl[52] br[52] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_55 
+ bl[53] br[53] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_56 
+ bl[54] br[54] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_57 
+ bl[55] br[55] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_58 
+ bl[56] br[56] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_59 
+ bl[57] br[57] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_60 
+ bl[58] br[58] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_61 
+ bl[59] br[59] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_62 
+ bl[60] br[60] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_63 
+ bl[61] br[61] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_64 
+ bl[62] br[62] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_65 
+ bl[63] br[63] vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_66 
+ vdd vdd vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_324_67 
+ vdd vdd vdd vss wl[322] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_0 
+ vdd vdd vss vdd vpb vnb wl[323] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_325_1 
+ rbl rbr vss vdd vpb vnb wl[323] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_325_2 
+ bl[0] br[0] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_3 
+ bl[1] br[1] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_4 
+ bl[2] br[2] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_5 
+ bl[3] br[3] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_6 
+ bl[4] br[4] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_7 
+ bl[5] br[5] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_8 
+ bl[6] br[6] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_9 
+ bl[7] br[7] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_10 
+ bl[8] br[8] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_11 
+ bl[9] br[9] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_12 
+ bl[10] br[10] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_13 
+ bl[11] br[11] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_14 
+ bl[12] br[12] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_15 
+ bl[13] br[13] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_16 
+ bl[14] br[14] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_17 
+ bl[15] br[15] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_18 
+ bl[16] br[16] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_19 
+ bl[17] br[17] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_20 
+ bl[18] br[18] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_21 
+ bl[19] br[19] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_22 
+ bl[20] br[20] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_23 
+ bl[21] br[21] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_24 
+ bl[22] br[22] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_25 
+ bl[23] br[23] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_26 
+ bl[24] br[24] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_27 
+ bl[25] br[25] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_28 
+ bl[26] br[26] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_29 
+ bl[27] br[27] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_30 
+ bl[28] br[28] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_31 
+ bl[29] br[29] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_32 
+ bl[30] br[30] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_33 
+ bl[31] br[31] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_34 
+ bl[32] br[32] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_35 
+ bl[33] br[33] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_36 
+ bl[34] br[34] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_37 
+ bl[35] br[35] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_38 
+ bl[36] br[36] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_39 
+ bl[37] br[37] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_40 
+ bl[38] br[38] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_41 
+ bl[39] br[39] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_42 
+ bl[40] br[40] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_43 
+ bl[41] br[41] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_44 
+ bl[42] br[42] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_45 
+ bl[43] br[43] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_46 
+ bl[44] br[44] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_47 
+ bl[45] br[45] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_48 
+ bl[46] br[46] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_49 
+ bl[47] br[47] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_50 
+ bl[48] br[48] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_51 
+ bl[49] br[49] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_52 
+ bl[50] br[50] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_53 
+ bl[51] br[51] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_54 
+ bl[52] br[52] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_55 
+ bl[53] br[53] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_56 
+ bl[54] br[54] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_57 
+ bl[55] br[55] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_58 
+ bl[56] br[56] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_59 
+ bl[57] br[57] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_60 
+ bl[58] br[58] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_61 
+ bl[59] br[59] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_62 
+ bl[60] br[60] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_63 
+ bl[61] br[61] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_64 
+ bl[62] br[62] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_65 
+ bl[63] br[63] vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_66 
+ vdd vdd vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_325_67 
+ vdd vdd vdd vss wl[323] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_0 
+ vdd vdd vss vdd vpb vnb wl[324] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_326_1 
+ rbl rbr vss vdd vpb vnb wl[324] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_326_2 
+ bl[0] br[0] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_3 
+ bl[1] br[1] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_4 
+ bl[2] br[2] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_5 
+ bl[3] br[3] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_6 
+ bl[4] br[4] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_7 
+ bl[5] br[5] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_8 
+ bl[6] br[6] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_9 
+ bl[7] br[7] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_10 
+ bl[8] br[8] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_11 
+ bl[9] br[9] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_12 
+ bl[10] br[10] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_13 
+ bl[11] br[11] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_14 
+ bl[12] br[12] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_15 
+ bl[13] br[13] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_16 
+ bl[14] br[14] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_17 
+ bl[15] br[15] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_18 
+ bl[16] br[16] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_19 
+ bl[17] br[17] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_20 
+ bl[18] br[18] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_21 
+ bl[19] br[19] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_22 
+ bl[20] br[20] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_23 
+ bl[21] br[21] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_24 
+ bl[22] br[22] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_25 
+ bl[23] br[23] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_26 
+ bl[24] br[24] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_27 
+ bl[25] br[25] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_28 
+ bl[26] br[26] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_29 
+ bl[27] br[27] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_30 
+ bl[28] br[28] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_31 
+ bl[29] br[29] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_32 
+ bl[30] br[30] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_33 
+ bl[31] br[31] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_34 
+ bl[32] br[32] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_35 
+ bl[33] br[33] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_36 
+ bl[34] br[34] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_37 
+ bl[35] br[35] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_38 
+ bl[36] br[36] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_39 
+ bl[37] br[37] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_40 
+ bl[38] br[38] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_41 
+ bl[39] br[39] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_42 
+ bl[40] br[40] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_43 
+ bl[41] br[41] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_44 
+ bl[42] br[42] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_45 
+ bl[43] br[43] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_46 
+ bl[44] br[44] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_47 
+ bl[45] br[45] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_48 
+ bl[46] br[46] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_49 
+ bl[47] br[47] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_50 
+ bl[48] br[48] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_51 
+ bl[49] br[49] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_52 
+ bl[50] br[50] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_53 
+ bl[51] br[51] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_54 
+ bl[52] br[52] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_55 
+ bl[53] br[53] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_56 
+ bl[54] br[54] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_57 
+ bl[55] br[55] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_58 
+ bl[56] br[56] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_59 
+ bl[57] br[57] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_60 
+ bl[58] br[58] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_61 
+ bl[59] br[59] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_62 
+ bl[60] br[60] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_63 
+ bl[61] br[61] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_64 
+ bl[62] br[62] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_65 
+ bl[63] br[63] vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_66 
+ vdd vdd vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_326_67 
+ vdd vdd vdd vss wl[324] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_0 
+ vdd vdd vss vdd vpb vnb wl[325] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_327_1 
+ rbl rbr vss vdd vpb vnb wl[325] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_327_2 
+ bl[0] br[0] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_3 
+ bl[1] br[1] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_4 
+ bl[2] br[2] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_5 
+ bl[3] br[3] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_6 
+ bl[4] br[4] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_7 
+ bl[5] br[5] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_8 
+ bl[6] br[6] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_9 
+ bl[7] br[7] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_10 
+ bl[8] br[8] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_11 
+ bl[9] br[9] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_12 
+ bl[10] br[10] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_13 
+ bl[11] br[11] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_14 
+ bl[12] br[12] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_15 
+ bl[13] br[13] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_16 
+ bl[14] br[14] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_17 
+ bl[15] br[15] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_18 
+ bl[16] br[16] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_19 
+ bl[17] br[17] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_20 
+ bl[18] br[18] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_21 
+ bl[19] br[19] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_22 
+ bl[20] br[20] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_23 
+ bl[21] br[21] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_24 
+ bl[22] br[22] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_25 
+ bl[23] br[23] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_26 
+ bl[24] br[24] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_27 
+ bl[25] br[25] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_28 
+ bl[26] br[26] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_29 
+ bl[27] br[27] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_30 
+ bl[28] br[28] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_31 
+ bl[29] br[29] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_32 
+ bl[30] br[30] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_33 
+ bl[31] br[31] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_34 
+ bl[32] br[32] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_35 
+ bl[33] br[33] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_36 
+ bl[34] br[34] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_37 
+ bl[35] br[35] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_38 
+ bl[36] br[36] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_39 
+ bl[37] br[37] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_40 
+ bl[38] br[38] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_41 
+ bl[39] br[39] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_42 
+ bl[40] br[40] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_43 
+ bl[41] br[41] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_44 
+ bl[42] br[42] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_45 
+ bl[43] br[43] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_46 
+ bl[44] br[44] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_47 
+ bl[45] br[45] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_48 
+ bl[46] br[46] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_49 
+ bl[47] br[47] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_50 
+ bl[48] br[48] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_51 
+ bl[49] br[49] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_52 
+ bl[50] br[50] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_53 
+ bl[51] br[51] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_54 
+ bl[52] br[52] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_55 
+ bl[53] br[53] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_56 
+ bl[54] br[54] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_57 
+ bl[55] br[55] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_58 
+ bl[56] br[56] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_59 
+ bl[57] br[57] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_60 
+ bl[58] br[58] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_61 
+ bl[59] br[59] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_62 
+ bl[60] br[60] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_63 
+ bl[61] br[61] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_64 
+ bl[62] br[62] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_65 
+ bl[63] br[63] vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_66 
+ vdd vdd vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_327_67 
+ vdd vdd vdd vss wl[325] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_0 
+ vdd vdd vss vdd vpb vnb wl[326] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_328_1 
+ rbl rbr vss vdd vpb vnb wl[326] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_328_2 
+ bl[0] br[0] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_3 
+ bl[1] br[1] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_4 
+ bl[2] br[2] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_5 
+ bl[3] br[3] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_6 
+ bl[4] br[4] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_7 
+ bl[5] br[5] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_8 
+ bl[6] br[6] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_9 
+ bl[7] br[7] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_10 
+ bl[8] br[8] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_11 
+ bl[9] br[9] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_12 
+ bl[10] br[10] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_13 
+ bl[11] br[11] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_14 
+ bl[12] br[12] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_15 
+ bl[13] br[13] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_16 
+ bl[14] br[14] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_17 
+ bl[15] br[15] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_18 
+ bl[16] br[16] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_19 
+ bl[17] br[17] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_20 
+ bl[18] br[18] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_21 
+ bl[19] br[19] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_22 
+ bl[20] br[20] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_23 
+ bl[21] br[21] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_24 
+ bl[22] br[22] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_25 
+ bl[23] br[23] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_26 
+ bl[24] br[24] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_27 
+ bl[25] br[25] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_28 
+ bl[26] br[26] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_29 
+ bl[27] br[27] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_30 
+ bl[28] br[28] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_31 
+ bl[29] br[29] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_32 
+ bl[30] br[30] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_33 
+ bl[31] br[31] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_34 
+ bl[32] br[32] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_35 
+ bl[33] br[33] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_36 
+ bl[34] br[34] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_37 
+ bl[35] br[35] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_38 
+ bl[36] br[36] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_39 
+ bl[37] br[37] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_40 
+ bl[38] br[38] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_41 
+ bl[39] br[39] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_42 
+ bl[40] br[40] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_43 
+ bl[41] br[41] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_44 
+ bl[42] br[42] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_45 
+ bl[43] br[43] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_46 
+ bl[44] br[44] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_47 
+ bl[45] br[45] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_48 
+ bl[46] br[46] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_49 
+ bl[47] br[47] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_50 
+ bl[48] br[48] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_51 
+ bl[49] br[49] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_52 
+ bl[50] br[50] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_53 
+ bl[51] br[51] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_54 
+ bl[52] br[52] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_55 
+ bl[53] br[53] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_56 
+ bl[54] br[54] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_57 
+ bl[55] br[55] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_58 
+ bl[56] br[56] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_59 
+ bl[57] br[57] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_60 
+ bl[58] br[58] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_61 
+ bl[59] br[59] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_62 
+ bl[60] br[60] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_63 
+ bl[61] br[61] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_64 
+ bl[62] br[62] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_65 
+ bl[63] br[63] vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_66 
+ vdd vdd vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_328_67 
+ vdd vdd vdd vss wl[326] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_0 
+ vdd vdd vss vdd vpb vnb wl[327] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_329_1 
+ rbl rbr vss vdd vpb vnb wl[327] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_329_2 
+ bl[0] br[0] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_3 
+ bl[1] br[1] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_4 
+ bl[2] br[2] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_5 
+ bl[3] br[3] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_6 
+ bl[4] br[4] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_7 
+ bl[5] br[5] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_8 
+ bl[6] br[6] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_9 
+ bl[7] br[7] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_10 
+ bl[8] br[8] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_11 
+ bl[9] br[9] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_12 
+ bl[10] br[10] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_13 
+ bl[11] br[11] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_14 
+ bl[12] br[12] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_15 
+ bl[13] br[13] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_16 
+ bl[14] br[14] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_17 
+ bl[15] br[15] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_18 
+ bl[16] br[16] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_19 
+ bl[17] br[17] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_20 
+ bl[18] br[18] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_21 
+ bl[19] br[19] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_22 
+ bl[20] br[20] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_23 
+ bl[21] br[21] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_24 
+ bl[22] br[22] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_25 
+ bl[23] br[23] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_26 
+ bl[24] br[24] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_27 
+ bl[25] br[25] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_28 
+ bl[26] br[26] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_29 
+ bl[27] br[27] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_30 
+ bl[28] br[28] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_31 
+ bl[29] br[29] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_32 
+ bl[30] br[30] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_33 
+ bl[31] br[31] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_34 
+ bl[32] br[32] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_35 
+ bl[33] br[33] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_36 
+ bl[34] br[34] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_37 
+ bl[35] br[35] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_38 
+ bl[36] br[36] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_39 
+ bl[37] br[37] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_40 
+ bl[38] br[38] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_41 
+ bl[39] br[39] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_42 
+ bl[40] br[40] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_43 
+ bl[41] br[41] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_44 
+ bl[42] br[42] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_45 
+ bl[43] br[43] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_46 
+ bl[44] br[44] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_47 
+ bl[45] br[45] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_48 
+ bl[46] br[46] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_49 
+ bl[47] br[47] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_50 
+ bl[48] br[48] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_51 
+ bl[49] br[49] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_52 
+ bl[50] br[50] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_53 
+ bl[51] br[51] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_54 
+ bl[52] br[52] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_55 
+ bl[53] br[53] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_56 
+ bl[54] br[54] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_57 
+ bl[55] br[55] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_58 
+ bl[56] br[56] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_59 
+ bl[57] br[57] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_60 
+ bl[58] br[58] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_61 
+ bl[59] br[59] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_62 
+ bl[60] br[60] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_63 
+ bl[61] br[61] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_64 
+ bl[62] br[62] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_65 
+ bl[63] br[63] vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_66 
+ vdd vdd vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_329_67 
+ vdd vdd vdd vss wl[327] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_0 
+ vdd vdd vss vdd vpb vnb wl[328] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_330_1 
+ rbl rbr vss vdd vpb vnb wl[328] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_330_2 
+ bl[0] br[0] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_3 
+ bl[1] br[1] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_4 
+ bl[2] br[2] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_5 
+ bl[3] br[3] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_6 
+ bl[4] br[4] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_7 
+ bl[5] br[5] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_8 
+ bl[6] br[6] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_9 
+ bl[7] br[7] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_10 
+ bl[8] br[8] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_11 
+ bl[9] br[9] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_12 
+ bl[10] br[10] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_13 
+ bl[11] br[11] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_14 
+ bl[12] br[12] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_15 
+ bl[13] br[13] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_16 
+ bl[14] br[14] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_17 
+ bl[15] br[15] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_18 
+ bl[16] br[16] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_19 
+ bl[17] br[17] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_20 
+ bl[18] br[18] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_21 
+ bl[19] br[19] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_22 
+ bl[20] br[20] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_23 
+ bl[21] br[21] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_24 
+ bl[22] br[22] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_25 
+ bl[23] br[23] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_26 
+ bl[24] br[24] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_27 
+ bl[25] br[25] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_28 
+ bl[26] br[26] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_29 
+ bl[27] br[27] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_30 
+ bl[28] br[28] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_31 
+ bl[29] br[29] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_32 
+ bl[30] br[30] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_33 
+ bl[31] br[31] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_34 
+ bl[32] br[32] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_35 
+ bl[33] br[33] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_36 
+ bl[34] br[34] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_37 
+ bl[35] br[35] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_38 
+ bl[36] br[36] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_39 
+ bl[37] br[37] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_40 
+ bl[38] br[38] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_41 
+ bl[39] br[39] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_42 
+ bl[40] br[40] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_43 
+ bl[41] br[41] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_44 
+ bl[42] br[42] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_45 
+ bl[43] br[43] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_46 
+ bl[44] br[44] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_47 
+ bl[45] br[45] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_48 
+ bl[46] br[46] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_49 
+ bl[47] br[47] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_50 
+ bl[48] br[48] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_51 
+ bl[49] br[49] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_52 
+ bl[50] br[50] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_53 
+ bl[51] br[51] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_54 
+ bl[52] br[52] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_55 
+ bl[53] br[53] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_56 
+ bl[54] br[54] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_57 
+ bl[55] br[55] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_58 
+ bl[56] br[56] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_59 
+ bl[57] br[57] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_60 
+ bl[58] br[58] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_61 
+ bl[59] br[59] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_62 
+ bl[60] br[60] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_63 
+ bl[61] br[61] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_64 
+ bl[62] br[62] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_65 
+ bl[63] br[63] vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_66 
+ vdd vdd vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_330_67 
+ vdd vdd vdd vss wl[328] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_0 
+ vdd vdd vss vdd vpb vnb wl[329] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_331_1 
+ rbl rbr vss vdd vpb vnb wl[329] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_331_2 
+ bl[0] br[0] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_3 
+ bl[1] br[1] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_4 
+ bl[2] br[2] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_5 
+ bl[3] br[3] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_6 
+ bl[4] br[4] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_7 
+ bl[5] br[5] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_8 
+ bl[6] br[6] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_9 
+ bl[7] br[7] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_10 
+ bl[8] br[8] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_11 
+ bl[9] br[9] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_12 
+ bl[10] br[10] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_13 
+ bl[11] br[11] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_14 
+ bl[12] br[12] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_15 
+ bl[13] br[13] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_16 
+ bl[14] br[14] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_17 
+ bl[15] br[15] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_18 
+ bl[16] br[16] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_19 
+ bl[17] br[17] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_20 
+ bl[18] br[18] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_21 
+ bl[19] br[19] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_22 
+ bl[20] br[20] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_23 
+ bl[21] br[21] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_24 
+ bl[22] br[22] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_25 
+ bl[23] br[23] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_26 
+ bl[24] br[24] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_27 
+ bl[25] br[25] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_28 
+ bl[26] br[26] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_29 
+ bl[27] br[27] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_30 
+ bl[28] br[28] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_31 
+ bl[29] br[29] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_32 
+ bl[30] br[30] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_33 
+ bl[31] br[31] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_34 
+ bl[32] br[32] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_35 
+ bl[33] br[33] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_36 
+ bl[34] br[34] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_37 
+ bl[35] br[35] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_38 
+ bl[36] br[36] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_39 
+ bl[37] br[37] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_40 
+ bl[38] br[38] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_41 
+ bl[39] br[39] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_42 
+ bl[40] br[40] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_43 
+ bl[41] br[41] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_44 
+ bl[42] br[42] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_45 
+ bl[43] br[43] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_46 
+ bl[44] br[44] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_47 
+ bl[45] br[45] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_48 
+ bl[46] br[46] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_49 
+ bl[47] br[47] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_50 
+ bl[48] br[48] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_51 
+ bl[49] br[49] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_52 
+ bl[50] br[50] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_53 
+ bl[51] br[51] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_54 
+ bl[52] br[52] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_55 
+ bl[53] br[53] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_56 
+ bl[54] br[54] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_57 
+ bl[55] br[55] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_58 
+ bl[56] br[56] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_59 
+ bl[57] br[57] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_60 
+ bl[58] br[58] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_61 
+ bl[59] br[59] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_62 
+ bl[60] br[60] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_63 
+ bl[61] br[61] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_64 
+ bl[62] br[62] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_65 
+ bl[63] br[63] vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_66 
+ vdd vdd vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_331_67 
+ vdd vdd vdd vss wl[329] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_0 
+ vdd vdd vss vdd vpb vnb wl[330] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_332_1 
+ rbl rbr vss vdd vpb vnb wl[330] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_332_2 
+ bl[0] br[0] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_3 
+ bl[1] br[1] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_4 
+ bl[2] br[2] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_5 
+ bl[3] br[3] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_6 
+ bl[4] br[4] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_7 
+ bl[5] br[5] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_8 
+ bl[6] br[6] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_9 
+ bl[7] br[7] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_10 
+ bl[8] br[8] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_11 
+ bl[9] br[9] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_12 
+ bl[10] br[10] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_13 
+ bl[11] br[11] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_14 
+ bl[12] br[12] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_15 
+ bl[13] br[13] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_16 
+ bl[14] br[14] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_17 
+ bl[15] br[15] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_18 
+ bl[16] br[16] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_19 
+ bl[17] br[17] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_20 
+ bl[18] br[18] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_21 
+ bl[19] br[19] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_22 
+ bl[20] br[20] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_23 
+ bl[21] br[21] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_24 
+ bl[22] br[22] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_25 
+ bl[23] br[23] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_26 
+ bl[24] br[24] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_27 
+ bl[25] br[25] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_28 
+ bl[26] br[26] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_29 
+ bl[27] br[27] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_30 
+ bl[28] br[28] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_31 
+ bl[29] br[29] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_32 
+ bl[30] br[30] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_33 
+ bl[31] br[31] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_34 
+ bl[32] br[32] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_35 
+ bl[33] br[33] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_36 
+ bl[34] br[34] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_37 
+ bl[35] br[35] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_38 
+ bl[36] br[36] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_39 
+ bl[37] br[37] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_40 
+ bl[38] br[38] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_41 
+ bl[39] br[39] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_42 
+ bl[40] br[40] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_43 
+ bl[41] br[41] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_44 
+ bl[42] br[42] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_45 
+ bl[43] br[43] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_46 
+ bl[44] br[44] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_47 
+ bl[45] br[45] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_48 
+ bl[46] br[46] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_49 
+ bl[47] br[47] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_50 
+ bl[48] br[48] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_51 
+ bl[49] br[49] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_52 
+ bl[50] br[50] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_53 
+ bl[51] br[51] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_54 
+ bl[52] br[52] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_55 
+ bl[53] br[53] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_56 
+ bl[54] br[54] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_57 
+ bl[55] br[55] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_58 
+ bl[56] br[56] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_59 
+ bl[57] br[57] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_60 
+ bl[58] br[58] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_61 
+ bl[59] br[59] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_62 
+ bl[60] br[60] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_63 
+ bl[61] br[61] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_64 
+ bl[62] br[62] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_65 
+ bl[63] br[63] vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_66 
+ vdd vdd vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_332_67 
+ vdd vdd vdd vss wl[330] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_0 
+ vdd vdd vss vdd vpb vnb wl[331] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_333_1 
+ rbl rbr vss vdd vpb vnb wl[331] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_333_2 
+ bl[0] br[0] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_3 
+ bl[1] br[1] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_4 
+ bl[2] br[2] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_5 
+ bl[3] br[3] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_6 
+ bl[4] br[4] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_7 
+ bl[5] br[5] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_8 
+ bl[6] br[6] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_9 
+ bl[7] br[7] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_10 
+ bl[8] br[8] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_11 
+ bl[9] br[9] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_12 
+ bl[10] br[10] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_13 
+ bl[11] br[11] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_14 
+ bl[12] br[12] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_15 
+ bl[13] br[13] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_16 
+ bl[14] br[14] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_17 
+ bl[15] br[15] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_18 
+ bl[16] br[16] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_19 
+ bl[17] br[17] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_20 
+ bl[18] br[18] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_21 
+ bl[19] br[19] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_22 
+ bl[20] br[20] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_23 
+ bl[21] br[21] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_24 
+ bl[22] br[22] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_25 
+ bl[23] br[23] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_26 
+ bl[24] br[24] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_27 
+ bl[25] br[25] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_28 
+ bl[26] br[26] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_29 
+ bl[27] br[27] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_30 
+ bl[28] br[28] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_31 
+ bl[29] br[29] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_32 
+ bl[30] br[30] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_33 
+ bl[31] br[31] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_34 
+ bl[32] br[32] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_35 
+ bl[33] br[33] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_36 
+ bl[34] br[34] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_37 
+ bl[35] br[35] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_38 
+ bl[36] br[36] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_39 
+ bl[37] br[37] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_40 
+ bl[38] br[38] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_41 
+ bl[39] br[39] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_42 
+ bl[40] br[40] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_43 
+ bl[41] br[41] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_44 
+ bl[42] br[42] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_45 
+ bl[43] br[43] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_46 
+ bl[44] br[44] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_47 
+ bl[45] br[45] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_48 
+ bl[46] br[46] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_49 
+ bl[47] br[47] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_50 
+ bl[48] br[48] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_51 
+ bl[49] br[49] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_52 
+ bl[50] br[50] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_53 
+ bl[51] br[51] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_54 
+ bl[52] br[52] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_55 
+ bl[53] br[53] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_56 
+ bl[54] br[54] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_57 
+ bl[55] br[55] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_58 
+ bl[56] br[56] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_59 
+ bl[57] br[57] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_60 
+ bl[58] br[58] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_61 
+ bl[59] br[59] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_62 
+ bl[60] br[60] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_63 
+ bl[61] br[61] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_64 
+ bl[62] br[62] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_65 
+ bl[63] br[63] vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_66 
+ vdd vdd vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_333_67 
+ vdd vdd vdd vss wl[331] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_0 
+ vdd vdd vss vdd vpb vnb wl[332] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_334_1 
+ rbl rbr vss vdd vpb vnb wl[332] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_334_2 
+ bl[0] br[0] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_3 
+ bl[1] br[1] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_4 
+ bl[2] br[2] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_5 
+ bl[3] br[3] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_6 
+ bl[4] br[4] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_7 
+ bl[5] br[5] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_8 
+ bl[6] br[6] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_9 
+ bl[7] br[7] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_10 
+ bl[8] br[8] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_11 
+ bl[9] br[9] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_12 
+ bl[10] br[10] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_13 
+ bl[11] br[11] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_14 
+ bl[12] br[12] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_15 
+ bl[13] br[13] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_16 
+ bl[14] br[14] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_17 
+ bl[15] br[15] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_18 
+ bl[16] br[16] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_19 
+ bl[17] br[17] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_20 
+ bl[18] br[18] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_21 
+ bl[19] br[19] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_22 
+ bl[20] br[20] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_23 
+ bl[21] br[21] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_24 
+ bl[22] br[22] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_25 
+ bl[23] br[23] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_26 
+ bl[24] br[24] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_27 
+ bl[25] br[25] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_28 
+ bl[26] br[26] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_29 
+ bl[27] br[27] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_30 
+ bl[28] br[28] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_31 
+ bl[29] br[29] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_32 
+ bl[30] br[30] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_33 
+ bl[31] br[31] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_34 
+ bl[32] br[32] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_35 
+ bl[33] br[33] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_36 
+ bl[34] br[34] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_37 
+ bl[35] br[35] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_38 
+ bl[36] br[36] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_39 
+ bl[37] br[37] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_40 
+ bl[38] br[38] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_41 
+ bl[39] br[39] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_42 
+ bl[40] br[40] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_43 
+ bl[41] br[41] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_44 
+ bl[42] br[42] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_45 
+ bl[43] br[43] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_46 
+ bl[44] br[44] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_47 
+ bl[45] br[45] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_48 
+ bl[46] br[46] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_49 
+ bl[47] br[47] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_50 
+ bl[48] br[48] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_51 
+ bl[49] br[49] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_52 
+ bl[50] br[50] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_53 
+ bl[51] br[51] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_54 
+ bl[52] br[52] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_55 
+ bl[53] br[53] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_56 
+ bl[54] br[54] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_57 
+ bl[55] br[55] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_58 
+ bl[56] br[56] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_59 
+ bl[57] br[57] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_60 
+ bl[58] br[58] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_61 
+ bl[59] br[59] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_62 
+ bl[60] br[60] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_63 
+ bl[61] br[61] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_64 
+ bl[62] br[62] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_65 
+ bl[63] br[63] vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_66 
+ vdd vdd vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_334_67 
+ vdd vdd vdd vss wl[332] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_0 
+ vdd vdd vss vdd vpb vnb wl[333] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_335_1 
+ rbl rbr vss vdd vpb vnb wl[333] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_335_2 
+ bl[0] br[0] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_3 
+ bl[1] br[1] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_4 
+ bl[2] br[2] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_5 
+ bl[3] br[3] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_6 
+ bl[4] br[4] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_7 
+ bl[5] br[5] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_8 
+ bl[6] br[6] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_9 
+ bl[7] br[7] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_10 
+ bl[8] br[8] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_11 
+ bl[9] br[9] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_12 
+ bl[10] br[10] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_13 
+ bl[11] br[11] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_14 
+ bl[12] br[12] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_15 
+ bl[13] br[13] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_16 
+ bl[14] br[14] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_17 
+ bl[15] br[15] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_18 
+ bl[16] br[16] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_19 
+ bl[17] br[17] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_20 
+ bl[18] br[18] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_21 
+ bl[19] br[19] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_22 
+ bl[20] br[20] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_23 
+ bl[21] br[21] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_24 
+ bl[22] br[22] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_25 
+ bl[23] br[23] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_26 
+ bl[24] br[24] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_27 
+ bl[25] br[25] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_28 
+ bl[26] br[26] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_29 
+ bl[27] br[27] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_30 
+ bl[28] br[28] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_31 
+ bl[29] br[29] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_32 
+ bl[30] br[30] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_33 
+ bl[31] br[31] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_34 
+ bl[32] br[32] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_35 
+ bl[33] br[33] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_36 
+ bl[34] br[34] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_37 
+ bl[35] br[35] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_38 
+ bl[36] br[36] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_39 
+ bl[37] br[37] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_40 
+ bl[38] br[38] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_41 
+ bl[39] br[39] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_42 
+ bl[40] br[40] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_43 
+ bl[41] br[41] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_44 
+ bl[42] br[42] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_45 
+ bl[43] br[43] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_46 
+ bl[44] br[44] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_47 
+ bl[45] br[45] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_48 
+ bl[46] br[46] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_49 
+ bl[47] br[47] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_50 
+ bl[48] br[48] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_51 
+ bl[49] br[49] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_52 
+ bl[50] br[50] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_53 
+ bl[51] br[51] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_54 
+ bl[52] br[52] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_55 
+ bl[53] br[53] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_56 
+ bl[54] br[54] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_57 
+ bl[55] br[55] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_58 
+ bl[56] br[56] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_59 
+ bl[57] br[57] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_60 
+ bl[58] br[58] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_61 
+ bl[59] br[59] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_62 
+ bl[60] br[60] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_63 
+ bl[61] br[61] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_64 
+ bl[62] br[62] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_65 
+ bl[63] br[63] vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_66 
+ vdd vdd vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_335_67 
+ vdd vdd vdd vss wl[333] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_0 
+ vdd vdd vss vdd vpb vnb wl[334] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_336_1 
+ rbl rbr vss vdd vpb vnb wl[334] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_336_2 
+ bl[0] br[0] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_3 
+ bl[1] br[1] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_4 
+ bl[2] br[2] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_5 
+ bl[3] br[3] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_6 
+ bl[4] br[4] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_7 
+ bl[5] br[5] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_8 
+ bl[6] br[6] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_9 
+ bl[7] br[7] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_10 
+ bl[8] br[8] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_11 
+ bl[9] br[9] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_12 
+ bl[10] br[10] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_13 
+ bl[11] br[11] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_14 
+ bl[12] br[12] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_15 
+ bl[13] br[13] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_16 
+ bl[14] br[14] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_17 
+ bl[15] br[15] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_18 
+ bl[16] br[16] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_19 
+ bl[17] br[17] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_20 
+ bl[18] br[18] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_21 
+ bl[19] br[19] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_22 
+ bl[20] br[20] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_23 
+ bl[21] br[21] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_24 
+ bl[22] br[22] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_25 
+ bl[23] br[23] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_26 
+ bl[24] br[24] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_27 
+ bl[25] br[25] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_28 
+ bl[26] br[26] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_29 
+ bl[27] br[27] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_30 
+ bl[28] br[28] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_31 
+ bl[29] br[29] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_32 
+ bl[30] br[30] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_33 
+ bl[31] br[31] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_34 
+ bl[32] br[32] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_35 
+ bl[33] br[33] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_36 
+ bl[34] br[34] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_37 
+ bl[35] br[35] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_38 
+ bl[36] br[36] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_39 
+ bl[37] br[37] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_40 
+ bl[38] br[38] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_41 
+ bl[39] br[39] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_42 
+ bl[40] br[40] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_43 
+ bl[41] br[41] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_44 
+ bl[42] br[42] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_45 
+ bl[43] br[43] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_46 
+ bl[44] br[44] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_47 
+ bl[45] br[45] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_48 
+ bl[46] br[46] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_49 
+ bl[47] br[47] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_50 
+ bl[48] br[48] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_51 
+ bl[49] br[49] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_52 
+ bl[50] br[50] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_53 
+ bl[51] br[51] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_54 
+ bl[52] br[52] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_55 
+ bl[53] br[53] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_56 
+ bl[54] br[54] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_57 
+ bl[55] br[55] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_58 
+ bl[56] br[56] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_59 
+ bl[57] br[57] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_60 
+ bl[58] br[58] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_61 
+ bl[59] br[59] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_62 
+ bl[60] br[60] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_63 
+ bl[61] br[61] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_64 
+ bl[62] br[62] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_65 
+ bl[63] br[63] vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_66 
+ vdd vdd vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_336_67 
+ vdd vdd vdd vss wl[334] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_0 
+ vdd vdd vss vdd vpb vnb wl[335] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_337_1 
+ rbl rbr vss vdd vpb vnb wl[335] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_337_2 
+ bl[0] br[0] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_3 
+ bl[1] br[1] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_4 
+ bl[2] br[2] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_5 
+ bl[3] br[3] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_6 
+ bl[4] br[4] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_7 
+ bl[5] br[5] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_8 
+ bl[6] br[6] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_9 
+ bl[7] br[7] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_10 
+ bl[8] br[8] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_11 
+ bl[9] br[9] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_12 
+ bl[10] br[10] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_13 
+ bl[11] br[11] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_14 
+ bl[12] br[12] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_15 
+ bl[13] br[13] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_16 
+ bl[14] br[14] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_17 
+ bl[15] br[15] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_18 
+ bl[16] br[16] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_19 
+ bl[17] br[17] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_20 
+ bl[18] br[18] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_21 
+ bl[19] br[19] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_22 
+ bl[20] br[20] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_23 
+ bl[21] br[21] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_24 
+ bl[22] br[22] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_25 
+ bl[23] br[23] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_26 
+ bl[24] br[24] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_27 
+ bl[25] br[25] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_28 
+ bl[26] br[26] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_29 
+ bl[27] br[27] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_30 
+ bl[28] br[28] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_31 
+ bl[29] br[29] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_32 
+ bl[30] br[30] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_33 
+ bl[31] br[31] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_34 
+ bl[32] br[32] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_35 
+ bl[33] br[33] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_36 
+ bl[34] br[34] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_37 
+ bl[35] br[35] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_38 
+ bl[36] br[36] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_39 
+ bl[37] br[37] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_40 
+ bl[38] br[38] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_41 
+ bl[39] br[39] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_42 
+ bl[40] br[40] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_43 
+ bl[41] br[41] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_44 
+ bl[42] br[42] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_45 
+ bl[43] br[43] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_46 
+ bl[44] br[44] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_47 
+ bl[45] br[45] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_48 
+ bl[46] br[46] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_49 
+ bl[47] br[47] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_50 
+ bl[48] br[48] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_51 
+ bl[49] br[49] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_52 
+ bl[50] br[50] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_53 
+ bl[51] br[51] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_54 
+ bl[52] br[52] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_55 
+ bl[53] br[53] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_56 
+ bl[54] br[54] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_57 
+ bl[55] br[55] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_58 
+ bl[56] br[56] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_59 
+ bl[57] br[57] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_60 
+ bl[58] br[58] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_61 
+ bl[59] br[59] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_62 
+ bl[60] br[60] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_63 
+ bl[61] br[61] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_64 
+ bl[62] br[62] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_65 
+ bl[63] br[63] vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_66 
+ vdd vdd vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_337_67 
+ vdd vdd vdd vss wl[335] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_0 
+ vdd vdd vss vdd vpb vnb wl[336] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_338_1 
+ rbl rbr vss vdd vpb vnb wl[336] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_338_2 
+ bl[0] br[0] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_3 
+ bl[1] br[1] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_4 
+ bl[2] br[2] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_5 
+ bl[3] br[3] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_6 
+ bl[4] br[4] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_7 
+ bl[5] br[5] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_8 
+ bl[6] br[6] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_9 
+ bl[7] br[7] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_10 
+ bl[8] br[8] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_11 
+ bl[9] br[9] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_12 
+ bl[10] br[10] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_13 
+ bl[11] br[11] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_14 
+ bl[12] br[12] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_15 
+ bl[13] br[13] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_16 
+ bl[14] br[14] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_17 
+ bl[15] br[15] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_18 
+ bl[16] br[16] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_19 
+ bl[17] br[17] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_20 
+ bl[18] br[18] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_21 
+ bl[19] br[19] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_22 
+ bl[20] br[20] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_23 
+ bl[21] br[21] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_24 
+ bl[22] br[22] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_25 
+ bl[23] br[23] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_26 
+ bl[24] br[24] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_27 
+ bl[25] br[25] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_28 
+ bl[26] br[26] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_29 
+ bl[27] br[27] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_30 
+ bl[28] br[28] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_31 
+ bl[29] br[29] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_32 
+ bl[30] br[30] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_33 
+ bl[31] br[31] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_34 
+ bl[32] br[32] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_35 
+ bl[33] br[33] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_36 
+ bl[34] br[34] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_37 
+ bl[35] br[35] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_38 
+ bl[36] br[36] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_39 
+ bl[37] br[37] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_40 
+ bl[38] br[38] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_41 
+ bl[39] br[39] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_42 
+ bl[40] br[40] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_43 
+ bl[41] br[41] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_44 
+ bl[42] br[42] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_45 
+ bl[43] br[43] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_46 
+ bl[44] br[44] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_47 
+ bl[45] br[45] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_48 
+ bl[46] br[46] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_49 
+ bl[47] br[47] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_50 
+ bl[48] br[48] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_51 
+ bl[49] br[49] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_52 
+ bl[50] br[50] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_53 
+ bl[51] br[51] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_54 
+ bl[52] br[52] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_55 
+ bl[53] br[53] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_56 
+ bl[54] br[54] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_57 
+ bl[55] br[55] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_58 
+ bl[56] br[56] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_59 
+ bl[57] br[57] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_60 
+ bl[58] br[58] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_61 
+ bl[59] br[59] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_62 
+ bl[60] br[60] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_63 
+ bl[61] br[61] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_64 
+ bl[62] br[62] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_65 
+ bl[63] br[63] vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_66 
+ vdd vdd vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_338_67 
+ vdd vdd vdd vss wl[336] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_0 
+ vdd vdd vss vdd vpb vnb wl[337] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_339_1 
+ rbl rbr vss vdd vpb vnb wl[337] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_339_2 
+ bl[0] br[0] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_3 
+ bl[1] br[1] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_4 
+ bl[2] br[2] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_5 
+ bl[3] br[3] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_6 
+ bl[4] br[4] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_7 
+ bl[5] br[5] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_8 
+ bl[6] br[6] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_9 
+ bl[7] br[7] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_10 
+ bl[8] br[8] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_11 
+ bl[9] br[9] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_12 
+ bl[10] br[10] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_13 
+ bl[11] br[11] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_14 
+ bl[12] br[12] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_15 
+ bl[13] br[13] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_16 
+ bl[14] br[14] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_17 
+ bl[15] br[15] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_18 
+ bl[16] br[16] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_19 
+ bl[17] br[17] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_20 
+ bl[18] br[18] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_21 
+ bl[19] br[19] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_22 
+ bl[20] br[20] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_23 
+ bl[21] br[21] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_24 
+ bl[22] br[22] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_25 
+ bl[23] br[23] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_26 
+ bl[24] br[24] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_27 
+ bl[25] br[25] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_28 
+ bl[26] br[26] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_29 
+ bl[27] br[27] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_30 
+ bl[28] br[28] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_31 
+ bl[29] br[29] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_32 
+ bl[30] br[30] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_33 
+ bl[31] br[31] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_34 
+ bl[32] br[32] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_35 
+ bl[33] br[33] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_36 
+ bl[34] br[34] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_37 
+ bl[35] br[35] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_38 
+ bl[36] br[36] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_39 
+ bl[37] br[37] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_40 
+ bl[38] br[38] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_41 
+ bl[39] br[39] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_42 
+ bl[40] br[40] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_43 
+ bl[41] br[41] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_44 
+ bl[42] br[42] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_45 
+ bl[43] br[43] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_46 
+ bl[44] br[44] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_47 
+ bl[45] br[45] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_48 
+ bl[46] br[46] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_49 
+ bl[47] br[47] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_50 
+ bl[48] br[48] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_51 
+ bl[49] br[49] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_52 
+ bl[50] br[50] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_53 
+ bl[51] br[51] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_54 
+ bl[52] br[52] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_55 
+ bl[53] br[53] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_56 
+ bl[54] br[54] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_57 
+ bl[55] br[55] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_58 
+ bl[56] br[56] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_59 
+ bl[57] br[57] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_60 
+ bl[58] br[58] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_61 
+ bl[59] br[59] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_62 
+ bl[60] br[60] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_63 
+ bl[61] br[61] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_64 
+ bl[62] br[62] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_65 
+ bl[63] br[63] vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_66 
+ vdd vdd vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_339_67 
+ vdd vdd vdd vss wl[337] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_0 
+ vdd vdd vss vdd vpb vnb wl[338] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_340_1 
+ rbl rbr vss vdd vpb vnb wl[338] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_340_2 
+ bl[0] br[0] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_3 
+ bl[1] br[1] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_4 
+ bl[2] br[2] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_5 
+ bl[3] br[3] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_6 
+ bl[4] br[4] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_7 
+ bl[5] br[5] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_8 
+ bl[6] br[6] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_9 
+ bl[7] br[7] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_10 
+ bl[8] br[8] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_11 
+ bl[9] br[9] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_12 
+ bl[10] br[10] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_13 
+ bl[11] br[11] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_14 
+ bl[12] br[12] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_15 
+ bl[13] br[13] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_16 
+ bl[14] br[14] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_17 
+ bl[15] br[15] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_18 
+ bl[16] br[16] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_19 
+ bl[17] br[17] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_20 
+ bl[18] br[18] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_21 
+ bl[19] br[19] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_22 
+ bl[20] br[20] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_23 
+ bl[21] br[21] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_24 
+ bl[22] br[22] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_25 
+ bl[23] br[23] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_26 
+ bl[24] br[24] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_27 
+ bl[25] br[25] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_28 
+ bl[26] br[26] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_29 
+ bl[27] br[27] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_30 
+ bl[28] br[28] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_31 
+ bl[29] br[29] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_32 
+ bl[30] br[30] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_33 
+ bl[31] br[31] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_34 
+ bl[32] br[32] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_35 
+ bl[33] br[33] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_36 
+ bl[34] br[34] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_37 
+ bl[35] br[35] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_38 
+ bl[36] br[36] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_39 
+ bl[37] br[37] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_40 
+ bl[38] br[38] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_41 
+ bl[39] br[39] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_42 
+ bl[40] br[40] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_43 
+ bl[41] br[41] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_44 
+ bl[42] br[42] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_45 
+ bl[43] br[43] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_46 
+ bl[44] br[44] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_47 
+ bl[45] br[45] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_48 
+ bl[46] br[46] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_49 
+ bl[47] br[47] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_50 
+ bl[48] br[48] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_51 
+ bl[49] br[49] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_52 
+ bl[50] br[50] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_53 
+ bl[51] br[51] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_54 
+ bl[52] br[52] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_55 
+ bl[53] br[53] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_56 
+ bl[54] br[54] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_57 
+ bl[55] br[55] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_58 
+ bl[56] br[56] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_59 
+ bl[57] br[57] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_60 
+ bl[58] br[58] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_61 
+ bl[59] br[59] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_62 
+ bl[60] br[60] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_63 
+ bl[61] br[61] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_64 
+ bl[62] br[62] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_65 
+ bl[63] br[63] vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_66 
+ vdd vdd vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_340_67 
+ vdd vdd vdd vss wl[338] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_0 
+ vdd vdd vss vdd vpb vnb wl[339] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_341_1 
+ rbl rbr vss vdd vpb vnb wl[339] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_341_2 
+ bl[0] br[0] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_3 
+ bl[1] br[1] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_4 
+ bl[2] br[2] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_5 
+ bl[3] br[3] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_6 
+ bl[4] br[4] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_7 
+ bl[5] br[5] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_8 
+ bl[6] br[6] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_9 
+ bl[7] br[7] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_10 
+ bl[8] br[8] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_11 
+ bl[9] br[9] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_12 
+ bl[10] br[10] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_13 
+ bl[11] br[11] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_14 
+ bl[12] br[12] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_15 
+ bl[13] br[13] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_16 
+ bl[14] br[14] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_17 
+ bl[15] br[15] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_18 
+ bl[16] br[16] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_19 
+ bl[17] br[17] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_20 
+ bl[18] br[18] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_21 
+ bl[19] br[19] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_22 
+ bl[20] br[20] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_23 
+ bl[21] br[21] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_24 
+ bl[22] br[22] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_25 
+ bl[23] br[23] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_26 
+ bl[24] br[24] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_27 
+ bl[25] br[25] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_28 
+ bl[26] br[26] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_29 
+ bl[27] br[27] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_30 
+ bl[28] br[28] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_31 
+ bl[29] br[29] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_32 
+ bl[30] br[30] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_33 
+ bl[31] br[31] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_34 
+ bl[32] br[32] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_35 
+ bl[33] br[33] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_36 
+ bl[34] br[34] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_37 
+ bl[35] br[35] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_38 
+ bl[36] br[36] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_39 
+ bl[37] br[37] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_40 
+ bl[38] br[38] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_41 
+ bl[39] br[39] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_42 
+ bl[40] br[40] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_43 
+ bl[41] br[41] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_44 
+ bl[42] br[42] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_45 
+ bl[43] br[43] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_46 
+ bl[44] br[44] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_47 
+ bl[45] br[45] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_48 
+ bl[46] br[46] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_49 
+ bl[47] br[47] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_50 
+ bl[48] br[48] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_51 
+ bl[49] br[49] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_52 
+ bl[50] br[50] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_53 
+ bl[51] br[51] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_54 
+ bl[52] br[52] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_55 
+ bl[53] br[53] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_56 
+ bl[54] br[54] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_57 
+ bl[55] br[55] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_58 
+ bl[56] br[56] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_59 
+ bl[57] br[57] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_60 
+ bl[58] br[58] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_61 
+ bl[59] br[59] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_62 
+ bl[60] br[60] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_63 
+ bl[61] br[61] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_64 
+ bl[62] br[62] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_65 
+ bl[63] br[63] vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_66 
+ vdd vdd vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_341_67 
+ vdd vdd vdd vss wl[339] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_0 
+ vdd vdd vss vdd vpb vnb wl[340] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_342_1 
+ rbl rbr vss vdd vpb vnb wl[340] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_342_2 
+ bl[0] br[0] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_3 
+ bl[1] br[1] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_4 
+ bl[2] br[2] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_5 
+ bl[3] br[3] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_6 
+ bl[4] br[4] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_7 
+ bl[5] br[5] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_8 
+ bl[6] br[6] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_9 
+ bl[7] br[7] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_10 
+ bl[8] br[8] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_11 
+ bl[9] br[9] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_12 
+ bl[10] br[10] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_13 
+ bl[11] br[11] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_14 
+ bl[12] br[12] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_15 
+ bl[13] br[13] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_16 
+ bl[14] br[14] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_17 
+ bl[15] br[15] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_18 
+ bl[16] br[16] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_19 
+ bl[17] br[17] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_20 
+ bl[18] br[18] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_21 
+ bl[19] br[19] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_22 
+ bl[20] br[20] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_23 
+ bl[21] br[21] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_24 
+ bl[22] br[22] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_25 
+ bl[23] br[23] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_26 
+ bl[24] br[24] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_27 
+ bl[25] br[25] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_28 
+ bl[26] br[26] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_29 
+ bl[27] br[27] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_30 
+ bl[28] br[28] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_31 
+ bl[29] br[29] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_32 
+ bl[30] br[30] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_33 
+ bl[31] br[31] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_34 
+ bl[32] br[32] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_35 
+ bl[33] br[33] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_36 
+ bl[34] br[34] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_37 
+ bl[35] br[35] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_38 
+ bl[36] br[36] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_39 
+ bl[37] br[37] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_40 
+ bl[38] br[38] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_41 
+ bl[39] br[39] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_42 
+ bl[40] br[40] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_43 
+ bl[41] br[41] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_44 
+ bl[42] br[42] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_45 
+ bl[43] br[43] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_46 
+ bl[44] br[44] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_47 
+ bl[45] br[45] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_48 
+ bl[46] br[46] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_49 
+ bl[47] br[47] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_50 
+ bl[48] br[48] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_51 
+ bl[49] br[49] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_52 
+ bl[50] br[50] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_53 
+ bl[51] br[51] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_54 
+ bl[52] br[52] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_55 
+ bl[53] br[53] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_56 
+ bl[54] br[54] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_57 
+ bl[55] br[55] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_58 
+ bl[56] br[56] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_59 
+ bl[57] br[57] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_60 
+ bl[58] br[58] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_61 
+ bl[59] br[59] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_62 
+ bl[60] br[60] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_63 
+ bl[61] br[61] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_64 
+ bl[62] br[62] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_65 
+ bl[63] br[63] vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_66 
+ vdd vdd vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_342_67 
+ vdd vdd vdd vss wl[340] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_0 
+ vdd vdd vss vdd vpb vnb wl[341] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_343_1 
+ rbl rbr vss vdd vpb vnb wl[341] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_343_2 
+ bl[0] br[0] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_3 
+ bl[1] br[1] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_4 
+ bl[2] br[2] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_5 
+ bl[3] br[3] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_6 
+ bl[4] br[4] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_7 
+ bl[5] br[5] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_8 
+ bl[6] br[6] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_9 
+ bl[7] br[7] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_10 
+ bl[8] br[8] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_11 
+ bl[9] br[9] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_12 
+ bl[10] br[10] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_13 
+ bl[11] br[11] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_14 
+ bl[12] br[12] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_15 
+ bl[13] br[13] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_16 
+ bl[14] br[14] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_17 
+ bl[15] br[15] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_18 
+ bl[16] br[16] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_19 
+ bl[17] br[17] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_20 
+ bl[18] br[18] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_21 
+ bl[19] br[19] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_22 
+ bl[20] br[20] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_23 
+ bl[21] br[21] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_24 
+ bl[22] br[22] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_25 
+ bl[23] br[23] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_26 
+ bl[24] br[24] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_27 
+ bl[25] br[25] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_28 
+ bl[26] br[26] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_29 
+ bl[27] br[27] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_30 
+ bl[28] br[28] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_31 
+ bl[29] br[29] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_32 
+ bl[30] br[30] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_33 
+ bl[31] br[31] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_34 
+ bl[32] br[32] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_35 
+ bl[33] br[33] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_36 
+ bl[34] br[34] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_37 
+ bl[35] br[35] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_38 
+ bl[36] br[36] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_39 
+ bl[37] br[37] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_40 
+ bl[38] br[38] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_41 
+ bl[39] br[39] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_42 
+ bl[40] br[40] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_43 
+ bl[41] br[41] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_44 
+ bl[42] br[42] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_45 
+ bl[43] br[43] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_46 
+ bl[44] br[44] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_47 
+ bl[45] br[45] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_48 
+ bl[46] br[46] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_49 
+ bl[47] br[47] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_50 
+ bl[48] br[48] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_51 
+ bl[49] br[49] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_52 
+ bl[50] br[50] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_53 
+ bl[51] br[51] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_54 
+ bl[52] br[52] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_55 
+ bl[53] br[53] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_56 
+ bl[54] br[54] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_57 
+ bl[55] br[55] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_58 
+ bl[56] br[56] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_59 
+ bl[57] br[57] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_60 
+ bl[58] br[58] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_61 
+ bl[59] br[59] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_62 
+ bl[60] br[60] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_63 
+ bl[61] br[61] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_64 
+ bl[62] br[62] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_65 
+ bl[63] br[63] vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_66 
+ vdd vdd vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_343_67 
+ vdd vdd vdd vss wl[341] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_0 
+ vdd vdd vss vdd vpb vnb wl[342] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_344_1 
+ rbl rbr vss vdd vpb vnb wl[342] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_344_2 
+ bl[0] br[0] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_3 
+ bl[1] br[1] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_4 
+ bl[2] br[2] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_5 
+ bl[3] br[3] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_6 
+ bl[4] br[4] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_7 
+ bl[5] br[5] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_8 
+ bl[6] br[6] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_9 
+ bl[7] br[7] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_10 
+ bl[8] br[8] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_11 
+ bl[9] br[9] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_12 
+ bl[10] br[10] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_13 
+ bl[11] br[11] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_14 
+ bl[12] br[12] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_15 
+ bl[13] br[13] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_16 
+ bl[14] br[14] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_17 
+ bl[15] br[15] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_18 
+ bl[16] br[16] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_19 
+ bl[17] br[17] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_20 
+ bl[18] br[18] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_21 
+ bl[19] br[19] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_22 
+ bl[20] br[20] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_23 
+ bl[21] br[21] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_24 
+ bl[22] br[22] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_25 
+ bl[23] br[23] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_26 
+ bl[24] br[24] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_27 
+ bl[25] br[25] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_28 
+ bl[26] br[26] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_29 
+ bl[27] br[27] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_30 
+ bl[28] br[28] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_31 
+ bl[29] br[29] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_32 
+ bl[30] br[30] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_33 
+ bl[31] br[31] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_34 
+ bl[32] br[32] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_35 
+ bl[33] br[33] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_36 
+ bl[34] br[34] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_37 
+ bl[35] br[35] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_38 
+ bl[36] br[36] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_39 
+ bl[37] br[37] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_40 
+ bl[38] br[38] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_41 
+ bl[39] br[39] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_42 
+ bl[40] br[40] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_43 
+ bl[41] br[41] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_44 
+ bl[42] br[42] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_45 
+ bl[43] br[43] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_46 
+ bl[44] br[44] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_47 
+ bl[45] br[45] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_48 
+ bl[46] br[46] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_49 
+ bl[47] br[47] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_50 
+ bl[48] br[48] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_51 
+ bl[49] br[49] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_52 
+ bl[50] br[50] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_53 
+ bl[51] br[51] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_54 
+ bl[52] br[52] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_55 
+ bl[53] br[53] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_56 
+ bl[54] br[54] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_57 
+ bl[55] br[55] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_58 
+ bl[56] br[56] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_59 
+ bl[57] br[57] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_60 
+ bl[58] br[58] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_61 
+ bl[59] br[59] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_62 
+ bl[60] br[60] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_63 
+ bl[61] br[61] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_64 
+ bl[62] br[62] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_65 
+ bl[63] br[63] vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_66 
+ vdd vdd vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_344_67 
+ vdd vdd vdd vss wl[342] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_0 
+ vdd vdd vss vdd vpb vnb wl[343] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_345_1 
+ rbl rbr vss vdd vpb vnb wl[343] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_345_2 
+ bl[0] br[0] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_3 
+ bl[1] br[1] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_4 
+ bl[2] br[2] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_5 
+ bl[3] br[3] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_6 
+ bl[4] br[4] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_7 
+ bl[5] br[5] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_8 
+ bl[6] br[6] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_9 
+ bl[7] br[7] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_10 
+ bl[8] br[8] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_11 
+ bl[9] br[9] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_12 
+ bl[10] br[10] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_13 
+ bl[11] br[11] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_14 
+ bl[12] br[12] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_15 
+ bl[13] br[13] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_16 
+ bl[14] br[14] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_17 
+ bl[15] br[15] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_18 
+ bl[16] br[16] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_19 
+ bl[17] br[17] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_20 
+ bl[18] br[18] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_21 
+ bl[19] br[19] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_22 
+ bl[20] br[20] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_23 
+ bl[21] br[21] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_24 
+ bl[22] br[22] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_25 
+ bl[23] br[23] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_26 
+ bl[24] br[24] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_27 
+ bl[25] br[25] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_28 
+ bl[26] br[26] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_29 
+ bl[27] br[27] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_30 
+ bl[28] br[28] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_31 
+ bl[29] br[29] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_32 
+ bl[30] br[30] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_33 
+ bl[31] br[31] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_34 
+ bl[32] br[32] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_35 
+ bl[33] br[33] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_36 
+ bl[34] br[34] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_37 
+ bl[35] br[35] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_38 
+ bl[36] br[36] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_39 
+ bl[37] br[37] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_40 
+ bl[38] br[38] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_41 
+ bl[39] br[39] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_42 
+ bl[40] br[40] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_43 
+ bl[41] br[41] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_44 
+ bl[42] br[42] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_45 
+ bl[43] br[43] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_46 
+ bl[44] br[44] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_47 
+ bl[45] br[45] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_48 
+ bl[46] br[46] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_49 
+ bl[47] br[47] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_50 
+ bl[48] br[48] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_51 
+ bl[49] br[49] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_52 
+ bl[50] br[50] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_53 
+ bl[51] br[51] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_54 
+ bl[52] br[52] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_55 
+ bl[53] br[53] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_56 
+ bl[54] br[54] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_57 
+ bl[55] br[55] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_58 
+ bl[56] br[56] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_59 
+ bl[57] br[57] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_60 
+ bl[58] br[58] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_61 
+ bl[59] br[59] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_62 
+ bl[60] br[60] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_63 
+ bl[61] br[61] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_64 
+ bl[62] br[62] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_65 
+ bl[63] br[63] vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_66 
+ vdd vdd vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_345_67 
+ vdd vdd vdd vss wl[343] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_0 
+ vdd vdd vss vdd vpb vnb wl[344] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_346_1 
+ rbl rbr vss vdd vpb vnb wl[344] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_346_2 
+ bl[0] br[0] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_3 
+ bl[1] br[1] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_4 
+ bl[2] br[2] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_5 
+ bl[3] br[3] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_6 
+ bl[4] br[4] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_7 
+ bl[5] br[5] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_8 
+ bl[6] br[6] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_9 
+ bl[7] br[7] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_10 
+ bl[8] br[8] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_11 
+ bl[9] br[9] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_12 
+ bl[10] br[10] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_13 
+ bl[11] br[11] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_14 
+ bl[12] br[12] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_15 
+ bl[13] br[13] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_16 
+ bl[14] br[14] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_17 
+ bl[15] br[15] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_18 
+ bl[16] br[16] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_19 
+ bl[17] br[17] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_20 
+ bl[18] br[18] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_21 
+ bl[19] br[19] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_22 
+ bl[20] br[20] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_23 
+ bl[21] br[21] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_24 
+ bl[22] br[22] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_25 
+ bl[23] br[23] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_26 
+ bl[24] br[24] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_27 
+ bl[25] br[25] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_28 
+ bl[26] br[26] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_29 
+ bl[27] br[27] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_30 
+ bl[28] br[28] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_31 
+ bl[29] br[29] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_32 
+ bl[30] br[30] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_33 
+ bl[31] br[31] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_34 
+ bl[32] br[32] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_35 
+ bl[33] br[33] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_36 
+ bl[34] br[34] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_37 
+ bl[35] br[35] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_38 
+ bl[36] br[36] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_39 
+ bl[37] br[37] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_40 
+ bl[38] br[38] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_41 
+ bl[39] br[39] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_42 
+ bl[40] br[40] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_43 
+ bl[41] br[41] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_44 
+ bl[42] br[42] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_45 
+ bl[43] br[43] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_46 
+ bl[44] br[44] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_47 
+ bl[45] br[45] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_48 
+ bl[46] br[46] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_49 
+ bl[47] br[47] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_50 
+ bl[48] br[48] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_51 
+ bl[49] br[49] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_52 
+ bl[50] br[50] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_53 
+ bl[51] br[51] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_54 
+ bl[52] br[52] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_55 
+ bl[53] br[53] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_56 
+ bl[54] br[54] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_57 
+ bl[55] br[55] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_58 
+ bl[56] br[56] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_59 
+ bl[57] br[57] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_60 
+ bl[58] br[58] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_61 
+ bl[59] br[59] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_62 
+ bl[60] br[60] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_63 
+ bl[61] br[61] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_64 
+ bl[62] br[62] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_65 
+ bl[63] br[63] vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_66 
+ vdd vdd vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_346_67 
+ vdd vdd vdd vss wl[344] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_0 
+ vdd vdd vss vdd vpb vnb wl[345] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_347_1 
+ rbl rbr vss vdd vpb vnb wl[345] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_347_2 
+ bl[0] br[0] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_3 
+ bl[1] br[1] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_4 
+ bl[2] br[2] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_5 
+ bl[3] br[3] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_6 
+ bl[4] br[4] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_7 
+ bl[5] br[5] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_8 
+ bl[6] br[6] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_9 
+ bl[7] br[7] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_10 
+ bl[8] br[8] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_11 
+ bl[9] br[9] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_12 
+ bl[10] br[10] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_13 
+ bl[11] br[11] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_14 
+ bl[12] br[12] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_15 
+ bl[13] br[13] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_16 
+ bl[14] br[14] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_17 
+ bl[15] br[15] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_18 
+ bl[16] br[16] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_19 
+ bl[17] br[17] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_20 
+ bl[18] br[18] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_21 
+ bl[19] br[19] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_22 
+ bl[20] br[20] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_23 
+ bl[21] br[21] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_24 
+ bl[22] br[22] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_25 
+ bl[23] br[23] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_26 
+ bl[24] br[24] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_27 
+ bl[25] br[25] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_28 
+ bl[26] br[26] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_29 
+ bl[27] br[27] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_30 
+ bl[28] br[28] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_31 
+ bl[29] br[29] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_32 
+ bl[30] br[30] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_33 
+ bl[31] br[31] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_34 
+ bl[32] br[32] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_35 
+ bl[33] br[33] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_36 
+ bl[34] br[34] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_37 
+ bl[35] br[35] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_38 
+ bl[36] br[36] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_39 
+ bl[37] br[37] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_40 
+ bl[38] br[38] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_41 
+ bl[39] br[39] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_42 
+ bl[40] br[40] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_43 
+ bl[41] br[41] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_44 
+ bl[42] br[42] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_45 
+ bl[43] br[43] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_46 
+ bl[44] br[44] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_47 
+ bl[45] br[45] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_48 
+ bl[46] br[46] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_49 
+ bl[47] br[47] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_50 
+ bl[48] br[48] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_51 
+ bl[49] br[49] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_52 
+ bl[50] br[50] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_53 
+ bl[51] br[51] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_54 
+ bl[52] br[52] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_55 
+ bl[53] br[53] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_56 
+ bl[54] br[54] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_57 
+ bl[55] br[55] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_58 
+ bl[56] br[56] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_59 
+ bl[57] br[57] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_60 
+ bl[58] br[58] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_61 
+ bl[59] br[59] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_62 
+ bl[60] br[60] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_63 
+ bl[61] br[61] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_64 
+ bl[62] br[62] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_65 
+ bl[63] br[63] vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_66 
+ vdd vdd vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_347_67 
+ vdd vdd vdd vss wl[345] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_0 
+ vdd vdd vss vdd vpb vnb wl[346] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_348_1 
+ rbl rbr vss vdd vpb vnb wl[346] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_348_2 
+ bl[0] br[0] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_3 
+ bl[1] br[1] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_4 
+ bl[2] br[2] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_5 
+ bl[3] br[3] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_6 
+ bl[4] br[4] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_7 
+ bl[5] br[5] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_8 
+ bl[6] br[6] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_9 
+ bl[7] br[7] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_10 
+ bl[8] br[8] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_11 
+ bl[9] br[9] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_12 
+ bl[10] br[10] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_13 
+ bl[11] br[11] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_14 
+ bl[12] br[12] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_15 
+ bl[13] br[13] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_16 
+ bl[14] br[14] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_17 
+ bl[15] br[15] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_18 
+ bl[16] br[16] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_19 
+ bl[17] br[17] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_20 
+ bl[18] br[18] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_21 
+ bl[19] br[19] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_22 
+ bl[20] br[20] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_23 
+ bl[21] br[21] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_24 
+ bl[22] br[22] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_25 
+ bl[23] br[23] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_26 
+ bl[24] br[24] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_27 
+ bl[25] br[25] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_28 
+ bl[26] br[26] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_29 
+ bl[27] br[27] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_30 
+ bl[28] br[28] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_31 
+ bl[29] br[29] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_32 
+ bl[30] br[30] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_33 
+ bl[31] br[31] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_34 
+ bl[32] br[32] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_35 
+ bl[33] br[33] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_36 
+ bl[34] br[34] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_37 
+ bl[35] br[35] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_38 
+ bl[36] br[36] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_39 
+ bl[37] br[37] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_40 
+ bl[38] br[38] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_41 
+ bl[39] br[39] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_42 
+ bl[40] br[40] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_43 
+ bl[41] br[41] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_44 
+ bl[42] br[42] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_45 
+ bl[43] br[43] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_46 
+ bl[44] br[44] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_47 
+ bl[45] br[45] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_48 
+ bl[46] br[46] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_49 
+ bl[47] br[47] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_50 
+ bl[48] br[48] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_51 
+ bl[49] br[49] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_52 
+ bl[50] br[50] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_53 
+ bl[51] br[51] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_54 
+ bl[52] br[52] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_55 
+ bl[53] br[53] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_56 
+ bl[54] br[54] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_57 
+ bl[55] br[55] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_58 
+ bl[56] br[56] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_59 
+ bl[57] br[57] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_60 
+ bl[58] br[58] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_61 
+ bl[59] br[59] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_62 
+ bl[60] br[60] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_63 
+ bl[61] br[61] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_64 
+ bl[62] br[62] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_65 
+ bl[63] br[63] vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_66 
+ vdd vdd vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_348_67 
+ vdd vdd vdd vss wl[346] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_0 
+ vdd vdd vss vdd vpb vnb wl[347] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_349_1 
+ rbl rbr vss vdd vpb vnb wl[347] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_349_2 
+ bl[0] br[0] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_3 
+ bl[1] br[1] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_4 
+ bl[2] br[2] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_5 
+ bl[3] br[3] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_6 
+ bl[4] br[4] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_7 
+ bl[5] br[5] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_8 
+ bl[6] br[6] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_9 
+ bl[7] br[7] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_10 
+ bl[8] br[8] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_11 
+ bl[9] br[9] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_12 
+ bl[10] br[10] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_13 
+ bl[11] br[11] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_14 
+ bl[12] br[12] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_15 
+ bl[13] br[13] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_16 
+ bl[14] br[14] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_17 
+ bl[15] br[15] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_18 
+ bl[16] br[16] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_19 
+ bl[17] br[17] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_20 
+ bl[18] br[18] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_21 
+ bl[19] br[19] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_22 
+ bl[20] br[20] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_23 
+ bl[21] br[21] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_24 
+ bl[22] br[22] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_25 
+ bl[23] br[23] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_26 
+ bl[24] br[24] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_27 
+ bl[25] br[25] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_28 
+ bl[26] br[26] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_29 
+ bl[27] br[27] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_30 
+ bl[28] br[28] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_31 
+ bl[29] br[29] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_32 
+ bl[30] br[30] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_33 
+ bl[31] br[31] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_34 
+ bl[32] br[32] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_35 
+ bl[33] br[33] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_36 
+ bl[34] br[34] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_37 
+ bl[35] br[35] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_38 
+ bl[36] br[36] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_39 
+ bl[37] br[37] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_40 
+ bl[38] br[38] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_41 
+ bl[39] br[39] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_42 
+ bl[40] br[40] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_43 
+ bl[41] br[41] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_44 
+ bl[42] br[42] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_45 
+ bl[43] br[43] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_46 
+ bl[44] br[44] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_47 
+ bl[45] br[45] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_48 
+ bl[46] br[46] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_49 
+ bl[47] br[47] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_50 
+ bl[48] br[48] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_51 
+ bl[49] br[49] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_52 
+ bl[50] br[50] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_53 
+ bl[51] br[51] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_54 
+ bl[52] br[52] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_55 
+ bl[53] br[53] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_56 
+ bl[54] br[54] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_57 
+ bl[55] br[55] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_58 
+ bl[56] br[56] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_59 
+ bl[57] br[57] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_60 
+ bl[58] br[58] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_61 
+ bl[59] br[59] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_62 
+ bl[60] br[60] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_63 
+ bl[61] br[61] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_64 
+ bl[62] br[62] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_65 
+ bl[63] br[63] vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_66 
+ vdd vdd vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_349_67 
+ vdd vdd vdd vss wl[347] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_0 
+ vdd vdd vss vdd vpb vnb wl[348] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_350_1 
+ rbl rbr vss vdd vpb vnb wl[348] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_350_2 
+ bl[0] br[0] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_3 
+ bl[1] br[1] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_4 
+ bl[2] br[2] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_5 
+ bl[3] br[3] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_6 
+ bl[4] br[4] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_7 
+ bl[5] br[5] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_8 
+ bl[6] br[6] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_9 
+ bl[7] br[7] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_10 
+ bl[8] br[8] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_11 
+ bl[9] br[9] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_12 
+ bl[10] br[10] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_13 
+ bl[11] br[11] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_14 
+ bl[12] br[12] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_15 
+ bl[13] br[13] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_16 
+ bl[14] br[14] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_17 
+ bl[15] br[15] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_18 
+ bl[16] br[16] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_19 
+ bl[17] br[17] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_20 
+ bl[18] br[18] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_21 
+ bl[19] br[19] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_22 
+ bl[20] br[20] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_23 
+ bl[21] br[21] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_24 
+ bl[22] br[22] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_25 
+ bl[23] br[23] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_26 
+ bl[24] br[24] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_27 
+ bl[25] br[25] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_28 
+ bl[26] br[26] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_29 
+ bl[27] br[27] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_30 
+ bl[28] br[28] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_31 
+ bl[29] br[29] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_32 
+ bl[30] br[30] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_33 
+ bl[31] br[31] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_34 
+ bl[32] br[32] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_35 
+ bl[33] br[33] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_36 
+ bl[34] br[34] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_37 
+ bl[35] br[35] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_38 
+ bl[36] br[36] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_39 
+ bl[37] br[37] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_40 
+ bl[38] br[38] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_41 
+ bl[39] br[39] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_42 
+ bl[40] br[40] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_43 
+ bl[41] br[41] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_44 
+ bl[42] br[42] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_45 
+ bl[43] br[43] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_46 
+ bl[44] br[44] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_47 
+ bl[45] br[45] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_48 
+ bl[46] br[46] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_49 
+ bl[47] br[47] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_50 
+ bl[48] br[48] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_51 
+ bl[49] br[49] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_52 
+ bl[50] br[50] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_53 
+ bl[51] br[51] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_54 
+ bl[52] br[52] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_55 
+ bl[53] br[53] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_56 
+ bl[54] br[54] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_57 
+ bl[55] br[55] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_58 
+ bl[56] br[56] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_59 
+ bl[57] br[57] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_60 
+ bl[58] br[58] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_61 
+ bl[59] br[59] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_62 
+ bl[60] br[60] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_63 
+ bl[61] br[61] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_64 
+ bl[62] br[62] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_65 
+ bl[63] br[63] vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_66 
+ vdd vdd vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_350_67 
+ vdd vdd vdd vss wl[348] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_0 
+ vdd vdd vss vdd vpb vnb wl[349] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_351_1 
+ rbl rbr vss vdd vpb vnb wl[349] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_351_2 
+ bl[0] br[0] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_3 
+ bl[1] br[1] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_4 
+ bl[2] br[2] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_5 
+ bl[3] br[3] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_6 
+ bl[4] br[4] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_7 
+ bl[5] br[5] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_8 
+ bl[6] br[6] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_9 
+ bl[7] br[7] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_10 
+ bl[8] br[8] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_11 
+ bl[9] br[9] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_12 
+ bl[10] br[10] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_13 
+ bl[11] br[11] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_14 
+ bl[12] br[12] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_15 
+ bl[13] br[13] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_16 
+ bl[14] br[14] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_17 
+ bl[15] br[15] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_18 
+ bl[16] br[16] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_19 
+ bl[17] br[17] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_20 
+ bl[18] br[18] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_21 
+ bl[19] br[19] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_22 
+ bl[20] br[20] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_23 
+ bl[21] br[21] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_24 
+ bl[22] br[22] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_25 
+ bl[23] br[23] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_26 
+ bl[24] br[24] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_27 
+ bl[25] br[25] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_28 
+ bl[26] br[26] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_29 
+ bl[27] br[27] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_30 
+ bl[28] br[28] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_31 
+ bl[29] br[29] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_32 
+ bl[30] br[30] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_33 
+ bl[31] br[31] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_34 
+ bl[32] br[32] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_35 
+ bl[33] br[33] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_36 
+ bl[34] br[34] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_37 
+ bl[35] br[35] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_38 
+ bl[36] br[36] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_39 
+ bl[37] br[37] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_40 
+ bl[38] br[38] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_41 
+ bl[39] br[39] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_42 
+ bl[40] br[40] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_43 
+ bl[41] br[41] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_44 
+ bl[42] br[42] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_45 
+ bl[43] br[43] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_46 
+ bl[44] br[44] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_47 
+ bl[45] br[45] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_48 
+ bl[46] br[46] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_49 
+ bl[47] br[47] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_50 
+ bl[48] br[48] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_51 
+ bl[49] br[49] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_52 
+ bl[50] br[50] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_53 
+ bl[51] br[51] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_54 
+ bl[52] br[52] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_55 
+ bl[53] br[53] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_56 
+ bl[54] br[54] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_57 
+ bl[55] br[55] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_58 
+ bl[56] br[56] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_59 
+ bl[57] br[57] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_60 
+ bl[58] br[58] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_61 
+ bl[59] br[59] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_62 
+ bl[60] br[60] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_63 
+ bl[61] br[61] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_64 
+ bl[62] br[62] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_65 
+ bl[63] br[63] vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_66 
+ vdd vdd vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_351_67 
+ vdd vdd vdd vss wl[349] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_0 
+ vdd vdd vss vdd vpb vnb wl[350] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_352_1 
+ rbl rbr vss vdd vpb vnb wl[350] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_352_2 
+ bl[0] br[0] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_3 
+ bl[1] br[1] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_4 
+ bl[2] br[2] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_5 
+ bl[3] br[3] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_6 
+ bl[4] br[4] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_7 
+ bl[5] br[5] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_8 
+ bl[6] br[6] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_9 
+ bl[7] br[7] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_10 
+ bl[8] br[8] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_11 
+ bl[9] br[9] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_12 
+ bl[10] br[10] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_13 
+ bl[11] br[11] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_14 
+ bl[12] br[12] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_15 
+ bl[13] br[13] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_16 
+ bl[14] br[14] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_17 
+ bl[15] br[15] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_18 
+ bl[16] br[16] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_19 
+ bl[17] br[17] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_20 
+ bl[18] br[18] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_21 
+ bl[19] br[19] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_22 
+ bl[20] br[20] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_23 
+ bl[21] br[21] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_24 
+ bl[22] br[22] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_25 
+ bl[23] br[23] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_26 
+ bl[24] br[24] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_27 
+ bl[25] br[25] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_28 
+ bl[26] br[26] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_29 
+ bl[27] br[27] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_30 
+ bl[28] br[28] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_31 
+ bl[29] br[29] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_32 
+ bl[30] br[30] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_33 
+ bl[31] br[31] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_34 
+ bl[32] br[32] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_35 
+ bl[33] br[33] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_36 
+ bl[34] br[34] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_37 
+ bl[35] br[35] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_38 
+ bl[36] br[36] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_39 
+ bl[37] br[37] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_40 
+ bl[38] br[38] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_41 
+ bl[39] br[39] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_42 
+ bl[40] br[40] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_43 
+ bl[41] br[41] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_44 
+ bl[42] br[42] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_45 
+ bl[43] br[43] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_46 
+ bl[44] br[44] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_47 
+ bl[45] br[45] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_48 
+ bl[46] br[46] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_49 
+ bl[47] br[47] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_50 
+ bl[48] br[48] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_51 
+ bl[49] br[49] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_52 
+ bl[50] br[50] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_53 
+ bl[51] br[51] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_54 
+ bl[52] br[52] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_55 
+ bl[53] br[53] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_56 
+ bl[54] br[54] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_57 
+ bl[55] br[55] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_58 
+ bl[56] br[56] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_59 
+ bl[57] br[57] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_60 
+ bl[58] br[58] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_61 
+ bl[59] br[59] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_62 
+ bl[60] br[60] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_63 
+ bl[61] br[61] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_64 
+ bl[62] br[62] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_65 
+ bl[63] br[63] vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_66 
+ vdd vdd vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_352_67 
+ vdd vdd vdd vss wl[350] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_0 
+ vdd vdd vss vdd vpb vnb wl[351] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_353_1 
+ rbl rbr vss vdd vpb vnb wl[351] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_353_2 
+ bl[0] br[0] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_3 
+ bl[1] br[1] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_4 
+ bl[2] br[2] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_5 
+ bl[3] br[3] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_6 
+ bl[4] br[4] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_7 
+ bl[5] br[5] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_8 
+ bl[6] br[6] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_9 
+ bl[7] br[7] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_10 
+ bl[8] br[8] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_11 
+ bl[9] br[9] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_12 
+ bl[10] br[10] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_13 
+ bl[11] br[11] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_14 
+ bl[12] br[12] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_15 
+ bl[13] br[13] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_16 
+ bl[14] br[14] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_17 
+ bl[15] br[15] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_18 
+ bl[16] br[16] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_19 
+ bl[17] br[17] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_20 
+ bl[18] br[18] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_21 
+ bl[19] br[19] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_22 
+ bl[20] br[20] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_23 
+ bl[21] br[21] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_24 
+ bl[22] br[22] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_25 
+ bl[23] br[23] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_26 
+ bl[24] br[24] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_27 
+ bl[25] br[25] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_28 
+ bl[26] br[26] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_29 
+ bl[27] br[27] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_30 
+ bl[28] br[28] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_31 
+ bl[29] br[29] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_32 
+ bl[30] br[30] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_33 
+ bl[31] br[31] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_34 
+ bl[32] br[32] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_35 
+ bl[33] br[33] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_36 
+ bl[34] br[34] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_37 
+ bl[35] br[35] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_38 
+ bl[36] br[36] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_39 
+ bl[37] br[37] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_40 
+ bl[38] br[38] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_41 
+ bl[39] br[39] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_42 
+ bl[40] br[40] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_43 
+ bl[41] br[41] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_44 
+ bl[42] br[42] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_45 
+ bl[43] br[43] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_46 
+ bl[44] br[44] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_47 
+ bl[45] br[45] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_48 
+ bl[46] br[46] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_49 
+ bl[47] br[47] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_50 
+ bl[48] br[48] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_51 
+ bl[49] br[49] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_52 
+ bl[50] br[50] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_53 
+ bl[51] br[51] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_54 
+ bl[52] br[52] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_55 
+ bl[53] br[53] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_56 
+ bl[54] br[54] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_57 
+ bl[55] br[55] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_58 
+ bl[56] br[56] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_59 
+ bl[57] br[57] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_60 
+ bl[58] br[58] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_61 
+ bl[59] br[59] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_62 
+ bl[60] br[60] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_63 
+ bl[61] br[61] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_64 
+ bl[62] br[62] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_65 
+ bl[63] br[63] vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_66 
+ vdd vdd vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_353_67 
+ vdd vdd vdd vss wl[351] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_0 
+ vdd vdd vss vdd vpb vnb wl[352] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_354_1 
+ rbl rbr vss vdd vpb vnb wl[352] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_354_2 
+ bl[0] br[0] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_3 
+ bl[1] br[1] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_4 
+ bl[2] br[2] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_5 
+ bl[3] br[3] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_6 
+ bl[4] br[4] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_7 
+ bl[5] br[5] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_8 
+ bl[6] br[6] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_9 
+ bl[7] br[7] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_10 
+ bl[8] br[8] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_11 
+ bl[9] br[9] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_12 
+ bl[10] br[10] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_13 
+ bl[11] br[11] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_14 
+ bl[12] br[12] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_15 
+ bl[13] br[13] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_16 
+ bl[14] br[14] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_17 
+ bl[15] br[15] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_18 
+ bl[16] br[16] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_19 
+ bl[17] br[17] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_20 
+ bl[18] br[18] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_21 
+ bl[19] br[19] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_22 
+ bl[20] br[20] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_23 
+ bl[21] br[21] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_24 
+ bl[22] br[22] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_25 
+ bl[23] br[23] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_26 
+ bl[24] br[24] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_27 
+ bl[25] br[25] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_28 
+ bl[26] br[26] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_29 
+ bl[27] br[27] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_30 
+ bl[28] br[28] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_31 
+ bl[29] br[29] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_32 
+ bl[30] br[30] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_33 
+ bl[31] br[31] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_34 
+ bl[32] br[32] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_35 
+ bl[33] br[33] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_36 
+ bl[34] br[34] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_37 
+ bl[35] br[35] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_38 
+ bl[36] br[36] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_39 
+ bl[37] br[37] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_40 
+ bl[38] br[38] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_41 
+ bl[39] br[39] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_42 
+ bl[40] br[40] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_43 
+ bl[41] br[41] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_44 
+ bl[42] br[42] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_45 
+ bl[43] br[43] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_46 
+ bl[44] br[44] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_47 
+ bl[45] br[45] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_48 
+ bl[46] br[46] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_49 
+ bl[47] br[47] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_50 
+ bl[48] br[48] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_51 
+ bl[49] br[49] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_52 
+ bl[50] br[50] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_53 
+ bl[51] br[51] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_54 
+ bl[52] br[52] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_55 
+ bl[53] br[53] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_56 
+ bl[54] br[54] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_57 
+ bl[55] br[55] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_58 
+ bl[56] br[56] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_59 
+ bl[57] br[57] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_60 
+ bl[58] br[58] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_61 
+ bl[59] br[59] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_62 
+ bl[60] br[60] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_63 
+ bl[61] br[61] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_64 
+ bl[62] br[62] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_65 
+ bl[63] br[63] vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_66 
+ vdd vdd vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_354_67 
+ vdd vdd vdd vss wl[352] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_0 
+ vdd vdd vss vdd vpb vnb wl[353] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_355_1 
+ rbl rbr vss vdd vpb vnb wl[353] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_355_2 
+ bl[0] br[0] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_3 
+ bl[1] br[1] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_4 
+ bl[2] br[2] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_5 
+ bl[3] br[3] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_6 
+ bl[4] br[4] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_7 
+ bl[5] br[5] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_8 
+ bl[6] br[6] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_9 
+ bl[7] br[7] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_10 
+ bl[8] br[8] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_11 
+ bl[9] br[9] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_12 
+ bl[10] br[10] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_13 
+ bl[11] br[11] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_14 
+ bl[12] br[12] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_15 
+ bl[13] br[13] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_16 
+ bl[14] br[14] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_17 
+ bl[15] br[15] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_18 
+ bl[16] br[16] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_19 
+ bl[17] br[17] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_20 
+ bl[18] br[18] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_21 
+ bl[19] br[19] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_22 
+ bl[20] br[20] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_23 
+ bl[21] br[21] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_24 
+ bl[22] br[22] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_25 
+ bl[23] br[23] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_26 
+ bl[24] br[24] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_27 
+ bl[25] br[25] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_28 
+ bl[26] br[26] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_29 
+ bl[27] br[27] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_30 
+ bl[28] br[28] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_31 
+ bl[29] br[29] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_32 
+ bl[30] br[30] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_33 
+ bl[31] br[31] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_34 
+ bl[32] br[32] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_35 
+ bl[33] br[33] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_36 
+ bl[34] br[34] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_37 
+ bl[35] br[35] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_38 
+ bl[36] br[36] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_39 
+ bl[37] br[37] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_40 
+ bl[38] br[38] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_41 
+ bl[39] br[39] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_42 
+ bl[40] br[40] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_43 
+ bl[41] br[41] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_44 
+ bl[42] br[42] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_45 
+ bl[43] br[43] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_46 
+ bl[44] br[44] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_47 
+ bl[45] br[45] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_48 
+ bl[46] br[46] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_49 
+ bl[47] br[47] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_50 
+ bl[48] br[48] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_51 
+ bl[49] br[49] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_52 
+ bl[50] br[50] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_53 
+ bl[51] br[51] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_54 
+ bl[52] br[52] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_55 
+ bl[53] br[53] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_56 
+ bl[54] br[54] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_57 
+ bl[55] br[55] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_58 
+ bl[56] br[56] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_59 
+ bl[57] br[57] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_60 
+ bl[58] br[58] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_61 
+ bl[59] br[59] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_62 
+ bl[60] br[60] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_63 
+ bl[61] br[61] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_64 
+ bl[62] br[62] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_65 
+ bl[63] br[63] vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_66 
+ vdd vdd vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_355_67 
+ vdd vdd vdd vss wl[353] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_0 
+ vdd vdd vss vdd vpb vnb wl[354] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_356_1 
+ rbl rbr vss vdd vpb vnb wl[354] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_356_2 
+ bl[0] br[0] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_3 
+ bl[1] br[1] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_4 
+ bl[2] br[2] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_5 
+ bl[3] br[3] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_6 
+ bl[4] br[4] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_7 
+ bl[5] br[5] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_8 
+ bl[6] br[6] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_9 
+ bl[7] br[7] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_10 
+ bl[8] br[8] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_11 
+ bl[9] br[9] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_12 
+ bl[10] br[10] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_13 
+ bl[11] br[11] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_14 
+ bl[12] br[12] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_15 
+ bl[13] br[13] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_16 
+ bl[14] br[14] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_17 
+ bl[15] br[15] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_18 
+ bl[16] br[16] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_19 
+ bl[17] br[17] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_20 
+ bl[18] br[18] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_21 
+ bl[19] br[19] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_22 
+ bl[20] br[20] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_23 
+ bl[21] br[21] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_24 
+ bl[22] br[22] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_25 
+ bl[23] br[23] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_26 
+ bl[24] br[24] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_27 
+ bl[25] br[25] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_28 
+ bl[26] br[26] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_29 
+ bl[27] br[27] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_30 
+ bl[28] br[28] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_31 
+ bl[29] br[29] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_32 
+ bl[30] br[30] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_33 
+ bl[31] br[31] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_34 
+ bl[32] br[32] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_35 
+ bl[33] br[33] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_36 
+ bl[34] br[34] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_37 
+ bl[35] br[35] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_38 
+ bl[36] br[36] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_39 
+ bl[37] br[37] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_40 
+ bl[38] br[38] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_41 
+ bl[39] br[39] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_42 
+ bl[40] br[40] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_43 
+ bl[41] br[41] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_44 
+ bl[42] br[42] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_45 
+ bl[43] br[43] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_46 
+ bl[44] br[44] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_47 
+ bl[45] br[45] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_48 
+ bl[46] br[46] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_49 
+ bl[47] br[47] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_50 
+ bl[48] br[48] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_51 
+ bl[49] br[49] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_52 
+ bl[50] br[50] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_53 
+ bl[51] br[51] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_54 
+ bl[52] br[52] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_55 
+ bl[53] br[53] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_56 
+ bl[54] br[54] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_57 
+ bl[55] br[55] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_58 
+ bl[56] br[56] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_59 
+ bl[57] br[57] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_60 
+ bl[58] br[58] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_61 
+ bl[59] br[59] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_62 
+ bl[60] br[60] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_63 
+ bl[61] br[61] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_64 
+ bl[62] br[62] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_65 
+ bl[63] br[63] vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_66 
+ vdd vdd vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_356_67 
+ vdd vdd vdd vss wl[354] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_0 
+ vdd vdd vss vdd vpb vnb wl[355] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_357_1 
+ rbl rbr vss vdd vpb vnb wl[355] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_357_2 
+ bl[0] br[0] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_3 
+ bl[1] br[1] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_4 
+ bl[2] br[2] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_5 
+ bl[3] br[3] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_6 
+ bl[4] br[4] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_7 
+ bl[5] br[5] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_8 
+ bl[6] br[6] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_9 
+ bl[7] br[7] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_10 
+ bl[8] br[8] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_11 
+ bl[9] br[9] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_12 
+ bl[10] br[10] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_13 
+ bl[11] br[11] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_14 
+ bl[12] br[12] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_15 
+ bl[13] br[13] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_16 
+ bl[14] br[14] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_17 
+ bl[15] br[15] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_18 
+ bl[16] br[16] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_19 
+ bl[17] br[17] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_20 
+ bl[18] br[18] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_21 
+ bl[19] br[19] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_22 
+ bl[20] br[20] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_23 
+ bl[21] br[21] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_24 
+ bl[22] br[22] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_25 
+ bl[23] br[23] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_26 
+ bl[24] br[24] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_27 
+ bl[25] br[25] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_28 
+ bl[26] br[26] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_29 
+ bl[27] br[27] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_30 
+ bl[28] br[28] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_31 
+ bl[29] br[29] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_32 
+ bl[30] br[30] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_33 
+ bl[31] br[31] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_34 
+ bl[32] br[32] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_35 
+ bl[33] br[33] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_36 
+ bl[34] br[34] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_37 
+ bl[35] br[35] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_38 
+ bl[36] br[36] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_39 
+ bl[37] br[37] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_40 
+ bl[38] br[38] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_41 
+ bl[39] br[39] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_42 
+ bl[40] br[40] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_43 
+ bl[41] br[41] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_44 
+ bl[42] br[42] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_45 
+ bl[43] br[43] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_46 
+ bl[44] br[44] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_47 
+ bl[45] br[45] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_48 
+ bl[46] br[46] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_49 
+ bl[47] br[47] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_50 
+ bl[48] br[48] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_51 
+ bl[49] br[49] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_52 
+ bl[50] br[50] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_53 
+ bl[51] br[51] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_54 
+ bl[52] br[52] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_55 
+ bl[53] br[53] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_56 
+ bl[54] br[54] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_57 
+ bl[55] br[55] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_58 
+ bl[56] br[56] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_59 
+ bl[57] br[57] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_60 
+ bl[58] br[58] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_61 
+ bl[59] br[59] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_62 
+ bl[60] br[60] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_63 
+ bl[61] br[61] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_64 
+ bl[62] br[62] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_65 
+ bl[63] br[63] vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_66 
+ vdd vdd vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_357_67 
+ vdd vdd vdd vss wl[355] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_0 
+ vdd vdd vss vdd vpb vnb wl[356] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_358_1 
+ rbl rbr vss vdd vpb vnb wl[356] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_358_2 
+ bl[0] br[0] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_3 
+ bl[1] br[1] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_4 
+ bl[2] br[2] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_5 
+ bl[3] br[3] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_6 
+ bl[4] br[4] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_7 
+ bl[5] br[5] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_8 
+ bl[6] br[6] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_9 
+ bl[7] br[7] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_10 
+ bl[8] br[8] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_11 
+ bl[9] br[9] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_12 
+ bl[10] br[10] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_13 
+ bl[11] br[11] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_14 
+ bl[12] br[12] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_15 
+ bl[13] br[13] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_16 
+ bl[14] br[14] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_17 
+ bl[15] br[15] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_18 
+ bl[16] br[16] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_19 
+ bl[17] br[17] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_20 
+ bl[18] br[18] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_21 
+ bl[19] br[19] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_22 
+ bl[20] br[20] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_23 
+ bl[21] br[21] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_24 
+ bl[22] br[22] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_25 
+ bl[23] br[23] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_26 
+ bl[24] br[24] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_27 
+ bl[25] br[25] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_28 
+ bl[26] br[26] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_29 
+ bl[27] br[27] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_30 
+ bl[28] br[28] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_31 
+ bl[29] br[29] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_32 
+ bl[30] br[30] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_33 
+ bl[31] br[31] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_34 
+ bl[32] br[32] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_35 
+ bl[33] br[33] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_36 
+ bl[34] br[34] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_37 
+ bl[35] br[35] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_38 
+ bl[36] br[36] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_39 
+ bl[37] br[37] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_40 
+ bl[38] br[38] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_41 
+ bl[39] br[39] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_42 
+ bl[40] br[40] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_43 
+ bl[41] br[41] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_44 
+ bl[42] br[42] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_45 
+ bl[43] br[43] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_46 
+ bl[44] br[44] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_47 
+ bl[45] br[45] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_48 
+ bl[46] br[46] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_49 
+ bl[47] br[47] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_50 
+ bl[48] br[48] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_51 
+ bl[49] br[49] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_52 
+ bl[50] br[50] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_53 
+ bl[51] br[51] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_54 
+ bl[52] br[52] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_55 
+ bl[53] br[53] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_56 
+ bl[54] br[54] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_57 
+ bl[55] br[55] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_58 
+ bl[56] br[56] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_59 
+ bl[57] br[57] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_60 
+ bl[58] br[58] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_61 
+ bl[59] br[59] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_62 
+ bl[60] br[60] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_63 
+ bl[61] br[61] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_64 
+ bl[62] br[62] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_65 
+ bl[63] br[63] vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_66 
+ vdd vdd vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_358_67 
+ vdd vdd vdd vss wl[356] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_0 
+ vdd vdd vss vdd vpb vnb wl[357] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_359_1 
+ rbl rbr vss vdd vpb vnb wl[357] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_359_2 
+ bl[0] br[0] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_3 
+ bl[1] br[1] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_4 
+ bl[2] br[2] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_5 
+ bl[3] br[3] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_6 
+ bl[4] br[4] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_7 
+ bl[5] br[5] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_8 
+ bl[6] br[6] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_9 
+ bl[7] br[7] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_10 
+ bl[8] br[8] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_11 
+ bl[9] br[9] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_12 
+ bl[10] br[10] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_13 
+ bl[11] br[11] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_14 
+ bl[12] br[12] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_15 
+ bl[13] br[13] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_16 
+ bl[14] br[14] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_17 
+ bl[15] br[15] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_18 
+ bl[16] br[16] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_19 
+ bl[17] br[17] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_20 
+ bl[18] br[18] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_21 
+ bl[19] br[19] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_22 
+ bl[20] br[20] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_23 
+ bl[21] br[21] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_24 
+ bl[22] br[22] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_25 
+ bl[23] br[23] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_26 
+ bl[24] br[24] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_27 
+ bl[25] br[25] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_28 
+ bl[26] br[26] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_29 
+ bl[27] br[27] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_30 
+ bl[28] br[28] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_31 
+ bl[29] br[29] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_32 
+ bl[30] br[30] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_33 
+ bl[31] br[31] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_34 
+ bl[32] br[32] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_35 
+ bl[33] br[33] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_36 
+ bl[34] br[34] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_37 
+ bl[35] br[35] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_38 
+ bl[36] br[36] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_39 
+ bl[37] br[37] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_40 
+ bl[38] br[38] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_41 
+ bl[39] br[39] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_42 
+ bl[40] br[40] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_43 
+ bl[41] br[41] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_44 
+ bl[42] br[42] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_45 
+ bl[43] br[43] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_46 
+ bl[44] br[44] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_47 
+ bl[45] br[45] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_48 
+ bl[46] br[46] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_49 
+ bl[47] br[47] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_50 
+ bl[48] br[48] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_51 
+ bl[49] br[49] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_52 
+ bl[50] br[50] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_53 
+ bl[51] br[51] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_54 
+ bl[52] br[52] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_55 
+ bl[53] br[53] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_56 
+ bl[54] br[54] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_57 
+ bl[55] br[55] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_58 
+ bl[56] br[56] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_59 
+ bl[57] br[57] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_60 
+ bl[58] br[58] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_61 
+ bl[59] br[59] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_62 
+ bl[60] br[60] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_63 
+ bl[61] br[61] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_64 
+ bl[62] br[62] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_65 
+ bl[63] br[63] vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_66 
+ vdd vdd vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_359_67 
+ vdd vdd vdd vss wl[357] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_0 
+ vdd vdd vss vdd vpb vnb wl[358] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_360_1 
+ rbl rbr vss vdd vpb vnb wl[358] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_360_2 
+ bl[0] br[0] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_3 
+ bl[1] br[1] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_4 
+ bl[2] br[2] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_5 
+ bl[3] br[3] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_6 
+ bl[4] br[4] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_7 
+ bl[5] br[5] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_8 
+ bl[6] br[6] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_9 
+ bl[7] br[7] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_10 
+ bl[8] br[8] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_11 
+ bl[9] br[9] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_12 
+ bl[10] br[10] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_13 
+ bl[11] br[11] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_14 
+ bl[12] br[12] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_15 
+ bl[13] br[13] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_16 
+ bl[14] br[14] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_17 
+ bl[15] br[15] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_18 
+ bl[16] br[16] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_19 
+ bl[17] br[17] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_20 
+ bl[18] br[18] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_21 
+ bl[19] br[19] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_22 
+ bl[20] br[20] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_23 
+ bl[21] br[21] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_24 
+ bl[22] br[22] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_25 
+ bl[23] br[23] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_26 
+ bl[24] br[24] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_27 
+ bl[25] br[25] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_28 
+ bl[26] br[26] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_29 
+ bl[27] br[27] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_30 
+ bl[28] br[28] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_31 
+ bl[29] br[29] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_32 
+ bl[30] br[30] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_33 
+ bl[31] br[31] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_34 
+ bl[32] br[32] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_35 
+ bl[33] br[33] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_36 
+ bl[34] br[34] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_37 
+ bl[35] br[35] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_38 
+ bl[36] br[36] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_39 
+ bl[37] br[37] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_40 
+ bl[38] br[38] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_41 
+ bl[39] br[39] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_42 
+ bl[40] br[40] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_43 
+ bl[41] br[41] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_44 
+ bl[42] br[42] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_45 
+ bl[43] br[43] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_46 
+ bl[44] br[44] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_47 
+ bl[45] br[45] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_48 
+ bl[46] br[46] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_49 
+ bl[47] br[47] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_50 
+ bl[48] br[48] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_51 
+ bl[49] br[49] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_52 
+ bl[50] br[50] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_53 
+ bl[51] br[51] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_54 
+ bl[52] br[52] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_55 
+ bl[53] br[53] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_56 
+ bl[54] br[54] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_57 
+ bl[55] br[55] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_58 
+ bl[56] br[56] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_59 
+ bl[57] br[57] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_60 
+ bl[58] br[58] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_61 
+ bl[59] br[59] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_62 
+ bl[60] br[60] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_63 
+ bl[61] br[61] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_64 
+ bl[62] br[62] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_65 
+ bl[63] br[63] vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_66 
+ vdd vdd vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_360_67 
+ vdd vdd vdd vss wl[358] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_0 
+ vdd vdd vss vdd vpb vnb wl[359] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_361_1 
+ rbl rbr vss vdd vpb vnb wl[359] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_361_2 
+ bl[0] br[0] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_3 
+ bl[1] br[1] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_4 
+ bl[2] br[2] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_5 
+ bl[3] br[3] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_6 
+ bl[4] br[4] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_7 
+ bl[5] br[5] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_8 
+ bl[6] br[6] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_9 
+ bl[7] br[7] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_10 
+ bl[8] br[8] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_11 
+ bl[9] br[9] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_12 
+ bl[10] br[10] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_13 
+ bl[11] br[11] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_14 
+ bl[12] br[12] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_15 
+ bl[13] br[13] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_16 
+ bl[14] br[14] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_17 
+ bl[15] br[15] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_18 
+ bl[16] br[16] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_19 
+ bl[17] br[17] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_20 
+ bl[18] br[18] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_21 
+ bl[19] br[19] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_22 
+ bl[20] br[20] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_23 
+ bl[21] br[21] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_24 
+ bl[22] br[22] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_25 
+ bl[23] br[23] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_26 
+ bl[24] br[24] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_27 
+ bl[25] br[25] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_28 
+ bl[26] br[26] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_29 
+ bl[27] br[27] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_30 
+ bl[28] br[28] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_31 
+ bl[29] br[29] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_32 
+ bl[30] br[30] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_33 
+ bl[31] br[31] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_34 
+ bl[32] br[32] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_35 
+ bl[33] br[33] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_36 
+ bl[34] br[34] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_37 
+ bl[35] br[35] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_38 
+ bl[36] br[36] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_39 
+ bl[37] br[37] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_40 
+ bl[38] br[38] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_41 
+ bl[39] br[39] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_42 
+ bl[40] br[40] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_43 
+ bl[41] br[41] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_44 
+ bl[42] br[42] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_45 
+ bl[43] br[43] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_46 
+ bl[44] br[44] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_47 
+ bl[45] br[45] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_48 
+ bl[46] br[46] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_49 
+ bl[47] br[47] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_50 
+ bl[48] br[48] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_51 
+ bl[49] br[49] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_52 
+ bl[50] br[50] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_53 
+ bl[51] br[51] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_54 
+ bl[52] br[52] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_55 
+ bl[53] br[53] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_56 
+ bl[54] br[54] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_57 
+ bl[55] br[55] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_58 
+ bl[56] br[56] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_59 
+ bl[57] br[57] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_60 
+ bl[58] br[58] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_61 
+ bl[59] br[59] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_62 
+ bl[60] br[60] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_63 
+ bl[61] br[61] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_64 
+ bl[62] br[62] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_65 
+ bl[63] br[63] vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_66 
+ vdd vdd vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_361_67 
+ vdd vdd vdd vss wl[359] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_0 
+ vdd vdd vss vdd vpb vnb wl[360] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_362_1 
+ rbl rbr vss vdd vpb vnb wl[360] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_362_2 
+ bl[0] br[0] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_3 
+ bl[1] br[1] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_4 
+ bl[2] br[2] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_5 
+ bl[3] br[3] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_6 
+ bl[4] br[4] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_7 
+ bl[5] br[5] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_8 
+ bl[6] br[6] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_9 
+ bl[7] br[7] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_10 
+ bl[8] br[8] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_11 
+ bl[9] br[9] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_12 
+ bl[10] br[10] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_13 
+ bl[11] br[11] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_14 
+ bl[12] br[12] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_15 
+ bl[13] br[13] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_16 
+ bl[14] br[14] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_17 
+ bl[15] br[15] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_18 
+ bl[16] br[16] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_19 
+ bl[17] br[17] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_20 
+ bl[18] br[18] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_21 
+ bl[19] br[19] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_22 
+ bl[20] br[20] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_23 
+ bl[21] br[21] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_24 
+ bl[22] br[22] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_25 
+ bl[23] br[23] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_26 
+ bl[24] br[24] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_27 
+ bl[25] br[25] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_28 
+ bl[26] br[26] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_29 
+ bl[27] br[27] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_30 
+ bl[28] br[28] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_31 
+ bl[29] br[29] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_32 
+ bl[30] br[30] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_33 
+ bl[31] br[31] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_34 
+ bl[32] br[32] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_35 
+ bl[33] br[33] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_36 
+ bl[34] br[34] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_37 
+ bl[35] br[35] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_38 
+ bl[36] br[36] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_39 
+ bl[37] br[37] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_40 
+ bl[38] br[38] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_41 
+ bl[39] br[39] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_42 
+ bl[40] br[40] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_43 
+ bl[41] br[41] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_44 
+ bl[42] br[42] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_45 
+ bl[43] br[43] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_46 
+ bl[44] br[44] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_47 
+ bl[45] br[45] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_48 
+ bl[46] br[46] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_49 
+ bl[47] br[47] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_50 
+ bl[48] br[48] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_51 
+ bl[49] br[49] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_52 
+ bl[50] br[50] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_53 
+ bl[51] br[51] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_54 
+ bl[52] br[52] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_55 
+ bl[53] br[53] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_56 
+ bl[54] br[54] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_57 
+ bl[55] br[55] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_58 
+ bl[56] br[56] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_59 
+ bl[57] br[57] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_60 
+ bl[58] br[58] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_61 
+ bl[59] br[59] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_62 
+ bl[60] br[60] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_63 
+ bl[61] br[61] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_64 
+ bl[62] br[62] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_65 
+ bl[63] br[63] vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_66 
+ vdd vdd vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_362_67 
+ vdd vdd vdd vss wl[360] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_0 
+ vdd vdd vss vdd vpb vnb wl[361] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_363_1 
+ rbl rbr vss vdd vpb vnb wl[361] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_363_2 
+ bl[0] br[0] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_3 
+ bl[1] br[1] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_4 
+ bl[2] br[2] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_5 
+ bl[3] br[3] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_6 
+ bl[4] br[4] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_7 
+ bl[5] br[5] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_8 
+ bl[6] br[6] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_9 
+ bl[7] br[7] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_10 
+ bl[8] br[8] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_11 
+ bl[9] br[9] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_12 
+ bl[10] br[10] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_13 
+ bl[11] br[11] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_14 
+ bl[12] br[12] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_15 
+ bl[13] br[13] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_16 
+ bl[14] br[14] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_17 
+ bl[15] br[15] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_18 
+ bl[16] br[16] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_19 
+ bl[17] br[17] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_20 
+ bl[18] br[18] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_21 
+ bl[19] br[19] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_22 
+ bl[20] br[20] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_23 
+ bl[21] br[21] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_24 
+ bl[22] br[22] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_25 
+ bl[23] br[23] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_26 
+ bl[24] br[24] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_27 
+ bl[25] br[25] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_28 
+ bl[26] br[26] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_29 
+ bl[27] br[27] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_30 
+ bl[28] br[28] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_31 
+ bl[29] br[29] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_32 
+ bl[30] br[30] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_33 
+ bl[31] br[31] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_34 
+ bl[32] br[32] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_35 
+ bl[33] br[33] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_36 
+ bl[34] br[34] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_37 
+ bl[35] br[35] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_38 
+ bl[36] br[36] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_39 
+ bl[37] br[37] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_40 
+ bl[38] br[38] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_41 
+ bl[39] br[39] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_42 
+ bl[40] br[40] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_43 
+ bl[41] br[41] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_44 
+ bl[42] br[42] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_45 
+ bl[43] br[43] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_46 
+ bl[44] br[44] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_47 
+ bl[45] br[45] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_48 
+ bl[46] br[46] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_49 
+ bl[47] br[47] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_50 
+ bl[48] br[48] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_51 
+ bl[49] br[49] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_52 
+ bl[50] br[50] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_53 
+ bl[51] br[51] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_54 
+ bl[52] br[52] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_55 
+ bl[53] br[53] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_56 
+ bl[54] br[54] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_57 
+ bl[55] br[55] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_58 
+ bl[56] br[56] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_59 
+ bl[57] br[57] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_60 
+ bl[58] br[58] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_61 
+ bl[59] br[59] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_62 
+ bl[60] br[60] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_63 
+ bl[61] br[61] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_64 
+ bl[62] br[62] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_65 
+ bl[63] br[63] vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_66 
+ vdd vdd vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_363_67 
+ vdd vdd vdd vss wl[361] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_0 
+ vdd vdd vss vdd vpb vnb wl[362] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_364_1 
+ rbl rbr vss vdd vpb vnb wl[362] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_364_2 
+ bl[0] br[0] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_3 
+ bl[1] br[1] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_4 
+ bl[2] br[2] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_5 
+ bl[3] br[3] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_6 
+ bl[4] br[4] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_7 
+ bl[5] br[5] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_8 
+ bl[6] br[6] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_9 
+ bl[7] br[7] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_10 
+ bl[8] br[8] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_11 
+ bl[9] br[9] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_12 
+ bl[10] br[10] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_13 
+ bl[11] br[11] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_14 
+ bl[12] br[12] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_15 
+ bl[13] br[13] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_16 
+ bl[14] br[14] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_17 
+ bl[15] br[15] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_18 
+ bl[16] br[16] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_19 
+ bl[17] br[17] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_20 
+ bl[18] br[18] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_21 
+ bl[19] br[19] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_22 
+ bl[20] br[20] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_23 
+ bl[21] br[21] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_24 
+ bl[22] br[22] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_25 
+ bl[23] br[23] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_26 
+ bl[24] br[24] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_27 
+ bl[25] br[25] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_28 
+ bl[26] br[26] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_29 
+ bl[27] br[27] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_30 
+ bl[28] br[28] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_31 
+ bl[29] br[29] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_32 
+ bl[30] br[30] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_33 
+ bl[31] br[31] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_34 
+ bl[32] br[32] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_35 
+ bl[33] br[33] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_36 
+ bl[34] br[34] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_37 
+ bl[35] br[35] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_38 
+ bl[36] br[36] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_39 
+ bl[37] br[37] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_40 
+ bl[38] br[38] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_41 
+ bl[39] br[39] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_42 
+ bl[40] br[40] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_43 
+ bl[41] br[41] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_44 
+ bl[42] br[42] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_45 
+ bl[43] br[43] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_46 
+ bl[44] br[44] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_47 
+ bl[45] br[45] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_48 
+ bl[46] br[46] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_49 
+ bl[47] br[47] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_50 
+ bl[48] br[48] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_51 
+ bl[49] br[49] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_52 
+ bl[50] br[50] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_53 
+ bl[51] br[51] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_54 
+ bl[52] br[52] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_55 
+ bl[53] br[53] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_56 
+ bl[54] br[54] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_57 
+ bl[55] br[55] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_58 
+ bl[56] br[56] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_59 
+ bl[57] br[57] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_60 
+ bl[58] br[58] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_61 
+ bl[59] br[59] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_62 
+ bl[60] br[60] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_63 
+ bl[61] br[61] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_64 
+ bl[62] br[62] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_65 
+ bl[63] br[63] vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_66 
+ vdd vdd vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_364_67 
+ vdd vdd vdd vss wl[362] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_0 
+ vdd vdd vss vdd vpb vnb wl[363] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_365_1 
+ rbl rbr vss vdd vpb vnb wl[363] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_365_2 
+ bl[0] br[0] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_3 
+ bl[1] br[1] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_4 
+ bl[2] br[2] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_5 
+ bl[3] br[3] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_6 
+ bl[4] br[4] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_7 
+ bl[5] br[5] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_8 
+ bl[6] br[6] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_9 
+ bl[7] br[7] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_10 
+ bl[8] br[8] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_11 
+ bl[9] br[9] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_12 
+ bl[10] br[10] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_13 
+ bl[11] br[11] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_14 
+ bl[12] br[12] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_15 
+ bl[13] br[13] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_16 
+ bl[14] br[14] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_17 
+ bl[15] br[15] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_18 
+ bl[16] br[16] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_19 
+ bl[17] br[17] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_20 
+ bl[18] br[18] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_21 
+ bl[19] br[19] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_22 
+ bl[20] br[20] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_23 
+ bl[21] br[21] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_24 
+ bl[22] br[22] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_25 
+ bl[23] br[23] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_26 
+ bl[24] br[24] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_27 
+ bl[25] br[25] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_28 
+ bl[26] br[26] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_29 
+ bl[27] br[27] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_30 
+ bl[28] br[28] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_31 
+ bl[29] br[29] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_32 
+ bl[30] br[30] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_33 
+ bl[31] br[31] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_34 
+ bl[32] br[32] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_35 
+ bl[33] br[33] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_36 
+ bl[34] br[34] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_37 
+ bl[35] br[35] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_38 
+ bl[36] br[36] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_39 
+ bl[37] br[37] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_40 
+ bl[38] br[38] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_41 
+ bl[39] br[39] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_42 
+ bl[40] br[40] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_43 
+ bl[41] br[41] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_44 
+ bl[42] br[42] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_45 
+ bl[43] br[43] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_46 
+ bl[44] br[44] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_47 
+ bl[45] br[45] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_48 
+ bl[46] br[46] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_49 
+ bl[47] br[47] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_50 
+ bl[48] br[48] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_51 
+ bl[49] br[49] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_52 
+ bl[50] br[50] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_53 
+ bl[51] br[51] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_54 
+ bl[52] br[52] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_55 
+ bl[53] br[53] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_56 
+ bl[54] br[54] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_57 
+ bl[55] br[55] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_58 
+ bl[56] br[56] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_59 
+ bl[57] br[57] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_60 
+ bl[58] br[58] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_61 
+ bl[59] br[59] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_62 
+ bl[60] br[60] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_63 
+ bl[61] br[61] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_64 
+ bl[62] br[62] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_65 
+ bl[63] br[63] vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_66 
+ vdd vdd vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_365_67 
+ vdd vdd vdd vss wl[363] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_0 
+ vdd vdd vss vdd vpb vnb wl[364] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_366_1 
+ rbl rbr vss vdd vpb vnb wl[364] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_366_2 
+ bl[0] br[0] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_3 
+ bl[1] br[1] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_4 
+ bl[2] br[2] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_5 
+ bl[3] br[3] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_6 
+ bl[4] br[4] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_7 
+ bl[5] br[5] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_8 
+ bl[6] br[6] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_9 
+ bl[7] br[7] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_10 
+ bl[8] br[8] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_11 
+ bl[9] br[9] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_12 
+ bl[10] br[10] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_13 
+ bl[11] br[11] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_14 
+ bl[12] br[12] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_15 
+ bl[13] br[13] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_16 
+ bl[14] br[14] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_17 
+ bl[15] br[15] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_18 
+ bl[16] br[16] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_19 
+ bl[17] br[17] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_20 
+ bl[18] br[18] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_21 
+ bl[19] br[19] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_22 
+ bl[20] br[20] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_23 
+ bl[21] br[21] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_24 
+ bl[22] br[22] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_25 
+ bl[23] br[23] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_26 
+ bl[24] br[24] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_27 
+ bl[25] br[25] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_28 
+ bl[26] br[26] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_29 
+ bl[27] br[27] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_30 
+ bl[28] br[28] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_31 
+ bl[29] br[29] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_32 
+ bl[30] br[30] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_33 
+ bl[31] br[31] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_34 
+ bl[32] br[32] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_35 
+ bl[33] br[33] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_36 
+ bl[34] br[34] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_37 
+ bl[35] br[35] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_38 
+ bl[36] br[36] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_39 
+ bl[37] br[37] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_40 
+ bl[38] br[38] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_41 
+ bl[39] br[39] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_42 
+ bl[40] br[40] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_43 
+ bl[41] br[41] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_44 
+ bl[42] br[42] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_45 
+ bl[43] br[43] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_46 
+ bl[44] br[44] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_47 
+ bl[45] br[45] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_48 
+ bl[46] br[46] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_49 
+ bl[47] br[47] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_50 
+ bl[48] br[48] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_51 
+ bl[49] br[49] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_52 
+ bl[50] br[50] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_53 
+ bl[51] br[51] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_54 
+ bl[52] br[52] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_55 
+ bl[53] br[53] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_56 
+ bl[54] br[54] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_57 
+ bl[55] br[55] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_58 
+ bl[56] br[56] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_59 
+ bl[57] br[57] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_60 
+ bl[58] br[58] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_61 
+ bl[59] br[59] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_62 
+ bl[60] br[60] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_63 
+ bl[61] br[61] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_64 
+ bl[62] br[62] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_65 
+ bl[63] br[63] vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_66 
+ vdd vdd vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_366_67 
+ vdd vdd vdd vss wl[364] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_0 
+ vdd vdd vss vdd vpb vnb wl[365] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_367_1 
+ rbl rbr vss vdd vpb vnb wl[365] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_367_2 
+ bl[0] br[0] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_3 
+ bl[1] br[1] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_4 
+ bl[2] br[2] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_5 
+ bl[3] br[3] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_6 
+ bl[4] br[4] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_7 
+ bl[5] br[5] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_8 
+ bl[6] br[6] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_9 
+ bl[7] br[7] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_10 
+ bl[8] br[8] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_11 
+ bl[9] br[9] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_12 
+ bl[10] br[10] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_13 
+ bl[11] br[11] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_14 
+ bl[12] br[12] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_15 
+ bl[13] br[13] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_16 
+ bl[14] br[14] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_17 
+ bl[15] br[15] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_18 
+ bl[16] br[16] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_19 
+ bl[17] br[17] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_20 
+ bl[18] br[18] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_21 
+ bl[19] br[19] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_22 
+ bl[20] br[20] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_23 
+ bl[21] br[21] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_24 
+ bl[22] br[22] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_25 
+ bl[23] br[23] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_26 
+ bl[24] br[24] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_27 
+ bl[25] br[25] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_28 
+ bl[26] br[26] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_29 
+ bl[27] br[27] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_30 
+ bl[28] br[28] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_31 
+ bl[29] br[29] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_32 
+ bl[30] br[30] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_33 
+ bl[31] br[31] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_34 
+ bl[32] br[32] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_35 
+ bl[33] br[33] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_36 
+ bl[34] br[34] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_37 
+ bl[35] br[35] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_38 
+ bl[36] br[36] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_39 
+ bl[37] br[37] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_40 
+ bl[38] br[38] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_41 
+ bl[39] br[39] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_42 
+ bl[40] br[40] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_43 
+ bl[41] br[41] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_44 
+ bl[42] br[42] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_45 
+ bl[43] br[43] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_46 
+ bl[44] br[44] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_47 
+ bl[45] br[45] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_48 
+ bl[46] br[46] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_49 
+ bl[47] br[47] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_50 
+ bl[48] br[48] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_51 
+ bl[49] br[49] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_52 
+ bl[50] br[50] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_53 
+ bl[51] br[51] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_54 
+ bl[52] br[52] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_55 
+ bl[53] br[53] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_56 
+ bl[54] br[54] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_57 
+ bl[55] br[55] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_58 
+ bl[56] br[56] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_59 
+ bl[57] br[57] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_60 
+ bl[58] br[58] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_61 
+ bl[59] br[59] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_62 
+ bl[60] br[60] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_63 
+ bl[61] br[61] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_64 
+ bl[62] br[62] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_65 
+ bl[63] br[63] vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_66 
+ vdd vdd vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_367_67 
+ vdd vdd vdd vss wl[365] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_0 
+ vdd vdd vss vdd vpb vnb wl[366] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_368_1 
+ rbl rbr vss vdd vpb vnb wl[366] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_368_2 
+ bl[0] br[0] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_3 
+ bl[1] br[1] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_4 
+ bl[2] br[2] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_5 
+ bl[3] br[3] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_6 
+ bl[4] br[4] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_7 
+ bl[5] br[5] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_8 
+ bl[6] br[6] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_9 
+ bl[7] br[7] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_10 
+ bl[8] br[8] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_11 
+ bl[9] br[9] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_12 
+ bl[10] br[10] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_13 
+ bl[11] br[11] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_14 
+ bl[12] br[12] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_15 
+ bl[13] br[13] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_16 
+ bl[14] br[14] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_17 
+ bl[15] br[15] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_18 
+ bl[16] br[16] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_19 
+ bl[17] br[17] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_20 
+ bl[18] br[18] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_21 
+ bl[19] br[19] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_22 
+ bl[20] br[20] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_23 
+ bl[21] br[21] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_24 
+ bl[22] br[22] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_25 
+ bl[23] br[23] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_26 
+ bl[24] br[24] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_27 
+ bl[25] br[25] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_28 
+ bl[26] br[26] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_29 
+ bl[27] br[27] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_30 
+ bl[28] br[28] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_31 
+ bl[29] br[29] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_32 
+ bl[30] br[30] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_33 
+ bl[31] br[31] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_34 
+ bl[32] br[32] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_35 
+ bl[33] br[33] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_36 
+ bl[34] br[34] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_37 
+ bl[35] br[35] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_38 
+ bl[36] br[36] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_39 
+ bl[37] br[37] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_40 
+ bl[38] br[38] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_41 
+ bl[39] br[39] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_42 
+ bl[40] br[40] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_43 
+ bl[41] br[41] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_44 
+ bl[42] br[42] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_45 
+ bl[43] br[43] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_46 
+ bl[44] br[44] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_47 
+ bl[45] br[45] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_48 
+ bl[46] br[46] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_49 
+ bl[47] br[47] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_50 
+ bl[48] br[48] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_51 
+ bl[49] br[49] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_52 
+ bl[50] br[50] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_53 
+ bl[51] br[51] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_54 
+ bl[52] br[52] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_55 
+ bl[53] br[53] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_56 
+ bl[54] br[54] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_57 
+ bl[55] br[55] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_58 
+ bl[56] br[56] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_59 
+ bl[57] br[57] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_60 
+ bl[58] br[58] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_61 
+ bl[59] br[59] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_62 
+ bl[60] br[60] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_63 
+ bl[61] br[61] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_64 
+ bl[62] br[62] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_65 
+ bl[63] br[63] vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_66 
+ vdd vdd vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_368_67 
+ vdd vdd vdd vss wl[366] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_0 
+ vdd vdd vss vdd vpb vnb wl[367] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_369_1 
+ rbl rbr vss vdd vpb vnb wl[367] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_369_2 
+ bl[0] br[0] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_3 
+ bl[1] br[1] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_4 
+ bl[2] br[2] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_5 
+ bl[3] br[3] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_6 
+ bl[4] br[4] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_7 
+ bl[5] br[5] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_8 
+ bl[6] br[6] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_9 
+ bl[7] br[7] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_10 
+ bl[8] br[8] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_11 
+ bl[9] br[9] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_12 
+ bl[10] br[10] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_13 
+ bl[11] br[11] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_14 
+ bl[12] br[12] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_15 
+ bl[13] br[13] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_16 
+ bl[14] br[14] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_17 
+ bl[15] br[15] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_18 
+ bl[16] br[16] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_19 
+ bl[17] br[17] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_20 
+ bl[18] br[18] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_21 
+ bl[19] br[19] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_22 
+ bl[20] br[20] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_23 
+ bl[21] br[21] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_24 
+ bl[22] br[22] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_25 
+ bl[23] br[23] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_26 
+ bl[24] br[24] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_27 
+ bl[25] br[25] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_28 
+ bl[26] br[26] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_29 
+ bl[27] br[27] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_30 
+ bl[28] br[28] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_31 
+ bl[29] br[29] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_32 
+ bl[30] br[30] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_33 
+ bl[31] br[31] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_34 
+ bl[32] br[32] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_35 
+ bl[33] br[33] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_36 
+ bl[34] br[34] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_37 
+ bl[35] br[35] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_38 
+ bl[36] br[36] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_39 
+ bl[37] br[37] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_40 
+ bl[38] br[38] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_41 
+ bl[39] br[39] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_42 
+ bl[40] br[40] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_43 
+ bl[41] br[41] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_44 
+ bl[42] br[42] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_45 
+ bl[43] br[43] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_46 
+ bl[44] br[44] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_47 
+ bl[45] br[45] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_48 
+ bl[46] br[46] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_49 
+ bl[47] br[47] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_50 
+ bl[48] br[48] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_51 
+ bl[49] br[49] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_52 
+ bl[50] br[50] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_53 
+ bl[51] br[51] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_54 
+ bl[52] br[52] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_55 
+ bl[53] br[53] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_56 
+ bl[54] br[54] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_57 
+ bl[55] br[55] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_58 
+ bl[56] br[56] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_59 
+ bl[57] br[57] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_60 
+ bl[58] br[58] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_61 
+ bl[59] br[59] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_62 
+ bl[60] br[60] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_63 
+ bl[61] br[61] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_64 
+ bl[62] br[62] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_65 
+ bl[63] br[63] vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_66 
+ vdd vdd vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_369_67 
+ vdd vdd vdd vss wl[367] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_0 
+ vdd vdd vss vdd vpb vnb wl[368] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_370_1 
+ rbl rbr vss vdd vpb vnb wl[368] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_370_2 
+ bl[0] br[0] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_3 
+ bl[1] br[1] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_4 
+ bl[2] br[2] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_5 
+ bl[3] br[3] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_6 
+ bl[4] br[4] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_7 
+ bl[5] br[5] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_8 
+ bl[6] br[6] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_9 
+ bl[7] br[7] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_10 
+ bl[8] br[8] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_11 
+ bl[9] br[9] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_12 
+ bl[10] br[10] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_13 
+ bl[11] br[11] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_14 
+ bl[12] br[12] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_15 
+ bl[13] br[13] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_16 
+ bl[14] br[14] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_17 
+ bl[15] br[15] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_18 
+ bl[16] br[16] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_19 
+ bl[17] br[17] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_20 
+ bl[18] br[18] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_21 
+ bl[19] br[19] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_22 
+ bl[20] br[20] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_23 
+ bl[21] br[21] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_24 
+ bl[22] br[22] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_25 
+ bl[23] br[23] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_26 
+ bl[24] br[24] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_27 
+ bl[25] br[25] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_28 
+ bl[26] br[26] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_29 
+ bl[27] br[27] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_30 
+ bl[28] br[28] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_31 
+ bl[29] br[29] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_32 
+ bl[30] br[30] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_33 
+ bl[31] br[31] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_34 
+ bl[32] br[32] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_35 
+ bl[33] br[33] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_36 
+ bl[34] br[34] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_37 
+ bl[35] br[35] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_38 
+ bl[36] br[36] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_39 
+ bl[37] br[37] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_40 
+ bl[38] br[38] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_41 
+ bl[39] br[39] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_42 
+ bl[40] br[40] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_43 
+ bl[41] br[41] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_44 
+ bl[42] br[42] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_45 
+ bl[43] br[43] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_46 
+ bl[44] br[44] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_47 
+ bl[45] br[45] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_48 
+ bl[46] br[46] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_49 
+ bl[47] br[47] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_50 
+ bl[48] br[48] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_51 
+ bl[49] br[49] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_52 
+ bl[50] br[50] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_53 
+ bl[51] br[51] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_54 
+ bl[52] br[52] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_55 
+ bl[53] br[53] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_56 
+ bl[54] br[54] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_57 
+ bl[55] br[55] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_58 
+ bl[56] br[56] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_59 
+ bl[57] br[57] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_60 
+ bl[58] br[58] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_61 
+ bl[59] br[59] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_62 
+ bl[60] br[60] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_63 
+ bl[61] br[61] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_64 
+ bl[62] br[62] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_65 
+ bl[63] br[63] vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_66 
+ vdd vdd vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_370_67 
+ vdd vdd vdd vss wl[368] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_0 
+ vdd vdd vss vdd vpb vnb wl[369] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_371_1 
+ rbl rbr vss vdd vpb vnb wl[369] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_371_2 
+ bl[0] br[0] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_3 
+ bl[1] br[1] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_4 
+ bl[2] br[2] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_5 
+ bl[3] br[3] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_6 
+ bl[4] br[4] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_7 
+ bl[5] br[5] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_8 
+ bl[6] br[6] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_9 
+ bl[7] br[7] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_10 
+ bl[8] br[8] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_11 
+ bl[9] br[9] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_12 
+ bl[10] br[10] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_13 
+ bl[11] br[11] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_14 
+ bl[12] br[12] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_15 
+ bl[13] br[13] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_16 
+ bl[14] br[14] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_17 
+ bl[15] br[15] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_18 
+ bl[16] br[16] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_19 
+ bl[17] br[17] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_20 
+ bl[18] br[18] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_21 
+ bl[19] br[19] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_22 
+ bl[20] br[20] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_23 
+ bl[21] br[21] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_24 
+ bl[22] br[22] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_25 
+ bl[23] br[23] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_26 
+ bl[24] br[24] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_27 
+ bl[25] br[25] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_28 
+ bl[26] br[26] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_29 
+ bl[27] br[27] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_30 
+ bl[28] br[28] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_31 
+ bl[29] br[29] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_32 
+ bl[30] br[30] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_33 
+ bl[31] br[31] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_34 
+ bl[32] br[32] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_35 
+ bl[33] br[33] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_36 
+ bl[34] br[34] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_37 
+ bl[35] br[35] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_38 
+ bl[36] br[36] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_39 
+ bl[37] br[37] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_40 
+ bl[38] br[38] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_41 
+ bl[39] br[39] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_42 
+ bl[40] br[40] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_43 
+ bl[41] br[41] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_44 
+ bl[42] br[42] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_45 
+ bl[43] br[43] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_46 
+ bl[44] br[44] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_47 
+ bl[45] br[45] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_48 
+ bl[46] br[46] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_49 
+ bl[47] br[47] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_50 
+ bl[48] br[48] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_51 
+ bl[49] br[49] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_52 
+ bl[50] br[50] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_53 
+ bl[51] br[51] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_54 
+ bl[52] br[52] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_55 
+ bl[53] br[53] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_56 
+ bl[54] br[54] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_57 
+ bl[55] br[55] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_58 
+ bl[56] br[56] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_59 
+ bl[57] br[57] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_60 
+ bl[58] br[58] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_61 
+ bl[59] br[59] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_62 
+ bl[60] br[60] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_63 
+ bl[61] br[61] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_64 
+ bl[62] br[62] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_65 
+ bl[63] br[63] vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_66 
+ vdd vdd vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_371_67 
+ vdd vdd vdd vss wl[369] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_0 
+ vdd vdd vss vdd vpb vnb wl[370] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_372_1 
+ rbl rbr vss vdd vpb vnb wl[370] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_372_2 
+ bl[0] br[0] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_3 
+ bl[1] br[1] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_4 
+ bl[2] br[2] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_5 
+ bl[3] br[3] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_6 
+ bl[4] br[4] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_7 
+ bl[5] br[5] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_8 
+ bl[6] br[6] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_9 
+ bl[7] br[7] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_10 
+ bl[8] br[8] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_11 
+ bl[9] br[9] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_12 
+ bl[10] br[10] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_13 
+ bl[11] br[11] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_14 
+ bl[12] br[12] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_15 
+ bl[13] br[13] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_16 
+ bl[14] br[14] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_17 
+ bl[15] br[15] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_18 
+ bl[16] br[16] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_19 
+ bl[17] br[17] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_20 
+ bl[18] br[18] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_21 
+ bl[19] br[19] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_22 
+ bl[20] br[20] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_23 
+ bl[21] br[21] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_24 
+ bl[22] br[22] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_25 
+ bl[23] br[23] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_26 
+ bl[24] br[24] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_27 
+ bl[25] br[25] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_28 
+ bl[26] br[26] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_29 
+ bl[27] br[27] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_30 
+ bl[28] br[28] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_31 
+ bl[29] br[29] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_32 
+ bl[30] br[30] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_33 
+ bl[31] br[31] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_34 
+ bl[32] br[32] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_35 
+ bl[33] br[33] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_36 
+ bl[34] br[34] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_37 
+ bl[35] br[35] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_38 
+ bl[36] br[36] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_39 
+ bl[37] br[37] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_40 
+ bl[38] br[38] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_41 
+ bl[39] br[39] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_42 
+ bl[40] br[40] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_43 
+ bl[41] br[41] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_44 
+ bl[42] br[42] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_45 
+ bl[43] br[43] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_46 
+ bl[44] br[44] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_47 
+ bl[45] br[45] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_48 
+ bl[46] br[46] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_49 
+ bl[47] br[47] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_50 
+ bl[48] br[48] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_51 
+ bl[49] br[49] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_52 
+ bl[50] br[50] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_53 
+ bl[51] br[51] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_54 
+ bl[52] br[52] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_55 
+ bl[53] br[53] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_56 
+ bl[54] br[54] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_57 
+ bl[55] br[55] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_58 
+ bl[56] br[56] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_59 
+ bl[57] br[57] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_60 
+ bl[58] br[58] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_61 
+ bl[59] br[59] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_62 
+ bl[60] br[60] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_63 
+ bl[61] br[61] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_64 
+ bl[62] br[62] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_65 
+ bl[63] br[63] vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_66 
+ vdd vdd vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_372_67 
+ vdd vdd vdd vss wl[370] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_0 
+ vdd vdd vss vdd vpb vnb wl[371] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_373_1 
+ rbl rbr vss vdd vpb vnb wl[371] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_373_2 
+ bl[0] br[0] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_3 
+ bl[1] br[1] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_4 
+ bl[2] br[2] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_5 
+ bl[3] br[3] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_6 
+ bl[4] br[4] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_7 
+ bl[5] br[5] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_8 
+ bl[6] br[6] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_9 
+ bl[7] br[7] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_10 
+ bl[8] br[8] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_11 
+ bl[9] br[9] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_12 
+ bl[10] br[10] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_13 
+ bl[11] br[11] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_14 
+ bl[12] br[12] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_15 
+ bl[13] br[13] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_16 
+ bl[14] br[14] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_17 
+ bl[15] br[15] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_18 
+ bl[16] br[16] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_19 
+ bl[17] br[17] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_20 
+ bl[18] br[18] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_21 
+ bl[19] br[19] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_22 
+ bl[20] br[20] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_23 
+ bl[21] br[21] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_24 
+ bl[22] br[22] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_25 
+ bl[23] br[23] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_26 
+ bl[24] br[24] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_27 
+ bl[25] br[25] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_28 
+ bl[26] br[26] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_29 
+ bl[27] br[27] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_30 
+ bl[28] br[28] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_31 
+ bl[29] br[29] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_32 
+ bl[30] br[30] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_33 
+ bl[31] br[31] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_34 
+ bl[32] br[32] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_35 
+ bl[33] br[33] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_36 
+ bl[34] br[34] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_37 
+ bl[35] br[35] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_38 
+ bl[36] br[36] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_39 
+ bl[37] br[37] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_40 
+ bl[38] br[38] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_41 
+ bl[39] br[39] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_42 
+ bl[40] br[40] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_43 
+ bl[41] br[41] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_44 
+ bl[42] br[42] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_45 
+ bl[43] br[43] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_46 
+ bl[44] br[44] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_47 
+ bl[45] br[45] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_48 
+ bl[46] br[46] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_49 
+ bl[47] br[47] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_50 
+ bl[48] br[48] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_51 
+ bl[49] br[49] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_52 
+ bl[50] br[50] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_53 
+ bl[51] br[51] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_54 
+ bl[52] br[52] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_55 
+ bl[53] br[53] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_56 
+ bl[54] br[54] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_57 
+ bl[55] br[55] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_58 
+ bl[56] br[56] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_59 
+ bl[57] br[57] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_60 
+ bl[58] br[58] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_61 
+ bl[59] br[59] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_62 
+ bl[60] br[60] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_63 
+ bl[61] br[61] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_64 
+ bl[62] br[62] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_65 
+ bl[63] br[63] vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_66 
+ vdd vdd vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_373_67 
+ vdd vdd vdd vss wl[371] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_0 
+ vdd vdd vss vdd vpb vnb wl[372] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_374_1 
+ rbl rbr vss vdd vpb vnb wl[372] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_374_2 
+ bl[0] br[0] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_3 
+ bl[1] br[1] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_4 
+ bl[2] br[2] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_5 
+ bl[3] br[3] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_6 
+ bl[4] br[4] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_7 
+ bl[5] br[5] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_8 
+ bl[6] br[6] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_9 
+ bl[7] br[7] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_10 
+ bl[8] br[8] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_11 
+ bl[9] br[9] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_12 
+ bl[10] br[10] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_13 
+ bl[11] br[11] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_14 
+ bl[12] br[12] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_15 
+ bl[13] br[13] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_16 
+ bl[14] br[14] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_17 
+ bl[15] br[15] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_18 
+ bl[16] br[16] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_19 
+ bl[17] br[17] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_20 
+ bl[18] br[18] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_21 
+ bl[19] br[19] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_22 
+ bl[20] br[20] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_23 
+ bl[21] br[21] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_24 
+ bl[22] br[22] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_25 
+ bl[23] br[23] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_26 
+ bl[24] br[24] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_27 
+ bl[25] br[25] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_28 
+ bl[26] br[26] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_29 
+ bl[27] br[27] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_30 
+ bl[28] br[28] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_31 
+ bl[29] br[29] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_32 
+ bl[30] br[30] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_33 
+ bl[31] br[31] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_34 
+ bl[32] br[32] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_35 
+ bl[33] br[33] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_36 
+ bl[34] br[34] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_37 
+ bl[35] br[35] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_38 
+ bl[36] br[36] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_39 
+ bl[37] br[37] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_40 
+ bl[38] br[38] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_41 
+ bl[39] br[39] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_42 
+ bl[40] br[40] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_43 
+ bl[41] br[41] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_44 
+ bl[42] br[42] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_45 
+ bl[43] br[43] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_46 
+ bl[44] br[44] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_47 
+ bl[45] br[45] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_48 
+ bl[46] br[46] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_49 
+ bl[47] br[47] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_50 
+ bl[48] br[48] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_51 
+ bl[49] br[49] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_52 
+ bl[50] br[50] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_53 
+ bl[51] br[51] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_54 
+ bl[52] br[52] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_55 
+ bl[53] br[53] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_56 
+ bl[54] br[54] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_57 
+ bl[55] br[55] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_58 
+ bl[56] br[56] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_59 
+ bl[57] br[57] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_60 
+ bl[58] br[58] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_61 
+ bl[59] br[59] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_62 
+ bl[60] br[60] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_63 
+ bl[61] br[61] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_64 
+ bl[62] br[62] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_65 
+ bl[63] br[63] vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_66 
+ vdd vdd vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_374_67 
+ vdd vdd vdd vss wl[372] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_0 
+ vdd vdd vss vdd vpb vnb wl[373] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_375_1 
+ rbl rbr vss vdd vpb vnb wl[373] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_375_2 
+ bl[0] br[0] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_3 
+ bl[1] br[1] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_4 
+ bl[2] br[2] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_5 
+ bl[3] br[3] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_6 
+ bl[4] br[4] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_7 
+ bl[5] br[5] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_8 
+ bl[6] br[6] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_9 
+ bl[7] br[7] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_10 
+ bl[8] br[8] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_11 
+ bl[9] br[9] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_12 
+ bl[10] br[10] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_13 
+ bl[11] br[11] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_14 
+ bl[12] br[12] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_15 
+ bl[13] br[13] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_16 
+ bl[14] br[14] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_17 
+ bl[15] br[15] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_18 
+ bl[16] br[16] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_19 
+ bl[17] br[17] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_20 
+ bl[18] br[18] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_21 
+ bl[19] br[19] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_22 
+ bl[20] br[20] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_23 
+ bl[21] br[21] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_24 
+ bl[22] br[22] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_25 
+ bl[23] br[23] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_26 
+ bl[24] br[24] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_27 
+ bl[25] br[25] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_28 
+ bl[26] br[26] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_29 
+ bl[27] br[27] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_30 
+ bl[28] br[28] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_31 
+ bl[29] br[29] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_32 
+ bl[30] br[30] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_33 
+ bl[31] br[31] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_34 
+ bl[32] br[32] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_35 
+ bl[33] br[33] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_36 
+ bl[34] br[34] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_37 
+ bl[35] br[35] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_38 
+ bl[36] br[36] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_39 
+ bl[37] br[37] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_40 
+ bl[38] br[38] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_41 
+ bl[39] br[39] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_42 
+ bl[40] br[40] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_43 
+ bl[41] br[41] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_44 
+ bl[42] br[42] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_45 
+ bl[43] br[43] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_46 
+ bl[44] br[44] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_47 
+ bl[45] br[45] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_48 
+ bl[46] br[46] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_49 
+ bl[47] br[47] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_50 
+ bl[48] br[48] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_51 
+ bl[49] br[49] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_52 
+ bl[50] br[50] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_53 
+ bl[51] br[51] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_54 
+ bl[52] br[52] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_55 
+ bl[53] br[53] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_56 
+ bl[54] br[54] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_57 
+ bl[55] br[55] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_58 
+ bl[56] br[56] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_59 
+ bl[57] br[57] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_60 
+ bl[58] br[58] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_61 
+ bl[59] br[59] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_62 
+ bl[60] br[60] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_63 
+ bl[61] br[61] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_64 
+ bl[62] br[62] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_65 
+ bl[63] br[63] vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_66 
+ vdd vdd vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_375_67 
+ vdd vdd vdd vss wl[373] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_0 
+ vdd vdd vss vdd vpb vnb wl[374] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_376_1 
+ rbl rbr vss vdd vpb vnb wl[374] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_376_2 
+ bl[0] br[0] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_3 
+ bl[1] br[1] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_4 
+ bl[2] br[2] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_5 
+ bl[3] br[3] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_6 
+ bl[4] br[4] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_7 
+ bl[5] br[5] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_8 
+ bl[6] br[6] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_9 
+ bl[7] br[7] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_10 
+ bl[8] br[8] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_11 
+ bl[9] br[9] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_12 
+ bl[10] br[10] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_13 
+ bl[11] br[11] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_14 
+ bl[12] br[12] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_15 
+ bl[13] br[13] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_16 
+ bl[14] br[14] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_17 
+ bl[15] br[15] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_18 
+ bl[16] br[16] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_19 
+ bl[17] br[17] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_20 
+ bl[18] br[18] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_21 
+ bl[19] br[19] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_22 
+ bl[20] br[20] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_23 
+ bl[21] br[21] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_24 
+ bl[22] br[22] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_25 
+ bl[23] br[23] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_26 
+ bl[24] br[24] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_27 
+ bl[25] br[25] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_28 
+ bl[26] br[26] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_29 
+ bl[27] br[27] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_30 
+ bl[28] br[28] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_31 
+ bl[29] br[29] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_32 
+ bl[30] br[30] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_33 
+ bl[31] br[31] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_34 
+ bl[32] br[32] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_35 
+ bl[33] br[33] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_36 
+ bl[34] br[34] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_37 
+ bl[35] br[35] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_38 
+ bl[36] br[36] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_39 
+ bl[37] br[37] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_40 
+ bl[38] br[38] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_41 
+ bl[39] br[39] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_42 
+ bl[40] br[40] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_43 
+ bl[41] br[41] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_44 
+ bl[42] br[42] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_45 
+ bl[43] br[43] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_46 
+ bl[44] br[44] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_47 
+ bl[45] br[45] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_48 
+ bl[46] br[46] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_49 
+ bl[47] br[47] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_50 
+ bl[48] br[48] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_51 
+ bl[49] br[49] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_52 
+ bl[50] br[50] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_53 
+ bl[51] br[51] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_54 
+ bl[52] br[52] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_55 
+ bl[53] br[53] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_56 
+ bl[54] br[54] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_57 
+ bl[55] br[55] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_58 
+ bl[56] br[56] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_59 
+ bl[57] br[57] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_60 
+ bl[58] br[58] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_61 
+ bl[59] br[59] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_62 
+ bl[60] br[60] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_63 
+ bl[61] br[61] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_64 
+ bl[62] br[62] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_65 
+ bl[63] br[63] vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_66 
+ vdd vdd vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_376_67 
+ vdd vdd vdd vss wl[374] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_0 
+ vdd vdd vss vdd vpb vnb wl[375] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_377_1 
+ rbl rbr vss vdd vpb vnb wl[375] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_377_2 
+ bl[0] br[0] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_3 
+ bl[1] br[1] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_4 
+ bl[2] br[2] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_5 
+ bl[3] br[3] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_6 
+ bl[4] br[4] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_7 
+ bl[5] br[5] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_8 
+ bl[6] br[6] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_9 
+ bl[7] br[7] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_10 
+ bl[8] br[8] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_11 
+ bl[9] br[9] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_12 
+ bl[10] br[10] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_13 
+ bl[11] br[11] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_14 
+ bl[12] br[12] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_15 
+ bl[13] br[13] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_16 
+ bl[14] br[14] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_17 
+ bl[15] br[15] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_18 
+ bl[16] br[16] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_19 
+ bl[17] br[17] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_20 
+ bl[18] br[18] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_21 
+ bl[19] br[19] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_22 
+ bl[20] br[20] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_23 
+ bl[21] br[21] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_24 
+ bl[22] br[22] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_25 
+ bl[23] br[23] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_26 
+ bl[24] br[24] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_27 
+ bl[25] br[25] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_28 
+ bl[26] br[26] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_29 
+ bl[27] br[27] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_30 
+ bl[28] br[28] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_31 
+ bl[29] br[29] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_32 
+ bl[30] br[30] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_33 
+ bl[31] br[31] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_34 
+ bl[32] br[32] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_35 
+ bl[33] br[33] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_36 
+ bl[34] br[34] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_37 
+ bl[35] br[35] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_38 
+ bl[36] br[36] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_39 
+ bl[37] br[37] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_40 
+ bl[38] br[38] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_41 
+ bl[39] br[39] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_42 
+ bl[40] br[40] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_43 
+ bl[41] br[41] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_44 
+ bl[42] br[42] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_45 
+ bl[43] br[43] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_46 
+ bl[44] br[44] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_47 
+ bl[45] br[45] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_48 
+ bl[46] br[46] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_49 
+ bl[47] br[47] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_50 
+ bl[48] br[48] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_51 
+ bl[49] br[49] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_52 
+ bl[50] br[50] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_53 
+ bl[51] br[51] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_54 
+ bl[52] br[52] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_55 
+ bl[53] br[53] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_56 
+ bl[54] br[54] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_57 
+ bl[55] br[55] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_58 
+ bl[56] br[56] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_59 
+ bl[57] br[57] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_60 
+ bl[58] br[58] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_61 
+ bl[59] br[59] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_62 
+ bl[60] br[60] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_63 
+ bl[61] br[61] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_64 
+ bl[62] br[62] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_65 
+ bl[63] br[63] vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_66 
+ vdd vdd vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_377_67 
+ vdd vdd vdd vss wl[375] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_0 
+ vdd vdd vss vdd vpb vnb wl[376] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_378_1 
+ rbl rbr vss vdd vpb vnb wl[376] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_378_2 
+ bl[0] br[0] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_3 
+ bl[1] br[1] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_4 
+ bl[2] br[2] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_5 
+ bl[3] br[3] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_6 
+ bl[4] br[4] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_7 
+ bl[5] br[5] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_8 
+ bl[6] br[6] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_9 
+ bl[7] br[7] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_10 
+ bl[8] br[8] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_11 
+ bl[9] br[9] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_12 
+ bl[10] br[10] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_13 
+ bl[11] br[11] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_14 
+ bl[12] br[12] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_15 
+ bl[13] br[13] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_16 
+ bl[14] br[14] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_17 
+ bl[15] br[15] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_18 
+ bl[16] br[16] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_19 
+ bl[17] br[17] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_20 
+ bl[18] br[18] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_21 
+ bl[19] br[19] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_22 
+ bl[20] br[20] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_23 
+ bl[21] br[21] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_24 
+ bl[22] br[22] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_25 
+ bl[23] br[23] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_26 
+ bl[24] br[24] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_27 
+ bl[25] br[25] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_28 
+ bl[26] br[26] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_29 
+ bl[27] br[27] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_30 
+ bl[28] br[28] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_31 
+ bl[29] br[29] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_32 
+ bl[30] br[30] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_33 
+ bl[31] br[31] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_34 
+ bl[32] br[32] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_35 
+ bl[33] br[33] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_36 
+ bl[34] br[34] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_37 
+ bl[35] br[35] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_38 
+ bl[36] br[36] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_39 
+ bl[37] br[37] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_40 
+ bl[38] br[38] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_41 
+ bl[39] br[39] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_42 
+ bl[40] br[40] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_43 
+ bl[41] br[41] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_44 
+ bl[42] br[42] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_45 
+ bl[43] br[43] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_46 
+ bl[44] br[44] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_47 
+ bl[45] br[45] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_48 
+ bl[46] br[46] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_49 
+ bl[47] br[47] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_50 
+ bl[48] br[48] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_51 
+ bl[49] br[49] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_52 
+ bl[50] br[50] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_53 
+ bl[51] br[51] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_54 
+ bl[52] br[52] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_55 
+ bl[53] br[53] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_56 
+ bl[54] br[54] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_57 
+ bl[55] br[55] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_58 
+ bl[56] br[56] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_59 
+ bl[57] br[57] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_60 
+ bl[58] br[58] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_61 
+ bl[59] br[59] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_62 
+ bl[60] br[60] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_63 
+ bl[61] br[61] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_64 
+ bl[62] br[62] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_65 
+ bl[63] br[63] vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_66 
+ vdd vdd vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_378_67 
+ vdd vdd vdd vss wl[376] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_0 
+ vdd vdd vss vdd vpb vnb wl[377] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_379_1 
+ rbl rbr vss vdd vpb vnb wl[377] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_379_2 
+ bl[0] br[0] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_3 
+ bl[1] br[1] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_4 
+ bl[2] br[2] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_5 
+ bl[3] br[3] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_6 
+ bl[4] br[4] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_7 
+ bl[5] br[5] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_8 
+ bl[6] br[6] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_9 
+ bl[7] br[7] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_10 
+ bl[8] br[8] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_11 
+ bl[9] br[9] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_12 
+ bl[10] br[10] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_13 
+ bl[11] br[11] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_14 
+ bl[12] br[12] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_15 
+ bl[13] br[13] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_16 
+ bl[14] br[14] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_17 
+ bl[15] br[15] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_18 
+ bl[16] br[16] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_19 
+ bl[17] br[17] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_20 
+ bl[18] br[18] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_21 
+ bl[19] br[19] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_22 
+ bl[20] br[20] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_23 
+ bl[21] br[21] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_24 
+ bl[22] br[22] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_25 
+ bl[23] br[23] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_26 
+ bl[24] br[24] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_27 
+ bl[25] br[25] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_28 
+ bl[26] br[26] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_29 
+ bl[27] br[27] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_30 
+ bl[28] br[28] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_31 
+ bl[29] br[29] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_32 
+ bl[30] br[30] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_33 
+ bl[31] br[31] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_34 
+ bl[32] br[32] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_35 
+ bl[33] br[33] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_36 
+ bl[34] br[34] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_37 
+ bl[35] br[35] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_38 
+ bl[36] br[36] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_39 
+ bl[37] br[37] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_40 
+ bl[38] br[38] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_41 
+ bl[39] br[39] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_42 
+ bl[40] br[40] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_43 
+ bl[41] br[41] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_44 
+ bl[42] br[42] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_45 
+ bl[43] br[43] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_46 
+ bl[44] br[44] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_47 
+ bl[45] br[45] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_48 
+ bl[46] br[46] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_49 
+ bl[47] br[47] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_50 
+ bl[48] br[48] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_51 
+ bl[49] br[49] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_52 
+ bl[50] br[50] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_53 
+ bl[51] br[51] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_54 
+ bl[52] br[52] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_55 
+ bl[53] br[53] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_56 
+ bl[54] br[54] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_57 
+ bl[55] br[55] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_58 
+ bl[56] br[56] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_59 
+ bl[57] br[57] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_60 
+ bl[58] br[58] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_61 
+ bl[59] br[59] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_62 
+ bl[60] br[60] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_63 
+ bl[61] br[61] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_64 
+ bl[62] br[62] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_65 
+ bl[63] br[63] vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_66 
+ vdd vdd vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_379_67 
+ vdd vdd vdd vss wl[377] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_0 
+ vdd vdd vss vdd vpb vnb wl[378] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_380_1 
+ rbl rbr vss vdd vpb vnb wl[378] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_380_2 
+ bl[0] br[0] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_3 
+ bl[1] br[1] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_4 
+ bl[2] br[2] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_5 
+ bl[3] br[3] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_6 
+ bl[4] br[4] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_7 
+ bl[5] br[5] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_8 
+ bl[6] br[6] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_9 
+ bl[7] br[7] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_10 
+ bl[8] br[8] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_11 
+ bl[9] br[9] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_12 
+ bl[10] br[10] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_13 
+ bl[11] br[11] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_14 
+ bl[12] br[12] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_15 
+ bl[13] br[13] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_16 
+ bl[14] br[14] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_17 
+ bl[15] br[15] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_18 
+ bl[16] br[16] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_19 
+ bl[17] br[17] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_20 
+ bl[18] br[18] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_21 
+ bl[19] br[19] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_22 
+ bl[20] br[20] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_23 
+ bl[21] br[21] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_24 
+ bl[22] br[22] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_25 
+ bl[23] br[23] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_26 
+ bl[24] br[24] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_27 
+ bl[25] br[25] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_28 
+ bl[26] br[26] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_29 
+ bl[27] br[27] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_30 
+ bl[28] br[28] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_31 
+ bl[29] br[29] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_32 
+ bl[30] br[30] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_33 
+ bl[31] br[31] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_34 
+ bl[32] br[32] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_35 
+ bl[33] br[33] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_36 
+ bl[34] br[34] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_37 
+ bl[35] br[35] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_38 
+ bl[36] br[36] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_39 
+ bl[37] br[37] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_40 
+ bl[38] br[38] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_41 
+ bl[39] br[39] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_42 
+ bl[40] br[40] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_43 
+ bl[41] br[41] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_44 
+ bl[42] br[42] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_45 
+ bl[43] br[43] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_46 
+ bl[44] br[44] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_47 
+ bl[45] br[45] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_48 
+ bl[46] br[46] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_49 
+ bl[47] br[47] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_50 
+ bl[48] br[48] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_51 
+ bl[49] br[49] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_52 
+ bl[50] br[50] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_53 
+ bl[51] br[51] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_54 
+ bl[52] br[52] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_55 
+ bl[53] br[53] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_56 
+ bl[54] br[54] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_57 
+ bl[55] br[55] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_58 
+ bl[56] br[56] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_59 
+ bl[57] br[57] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_60 
+ bl[58] br[58] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_61 
+ bl[59] br[59] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_62 
+ bl[60] br[60] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_63 
+ bl[61] br[61] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_64 
+ bl[62] br[62] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_65 
+ bl[63] br[63] vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_66 
+ vdd vdd vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_380_67 
+ vdd vdd vdd vss wl[378] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_0 
+ vdd vdd vss vdd vpb vnb wl[379] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_381_1 
+ rbl rbr vss vdd vpb vnb wl[379] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_381_2 
+ bl[0] br[0] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_3 
+ bl[1] br[1] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_4 
+ bl[2] br[2] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_5 
+ bl[3] br[3] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_6 
+ bl[4] br[4] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_7 
+ bl[5] br[5] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_8 
+ bl[6] br[6] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_9 
+ bl[7] br[7] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_10 
+ bl[8] br[8] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_11 
+ bl[9] br[9] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_12 
+ bl[10] br[10] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_13 
+ bl[11] br[11] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_14 
+ bl[12] br[12] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_15 
+ bl[13] br[13] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_16 
+ bl[14] br[14] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_17 
+ bl[15] br[15] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_18 
+ bl[16] br[16] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_19 
+ bl[17] br[17] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_20 
+ bl[18] br[18] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_21 
+ bl[19] br[19] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_22 
+ bl[20] br[20] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_23 
+ bl[21] br[21] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_24 
+ bl[22] br[22] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_25 
+ bl[23] br[23] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_26 
+ bl[24] br[24] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_27 
+ bl[25] br[25] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_28 
+ bl[26] br[26] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_29 
+ bl[27] br[27] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_30 
+ bl[28] br[28] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_31 
+ bl[29] br[29] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_32 
+ bl[30] br[30] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_33 
+ bl[31] br[31] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_34 
+ bl[32] br[32] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_35 
+ bl[33] br[33] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_36 
+ bl[34] br[34] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_37 
+ bl[35] br[35] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_38 
+ bl[36] br[36] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_39 
+ bl[37] br[37] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_40 
+ bl[38] br[38] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_41 
+ bl[39] br[39] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_42 
+ bl[40] br[40] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_43 
+ bl[41] br[41] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_44 
+ bl[42] br[42] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_45 
+ bl[43] br[43] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_46 
+ bl[44] br[44] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_47 
+ bl[45] br[45] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_48 
+ bl[46] br[46] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_49 
+ bl[47] br[47] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_50 
+ bl[48] br[48] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_51 
+ bl[49] br[49] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_52 
+ bl[50] br[50] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_53 
+ bl[51] br[51] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_54 
+ bl[52] br[52] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_55 
+ bl[53] br[53] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_56 
+ bl[54] br[54] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_57 
+ bl[55] br[55] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_58 
+ bl[56] br[56] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_59 
+ bl[57] br[57] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_60 
+ bl[58] br[58] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_61 
+ bl[59] br[59] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_62 
+ bl[60] br[60] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_63 
+ bl[61] br[61] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_64 
+ bl[62] br[62] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_65 
+ bl[63] br[63] vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_66 
+ vdd vdd vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_381_67 
+ vdd vdd vdd vss wl[379] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_0 
+ vdd vdd vss vdd vpb vnb wl[380] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_382_1 
+ rbl rbr vss vdd vpb vnb wl[380] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_382_2 
+ bl[0] br[0] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_3 
+ bl[1] br[1] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_4 
+ bl[2] br[2] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_5 
+ bl[3] br[3] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_6 
+ bl[4] br[4] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_7 
+ bl[5] br[5] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_8 
+ bl[6] br[6] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_9 
+ bl[7] br[7] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_10 
+ bl[8] br[8] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_11 
+ bl[9] br[9] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_12 
+ bl[10] br[10] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_13 
+ bl[11] br[11] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_14 
+ bl[12] br[12] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_15 
+ bl[13] br[13] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_16 
+ bl[14] br[14] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_17 
+ bl[15] br[15] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_18 
+ bl[16] br[16] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_19 
+ bl[17] br[17] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_20 
+ bl[18] br[18] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_21 
+ bl[19] br[19] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_22 
+ bl[20] br[20] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_23 
+ bl[21] br[21] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_24 
+ bl[22] br[22] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_25 
+ bl[23] br[23] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_26 
+ bl[24] br[24] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_27 
+ bl[25] br[25] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_28 
+ bl[26] br[26] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_29 
+ bl[27] br[27] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_30 
+ bl[28] br[28] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_31 
+ bl[29] br[29] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_32 
+ bl[30] br[30] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_33 
+ bl[31] br[31] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_34 
+ bl[32] br[32] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_35 
+ bl[33] br[33] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_36 
+ bl[34] br[34] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_37 
+ bl[35] br[35] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_38 
+ bl[36] br[36] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_39 
+ bl[37] br[37] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_40 
+ bl[38] br[38] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_41 
+ bl[39] br[39] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_42 
+ bl[40] br[40] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_43 
+ bl[41] br[41] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_44 
+ bl[42] br[42] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_45 
+ bl[43] br[43] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_46 
+ bl[44] br[44] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_47 
+ bl[45] br[45] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_48 
+ bl[46] br[46] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_49 
+ bl[47] br[47] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_50 
+ bl[48] br[48] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_51 
+ bl[49] br[49] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_52 
+ bl[50] br[50] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_53 
+ bl[51] br[51] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_54 
+ bl[52] br[52] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_55 
+ bl[53] br[53] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_56 
+ bl[54] br[54] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_57 
+ bl[55] br[55] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_58 
+ bl[56] br[56] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_59 
+ bl[57] br[57] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_60 
+ bl[58] br[58] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_61 
+ bl[59] br[59] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_62 
+ bl[60] br[60] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_63 
+ bl[61] br[61] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_64 
+ bl[62] br[62] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_65 
+ bl[63] br[63] vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_66 
+ vdd vdd vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_382_67 
+ vdd vdd vdd vss wl[380] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_0 
+ vdd vdd vss vdd vpb vnb wl[381] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_383_1 
+ rbl rbr vss vdd vpb vnb wl[381] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_383_2 
+ bl[0] br[0] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_3 
+ bl[1] br[1] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_4 
+ bl[2] br[2] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_5 
+ bl[3] br[3] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_6 
+ bl[4] br[4] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_7 
+ bl[5] br[5] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_8 
+ bl[6] br[6] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_9 
+ bl[7] br[7] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_10 
+ bl[8] br[8] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_11 
+ bl[9] br[9] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_12 
+ bl[10] br[10] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_13 
+ bl[11] br[11] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_14 
+ bl[12] br[12] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_15 
+ bl[13] br[13] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_16 
+ bl[14] br[14] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_17 
+ bl[15] br[15] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_18 
+ bl[16] br[16] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_19 
+ bl[17] br[17] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_20 
+ bl[18] br[18] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_21 
+ bl[19] br[19] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_22 
+ bl[20] br[20] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_23 
+ bl[21] br[21] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_24 
+ bl[22] br[22] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_25 
+ bl[23] br[23] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_26 
+ bl[24] br[24] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_27 
+ bl[25] br[25] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_28 
+ bl[26] br[26] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_29 
+ bl[27] br[27] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_30 
+ bl[28] br[28] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_31 
+ bl[29] br[29] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_32 
+ bl[30] br[30] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_33 
+ bl[31] br[31] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_34 
+ bl[32] br[32] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_35 
+ bl[33] br[33] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_36 
+ bl[34] br[34] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_37 
+ bl[35] br[35] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_38 
+ bl[36] br[36] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_39 
+ bl[37] br[37] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_40 
+ bl[38] br[38] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_41 
+ bl[39] br[39] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_42 
+ bl[40] br[40] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_43 
+ bl[41] br[41] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_44 
+ bl[42] br[42] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_45 
+ bl[43] br[43] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_46 
+ bl[44] br[44] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_47 
+ bl[45] br[45] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_48 
+ bl[46] br[46] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_49 
+ bl[47] br[47] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_50 
+ bl[48] br[48] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_51 
+ bl[49] br[49] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_52 
+ bl[50] br[50] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_53 
+ bl[51] br[51] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_54 
+ bl[52] br[52] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_55 
+ bl[53] br[53] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_56 
+ bl[54] br[54] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_57 
+ bl[55] br[55] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_58 
+ bl[56] br[56] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_59 
+ bl[57] br[57] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_60 
+ bl[58] br[58] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_61 
+ bl[59] br[59] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_62 
+ bl[60] br[60] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_63 
+ bl[61] br[61] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_64 
+ bl[62] br[62] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_65 
+ bl[63] br[63] vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_66 
+ vdd vdd vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_383_67 
+ vdd vdd vdd vss wl[381] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_0 
+ vdd vdd vss vdd vpb vnb wl[382] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_384_1 
+ rbl rbr vss vdd vpb vnb wl[382] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_384_2 
+ bl[0] br[0] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_3 
+ bl[1] br[1] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_4 
+ bl[2] br[2] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_5 
+ bl[3] br[3] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_6 
+ bl[4] br[4] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_7 
+ bl[5] br[5] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_8 
+ bl[6] br[6] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_9 
+ bl[7] br[7] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_10 
+ bl[8] br[8] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_11 
+ bl[9] br[9] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_12 
+ bl[10] br[10] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_13 
+ bl[11] br[11] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_14 
+ bl[12] br[12] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_15 
+ bl[13] br[13] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_16 
+ bl[14] br[14] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_17 
+ bl[15] br[15] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_18 
+ bl[16] br[16] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_19 
+ bl[17] br[17] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_20 
+ bl[18] br[18] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_21 
+ bl[19] br[19] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_22 
+ bl[20] br[20] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_23 
+ bl[21] br[21] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_24 
+ bl[22] br[22] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_25 
+ bl[23] br[23] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_26 
+ bl[24] br[24] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_27 
+ bl[25] br[25] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_28 
+ bl[26] br[26] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_29 
+ bl[27] br[27] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_30 
+ bl[28] br[28] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_31 
+ bl[29] br[29] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_32 
+ bl[30] br[30] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_33 
+ bl[31] br[31] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_34 
+ bl[32] br[32] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_35 
+ bl[33] br[33] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_36 
+ bl[34] br[34] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_37 
+ bl[35] br[35] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_38 
+ bl[36] br[36] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_39 
+ bl[37] br[37] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_40 
+ bl[38] br[38] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_41 
+ bl[39] br[39] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_42 
+ bl[40] br[40] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_43 
+ bl[41] br[41] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_44 
+ bl[42] br[42] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_45 
+ bl[43] br[43] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_46 
+ bl[44] br[44] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_47 
+ bl[45] br[45] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_48 
+ bl[46] br[46] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_49 
+ bl[47] br[47] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_50 
+ bl[48] br[48] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_51 
+ bl[49] br[49] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_52 
+ bl[50] br[50] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_53 
+ bl[51] br[51] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_54 
+ bl[52] br[52] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_55 
+ bl[53] br[53] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_56 
+ bl[54] br[54] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_57 
+ bl[55] br[55] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_58 
+ bl[56] br[56] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_59 
+ bl[57] br[57] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_60 
+ bl[58] br[58] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_61 
+ bl[59] br[59] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_62 
+ bl[60] br[60] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_63 
+ bl[61] br[61] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_64 
+ bl[62] br[62] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_65 
+ bl[63] br[63] vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_66 
+ vdd vdd vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_384_67 
+ vdd vdd vdd vss wl[382] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_0 
+ vdd vdd vss vdd vpb vnb wl[383] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_385_1 
+ rbl rbr vss vdd vpb vnb wl[383] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_385_2 
+ bl[0] br[0] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_3 
+ bl[1] br[1] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_4 
+ bl[2] br[2] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_5 
+ bl[3] br[3] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_6 
+ bl[4] br[4] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_7 
+ bl[5] br[5] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_8 
+ bl[6] br[6] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_9 
+ bl[7] br[7] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_10 
+ bl[8] br[8] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_11 
+ bl[9] br[9] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_12 
+ bl[10] br[10] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_13 
+ bl[11] br[11] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_14 
+ bl[12] br[12] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_15 
+ bl[13] br[13] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_16 
+ bl[14] br[14] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_17 
+ bl[15] br[15] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_18 
+ bl[16] br[16] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_19 
+ bl[17] br[17] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_20 
+ bl[18] br[18] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_21 
+ bl[19] br[19] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_22 
+ bl[20] br[20] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_23 
+ bl[21] br[21] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_24 
+ bl[22] br[22] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_25 
+ bl[23] br[23] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_26 
+ bl[24] br[24] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_27 
+ bl[25] br[25] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_28 
+ bl[26] br[26] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_29 
+ bl[27] br[27] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_30 
+ bl[28] br[28] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_31 
+ bl[29] br[29] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_32 
+ bl[30] br[30] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_33 
+ bl[31] br[31] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_34 
+ bl[32] br[32] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_35 
+ bl[33] br[33] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_36 
+ bl[34] br[34] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_37 
+ bl[35] br[35] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_38 
+ bl[36] br[36] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_39 
+ bl[37] br[37] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_40 
+ bl[38] br[38] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_41 
+ bl[39] br[39] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_42 
+ bl[40] br[40] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_43 
+ bl[41] br[41] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_44 
+ bl[42] br[42] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_45 
+ bl[43] br[43] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_46 
+ bl[44] br[44] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_47 
+ bl[45] br[45] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_48 
+ bl[46] br[46] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_49 
+ bl[47] br[47] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_50 
+ bl[48] br[48] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_51 
+ bl[49] br[49] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_52 
+ bl[50] br[50] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_53 
+ bl[51] br[51] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_54 
+ bl[52] br[52] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_55 
+ bl[53] br[53] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_56 
+ bl[54] br[54] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_57 
+ bl[55] br[55] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_58 
+ bl[56] br[56] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_59 
+ bl[57] br[57] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_60 
+ bl[58] br[58] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_61 
+ bl[59] br[59] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_62 
+ bl[60] br[60] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_63 
+ bl[61] br[61] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_64 
+ bl[62] br[62] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_65 
+ bl[63] br[63] vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_66 
+ vdd vdd vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_385_67 
+ vdd vdd vdd vss wl[383] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_0 
+ vdd vdd vss vdd vpb vnb wl[384] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_386_1 
+ rbl rbr vss vdd vpb vnb wl[384] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_386_2 
+ bl[0] br[0] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_3 
+ bl[1] br[1] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_4 
+ bl[2] br[2] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_5 
+ bl[3] br[3] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_6 
+ bl[4] br[4] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_7 
+ bl[5] br[5] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_8 
+ bl[6] br[6] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_9 
+ bl[7] br[7] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_10 
+ bl[8] br[8] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_11 
+ bl[9] br[9] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_12 
+ bl[10] br[10] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_13 
+ bl[11] br[11] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_14 
+ bl[12] br[12] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_15 
+ bl[13] br[13] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_16 
+ bl[14] br[14] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_17 
+ bl[15] br[15] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_18 
+ bl[16] br[16] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_19 
+ bl[17] br[17] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_20 
+ bl[18] br[18] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_21 
+ bl[19] br[19] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_22 
+ bl[20] br[20] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_23 
+ bl[21] br[21] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_24 
+ bl[22] br[22] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_25 
+ bl[23] br[23] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_26 
+ bl[24] br[24] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_27 
+ bl[25] br[25] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_28 
+ bl[26] br[26] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_29 
+ bl[27] br[27] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_30 
+ bl[28] br[28] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_31 
+ bl[29] br[29] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_32 
+ bl[30] br[30] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_33 
+ bl[31] br[31] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_34 
+ bl[32] br[32] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_35 
+ bl[33] br[33] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_36 
+ bl[34] br[34] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_37 
+ bl[35] br[35] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_38 
+ bl[36] br[36] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_39 
+ bl[37] br[37] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_40 
+ bl[38] br[38] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_41 
+ bl[39] br[39] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_42 
+ bl[40] br[40] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_43 
+ bl[41] br[41] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_44 
+ bl[42] br[42] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_45 
+ bl[43] br[43] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_46 
+ bl[44] br[44] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_47 
+ bl[45] br[45] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_48 
+ bl[46] br[46] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_49 
+ bl[47] br[47] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_50 
+ bl[48] br[48] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_51 
+ bl[49] br[49] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_52 
+ bl[50] br[50] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_53 
+ bl[51] br[51] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_54 
+ bl[52] br[52] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_55 
+ bl[53] br[53] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_56 
+ bl[54] br[54] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_57 
+ bl[55] br[55] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_58 
+ bl[56] br[56] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_59 
+ bl[57] br[57] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_60 
+ bl[58] br[58] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_61 
+ bl[59] br[59] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_62 
+ bl[60] br[60] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_63 
+ bl[61] br[61] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_64 
+ bl[62] br[62] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_65 
+ bl[63] br[63] vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_66 
+ vdd vdd vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_386_67 
+ vdd vdd vdd vss wl[384] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_0 
+ vdd vdd vss vdd vpb vnb wl[385] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_387_1 
+ rbl rbr vss vdd vpb vnb wl[385] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_387_2 
+ bl[0] br[0] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_3 
+ bl[1] br[1] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_4 
+ bl[2] br[2] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_5 
+ bl[3] br[3] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_6 
+ bl[4] br[4] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_7 
+ bl[5] br[5] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_8 
+ bl[6] br[6] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_9 
+ bl[7] br[7] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_10 
+ bl[8] br[8] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_11 
+ bl[9] br[9] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_12 
+ bl[10] br[10] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_13 
+ bl[11] br[11] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_14 
+ bl[12] br[12] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_15 
+ bl[13] br[13] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_16 
+ bl[14] br[14] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_17 
+ bl[15] br[15] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_18 
+ bl[16] br[16] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_19 
+ bl[17] br[17] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_20 
+ bl[18] br[18] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_21 
+ bl[19] br[19] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_22 
+ bl[20] br[20] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_23 
+ bl[21] br[21] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_24 
+ bl[22] br[22] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_25 
+ bl[23] br[23] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_26 
+ bl[24] br[24] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_27 
+ bl[25] br[25] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_28 
+ bl[26] br[26] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_29 
+ bl[27] br[27] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_30 
+ bl[28] br[28] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_31 
+ bl[29] br[29] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_32 
+ bl[30] br[30] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_33 
+ bl[31] br[31] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_34 
+ bl[32] br[32] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_35 
+ bl[33] br[33] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_36 
+ bl[34] br[34] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_37 
+ bl[35] br[35] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_38 
+ bl[36] br[36] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_39 
+ bl[37] br[37] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_40 
+ bl[38] br[38] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_41 
+ bl[39] br[39] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_42 
+ bl[40] br[40] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_43 
+ bl[41] br[41] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_44 
+ bl[42] br[42] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_45 
+ bl[43] br[43] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_46 
+ bl[44] br[44] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_47 
+ bl[45] br[45] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_48 
+ bl[46] br[46] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_49 
+ bl[47] br[47] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_50 
+ bl[48] br[48] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_51 
+ bl[49] br[49] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_52 
+ bl[50] br[50] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_53 
+ bl[51] br[51] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_54 
+ bl[52] br[52] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_55 
+ bl[53] br[53] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_56 
+ bl[54] br[54] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_57 
+ bl[55] br[55] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_58 
+ bl[56] br[56] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_59 
+ bl[57] br[57] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_60 
+ bl[58] br[58] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_61 
+ bl[59] br[59] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_62 
+ bl[60] br[60] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_63 
+ bl[61] br[61] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_64 
+ bl[62] br[62] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_65 
+ bl[63] br[63] vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_66 
+ vdd vdd vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_387_67 
+ vdd vdd vdd vss wl[385] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_0 
+ vdd vdd vss vdd vpb vnb wl[386] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_388_1 
+ rbl rbr vss vdd vpb vnb wl[386] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_388_2 
+ bl[0] br[0] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_3 
+ bl[1] br[1] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_4 
+ bl[2] br[2] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_5 
+ bl[3] br[3] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_6 
+ bl[4] br[4] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_7 
+ bl[5] br[5] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_8 
+ bl[6] br[6] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_9 
+ bl[7] br[7] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_10 
+ bl[8] br[8] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_11 
+ bl[9] br[9] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_12 
+ bl[10] br[10] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_13 
+ bl[11] br[11] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_14 
+ bl[12] br[12] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_15 
+ bl[13] br[13] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_16 
+ bl[14] br[14] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_17 
+ bl[15] br[15] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_18 
+ bl[16] br[16] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_19 
+ bl[17] br[17] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_20 
+ bl[18] br[18] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_21 
+ bl[19] br[19] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_22 
+ bl[20] br[20] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_23 
+ bl[21] br[21] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_24 
+ bl[22] br[22] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_25 
+ bl[23] br[23] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_26 
+ bl[24] br[24] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_27 
+ bl[25] br[25] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_28 
+ bl[26] br[26] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_29 
+ bl[27] br[27] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_30 
+ bl[28] br[28] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_31 
+ bl[29] br[29] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_32 
+ bl[30] br[30] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_33 
+ bl[31] br[31] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_34 
+ bl[32] br[32] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_35 
+ bl[33] br[33] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_36 
+ bl[34] br[34] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_37 
+ bl[35] br[35] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_38 
+ bl[36] br[36] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_39 
+ bl[37] br[37] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_40 
+ bl[38] br[38] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_41 
+ bl[39] br[39] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_42 
+ bl[40] br[40] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_43 
+ bl[41] br[41] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_44 
+ bl[42] br[42] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_45 
+ bl[43] br[43] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_46 
+ bl[44] br[44] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_47 
+ bl[45] br[45] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_48 
+ bl[46] br[46] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_49 
+ bl[47] br[47] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_50 
+ bl[48] br[48] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_51 
+ bl[49] br[49] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_52 
+ bl[50] br[50] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_53 
+ bl[51] br[51] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_54 
+ bl[52] br[52] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_55 
+ bl[53] br[53] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_56 
+ bl[54] br[54] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_57 
+ bl[55] br[55] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_58 
+ bl[56] br[56] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_59 
+ bl[57] br[57] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_60 
+ bl[58] br[58] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_61 
+ bl[59] br[59] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_62 
+ bl[60] br[60] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_63 
+ bl[61] br[61] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_64 
+ bl[62] br[62] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_65 
+ bl[63] br[63] vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_66 
+ vdd vdd vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_388_67 
+ vdd vdd vdd vss wl[386] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_0 
+ vdd vdd vss vdd vpb vnb wl[387] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_389_1 
+ rbl rbr vss vdd vpb vnb wl[387] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_389_2 
+ bl[0] br[0] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_3 
+ bl[1] br[1] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_4 
+ bl[2] br[2] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_5 
+ bl[3] br[3] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_6 
+ bl[4] br[4] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_7 
+ bl[5] br[5] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_8 
+ bl[6] br[6] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_9 
+ bl[7] br[7] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_10 
+ bl[8] br[8] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_11 
+ bl[9] br[9] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_12 
+ bl[10] br[10] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_13 
+ bl[11] br[11] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_14 
+ bl[12] br[12] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_15 
+ bl[13] br[13] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_16 
+ bl[14] br[14] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_17 
+ bl[15] br[15] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_18 
+ bl[16] br[16] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_19 
+ bl[17] br[17] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_20 
+ bl[18] br[18] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_21 
+ bl[19] br[19] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_22 
+ bl[20] br[20] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_23 
+ bl[21] br[21] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_24 
+ bl[22] br[22] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_25 
+ bl[23] br[23] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_26 
+ bl[24] br[24] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_27 
+ bl[25] br[25] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_28 
+ bl[26] br[26] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_29 
+ bl[27] br[27] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_30 
+ bl[28] br[28] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_31 
+ bl[29] br[29] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_32 
+ bl[30] br[30] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_33 
+ bl[31] br[31] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_34 
+ bl[32] br[32] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_35 
+ bl[33] br[33] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_36 
+ bl[34] br[34] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_37 
+ bl[35] br[35] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_38 
+ bl[36] br[36] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_39 
+ bl[37] br[37] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_40 
+ bl[38] br[38] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_41 
+ bl[39] br[39] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_42 
+ bl[40] br[40] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_43 
+ bl[41] br[41] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_44 
+ bl[42] br[42] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_45 
+ bl[43] br[43] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_46 
+ bl[44] br[44] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_47 
+ bl[45] br[45] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_48 
+ bl[46] br[46] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_49 
+ bl[47] br[47] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_50 
+ bl[48] br[48] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_51 
+ bl[49] br[49] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_52 
+ bl[50] br[50] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_53 
+ bl[51] br[51] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_54 
+ bl[52] br[52] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_55 
+ bl[53] br[53] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_56 
+ bl[54] br[54] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_57 
+ bl[55] br[55] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_58 
+ bl[56] br[56] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_59 
+ bl[57] br[57] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_60 
+ bl[58] br[58] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_61 
+ bl[59] br[59] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_62 
+ bl[60] br[60] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_63 
+ bl[61] br[61] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_64 
+ bl[62] br[62] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_65 
+ bl[63] br[63] vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_66 
+ vdd vdd vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_389_67 
+ vdd vdd vdd vss wl[387] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_0 
+ vdd vdd vss vdd vpb vnb wl[388] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_390_1 
+ rbl rbr vss vdd vpb vnb wl[388] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_390_2 
+ bl[0] br[0] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_3 
+ bl[1] br[1] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_4 
+ bl[2] br[2] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_5 
+ bl[3] br[3] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_6 
+ bl[4] br[4] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_7 
+ bl[5] br[5] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_8 
+ bl[6] br[6] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_9 
+ bl[7] br[7] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_10 
+ bl[8] br[8] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_11 
+ bl[9] br[9] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_12 
+ bl[10] br[10] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_13 
+ bl[11] br[11] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_14 
+ bl[12] br[12] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_15 
+ bl[13] br[13] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_16 
+ bl[14] br[14] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_17 
+ bl[15] br[15] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_18 
+ bl[16] br[16] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_19 
+ bl[17] br[17] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_20 
+ bl[18] br[18] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_21 
+ bl[19] br[19] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_22 
+ bl[20] br[20] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_23 
+ bl[21] br[21] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_24 
+ bl[22] br[22] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_25 
+ bl[23] br[23] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_26 
+ bl[24] br[24] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_27 
+ bl[25] br[25] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_28 
+ bl[26] br[26] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_29 
+ bl[27] br[27] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_30 
+ bl[28] br[28] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_31 
+ bl[29] br[29] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_32 
+ bl[30] br[30] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_33 
+ bl[31] br[31] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_34 
+ bl[32] br[32] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_35 
+ bl[33] br[33] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_36 
+ bl[34] br[34] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_37 
+ bl[35] br[35] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_38 
+ bl[36] br[36] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_39 
+ bl[37] br[37] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_40 
+ bl[38] br[38] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_41 
+ bl[39] br[39] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_42 
+ bl[40] br[40] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_43 
+ bl[41] br[41] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_44 
+ bl[42] br[42] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_45 
+ bl[43] br[43] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_46 
+ bl[44] br[44] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_47 
+ bl[45] br[45] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_48 
+ bl[46] br[46] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_49 
+ bl[47] br[47] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_50 
+ bl[48] br[48] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_51 
+ bl[49] br[49] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_52 
+ bl[50] br[50] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_53 
+ bl[51] br[51] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_54 
+ bl[52] br[52] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_55 
+ bl[53] br[53] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_56 
+ bl[54] br[54] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_57 
+ bl[55] br[55] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_58 
+ bl[56] br[56] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_59 
+ bl[57] br[57] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_60 
+ bl[58] br[58] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_61 
+ bl[59] br[59] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_62 
+ bl[60] br[60] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_63 
+ bl[61] br[61] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_64 
+ bl[62] br[62] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_65 
+ bl[63] br[63] vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_66 
+ vdd vdd vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_390_67 
+ vdd vdd vdd vss wl[388] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_0 
+ vdd vdd vss vdd vpb vnb wl[389] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_391_1 
+ rbl rbr vss vdd vpb vnb wl[389] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_391_2 
+ bl[0] br[0] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_3 
+ bl[1] br[1] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_4 
+ bl[2] br[2] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_5 
+ bl[3] br[3] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_6 
+ bl[4] br[4] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_7 
+ bl[5] br[5] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_8 
+ bl[6] br[6] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_9 
+ bl[7] br[7] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_10 
+ bl[8] br[8] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_11 
+ bl[9] br[9] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_12 
+ bl[10] br[10] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_13 
+ bl[11] br[11] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_14 
+ bl[12] br[12] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_15 
+ bl[13] br[13] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_16 
+ bl[14] br[14] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_17 
+ bl[15] br[15] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_18 
+ bl[16] br[16] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_19 
+ bl[17] br[17] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_20 
+ bl[18] br[18] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_21 
+ bl[19] br[19] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_22 
+ bl[20] br[20] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_23 
+ bl[21] br[21] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_24 
+ bl[22] br[22] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_25 
+ bl[23] br[23] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_26 
+ bl[24] br[24] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_27 
+ bl[25] br[25] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_28 
+ bl[26] br[26] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_29 
+ bl[27] br[27] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_30 
+ bl[28] br[28] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_31 
+ bl[29] br[29] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_32 
+ bl[30] br[30] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_33 
+ bl[31] br[31] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_34 
+ bl[32] br[32] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_35 
+ bl[33] br[33] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_36 
+ bl[34] br[34] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_37 
+ bl[35] br[35] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_38 
+ bl[36] br[36] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_39 
+ bl[37] br[37] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_40 
+ bl[38] br[38] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_41 
+ bl[39] br[39] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_42 
+ bl[40] br[40] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_43 
+ bl[41] br[41] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_44 
+ bl[42] br[42] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_45 
+ bl[43] br[43] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_46 
+ bl[44] br[44] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_47 
+ bl[45] br[45] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_48 
+ bl[46] br[46] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_49 
+ bl[47] br[47] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_50 
+ bl[48] br[48] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_51 
+ bl[49] br[49] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_52 
+ bl[50] br[50] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_53 
+ bl[51] br[51] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_54 
+ bl[52] br[52] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_55 
+ bl[53] br[53] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_56 
+ bl[54] br[54] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_57 
+ bl[55] br[55] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_58 
+ bl[56] br[56] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_59 
+ bl[57] br[57] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_60 
+ bl[58] br[58] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_61 
+ bl[59] br[59] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_62 
+ bl[60] br[60] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_63 
+ bl[61] br[61] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_64 
+ bl[62] br[62] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_65 
+ bl[63] br[63] vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_66 
+ vdd vdd vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_391_67 
+ vdd vdd vdd vss wl[389] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_0 
+ vdd vdd vss vdd vpb vnb wl[390] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_392_1 
+ rbl rbr vss vdd vpb vnb wl[390] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_392_2 
+ bl[0] br[0] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_3 
+ bl[1] br[1] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_4 
+ bl[2] br[2] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_5 
+ bl[3] br[3] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_6 
+ bl[4] br[4] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_7 
+ bl[5] br[5] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_8 
+ bl[6] br[6] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_9 
+ bl[7] br[7] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_10 
+ bl[8] br[8] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_11 
+ bl[9] br[9] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_12 
+ bl[10] br[10] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_13 
+ bl[11] br[11] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_14 
+ bl[12] br[12] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_15 
+ bl[13] br[13] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_16 
+ bl[14] br[14] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_17 
+ bl[15] br[15] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_18 
+ bl[16] br[16] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_19 
+ bl[17] br[17] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_20 
+ bl[18] br[18] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_21 
+ bl[19] br[19] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_22 
+ bl[20] br[20] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_23 
+ bl[21] br[21] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_24 
+ bl[22] br[22] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_25 
+ bl[23] br[23] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_26 
+ bl[24] br[24] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_27 
+ bl[25] br[25] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_28 
+ bl[26] br[26] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_29 
+ bl[27] br[27] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_30 
+ bl[28] br[28] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_31 
+ bl[29] br[29] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_32 
+ bl[30] br[30] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_33 
+ bl[31] br[31] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_34 
+ bl[32] br[32] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_35 
+ bl[33] br[33] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_36 
+ bl[34] br[34] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_37 
+ bl[35] br[35] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_38 
+ bl[36] br[36] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_39 
+ bl[37] br[37] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_40 
+ bl[38] br[38] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_41 
+ bl[39] br[39] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_42 
+ bl[40] br[40] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_43 
+ bl[41] br[41] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_44 
+ bl[42] br[42] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_45 
+ bl[43] br[43] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_46 
+ bl[44] br[44] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_47 
+ bl[45] br[45] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_48 
+ bl[46] br[46] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_49 
+ bl[47] br[47] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_50 
+ bl[48] br[48] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_51 
+ bl[49] br[49] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_52 
+ bl[50] br[50] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_53 
+ bl[51] br[51] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_54 
+ bl[52] br[52] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_55 
+ bl[53] br[53] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_56 
+ bl[54] br[54] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_57 
+ bl[55] br[55] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_58 
+ bl[56] br[56] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_59 
+ bl[57] br[57] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_60 
+ bl[58] br[58] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_61 
+ bl[59] br[59] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_62 
+ bl[60] br[60] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_63 
+ bl[61] br[61] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_64 
+ bl[62] br[62] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_65 
+ bl[63] br[63] vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_66 
+ vdd vdd vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_392_67 
+ vdd vdd vdd vss wl[390] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_0 
+ vdd vdd vss vdd vpb vnb wl[391] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_393_1 
+ rbl rbr vss vdd vpb vnb wl[391] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_393_2 
+ bl[0] br[0] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_3 
+ bl[1] br[1] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_4 
+ bl[2] br[2] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_5 
+ bl[3] br[3] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_6 
+ bl[4] br[4] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_7 
+ bl[5] br[5] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_8 
+ bl[6] br[6] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_9 
+ bl[7] br[7] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_10 
+ bl[8] br[8] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_11 
+ bl[9] br[9] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_12 
+ bl[10] br[10] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_13 
+ bl[11] br[11] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_14 
+ bl[12] br[12] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_15 
+ bl[13] br[13] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_16 
+ bl[14] br[14] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_17 
+ bl[15] br[15] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_18 
+ bl[16] br[16] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_19 
+ bl[17] br[17] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_20 
+ bl[18] br[18] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_21 
+ bl[19] br[19] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_22 
+ bl[20] br[20] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_23 
+ bl[21] br[21] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_24 
+ bl[22] br[22] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_25 
+ bl[23] br[23] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_26 
+ bl[24] br[24] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_27 
+ bl[25] br[25] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_28 
+ bl[26] br[26] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_29 
+ bl[27] br[27] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_30 
+ bl[28] br[28] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_31 
+ bl[29] br[29] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_32 
+ bl[30] br[30] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_33 
+ bl[31] br[31] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_34 
+ bl[32] br[32] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_35 
+ bl[33] br[33] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_36 
+ bl[34] br[34] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_37 
+ bl[35] br[35] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_38 
+ bl[36] br[36] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_39 
+ bl[37] br[37] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_40 
+ bl[38] br[38] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_41 
+ bl[39] br[39] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_42 
+ bl[40] br[40] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_43 
+ bl[41] br[41] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_44 
+ bl[42] br[42] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_45 
+ bl[43] br[43] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_46 
+ bl[44] br[44] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_47 
+ bl[45] br[45] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_48 
+ bl[46] br[46] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_49 
+ bl[47] br[47] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_50 
+ bl[48] br[48] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_51 
+ bl[49] br[49] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_52 
+ bl[50] br[50] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_53 
+ bl[51] br[51] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_54 
+ bl[52] br[52] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_55 
+ bl[53] br[53] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_56 
+ bl[54] br[54] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_57 
+ bl[55] br[55] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_58 
+ bl[56] br[56] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_59 
+ bl[57] br[57] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_60 
+ bl[58] br[58] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_61 
+ bl[59] br[59] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_62 
+ bl[60] br[60] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_63 
+ bl[61] br[61] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_64 
+ bl[62] br[62] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_65 
+ bl[63] br[63] vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_66 
+ vdd vdd vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_393_67 
+ vdd vdd vdd vss wl[391] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_0 
+ vdd vdd vss vdd vpb vnb wl[392] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_394_1 
+ rbl rbr vss vdd vpb vnb wl[392] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_394_2 
+ bl[0] br[0] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_3 
+ bl[1] br[1] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_4 
+ bl[2] br[2] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_5 
+ bl[3] br[3] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_6 
+ bl[4] br[4] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_7 
+ bl[5] br[5] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_8 
+ bl[6] br[6] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_9 
+ bl[7] br[7] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_10 
+ bl[8] br[8] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_11 
+ bl[9] br[9] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_12 
+ bl[10] br[10] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_13 
+ bl[11] br[11] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_14 
+ bl[12] br[12] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_15 
+ bl[13] br[13] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_16 
+ bl[14] br[14] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_17 
+ bl[15] br[15] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_18 
+ bl[16] br[16] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_19 
+ bl[17] br[17] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_20 
+ bl[18] br[18] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_21 
+ bl[19] br[19] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_22 
+ bl[20] br[20] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_23 
+ bl[21] br[21] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_24 
+ bl[22] br[22] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_25 
+ bl[23] br[23] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_26 
+ bl[24] br[24] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_27 
+ bl[25] br[25] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_28 
+ bl[26] br[26] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_29 
+ bl[27] br[27] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_30 
+ bl[28] br[28] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_31 
+ bl[29] br[29] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_32 
+ bl[30] br[30] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_33 
+ bl[31] br[31] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_34 
+ bl[32] br[32] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_35 
+ bl[33] br[33] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_36 
+ bl[34] br[34] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_37 
+ bl[35] br[35] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_38 
+ bl[36] br[36] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_39 
+ bl[37] br[37] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_40 
+ bl[38] br[38] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_41 
+ bl[39] br[39] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_42 
+ bl[40] br[40] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_43 
+ bl[41] br[41] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_44 
+ bl[42] br[42] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_45 
+ bl[43] br[43] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_46 
+ bl[44] br[44] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_47 
+ bl[45] br[45] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_48 
+ bl[46] br[46] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_49 
+ bl[47] br[47] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_50 
+ bl[48] br[48] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_51 
+ bl[49] br[49] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_52 
+ bl[50] br[50] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_53 
+ bl[51] br[51] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_54 
+ bl[52] br[52] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_55 
+ bl[53] br[53] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_56 
+ bl[54] br[54] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_57 
+ bl[55] br[55] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_58 
+ bl[56] br[56] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_59 
+ bl[57] br[57] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_60 
+ bl[58] br[58] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_61 
+ bl[59] br[59] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_62 
+ bl[60] br[60] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_63 
+ bl[61] br[61] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_64 
+ bl[62] br[62] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_65 
+ bl[63] br[63] vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_66 
+ vdd vdd vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_394_67 
+ vdd vdd vdd vss wl[392] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_0 
+ vdd vdd vss vdd vpb vnb wl[393] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_395_1 
+ rbl rbr vss vdd vpb vnb wl[393] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_395_2 
+ bl[0] br[0] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_3 
+ bl[1] br[1] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_4 
+ bl[2] br[2] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_5 
+ bl[3] br[3] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_6 
+ bl[4] br[4] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_7 
+ bl[5] br[5] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_8 
+ bl[6] br[6] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_9 
+ bl[7] br[7] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_10 
+ bl[8] br[8] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_11 
+ bl[9] br[9] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_12 
+ bl[10] br[10] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_13 
+ bl[11] br[11] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_14 
+ bl[12] br[12] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_15 
+ bl[13] br[13] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_16 
+ bl[14] br[14] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_17 
+ bl[15] br[15] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_18 
+ bl[16] br[16] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_19 
+ bl[17] br[17] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_20 
+ bl[18] br[18] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_21 
+ bl[19] br[19] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_22 
+ bl[20] br[20] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_23 
+ bl[21] br[21] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_24 
+ bl[22] br[22] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_25 
+ bl[23] br[23] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_26 
+ bl[24] br[24] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_27 
+ bl[25] br[25] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_28 
+ bl[26] br[26] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_29 
+ bl[27] br[27] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_30 
+ bl[28] br[28] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_31 
+ bl[29] br[29] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_32 
+ bl[30] br[30] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_33 
+ bl[31] br[31] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_34 
+ bl[32] br[32] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_35 
+ bl[33] br[33] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_36 
+ bl[34] br[34] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_37 
+ bl[35] br[35] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_38 
+ bl[36] br[36] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_39 
+ bl[37] br[37] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_40 
+ bl[38] br[38] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_41 
+ bl[39] br[39] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_42 
+ bl[40] br[40] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_43 
+ bl[41] br[41] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_44 
+ bl[42] br[42] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_45 
+ bl[43] br[43] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_46 
+ bl[44] br[44] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_47 
+ bl[45] br[45] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_48 
+ bl[46] br[46] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_49 
+ bl[47] br[47] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_50 
+ bl[48] br[48] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_51 
+ bl[49] br[49] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_52 
+ bl[50] br[50] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_53 
+ bl[51] br[51] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_54 
+ bl[52] br[52] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_55 
+ bl[53] br[53] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_56 
+ bl[54] br[54] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_57 
+ bl[55] br[55] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_58 
+ bl[56] br[56] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_59 
+ bl[57] br[57] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_60 
+ bl[58] br[58] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_61 
+ bl[59] br[59] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_62 
+ bl[60] br[60] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_63 
+ bl[61] br[61] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_64 
+ bl[62] br[62] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_65 
+ bl[63] br[63] vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_66 
+ vdd vdd vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_395_67 
+ vdd vdd vdd vss wl[393] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_0 
+ vdd vdd vss vdd vpb vnb wl[394] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_396_1 
+ rbl rbr vss vdd vpb vnb wl[394] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_396_2 
+ bl[0] br[0] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_3 
+ bl[1] br[1] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_4 
+ bl[2] br[2] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_5 
+ bl[3] br[3] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_6 
+ bl[4] br[4] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_7 
+ bl[5] br[5] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_8 
+ bl[6] br[6] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_9 
+ bl[7] br[7] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_10 
+ bl[8] br[8] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_11 
+ bl[9] br[9] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_12 
+ bl[10] br[10] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_13 
+ bl[11] br[11] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_14 
+ bl[12] br[12] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_15 
+ bl[13] br[13] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_16 
+ bl[14] br[14] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_17 
+ bl[15] br[15] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_18 
+ bl[16] br[16] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_19 
+ bl[17] br[17] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_20 
+ bl[18] br[18] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_21 
+ bl[19] br[19] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_22 
+ bl[20] br[20] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_23 
+ bl[21] br[21] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_24 
+ bl[22] br[22] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_25 
+ bl[23] br[23] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_26 
+ bl[24] br[24] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_27 
+ bl[25] br[25] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_28 
+ bl[26] br[26] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_29 
+ bl[27] br[27] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_30 
+ bl[28] br[28] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_31 
+ bl[29] br[29] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_32 
+ bl[30] br[30] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_33 
+ bl[31] br[31] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_34 
+ bl[32] br[32] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_35 
+ bl[33] br[33] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_36 
+ bl[34] br[34] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_37 
+ bl[35] br[35] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_38 
+ bl[36] br[36] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_39 
+ bl[37] br[37] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_40 
+ bl[38] br[38] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_41 
+ bl[39] br[39] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_42 
+ bl[40] br[40] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_43 
+ bl[41] br[41] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_44 
+ bl[42] br[42] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_45 
+ bl[43] br[43] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_46 
+ bl[44] br[44] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_47 
+ bl[45] br[45] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_48 
+ bl[46] br[46] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_49 
+ bl[47] br[47] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_50 
+ bl[48] br[48] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_51 
+ bl[49] br[49] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_52 
+ bl[50] br[50] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_53 
+ bl[51] br[51] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_54 
+ bl[52] br[52] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_55 
+ bl[53] br[53] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_56 
+ bl[54] br[54] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_57 
+ bl[55] br[55] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_58 
+ bl[56] br[56] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_59 
+ bl[57] br[57] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_60 
+ bl[58] br[58] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_61 
+ bl[59] br[59] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_62 
+ bl[60] br[60] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_63 
+ bl[61] br[61] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_64 
+ bl[62] br[62] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_65 
+ bl[63] br[63] vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_66 
+ vdd vdd vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_396_67 
+ vdd vdd vdd vss wl[394] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_0 
+ vdd vdd vss vdd vpb vnb wl[395] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_397_1 
+ rbl rbr vss vdd vpb vnb wl[395] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_397_2 
+ bl[0] br[0] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_3 
+ bl[1] br[1] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_4 
+ bl[2] br[2] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_5 
+ bl[3] br[3] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_6 
+ bl[4] br[4] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_7 
+ bl[5] br[5] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_8 
+ bl[6] br[6] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_9 
+ bl[7] br[7] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_10 
+ bl[8] br[8] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_11 
+ bl[9] br[9] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_12 
+ bl[10] br[10] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_13 
+ bl[11] br[11] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_14 
+ bl[12] br[12] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_15 
+ bl[13] br[13] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_16 
+ bl[14] br[14] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_17 
+ bl[15] br[15] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_18 
+ bl[16] br[16] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_19 
+ bl[17] br[17] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_20 
+ bl[18] br[18] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_21 
+ bl[19] br[19] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_22 
+ bl[20] br[20] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_23 
+ bl[21] br[21] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_24 
+ bl[22] br[22] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_25 
+ bl[23] br[23] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_26 
+ bl[24] br[24] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_27 
+ bl[25] br[25] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_28 
+ bl[26] br[26] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_29 
+ bl[27] br[27] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_30 
+ bl[28] br[28] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_31 
+ bl[29] br[29] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_32 
+ bl[30] br[30] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_33 
+ bl[31] br[31] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_34 
+ bl[32] br[32] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_35 
+ bl[33] br[33] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_36 
+ bl[34] br[34] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_37 
+ bl[35] br[35] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_38 
+ bl[36] br[36] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_39 
+ bl[37] br[37] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_40 
+ bl[38] br[38] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_41 
+ bl[39] br[39] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_42 
+ bl[40] br[40] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_43 
+ bl[41] br[41] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_44 
+ bl[42] br[42] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_45 
+ bl[43] br[43] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_46 
+ bl[44] br[44] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_47 
+ bl[45] br[45] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_48 
+ bl[46] br[46] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_49 
+ bl[47] br[47] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_50 
+ bl[48] br[48] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_51 
+ bl[49] br[49] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_52 
+ bl[50] br[50] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_53 
+ bl[51] br[51] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_54 
+ bl[52] br[52] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_55 
+ bl[53] br[53] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_56 
+ bl[54] br[54] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_57 
+ bl[55] br[55] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_58 
+ bl[56] br[56] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_59 
+ bl[57] br[57] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_60 
+ bl[58] br[58] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_61 
+ bl[59] br[59] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_62 
+ bl[60] br[60] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_63 
+ bl[61] br[61] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_64 
+ bl[62] br[62] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_65 
+ bl[63] br[63] vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_66 
+ vdd vdd vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_397_67 
+ vdd vdd vdd vss wl[395] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_0 
+ vdd vdd vss vdd vpb vnb wl[396] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_398_1 
+ rbl rbr vss vdd vpb vnb wl[396] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_398_2 
+ bl[0] br[0] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_3 
+ bl[1] br[1] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_4 
+ bl[2] br[2] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_5 
+ bl[3] br[3] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_6 
+ bl[4] br[4] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_7 
+ bl[5] br[5] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_8 
+ bl[6] br[6] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_9 
+ bl[7] br[7] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_10 
+ bl[8] br[8] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_11 
+ bl[9] br[9] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_12 
+ bl[10] br[10] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_13 
+ bl[11] br[11] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_14 
+ bl[12] br[12] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_15 
+ bl[13] br[13] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_16 
+ bl[14] br[14] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_17 
+ bl[15] br[15] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_18 
+ bl[16] br[16] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_19 
+ bl[17] br[17] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_20 
+ bl[18] br[18] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_21 
+ bl[19] br[19] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_22 
+ bl[20] br[20] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_23 
+ bl[21] br[21] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_24 
+ bl[22] br[22] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_25 
+ bl[23] br[23] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_26 
+ bl[24] br[24] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_27 
+ bl[25] br[25] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_28 
+ bl[26] br[26] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_29 
+ bl[27] br[27] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_30 
+ bl[28] br[28] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_31 
+ bl[29] br[29] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_32 
+ bl[30] br[30] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_33 
+ bl[31] br[31] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_34 
+ bl[32] br[32] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_35 
+ bl[33] br[33] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_36 
+ bl[34] br[34] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_37 
+ bl[35] br[35] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_38 
+ bl[36] br[36] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_39 
+ bl[37] br[37] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_40 
+ bl[38] br[38] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_41 
+ bl[39] br[39] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_42 
+ bl[40] br[40] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_43 
+ bl[41] br[41] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_44 
+ bl[42] br[42] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_45 
+ bl[43] br[43] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_46 
+ bl[44] br[44] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_47 
+ bl[45] br[45] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_48 
+ bl[46] br[46] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_49 
+ bl[47] br[47] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_50 
+ bl[48] br[48] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_51 
+ bl[49] br[49] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_52 
+ bl[50] br[50] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_53 
+ bl[51] br[51] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_54 
+ bl[52] br[52] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_55 
+ bl[53] br[53] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_56 
+ bl[54] br[54] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_57 
+ bl[55] br[55] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_58 
+ bl[56] br[56] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_59 
+ bl[57] br[57] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_60 
+ bl[58] br[58] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_61 
+ bl[59] br[59] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_62 
+ bl[60] br[60] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_63 
+ bl[61] br[61] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_64 
+ bl[62] br[62] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_65 
+ bl[63] br[63] vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_66 
+ vdd vdd vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_398_67 
+ vdd vdd vdd vss wl[396] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_0 
+ vdd vdd vss vdd vpb vnb wl[397] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_399_1 
+ rbl rbr vss vdd vpb vnb wl[397] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_399_2 
+ bl[0] br[0] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_3 
+ bl[1] br[1] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_4 
+ bl[2] br[2] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_5 
+ bl[3] br[3] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_6 
+ bl[4] br[4] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_7 
+ bl[5] br[5] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_8 
+ bl[6] br[6] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_9 
+ bl[7] br[7] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_10 
+ bl[8] br[8] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_11 
+ bl[9] br[9] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_12 
+ bl[10] br[10] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_13 
+ bl[11] br[11] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_14 
+ bl[12] br[12] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_15 
+ bl[13] br[13] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_16 
+ bl[14] br[14] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_17 
+ bl[15] br[15] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_18 
+ bl[16] br[16] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_19 
+ bl[17] br[17] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_20 
+ bl[18] br[18] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_21 
+ bl[19] br[19] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_22 
+ bl[20] br[20] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_23 
+ bl[21] br[21] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_24 
+ bl[22] br[22] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_25 
+ bl[23] br[23] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_26 
+ bl[24] br[24] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_27 
+ bl[25] br[25] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_28 
+ bl[26] br[26] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_29 
+ bl[27] br[27] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_30 
+ bl[28] br[28] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_31 
+ bl[29] br[29] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_32 
+ bl[30] br[30] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_33 
+ bl[31] br[31] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_34 
+ bl[32] br[32] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_35 
+ bl[33] br[33] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_36 
+ bl[34] br[34] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_37 
+ bl[35] br[35] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_38 
+ bl[36] br[36] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_39 
+ bl[37] br[37] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_40 
+ bl[38] br[38] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_41 
+ bl[39] br[39] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_42 
+ bl[40] br[40] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_43 
+ bl[41] br[41] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_44 
+ bl[42] br[42] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_45 
+ bl[43] br[43] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_46 
+ bl[44] br[44] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_47 
+ bl[45] br[45] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_48 
+ bl[46] br[46] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_49 
+ bl[47] br[47] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_50 
+ bl[48] br[48] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_51 
+ bl[49] br[49] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_52 
+ bl[50] br[50] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_53 
+ bl[51] br[51] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_54 
+ bl[52] br[52] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_55 
+ bl[53] br[53] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_56 
+ bl[54] br[54] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_57 
+ bl[55] br[55] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_58 
+ bl[56] br[56] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_59 
+ bl[57] br[57] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_60 
+ bl[58] br[58] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_61 
+ bl[59] br[59] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_62 
+ bl[60] br[60] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_63 
+ bl[61] br[61] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_64 
+ bl[62] br[62] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_65 
+ bl[63] br[63] vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_66 
+ vdd vdd vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_399_67 
+ vdd vdd vdd vss wl[397] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_0 
+ vdd vdd vss vdd vpb vnb wl[398] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_400_1 
+ rbl rbr vss vdd vpb vnb wl[398] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_400_2 
+ bl[0] br[0] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_3 
+ bl[1] br[1] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_4 
+ bl[2] br[2] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_5 
+ bl[3] br[3] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_6 
+ bl[4] br[4] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_7 
+ bl[5] br[5] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_8 
+ bl[6] br[6] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_9 
+ bl[7] br[7] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_10 
+ bl[8] br[8] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_11 
+ bl[9] br[9] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_12 
+ bl[10] br[10] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_13 
+ bl[11] br[11] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_14 
+ bl[12] br[12] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_15 
+ bl[13] br[13] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_16 
+ bl[14] br[14] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_17 
+ bl[15] br[15] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_18 
+ bl[16] br[16] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_19 
+ bl[17] br[17] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_20 
+ bl[18] br[18] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_21 
+ bl[19] br[19] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_22 
+ bl[20] br[20] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_23 
+ bl[21] br[21] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_24 
+ bl[22] br[22] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_25 
+ bl[23] br[23] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_26 
+ bl[24] br[24] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_27 
+ bl[25] br[25] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_28 
+ bl[26] br[26] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_29 
+ bl[27] br[27] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_30 
+ bl[28] br[28] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_31 
+ bl[29] br[29] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_32 
+ bl[30] br[30] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_33 
+ bl[31] br[31] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_34 
+ bl[32] br[32] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_35 
+ bl[33] br[33] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_36 
+ bl[34] br[34] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_37 
+ bl[35] br[35] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_38 
+ bl[36] br[36] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_39 
+ bl[37] br[37] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_40 
+ bl[38] br[38] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_41 
+ bl[39] br[39] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_42 
+ bl[40] br[40] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_43 
+ bl[41] br[41] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_44 
+ bl[42] br[42] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_45 
+ bl[43] br[43] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_46 
+ bl[44] br[44] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_47 
+ bl[45] br[45] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_48 
+ bl[46] br[46] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_49 
+ bl[47] br[47] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_50 
+ bl[48] br[48] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_51 
+ bl[49] br[49] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_52 
+ bl[50] br[50] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_53 
+ bl[51] br[51] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_54 
+ bl[52] br[52] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_55 
+ bl[53] br[53] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_56 
+ bl[54] br[54] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_57 
+ bl[55] br[55] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_58 
+ bl[56] br[56] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_59 
+ bl[57] br[57] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_60 
+ bl[58] br[58] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_61 
+ bl[59] br[59] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_62 
+ bl[60] br[60] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_63 
+ bl[61] br[61] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_64 
+ bl[62] br[62] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_65 
+ bl[63] br[63] vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_66 
+ vdd vdd vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_400_67 
+ vdd vdd vdd vss wl[398] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_0 
+ vdd vdd vss vdd vpb vnb wl[399] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_401_1 
+ rbl rbr vss vdd vpb vnb wl[399] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_401_2 
+ bl[0] br[0] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_3 
+ bl[1] br[1] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_4 
+ bl[2] br[2] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_5 
+ bl[3] br[3] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_6 
+ bl[4] br[4] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_7 
+ bl[5] br[5] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_8 
+ bl[6] br[6] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_9 
+ bl[7] br[7] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_10 
+ bl[8] br[8] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_11 
+ bl[9] br[9] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_12 
+ bl[10] br[10] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_13 
+ bl[11] br[11] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_14 
+ bl[12] br[12] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_15 
+ bl[13] br[13] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_16 
+ bl[14] br[14] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_17 
+ bl[15] br[15] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_18 
+ bl[16] br[16] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_19 
+ bl[17] br[17] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_20 
+ bl[18] br[18] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_21 
+ bl[19] br[19] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_22 
+ bl[20] br[20] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_23 
+ bl[21] br[21] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_24 
+ bl[22] br[22] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_25 
+ bl[23] br[23] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_26 
+ bl[24] br[24] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_27 
+ bl[25] br[25] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_28 
+ bl[26] br[26] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_29 
+ bl[27] br[27] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_30 
+ bl[28] br[28] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_31 
+ bl[29] br[29] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_32 
+ bl[30] br[30] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_33 
+ bl[31] br[31] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_34 
+ bl[32] br[32] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_35 
+ bl[33] br[33] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_36 
+ bl[34] br[34] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_37 
+ bl[35] br[35] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_38 
+ bl[36] br[36] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_39 
+ bl[37] br[37] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_40 
+ bl[38] br[38] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_41 
+ bl[39] br[39] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_42 
+ bl[40] br[40] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_43 
+ bl[41] br[41] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_44 
+ bl[42] br[42] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_45 
+ bl[43] br[43] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_46 
+ bl[44] br[44] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_47 
+ bl[45] br[45] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_48 
+ bl[46] br[46] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_49 
+ bl[47] br[47] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_50 
+ bl[48] br[48] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_51 
+ bl[49] br[49] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_52 
+ bl[50] br[50] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_53 
+ bl[51] br[51] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_54 
+ bl[52] br[52] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_55 
+ bl[53] br[53] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_56 
+ bl[54] br[54] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_57 
+ bl[55] br[55] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_58 
+ bl[56] br[56] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_59 
+ bl[57] br[57] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_60 
+ bl[58] br[58] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_61 
+ bl[59] br[59] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_62 
+ bl[60] br[60] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_63 
+ bl[61] br[61] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_64 
+ bl[62] br[62] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_65 
+ bl[63] br[63] vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_66 
+ vdd vdd vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_401_67 
+ vdd vdd vdd vss wl[399] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_0 
+ vdd vdd vss vdd vpb vnb wl[400] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_402_1 
+ rbl rbr vss vdd vpb vnb wl[400] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_402_2 
+ bl[0] br[0] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_3 
+ bl[1] br[1] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_4 
+ bl[2] br[2] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_5 
+ bl[3] br[3] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_6 
+ bl[4] br[4] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_7 
+ bl[5] br[5] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_8 
+ bl[6] br[6] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_9 
+ bl[7] br[7] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_10 
+ bl[8] br[8] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_11 
+ bl[9] br[9] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_12 
+ bl[10] br[10] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_13 
+ bl[11] br[11] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_14 
+ bl[12] br[12] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_15 
+ bl[13] br[13] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_16 
+ bl[14] br[14] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_17 
+ bl[15] br[15] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_18 
+ bl[16] br[16] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_19 
+ bl[17] br[17] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_20 
+ bl[18] br[18] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_21 
+ bl[19] br[19] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_22 
+ bl[20] br[20] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_23 
+ bl[21] br[21] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_24 
+ bl[22] br[22] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_25 
+ bl[23] br[23] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_26 
+ bl[24] br[24] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_27 
+ bl[25] br[25] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_28 
+ bl[26] br[26] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_29 
+ bl[27] br[27] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_30 
+ bl[28] br[28] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_31 
+ bl[29] br[29] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_32 
+ bl[30] br[30] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_33 
+ bl[31] br[31] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_34 
+ bl[32] br[32] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_35 
+ bl[33] br[33] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_36 
+ bl[34] br[34] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_37 
+ bl[35] br[35] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_38 
+ bl[36] br[36] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_39 
+ bl[37] br[37] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_40 
+ bl[38] br[38] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_41 
+ bl[39] br[39] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_42 
+ bl[40] br[40] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_43 
+ bl[41] br[41] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_44 
+ bl[42] br[42] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_45 
+ bl[43] br[43] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_46 
+ bl[44] br[44] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_47 
+ bl[45] br[45] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_48 
+ bl[46] br[46] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_49 
+ bl[47] br[47] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_50 
+ bl[48] br[48] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_51 
+ bl[49] br[49] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_52 
+ bl[50] br[50] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_53 
+ bl[51] br[51] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_54 
+ bl[52] br[52] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_55 
+ bl[53] br[53] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_56 
+ bl[54] br[54] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_57 
+ bl[55] br[55] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_58 
+ bl[56] br[56] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_59 
+ bl[57] br[57] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_60 
+ bl[58] br[58] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_61 
+ bl[59] br[59] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_62 
+ bl[60] br[60] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_63 
+ bl[61] br[61] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_64 
+ bl[62] br[62] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_65 
+ bl[63] br[63] vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_66 
+ vdd vdd vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_402_67 
+ vdd vdd vdd vss wl[400] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_0 
+ vdd vdd vss vdd vpb vnb wl[401] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_403_1 
+ rbl rbr vss vdd vpb vnb wl[401] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_403_2 
+ bl[0] br[0] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_3 
+ bl[1] br[1] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_4 
+ bl[2] br[2] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_5 
+ bl[3] br[3] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_6 
+ bl[4] br[4] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_7 
+ bl[5] br[5] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_8 
+ bl[6] br[6] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_9 
+ bl[7] br[7] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_10 
+ bl[8] br[8] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_11 
+ bl[9] br[9] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_12 
+ bl[10] br[10] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_13 
+ bl[11] br[11] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_14 
+ bl[12] br[12] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_15 
+ bl[13] br[13] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_16 
+ bl[14] br[14] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_17 
+ bl[15] br[15] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_18 
+ bl[16] br[16] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_19 
+ bl[17] br[17] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_20 
+ bl[18] br[18] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_21 
+ bl[19] br[19] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_22 
+ bl[20] br[20] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_23 
+ bl[21] br[21] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_24 
+ bl[22] br[22] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_25 
+ bl[23] br[23] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_26 
+ bl[24] br[24] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_27 
+ bl[25] br[25] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_28 
+ bl[26] br[26] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_29 
+ bl[27] br[27] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_30 
+ bl[28] br[28] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_31 
+ bl[29] br[29] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_32 
+ bl[30] br[30] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_33 
+ bl[31] br[31] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_34 
+ bl[32] br[32] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_35 
+ bl[33] br[33] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_36 
+ bl[34] br[34] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_37 
+ bl[35] br[35] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_38 
+ bl[36] br[36] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_39 
+ bl[37] br[37] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_40 
+ bl[38] br[38] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_41 
+ bl[39] br[39] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_42 
+ bl[40] br[40] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_43 
+ bl[41] br[41] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_44 
+ bl[42] br[42] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_45 
+ bl[43] br[43] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_46 
+ bl[44] br[44] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_47 
+ bl[45] br[45] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_48 
+ bl[46] br[46] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_49 
+ bl[47] br[47] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_50 
+ bl[48] br[48] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_51 
+ bl[49] br[49] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_52 
+ bl[50] br[50] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_53 
+ bl[51] br[51] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_54 
+ bl[52] br[52] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_55 
+ bl[53] br[53] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_56 
+ bl[54] br[54] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_57 
+ bl[55] br[55] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_58 
+ bl[56] br[56] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_59 
+ bl[57] br[57] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_60 
+ bl[58] br[58] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_61 
+ bl[59] br[59] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_62 
+ bl[60] br[60] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_63 
+ bl[61] br[61] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_64 
+ bl[62] br[62] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_65 
+ bl[63] br[63] vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_66 
+ vdd vdd vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_403_67 
+ vdd vdd vdd vss wl[401] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_0 
+ vdd vdd vss vdd vpb vnb wl[402] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_404_1 
+ rbl rbr vss vdd vpb vnb wl[402] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_404_2 
+ bl[0] br[0] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_3 
+ bl[1] br[1] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_4 
+ bl[2] br[2] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_5 
+ bl[3] br[3] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_6 
+ bl[4] br[4] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_7 
+ bl[5] br[5] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_8 
+ bl[6] br[6] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_9 
+ bl[7] br[7] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_10 
+ bl[8] br[8] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_11 
+ bl[9] br[9] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_12 
+ bl[10] br[10] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_13 
+ bl[11] br[11] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_14 
+ bl[12] br[12] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_15 
+ bl[13] br[13] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_16 
+ bl[14] br[14] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_17 
+ bl[15] br[15] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_18 
+ bl[16] br[16] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_19 
+ bl[17] br[17] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_20 
+ bl[18] br[18] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_21 
+ bl[19] br[19] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_22 
+ bl[20] br[20] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_23 
+ bl[21] br[21] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_24 
+ bl[22] br[22] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_25 
+ bl[23] br[23] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_26 
+ bl[24] br[24] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_27 
+ bl[25] br[25] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_28 
+ bl[26] br[26] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_29 
+ bl[27] br[27] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_30 
+ bl[28] br[28] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_31 
+ bl[29] br[29] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_32 
+ bl[30] br[30] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_33 
+ bl[31] br[31] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_34 
+ bl[32] br[32] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_35 
+ bl[33] br[33] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_36 
+ bl[34] br[34] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_37 
+ bl[35] br[35] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_38 
+ bl[36] br[36] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_39 
+ bl[37] br[37] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_40 
+ bl[38] br[38] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_41 
+ bl[39] br[39] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_42 
+ bl[40] br[40] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_43 
+ bl[41] br[41] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_44 
+ bl[42] br[42] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_45 
+ bl[43] br[43] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_46 
+ bl[44] br[44] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_47 
+ bl[45] br[45] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_48 
+ bl[46] br[46] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_49 
+ bl[47] br[47] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_50 
+ bl[48] br[48] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_51 
+ bl[49] br[49] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_52 
+ bl[50] br[50] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_53 
+ bl[51] br[51] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_54 
+ bl[52] br[52] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_55 
+ bl[53] br[53] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_56 
+ bl[54] br[54] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_57 
+ bl[55] br[55] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_58 
+ bl[56] br[56] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_59 
+ bl[57] br[57] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_60 
+ bl[58] br[58] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_61 
+ bl[59] br[59] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_62 
+ bl[60] br[60] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_63 
+ bl[61] br[61] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_64 
+ bl[62] br[62] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_65 
+ bl[63] br[63] vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_66 
+ vdd vdd vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_404_67 
+ vdd vdd vdd vss wl[402] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_0 
+ vdd vdd vss vdd vpb vnb wl[403] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_405_1 
+ rbl rbr vss vdd vpb vnb wl[403] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_405_2 
+ bl[0] br[0] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_3 
+ bl[1] br[1] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_4 
+ bl[2] br[2] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_5 
+ bl[3] br[3] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_6 
+ bl[4] br[4] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_7 
+ bl[5] br[5] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_8 
+ bl[6] br[6] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_9 
+ bl[7] br[7] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_10 
+ bl[8] br[8] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_11 
+ bl[9] br[9] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_12 
+ bl[10] br[10] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_13 
+ bl[11] br[11] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_14 
+ bl[12] br[12] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_15 
+ bl[13] br[13] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_16 
+ bl[14] br[14] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_17 
+ bl[15] br[15] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_18 
+ bl[16] br[16] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_19 
+ bl[17] br[17] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_20 
+ bl[18] br[18] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_21 
+ bl[19] br[19] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_22 
+ bl[20] br[20] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_23 
+ bl[21] br[21] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_24 
+ bl[22] br[22] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_25 
+ bl[23] br[23] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_26 
+ bl[24] br[24] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_27 
+ bl[25] br[25] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_28 
+ bl[26] br[26] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_29 
+ bl[27] br[27] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_30 
+ bl[28] br[28] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_31 
+ bl[29] br[29] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_32 
+ bl[30] br[30] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_33 
+ bl[31] br[31] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_34 
+ bl[32] br[32] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_35 
+ bl[33] br[33] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_36 
+ bl[34] br[34] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_37 
+ bl[35] br[35] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_38 
+ bl[36] br[36] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_39 
+ bl[37] br[37] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_40 
+ bl[38] br[38] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_41 
+ bl[39] br[39] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_42 
+ bl[40] br[40] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_43 
+ bl[41] br[41] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_44 
+ bl[42] br[42] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_45 
+ bl[43] br[43] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_46 
+ bl[44] br[44] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_47 
+ bl[45] br[45] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_48 
+ bl[46] br[46] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_49 
+ bl[47] br[47] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_50 
+ bl[48] br[48] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_51 
+ bl[49] br[49] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_52 
+ bl[50] br[50] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_53 
+ bl[51] br[51] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_54 
+ bl[52] br[52] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_55 
+ bl[53] br[53] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_56 
+ bl[54] br[54] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_57 
+ bl[55] br[55] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_58 
+ bl[56] br[56] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_59 
+ bl[57] br[57] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_60 
+ bl[58] br[58] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_61 
+ bl[59] br[59] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_62 
+ bl[60] br[60] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_63 
+ bl[61] br[61] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_64 
+ bl[62] br[62] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_65 
+ bl[63] br[63] vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_66 
+ vdd vdd vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_405_67 
+ vdd vdd vdd vss wl[403] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_0 
+ vdd vdd vss vdd vpb vnb wl[404] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_406_1 
+ rbl rbr vss vdd vpb vnb wl[404] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_406_2 
+ bl[0] br[0] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_3 
+ bl[1] br[1] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_4 
+ bl[2] br[2] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_5 
+ bl[3] br[3] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_6 
+ bl[4] br[4] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_7 
+ bl[5] br[5] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_8 
+ bl[6] br[6] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_9 
+ bl[7] br[7] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_10 
+ bl[8] br[8] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_11 
+ bl[9] br[9] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_12 
+ bl[10] br[10] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_13 
+ bl[11] br[11] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_14 
+ bl[12] br[12] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_15 
+ bl[13] br[13] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_16 
+ bl[14] br[14] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_17 
+ bl[15] br[15] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_18 
+ bl[16] br[16] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_19 
+ bl[17] br[17] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_20 
+ bl[18] br[18] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_21 
+ bl[19] br[19] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_22 
+ bl[20] br[20] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_23 
+ bl[21] br[21] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_24 
+ bl[22] br[22] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_25 
+ bl[23] br[23] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_26 
+ bl[24] br[24] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_27 
+ bl[25] br[25] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_28 
+ bl[26] br[26] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_29 
+ bl[27] br[27] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_30 
+ bl[28] br[28] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_31 
+ bl[29] br[29] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_32 
+ bl[30] br[30] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_33 
+ bl[31] br[31] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_34 
+ bl[32] br[32] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_35 
+ bl[33] br[33] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_36 
+ bl[34] br[34] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_37 
+ bl[35] br[35] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_38 
+ bl[36] br[36] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_39 
+ bl[37] br[37] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_40 
+ bl[38] br[38] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_41 
+ bl[39] br[39] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_42 
+ bl[40] br[40] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_43 
+ bl[41] br[41] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_44 
+ bl[42] br[42] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_45 
+ bl[43] br[43] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_46 
+ bl[44] br[44] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_47 
+ bl[45] br[45] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_48 
+ bl[46] br[46] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_49 
+ bl[47] br[47] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_50 
+ bl[48] br[48] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_51 
+ bl[49] br[49] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_52 
+ bl[50] br[50] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_53 
+ bl[51] br[51] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_54 
+ bl[52] br[52] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_55 
+ bl[53] br[53] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_56 
+ bl[54] br[54] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_57 
+ bl[55] br[55] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_58 
+ bl[56] br[56] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_59 
+ bl[57] br[57] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_60 
+ bl[58] br[58] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_61 
+ bl[59] br[59] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_62 
+ bl[60] br[60] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_63 
+ bl[61] br[61] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_64 
+ bl[62] br[62] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_65 
+ bl[63] br[63] vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_66 
+ vdd vdd vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_406_67 
+ vdd vdd vdd vss wl[404] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_0 
+ vdd vdd vss vdd vpb vnb wl[405] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_407_1 
+ rbl rbr vss vdd vpb vnb wl[405] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_407_2 
+ bl[0] br[0] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_3 
+ bl[1] br[1] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_4 
+ bl[2] br[2] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_5 
+ bl[3] br[3] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_6 
+ bl[4] br[4] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_7 
+ bl[5] br[5] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_8 
+ bl[6] br[6] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_9 
+ bl[7] br[7] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_10 
+ bl[8] br[8] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_11 
+ bl[9] br[9] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_12 
+ bl[10] br[10] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_13 
+ bl[11] br[11] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_14 
+ bl[12] br[12] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_15 
+ bl[13] br[13] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_16 
+ bl[14] br[14] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_17 
+ bl[15] br[15] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_18 
+ bl[16] br[16] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_19 
+ bl[17] br[17] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_20 
+ bl[18] br[18] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_21 
+ bl[19] br[19] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_22 
+ bl[20] br[20] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_23 
+ bl[21] br[21] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_24 
+ bl[22] br[22] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_25 
+ bl[23] br[23] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_26 
+ bl[24] br[24] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_27 
+ bl[25] br[25] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_28 
+ bl[26] br[26] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_29 
+ bl[27] br[27] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_30 
+ bl[28] br[28] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_31 
+ bl[29] br[29] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_32 
+ bl[30] br[30] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_33 
+ bl[31] br[31] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_34 
+ bl[32] br[32] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_35 
+ bl[33] br[33] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_36 
+ bl[34] br[34] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_37 
+ bl[35] br[35] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_38 
+ bl[36] br[36] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_39 
+ bl[37] br[37] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_40 
+ bl[38] br[38] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_41 
+ bl[39] br[39] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_42 
+ bl[40] br[40] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_43 
+ bl[41] br[41] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_44 
+ bl[42] br[42] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_45 
+ bl[43] br[43] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_46 
+ bl[44] br[44] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_47 
+ bl[45] br[45] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_48 
+ bl[46] br[46] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_49 
+ bl[47] br[47] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_50 
+ bl[48] br[48] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_51 
+ bl[49] br[49] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_52 
+ bl[50] br[50] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_53 
+ bl[51] br[51] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_54 
+ bl[52] br[52] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_55 
+ bl[53] br[53] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_56 
+ bl[54] br[54] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_57 
+ bl[55] br[55] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_58 
+ bl[56] br[56] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_59 
+ bl[57] br[57] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_60 
+ bl[58] br[58] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_61 
+ bl[59] br[59] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_62 
+ bl[60] br[60] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_63 
+ bl[61] br[61] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_64 
+ bl[62] br[62] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_65 
+ bl[63] br[63] vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_66 
+ vdd vdd vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_407_67 
+ vdd vdd vdd vss wl[405] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_0 
+ vdd vdd vss vdd vpb vnb wl[406] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_408_1 
+ rbl rbr vss vdd vpb vnb wl[406] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_408_2 
+ bl[0] br[0] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_3 
+ bl[1] br[1] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_4 
+ bl[2] br[2] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_5 
+ bl[3] br[3] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_6 
+ bl[4] br[4] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_7 
+ bl[5] br[5] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_8 
+ bl[6] br[6] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_9 
+ bl[7] br[7] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_10 
+ bl[8] br[8] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_11 
+ bl[9] br[9] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_12 
+ bl[10] br[10] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_13 
+ bl[11] br[11] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_14 
+ bl[12] br[12] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_15 
+ bl[13] br[13] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_16 
+ bl[14] br[14] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_17 
+ bl[15] br[15] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_18 
+ bl[16] br[16] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_19 
+ bl[17] br[17] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_20 
+ bl[18] br[18] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_21 
+ bl[19] br[19] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_22 
+ bl[20] br[20] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_23 
+ bl[21] br[21] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_24 
+ bl[22] br[22] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_25 
+ bl[23] br[23] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_26 
+ bl[24] br[24] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_27 
+ bl[25] br[25] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_28 
+ bl[26] br[26] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_29 
+ bl[27] br[27] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_30 
+ bl[28] br[28] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_31 
+ bl[29] br[29] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_32 
+ bl[30] br[30] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_33 
+ bl[31] br[31] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_34 
+ bl[32] br[32] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_35 
+ bl[33] br[33] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_36 
+ bl[34] br[34] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_37 
+ bl[35] br[35] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_38 
+ bl[36] br[36] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_39 
+ bl[37] br[37] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_40 
+ bl[38] br[38] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_41 
+ bl[39] br[39] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_42 
+ bl[40] br[40] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_43 
+ bl[41] br[41] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_44 
+ bl[42] br[42] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_45 
+ bl[43] br[43] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_46 
+ bl[44] br[44] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_47 
+ bl[45] br[45] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_48 
+ bl[46] br[46] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_49 
+ bl[47] br[47] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_50 
+ bl[48] br[48] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_51 
+ bl[49] br[49] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_52 
+ bl[50] br[50] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_53 
+ bl[51] br[51] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_54 
+ bl[52] br[52] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_55 
+ bl[53] br[53] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_56 
+ bl[54] br[54] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_57 
+ bl[55] br[55] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_58 
+ bl[56] br[56] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_59 
+ bl[57] br[57] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_60 
+ bl[58] br[58] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_61 
+ bl[59] br[59] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_62 
+ bl[60] br[60] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_63 
+ bl[61] br[61] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_64 
+ bl[62] br[62] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_65 
+ bl[63] br[63] vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_66 
+ vdd vdd vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_408_67 
+ vdd vdd vdd vss wl[406] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_0 
+ vdd vdd vss vdd vpb vnb wl[407] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_409_1 
+ rbl rbr vss vdd vpb vnb wl[407] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_409_2 
+ bl[0] br[0] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_3 
+ bl[1] br[1] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_4 
+ bl[2] br[2] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_5 
+ bl[3] br[3] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_6 
+ bl[4] br[4] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_7 
+ bl[5] br[5] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_8 
+ bl[6] br[6] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_9 
+ bl[7] br[7] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_10 
+ bl[8] br[8] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_11 
+ bl[9] br[9] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_12 
+ bl[10] br[10] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_13 
+ bl[11] br[11] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_14 
+ bl[12] br[12] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_15 
+ bl[13] br[13] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_16 
+ bl[14] br[14] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_17 
+ bl[15] br[15] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_18 
+ bl[16] br[16] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_19 
+ bl[17] br[17] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_20 
+ bl[18] br[18] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_21 
+ bl[19] br[19] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_22 
+ bl[20] br[20] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_23 
+ bl[21] br[21] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_24 
+ bl[22] br[22] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_25 
+ bl[23] br[23] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_26 
+ bl[24] br[24] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_27 
+ bl[25] br[25] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_28 
+ bl[26] br[26] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_29 
+ bl[27] br[27] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_30 
+ bl[28] br[28] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_31 
+ bl[29] br[29] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_32 
+ bl[30] br[30] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_33 
+ bl[31] br[31] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_34 
+ bl[32] br[32] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_35 
+ bl[33] br[33] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_36 
+ bl[34] br[34] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_37 
+ bl[35] br[35] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_38 
+ bl[36] br[36] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_39 
+ bl[37] br[37] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_40 
+ bl[38] br[38] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_41 
+ bl[39] br[39] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_42 
+ bl[40] br[40] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_43 
+ bl[41] br[41] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_44 
+ bl[42] br[42] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_45 
+ bl[43] br[43] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_46 
+ bl[44] br[44] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_47 
+ bl[45] br[45] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_48 
+ bl[46] br[46] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_49 
+ bl[47] br[47] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_50 
+ bl[48] br[48] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_51 
+ bl[49] br[49] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_52 
+ bl[50] br[50] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_53 
+ bl[51] br[51] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_54 
+ bl[52] br[52] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_55 
+ bl[53] br[53] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_56 
+ bl[54] br[54] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_57 
+ bl[55] br[55] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_58 
+ bl[56] br[56] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_59 
+ bl[57] br[57] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_60 
+ bl[58] br[58] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_61 
+ bl[59] br[59] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_62 
+ bl[60] br[60] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_63 
+ bl[61] br[61] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_64 
+ bl[62] br[62] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_65 
+ bl[63] br[63] vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_66 
+ vdd vdd vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_409_67 
+ vdd vdd vdd vss wl[407] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_0 
+ vdd vdd vss vdd vpb vnb wl[408] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_410_1 
+ rbl rbr vss vdd vpb vnb wl[408] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_410_2 
+ bl[0] br[0] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_3 
+ bl[1] br[1] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_4 
+ bl[2] br[2] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_5 
+ bl[3] br[3] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_6 
+ bl[4] br[4] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_7 
+ bl[5] br[5] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_8 
+ bl[6] br[6] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_9 
+ bl[7] br[7] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_10 
+ bl[8] br[8] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_11 
+ bl[9] br[9] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_12 
+ bl[10] br[10] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_13 
+ bl[11] br[11] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_14 
+ bl[12] br[12] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_15 
+ bl[13] br[13] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_16 
+ bl[14] br[14] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_17 
+ bl[15] br[15] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_18 
+ bl[16] br[16] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_19 
+ bl[17] br[17] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_20 
+ bl[18] br[18] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_21 
+ bl[19] br[19] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_22 
+ bl[20] br[20] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_23 
+ bl[21] br[21] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_24 
+ bl[22] br[22] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_25 
+ bl[23] br[23] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_26 
+ bl[24] br[24] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_27 
+ bl[25] br[25] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_28 
+ bl[26] br[26] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_29 
+ bl[27] br[27] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_30 
+ bl[28] br[28] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_31 
+ bl[29] br[29] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_32 
+ bl[30] br[30] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_33 
+ bl[31] br[31] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_34 
+ bl[32] br[32] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_35 
+ bl[33] br[33] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_36 
+ bl[34] br[34] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_37 
+ bl[35] br[35] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_38 
+ bl[36] br[36] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_39 
+ bl[37] br[37] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_40 
+ bl[38] br[38] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_41 
+ bl[39] br[39] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_42 
+ bl[40] br[40] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_43 
+ bl[41] br[41] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_44 
+ bl[42] br[42] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_45 
+ bl[43] br[43] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_46 
+ bl[44] br[44] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_47 
+ bl[45] br[45] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_48 
+ bl[46] br[46] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_49 
+ bl[47] br[47] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_50 
+ bl[48] br[48] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_51 
+ bl[49] br[49] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_52 
+ bl[50] br[50] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_53 
+ bl[51] br[51] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_54 
+ bl[52] br[52] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_55 
+ bl[53] br[53] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_56 
+ bl[54] br[54] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_57 
+ bl[55] br[55] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_58 
+ bl[56] br[56] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_59 
+ bl[57] br[57] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_60 
+ bl[58] br[58] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_61 
+ bl[59] br[59] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_62 
+ bl[60] br[60] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_63 
+ bl[61] br[61] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_64 
+ bl[62] br[62] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_65 
+ bl[63] br[63] vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_66 
+ vdd vdd vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_410_67 
+ vdd vdd vdd vss wl[408] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_0 
+ vdd vdd vss vdd vpb vnb wl[409] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_411_1 
+ rbl rbr vss vdd vpb vnb wl[409] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_411_2 
+ bl[0] br[0] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_3 
+ bl[1] br[1] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_4 
+ bl[2] br[2] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_5 
+ bl[3] br[3] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_6 
+ bl[4] br[4] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_7 
+ bl[5] br[5] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_8 
+ bl[6] br[6] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_9 
+ bl[7] br[7] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_10 
+ bl[8] br[8] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_11 
+ bl[9] br[9] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_12 
+ bl[10] br[10] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_13 
+ bl[11] br[11] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_14 
+ bl[12] br[12] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_15 
+ bl[13] br[13] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_16 
+ bl[14] br[14] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_17 
+ bl[15] br[15] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_18 
+ bl[16] br[16] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_19 
+ bl[17] br[17] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_20 
+ bl[18] br[18] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_21 
+ bl[19] br[19] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_22 
+ bl[20] br[20] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_23 
+ bl[21] br[21] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_24 
+ bl[22] br[22] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_25 
+ bl[23] br[23] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_26 
+ bl[24] br[24] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_27 
+ bl[25] br[25] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_28 
+ bl[26] br[26] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_29 
+ bl[27] br[27] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_30 
+ bl[28] br[28] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_31 
+ bl[29] br[29] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_32 
+ bl[30] br[30] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_33 
+ bl[31] br[31] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_34 
+ bl[32] br[32] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_35 
+ bl[33] br[33] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_36 
+ bl[34] br[34] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_37 
+ bl[35] br[35] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_38 
+ bl[36] br[36] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_39 
+ bl[37] br[37] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_40 
+ bl[38] br[38] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_41 
+ bl[39] br[39] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_42 
+ bl[40] br[40] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_43 
+ bl[41] br[41] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_44 
+ bl[42] br[42] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_45 
+ bl[43] br[43] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_46 
+ bl[44] br[44] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_47 
+ bl[45] br[45] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_48 
+ bl[46] br[46] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_49 
+ bl[47] br[47] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_50 
+ bl[48] br[48] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_51 
+ bl[49] br[49] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_52 
+ bl[50] br[50] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_53 
+ bl[51] br[51] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_54 
+ bl[52] br[52] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_55 
+ bl[53] br[53] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_56 
+ bl[54] br[54] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_57 
+ bl[55] br[55] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_58 
+ bl[56] br[56] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_59 
+ bl[57] br[57] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_60 
+ bl[58] br[58] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_61 
+ bl[59] br[59] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_62 
+ bl[60] br[60] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_63 
+ bl[61] br[61] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_64 
+ bl[62] br[62] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_65 
+ bl[63] br[63] vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_66 
+ vdd vdd vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_411_67 
+ vdd vdd vdd vss wl[409] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_0 
+ vdd vdd vss vdd vpb vnb wl[410] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_412_1 
+ rbl rbr vss vdd vpb vnb wl[410] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_412_2 
+ bl[0] br[0] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_3 
+ bl[1] br[1] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_4 
+ bl[2] br[2] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_5 
+ bl[3] br[3] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_6 
+ bl[4] br[4] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_7 
+ bl[5] br[5] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_8 
+ bl[6] br[6] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_9 
+ bl[7] br[7] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_10 
+ bl[8] br[8] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_11 
+ bl[9] br[9] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_12 
+ bl[10] br[10] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_13 
+ bl[11] br[11] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_14 
+ bl[12] br[12] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_15 
+ bl[13] br[13] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_16 
+ bl[14] br[14] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_17 
+ bl[15] br[15] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_18 
+ bl[16] br[16] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_19 
+ bl[17] br[17] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_20 
+ bl[18] br[18] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_21 
+ bl[19] br[19] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_22 
+ bl[20] br[20] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_23 
+ bl[21] br[21] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_24 
+ bl[22] br[22] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_25 
+ bl[23] br[23] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_26 
+ bl[24] br[24] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_27 
+ bl[25] br[25] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_28 
+ bl[26] br[26] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_29 
+ bl[27] br[27] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_30 
+ bl[28] br[28] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_31 
+ bl[29] br[29] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_32 
+ bl[30] br[30] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_33 
+ bl[31] br[31] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_34 
+ bl[32] br[32] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_35 
+ bl[33] br[33] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_36 
+ bl[34] br[34] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_37 
+ bl[35] br[35] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_38 
+ bl[36] br[36] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_39 
+ bl[37] br[37] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_40 
+ bl[38] br[38] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_41 
+ bl[39] br[39] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_42 
+ bl[40] br[40] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_43 
+ bl[41] br[41] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_44 
+ bl[42] br[42] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_45 
+ bl[43] br[43] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_46 
+ bl[44] br[44] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_47 
+ bl[45] br[45] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_48 
+ bl[46] br[46] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_49 
+ bl[47] br[47] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_50 
+ bl[48] br[48] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_51 
+ bl[49] br[49] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_52 
+ bl[50] br[50] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_53 
+ bl[51] br[51] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_54 
+ bl[52] br[52] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_55 
+ bl[53] br[53] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_56 
+ bl[54] br[54] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_57 
+ bl[55] br[55] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_58 
+ bl[56] br[56] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_59 
+ bl[57] br[57] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_60 
+ bl[58] br[58] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_61 
+ bl[59] br[59] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_62 
+ bl[60] br[60] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_63 
+ bl[61] br[61] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_64 
+ bl[62] br[62] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_65 
+ bl[63] br[63] vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_66 
+ vdd vdd vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_412_67 
+ vdd vdd vdd vss wl[410] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_0 
+ vdd vdd vss vdd vpb vnb wl[411] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_413_1 
+ rbl rbr vss vdd vpb vnb wl[411] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_413_2 
+ bl[0] br[0] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_3 
+ bl[1] br[1] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_4 
+ bl[2] br[2] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_5 
+ bl[3] br[3] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_6 
+ bl[4] br[4] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_7 
+ bl[5] br[5] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_8 
+ bl[6] br[6] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_9 
+ bl[7] br[7] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_10 
+ bl[8] br[8] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_11 
+ bl[9] br[9] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_12 
+ bl[10] br[10] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_13 
+ bl[11] br[11] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_14 
+ bl[12] br[12] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_15 
+ bl[13] br[13] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_16 
+ bl[14] br[14] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_17 
+ bl[15] br[15] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_18 
+ bl[16] br[16] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_19 
+ bl[17] br[17] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_20 
+ bl[18] br[18] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_21 
+ bl[19] br[19] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_22 
+ bl[20] br[20] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_23 
+ bl[21] br[21] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_24 
+ bl[22] br[22] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_25 
+ bl[23] br[23] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_26 
+ bl[24] br[24] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_27 
+ bl[25] br[25] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_28 
+ bl[26] br[26] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_29 
+ bl[27] br[27] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_30 
+ bl[28] br[28] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_31 
+ bl[29] br[29] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_32 
+ bl[30] br[30] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_33 
+ bl[31] br[31] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_34 
+ bl[32] br[32] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_35 
+ bl[33] br[33] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_36 
+ bl[34] br[34] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_37 
+ bl[35] br[35] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_38 
+ bl[36] br[36] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_39 
+ bl[37] br[37] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_40 
+ bl[38] br[38] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_41 
+ bl[39] br[39] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_42 
+ bl[40] br[40] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_43 
+ bl[41] br[41] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_44 
+ bl[42] br[42] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_45 
+ bl[43] br[43] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_46 
+ bl[44] br[44] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_47 
+ bl[45] br[45] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_48 
+ bl[46] br[46] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_49 
+ bl[47] br[47] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_50 
+ bl[48] br[48] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_51 
+ bl[49] br[49] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_52 
+ bl[50] br[50] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_53 
+ bl[51] br[51] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_54 
+ bl[52] br[52] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_55 
+ bl[53] br[53] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_56 
+ bl[54] br[54] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_57 
+ bl[55] br[55] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_58 
+ bl[56] br[56] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_59 
+ bl[57] br[57] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_60 
+ bl[58] br[58] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_61 
+ bl[59] br[59] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_62 
+ bl[60] br[60] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_63 
+ bl[61] br[61] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_64 
+ bl[62] br[62] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_65 
+ bl[63] br[63] vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_66 
+ vdd vdd vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_413_67 
+ vdd vdd vdd vss wl[411] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_0 
+ vdd vdd vss vdd vpb vnb wl[412] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_414_1 
+ rbl rbr vss vdd vpb vnb wl[412] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_414_2 
+ bl[0] br[0] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_3 
+ bl[1] br[1] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_4 
+ bl[2] br[2] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_5 
+ bl[3] br[3] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_6 
+ bl[4] br[4] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_7 
+ bl[5] br[5] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_8 
+ bl[6] br[6] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_9 
+ bl[7] br[7] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_10 
+ bl[8] br[8] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_11 
+ bl[9] br[9] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_12 
+ bl[10] br[10] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_13 
+ bl[11] br[11] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_14 
+ bl[12] br[12] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_15 
+ bl[13] br[13] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_16 
+ bl[14] br[14] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_17 
+ bl[15] br[15] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_18 
+ bl[16] br[16] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_19 
+ bl[17] br[17] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_20 
+ bl[18] br[18] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_21 
+ bl[19] br[19] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_22 
+ bl[20] br[20] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_23 
+ bl[21] br[21] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_24 
+ bl[22] br[22] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_25 
+ bl[23] br[23] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_26 
+ bl[24] br[24] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_27 
+ bl[25] br[25] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_28 
+ bl[26] br[26] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_29 
+ bl[27] br[27] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_30 
+ bl[28] br[28] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_31 
+ bl[29] br[29] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_32 
+ bl[30] br[30] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_33 
+ bl[31] br[31] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_34 
+ bl[32] br[32] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_35 
+ bl[33] br[33] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_36 
+ bl[34] br[34] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_37 
+ bl[35] br[35] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_38 
+ bl[36] br[36] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_39 
+ bl[37] br[37] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_40 
+ bl[38] br[38] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_41 
+ bl[39] br[39] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_42 
+ bl[40] br[40] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_43 
+ bl[41] br[41] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_44 
+ bl[42] br[42] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_45 
+ bl[43] br[43] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_46 
+ bl[44] br[44] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_47 
+ bl[45] br[45] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_48 
+ bl[46] br[46] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_49 
+ bl[47] br[47] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_50 
+ bl[48] br[48] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_51 
+ bl[49] br[49] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_52 
+ bl[50] br[50] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_53 
+ bl[51] br[51] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_54 
+ bl[52] br[52] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_55 
+ bl[53] br[53] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_56 
+ bl[54] br[54] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_57 
+ bl[55] br[55] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_58 
+ bl[56] br[56] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_59 
+ bl[57] br[57] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_60 
+ bl[58] br[58] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_61 
+ bl[59] br[59] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_62 
+ bl[60] br[60] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_63 
+ bl[61] br[61] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_64 
+ bl[62] br[62] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_65 
+ bl[63] br[63] vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_66 
+ vdd vdd vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_414_67 
+ vdd vdd vdd vss wl[412] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_0 
+ vdd vdd vss vdd vpb vnb wl[413] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_415_1 
+ rbl rbr vss vdd vpb vnb wl[413] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_415_2 
+ bl[0] br[0] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_3 
+ bl[1] br[1] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_4 
+ bl[2] br[2] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_5 
+ bl[3] br[3] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_6 
+ bl[4] br[4] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_7 
+ bl[5] br[5] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_8 
+ bl[6] br[6] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_9 
+ bl[7] br[7] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_10 
+ bl[8] br[8] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_11 
+ bl[9] br[9] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_12 
+ bl[10] br[10] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_13 
+ bl[11] br[11] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_14 
+ bl[12] br[12] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_15 
+ bl[13] br[13] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_16 
+ bl[14] br[14] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_17 
+ bl[15] br[15] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_18 
+ bl[16] br[16] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_19 
+ bl[17] br[17] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_20 
+ bl[18] br[18] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_21 
+ bl[19] br[19] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_22 
+ bl[20] br[20] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_23 
+ bl[21] br[21] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_24 
+ bl[22] br[22] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_25 
+ bl[23] br[23] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_26 
+ bl[24] br[24] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_27 
+ bl[25] br[25] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_28 
+ bl[26] br[26] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_29 
+ bl[27] br[27] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_30 
+ bl[28] br[28] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_31 
+ bl[29] br[29] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_32 
+ bl[30] br[30] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_33 
+ bl[31] br[31] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_34 
+ bl[32] br[32] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_35 
+ bl[33] br[33] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_36 
+ bl[34] br[34] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_37 
+ bl[35] br[35] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_38 
+ bl[36] br[36] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_39 
+ bl[37] br[37] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_40 
+ bl[38] br[38] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_41 
+ bl[39] br[39] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_42 
+ bl[40] br[40] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_43 
+ bl[41] br[41] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_44 
+ bl[42] br[42] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_45 
+ bl[43] br[43] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_46 
+ bl[44] br[44] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_47 
+ bl[45] br[45] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_48 
+ bl[46] br[46] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_49 
+ bl[47] br[47] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_50 
+ bl[48] br[48] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_51 
+ bl[49] br[49] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_52 
+ bl[50] br[50] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_53 
+ bl[51] br[51] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_54 
+ bl[52] br[52] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_55 
+ bl[53] br[53] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_56 
+ bl[54] br[54] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_57 
+ bl[55] br[55] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_58 
+ bl[56] br[56] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_59 
+ bl[57] br[57] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_60 
+ bl[58] br[58] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_61 
+ bl[59] br[59] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_62 
+ bl[60] br[60] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_63 
+ bl[61] br[61] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_64 
+ bl[62] br[62] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_65 
+ bl[63] br[63] vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_66 
+ vdd vdd vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_415_67 
+ vdd vdd vdd vss wl[413] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_0 
+ vdd vdd vss vdd vpb vnb wl[414] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_416_1 
+ rbl rbr vss vdd vpb vnb wl[414] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_416_2 
+ bl[0] br[0] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_3 
+ bl[1] br[1] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_4 
+ bl[2] br[2] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_5 
+ bl[3] br[3] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_6 
+ bl[4] br[4] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_7 
+ bl[5] br[5] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_8 
+ bl[6] br[6] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_9 
+ bl[7] br[7] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_10 
+ bl[8] br[8] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_11 
+ bl[9] br[9] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_12 
+ bl[10] br[10] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_13 
+ bl[11] br[11] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_14 
+ bl[12] br[12] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_15 
+ bl[13] br[13] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_16 
+ bl[14] br[14] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_17 
+ bl[15] br[15] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_18 
+ bl[16] br[16] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_19 
+ bl[17] br[17] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_20 
+ bl[18] br[18] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_21 
+ bl[19] br[19] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_22 
+ bl[20] br[20] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_23 
+ bl[21] br[21] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_24 
+ bl[22] br[22] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_25 
+ bl[23] br[23] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_26 
+ bl[24] br[24] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_27 
+ bl[25] br[25] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_28 
+ bl[26] br[26] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_29 
+ bl[27] br[27] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_30 
+ bl[28] br[28] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_31 
+ bl[29] br[29] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_32 
+ bl[30] br[30] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_33 
+ bl[31] br[31] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_34 
+ bl[32] br[32] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_35 
+ bl[33] br[33] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_36 
+ bl[34] br[34] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_37 
+ bl[35] br[35] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_38 
+ bl[36] br[36] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_39 
+ bl[37] br[37] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_40 
+ bl[38] br[38] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_41 
+ bl[39] br[39] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_42 
+ bl[40] br[40] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_43 
+ bl[41] br[41] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_44 
+ bl[42] br[42] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_45 
+ bl[43] br[43] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_46 
+ bl[44] br[44] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_47 
+ bl[45] br[45] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_48 
+ bl[46] br[46] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_49 
+ bl[47] br[47] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_50 
+ bl[48] br[48] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_51 
+ bl[49] br[49] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_52 
+ bl[50] br[50] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_53 
+ bl[51] br[51] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_54 
+ bl[52] br[52] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_55 
+ bl[53] br[53] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_56 
+ bl[54] br[54] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_57 
+ bl[55] br[55] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_58 
+ bl[56] br[56] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_59 
+ bl[57] br[57] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_60 
+ bl[58] br[58] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_61 
+ bl[59] br[59] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_62 
+ bl[60] br[60] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_63 
+ bl[61] br[61] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_64 
+ bl[62] br[62] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_65 
+ bl[63] br[63] vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_66 
+ vdd vdd vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_416_67 
+ vdd vdd vdd vss wl[414] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_0 
+ vdd vdd vss vdd vpb vnb wl[415] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_417_1 
+ rbl rbr vss vdd vpb vnb wl[415] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_417_2 
+ bl[0] br[0] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_3 
+ bl[1] br[1] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_4 
+ bl[2] br[2] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_5 
+ bl[3] br[3] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_6 
+ bl[4] br[4] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_7 
+ bl[5] br[5] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_8 
+ bl[6] br[6] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_9 
+ bl[7] br[7] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_10 
+ bl[8] br[8] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_11 
+ bl[9] br[9] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_12 
+ bl[10] br[10] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_13 
+ bl[11] br[11] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_14 
+ bl[12] br[12] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_15 
+ bl[13] br[13] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_16 
+ bl[14] br[14] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_17 
+ bl[15] br[15] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_18 
+ bl[16] br[16] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_19 
+ bl[17] br[17] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_20 
+ bl[18] br[18] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_21 
+ bl[19] br[19] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_22 
+ bl[20] br[20] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_23 
+ bl[21] br[21] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_24 
+ bl[22] br[22] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_25 
+ bl[23] br[23] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_26 
+ bl[24] br[24] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_27 
+ bl[25] br[25] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_28 
+ bl[26] br[26] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_29 
+ bl[27] br[27] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_30 
+ bl[28] br[28] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_31 
+ bl[29] br[29] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_32 
+ bl[30] br[30] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_33 
+ bl[31] br[31] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_34 
+ bl[32] br[32] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_35 
+ bl[33] br[33] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_36 
+ bl[34] br[34] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_37 
+ bl[35] br[35] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_38 
+ bl[36] br[36] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_39 
+ bl[37] br[37] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_40 
+ bl[38] br[38] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_41 
+ bl[39] br[39] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_42 
+ bl[40] br[40] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_43 
+ bl[41] br[41] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_44 
+ bl[42] br[42] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_45 
+ bl[43] br[43] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_46 
+ bl[44] br[44] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_47 
+ bl[45] br[45] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_48 
+ bl[46] br[46] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_49 
+ bl[47] br[47] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_50 
+ bl[48] br[48] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_51 
+ bl[49] br[49] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_52 
+ bl[50] br[50] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_53 
+ bl[51] br[51] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_54 
+ bl[52] br[52] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_55 
+ bl[53] br[53] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_56 
+ bl[54] br[54] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_57 
+ bl[55] br[55] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_58 
+ bl[56] br[56] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_59 
+ bl[57] br[57] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_60 
+ bl[58] br[58] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_61 
+ bl[59] br[59] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_62 
+ bl[60] br[60] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_63 
+ bl[61] br[61] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_64 
+ bl[62] br[62] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_65 
+ bl[63] br[63] vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_66 
+ vdd vdd vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_417_67 
+ vdd vdd vdd vss wl[415] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_0 
+ vdd vdd vss vdd vpb vnb wl[416] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_418_1 
+ rbl rbr vss vdd vpb vnb wl[416] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_418_2 
+ bl[0] br[0] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_3 
+ bl[1] br[1] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_4 
+ bl[2] br[2] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_5 
+ bl[3] br[3] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_6 
+ bl[4] br[4] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_7 
+ bl[5] br[5] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_8 
+ bl[6] br[6] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_9 
+ bl[7] br[7] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_10 
+ bl[8] br[8] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_11 
+ bl[9] br[9] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_12 
+ bl[10] br[10] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_13 
+ bl[11] br[11] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_14 
+ bl[12] br[12] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_15 
+ bl[13] br[13] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_16 
+ bl[14] br[14] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_17 
+ bl[15] br[15] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_18 
+ bl[16] br[16] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_19 
+ bl[17] br[17] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_20 
+ bl[18] br[18] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_21 
+ bl[19] br[19] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_22 
+ bl[20] br[20] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_23 
+ bl[21] br[21] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_24 
+ bl[22] br[22] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_25 
+ bl[23] br[23] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_26 
+ bl[24] br[24] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_27 
+ bl[25] br[25] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_28 
+ bl[26] br[26] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_29 
+ bl[27] br[27] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_30 
+ bl[28] br[28] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_31 
+ bl[29] br[29] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_32 
+ bl[30] br[30] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_33 
+ bl[31] br[31] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_34 
+ bl[32] br[32] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_35 
+ bl[33] br[33] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_36 
+ bl[34] br[34] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_37 
+ bl[35] br[35] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_38 
+ bl[36] br[36] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_39 
+ bl[37] br[37] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_40 
+ bl[38] br[38] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_41 
+ bl[39] br[39] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_42 
+ bl[40] br[40] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_43 
+ bl[41] br[41] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_44 
+ bl[42] br[42] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_45 
+ bl[43] br[43] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_46 
+ bl[44] br[44] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_47 
+ bl[45] br[45] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_48 
+ bl[46] br[46] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_49 
+ bl[47] br[47] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_50 
+ bl[48] br[48] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_51 
+ bl[49] br[49] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_52 
+ bl[50] br[50] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_53 
+ bl[51] br[51] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_54 
+ bl[52] br[52] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_55 
+ bl[53] br[53] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_56 
+ bl[54] br[54] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_57 
+ bl[55] br[55] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_58 
+ bl[56] br[56] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_59 
+ bl[57] br[57] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_60 
+ bl[58] br[58] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_61 
+ bl[59] br[59] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_62 
+ bl[60] br[60] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_63 
+ bl[61] br[61] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_64 
+ bl[62] br[62] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_65 
+ bl[63] br[63] vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_66 
+ vdd vdd vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_418_67 
+ vdd vdd vdd vss wl[416] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_0 
+ vdd vdd vss vdd vpb vnb wl[417] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_419_1 
+ rbl rbr vss vdd vpb vnb wl[417] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_419_2 
+ bl[0] br[0] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_3 
+ bl[1] br[1] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_4 
+ bl[2] br[2] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_5 
+ bl[3] br[3] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_6 
+ bl[4] br[4] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_7 
+ bl[5] br[5] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_8 
+ bl[6] br[6] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_9 
+ bl[7] br[7] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_10 
+ bl[8] br[8] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_11 
+ bl[9] br[9] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_12 
+ bl[10] br[10] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_13 
+ bl[11] br[11] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_14 
+ bl[12] br[12] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_15 
+ bl[13] br[13] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_16 
+ bl[14] br[14] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_17 
+ bl[15] br[15] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_18 
+ bl[16] br[16] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_19 
+ bl[17] br[17] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_20 
+ bl[18] br[18] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_21 
+ bl[19] br[19] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_22 
+ bl[20] br[20] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_23 
+ bl[21] br[21] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_24 
+ bl[22] br[22] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_25 
+ bl[23] br[23] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_26 
+ bl[24] br[24] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_27 
+ bl[25] br[25] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_28 
+ bl[26] br[26] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_29 
+ bl[27] br[27] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_30 
+ bl[28] br[28] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_31 
+ bl[29] br[29] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_32 
+ bl[30] br[30] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_33 
+ bl[31] br[31] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_34 
+ bl[32] br[32] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_35 
+ bl[33] br[33] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_36 
+ bl[34] br[34] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_37 
+ bl[35] br[35] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_38 
+ bl[36] br[36] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_39 
+ bl[37] br[37] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_40 
+ bl[38] br[38] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_41 
+ bl[39] br[39] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_42 
+ bl[40] br[40] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_43 
+ bl[41] br[41] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_44 
+ bl[42] br[42] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_45 
+ bl[43] br[43] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_46 
+ bl[44] br[44] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_47 
+ bl[45] br[45] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_48 
+ bl[46] br[46] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_49 
+ bl[47] br[47] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_50 
+ bl[48] br[48] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_51 
+ bl[49] br[49] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_52 
+ bl[50] br[50] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_53 
+ bl[51] br[51] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_54 
+ bl[52] br[52] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_55 
+ bl[53] br[53] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_56 
+ bl[54] br[54] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_57 
+ bl[55] br[55] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_58 
+ bl[56] br[56] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_59 
+ bl[57] br[57] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_60 
+ bl[58] br[58] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_61 
+ bl[59] br[59] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_62 
+ bl[60] br[60] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_63 
+ bl[61] br[61] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_64 
+ bl[62] br[62] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_65 
+ bl[63] br[63] vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_66 
+ vdd vdd vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_419_67 
+ vdd vdd vdd vss wl[417] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_0 
+ vdd vdd vss vdd vpb vnb wl[418] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_420_1 
+ rbl rbr vss vdd vpb vnb wl[418] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_420_2 
+ bl[0] br[0] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_3 
+ bl[1] br[1] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_4 
+ bl[2] br[2] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_5 
+ bl[3] br[3] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_6 
+ bl[4] br[4] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_7 
+ bl[5] br[5] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_8 
+ bl[6] br[6] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_9 
+ bl[7] br[7] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_10 
+ bl[8] br[8] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_11 
+ bl[9] br[9] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_12 
+ bl[10] br[10] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_13 
+ bl[11] br[11] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_14 
+ bl[12] br[12] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_15 
+ bl[13] br[13] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_16 
+ bl[14] br[14] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_17 
+ bl[15] br[15] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_18 
+ bl[16] br[16] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_19 
+ bl[17] br[17] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_20 
+ bl[18] br[18] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_21 
+ bl[19] br[19] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_22 
+ bl[20] br[20] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_23 
+ bl[21] br[21] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_24 
+ bl[22] br[22] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_25 
+ bl[23] br[23] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_26 
+ bl[24] br[24] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_27 
+ bl[25] br[25] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_28 
+ bl[26] br[26] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_29 
+ bl[27] br[27] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_30 
+ bl[28] br[28] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_31 
+ bl[29] br[29] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_32 
+ bl[30] br[30] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_33 
+ bl[31] br[31] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_34 
+ bl[32] br[32] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_35 
+ bl[33] br[33] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_36 
+ bl[34] br[34] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_37 
+ bl[35] br[35] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_38 
+ bl[36] br[36] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_39 
+ bl[37] br[37] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_40 
+ bl[38] br[38] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_41 
+ bl[39] br[39] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_42 
+ bl[40] br[40] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_43 
+ bl[41] br[41] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_44 
+ bl[42] br[42] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_45 
+ bl[43] br[43] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_46 
+ bl[44] br[44] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_47 
+ bl[45] br[45] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_48 
+ bl[46] br[46] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_49 
+ bl[47] br[47] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_50 
+ bl[48] br[48] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_51 
+ bl[49] br[49] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_52 
+ bl[50] br[50] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_53 
+ bl[51] br[51] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_54 
+ bl[52] br[52] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_55 
+ bl[53] br[53] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_56 
+ bl[54] br[54] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_57 
+ bl[55] br[55] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_58 
+ bl[56] br[56] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_59 
+ bl[57] br[57] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_60 
+ bl[58] br[58] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_61 
+ bl[59] br[59] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_62 
+ bl[60] br[60] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_63 
+ bl[61] br[61] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_64 
+ bl[62] br[62] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_65 
+ bl[63] br[63] vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_66 
+ vdd vdd vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_420_67 
+ vdd vdd vdd vss wl[418] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_0 
+ vdd vdd vss vdd vpb vnb wl[419] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_421_1 
+ rbl rbr vss vdd vpb vnb wl[419] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_421_2 
+ bl[0] br[0] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_3 
+ bl[1] br[1] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_4 
+ bl[2] br[2] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_5 
+ bl[3] br[3] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_6 
+ bl[4] br[4] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_7 
+ bl[5] br[5] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_8 
+ bl[6] br[6] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_9 
+ bl[7] br[7] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_10 
+ bl[8] br[8] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_11 
+ bl[9] br[9] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_12 
+ bl[10] br[10] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_13 
+ bl[11] br[11] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_14 
+ bl[12] br[12] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_15 
+ bl[13] br[13] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_16 
+ bl[14] br[14] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_17 
+ bl[15] br[15] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_18 
+ bl[16] br[16] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_19 
+ bl[17] br[17] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_20 
+ bl[18] br[18] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_21 
+ bl[19] br[19] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_22 
+ bl[20] br[20] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_23 
+ bl[21] br[21] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_24 
+ bl[22] br[22] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_25 
+ bl[23] br[23] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_26 
+ bl[24] br[24] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_27 
+ bl[25] br[25] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_28 
+ bl[26] br[26] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_29 
+ bl[27] br[27] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_30 
+ bl[28] br[28] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_31 
+ bl[29] br[29] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_32 
+ bl[30] br[30] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_33 
+ bl[31] br[31] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_34 
+ bl[32] br[32] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_35 
+ bl[33] br[33] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_36 
+ bl[34] br[34] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_37 
+ bl[35] br[35] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_38 
+ bl[36] br[36] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_39 
+ bl[37] br[37] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_40 
+ bl[38] br[38] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_41 
+ bl[39] br[39] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_42 
+ bl[40] br[40] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_43 
+ bl[41] br[41] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_44 
+ bl[42] br[42] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_45 
+ bl[43] br[43] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_46 
+ bl[44] br[44] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_47 
+ bl[45] br[45] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_48 
+ bl[46] br[46] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_49 
+ bl[47] br[47] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_50 
+ bl[48] br[48] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_51 
+ bl[49] br[49] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_52 
+ bl[50] br[50] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_53 
+ bl[51] br[51] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_54 
+ bl[52] br[52] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_55 
+ bl[53] br[53] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_56 
+ bl[54] br[54] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_57 
+ bl[55] br[55] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_58 
+ bl[56] br[56] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_59 
+ bl[57] br[57] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_60 
+ bl[58] br[58] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_61 
+ bl[59] br[59] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_62 
+ bl[60] br[60] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_63 
+ bl[61] br[61] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_64 
+ bl[62] br[62] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_65 
+ bl[63] br[63] vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_66 
+ vdd vdd vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_421_67 
+ vdd vdd vdd vss wl[419] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_0 
+ vdd vdd vss vdd vpb vnb wl[420] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_422_1 
+ rbl rbr vss vdd vpb vnb wl[420] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_422_2 
+ bl[0] br[0] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_3 
+ bl[1] br[1] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_4 
+ bl[2] br[2] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_5 
+ bl[3] br[3] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_6 
+ bl[4] br[4] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_7 
+ bl[5] br[5] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_8 
+ bl[6] br[6] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_9 
+ bl[7] br[7] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_10 
+ bl[8] br[8] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_11 
+ bl[9] br[9] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_12 
+ bl[10] br[10] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_13 
+ bl[11] br[11] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_14 
+ bl[12] br[12] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_15 
+ bl[13] br[13] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_16 
+ bl[14] br[14] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_17 
+ bl[15] br[15] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_18 
+ bl[16] br[16] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_19 
+ bl[17] br[17] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_20 
+ bl[18] br[18] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_21 
+ bl[19] br[19] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_22 
+ bl[20] br[20] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_23 
+ bl[21] br[21] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_24 
+ bl[22] br[22] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_25 
+ bl[23] br[23] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_26 
+ bl[24] br[24] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_27 
+ bl[25] br[25] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_28 
+ bl[26] br[26] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_29 
+ bl[27] br[27] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_30 
+ bl[28] br[28] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_31 
+ bl[29] br[29] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_32 
+ bl[30] br[30] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_33 
+ bl[31] br[31] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_34 
+ bl[32] br[32] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_35 
+ bl[33] br[33] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_36 
+ bl[34] br[34] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_37 
+ bl[35] br[35] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_38 
+ bl[36] br[36] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_39 
+ bl[37] br[37] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_40 
+ bl[38] br[38] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_41 
+ bl[39] br[39] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_42 
+ bl[40] br[40] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_43 
+ bl[41] br[41] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_44 
+ bl[42] br[42] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_45 
+ bl[43] br[43] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_46 
+ bl[44] br[44] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_47 
+ bl[45] br[45] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_48 
+ bl[46] br[46] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_49 
+ bl[47] br[47] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_50 
+ bl[48] br[48] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_51 
+ bl[49] br[49] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_52 
+ bl[50] br[50] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_53 
+ bl[51] br[51] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_54 
+ bl[52] br[52] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_55 
+ bl[53] br[53] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_56 
+ bl[54] br[54] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_57 
+ bl[55] br[55] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_58 
+ bl[56] br[56] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_59 
+ bl[57] br[57] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_60 
+ bl[58] br[58] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_61 
+ bl[59] br[59] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_62 
+ bl[60] br[60] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_63 
+ bl[61] br[61] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_64 
+ bl[62] br[62] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_65 
+ bl[63] br[63] vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_66 
+ vdd vdd vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_422_67 
+ vdd vdd vdd vss wl[420] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_0 
+ vdd vdd vss vdd vpb vnb wl[421] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_423_1 
+ rbl rbr vss vdd vpb vnb wl[421] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_423_2 
+ bl[0] br[0] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_3 
+ bl[1] br[1] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_4 
+ bl[2] br[2] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_5 
+ bl[3] br[3] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_6 
+ bl[4] br[4] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_7 
+ bl[5] br[5] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_8 
+ bl[6] br[6] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_9 
+ bl[7] br[7] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_10 
+ bl[8] br[8] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_11 
+ bl[9] br[9] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_12 
+ bl[10] br[10] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_13 
+ bl[11] br[11] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_14 
+ bl[12] br[12] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_15 
+ bl[13] br[13] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_16 
+ bl[14] br[14] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_17 
+ bl[15] br[15] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_18 
+ bl[16] br[16] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_19 
+ bl[17] br[17] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_20 
+ bl[18] br[18] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_21 
+ bl[19] br[19] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_22 
+ bl[20] br[20] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_23 
+ bl[21] br[21] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_24 
+ bl[22] br[22] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_25 
+ bl[23] br[23] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_26 
+ bl[24] br[24] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_27 
+ bl[25] br[25] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_28 
+ bl[26] br[26] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_29 
+ bl[27] br[27] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_30 
+ bl[28] br[28] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_31 
+ bl[29] br[29] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_32 
+ bl[30] br[30] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_33 
+ bl[31] br[31] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_34 
+ bl[32] br[32] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_35 
+ bl[33] br[33] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_36 
+ bl[34] br[34] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_37 
+ bl[35] br[35] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_38 
+ bl[36] br[36] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_39 
+ bl[37] br[37] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_40 
+ bl[38] br[38] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_41 
+ bl[39] br[39] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_42 
+ bl[40] br[40] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_43 
+ bl[41] br[41] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_44 
+ bl[42] br[42] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_45 
+ bl[43] br[43] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_46 
+ bl[44] br[44] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_47 
+ bl[45] br[45] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_48 
+ bl[46] br[46] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_49 
+ bl[47] br[47] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_50 
+ bl[48] br[48] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_51 
+ bl[49] br[49] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_52 
+ bl[50] br[50] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_53 
+ bl[51] br[51] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_54 
+ bl[52] br[52] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_55 
+ bl[53] br[53] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_56 
+ bl[54] br[54] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_57 
+ bl[55] br[55] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_58 
+ bl[56] br[56] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_59 
+ bl[57] br[57] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_60 
+ bl[58] br[58] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_61 
+ bl[59] br[59] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_62 
+ bl[60] br[60] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_63 
+ bl[61] br[61] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_64 
+ bl[62] br[62] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_65 
+ bl[63] br[63] vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_66 
+ vdd vdd vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_423_67 
+ vdd vdd vdd vss wl[421] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_0 
+ vdd vdd vss vdd vpb vnb wl[422] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_424_1 
+ rbl rbr vss vdd vpb vnb wl[422] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_424_2 
+ bl[0] br[0] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_3 
+ bl[1] br[1] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_4 
+ bl[2] br[2] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_5 
+ bl[3] br[3] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_6 
+ bl[4] br[4] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_7 
+ bl[5] br[5] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_8 
+ bl[6] br[6] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_9 
+ bl[7] br[7] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_10 
+ bl[8] br[8] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_11 
+ bl[9] br[9] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_12 
+ bl[10] br[10] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_13 
+ bl[11] br[11] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_14 
+ bl[12] br[12] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_15 
+ bl[13] br[13] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_16 
+ bl[14] br[14] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_17 
+ bl[15] br[15] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_18 
+ bl[16] br[16] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_19 
+ bl[17] br[17] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_20 
+ bl[18] br[18] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_21 
+ bl[19] br[19] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_22 
+ bl[20] br[20] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_23 
+ bl[21] br[21] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_24 
+ bl[22] br[22] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_25 
+ bl[23] br[23] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_26 
+ bl[24] br[24] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_27 
+ bl[25] br[25] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_28 
+ bl[26] br[26] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_29 
+ bl[27] br[27] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_30 
+ bl[28] br[28] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_31 
+ bl[29] br[29] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_32 
+ bl[30] br[30] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_33 
+ bl[31] br[31] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_34 
+ bl[32] br[32] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_35 
+ bl[33] br[33] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_36 
+ bl[34] br[34] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_37 
+ bl[35] br[35] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_38 
+ bl[36] br[36] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_39 
+ bl[37] br[37] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_40 
+ bl[38] br[38] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_41 
+ bl[39] br[39] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_42 
+ bl[40] br[40] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_43 
+ bl[41] br[41] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_44 
+ bl[42] br[42] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_45 
+ bl[43] br[43] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_46 
+ bl[44] br[44] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_47 
+ bl[45] br[45] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_48 
+ bl[46] br[46] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_49 
+ bl[47] br[47] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_50 
+ bl[48] br[48] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_51 
+ bl[49] br[49] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_52 
+ bl[50] br[50] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_53 
+ bl[51] br[51] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_54 
+ bl[52] br[52] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_55 
+ bl[53] br[53] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_56 
+ bl[54] br[54] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_57 
+ bl[55] br[55] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_58 
+ bl[56] br[56] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_59 
+ bl[57] br[57] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_60 
+ bl[58] br[58] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_61 
+ bl[59] br[59] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_62 
+ bl[60] br[60] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_63 
+ bl[61] br[61] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_64 
+ bl[62] br[62] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_65 
+ bl[63] br[63] vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_66 
+ vdd vdd vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_424_67 
+ vdd vdd vdd vss wl[422] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_0 
+ vdd vdd vss vdd vpb vnb wl[423] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_425_1 
+ rbl rbr vss vdd vpb vnb wl[423] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_425_2 
+ bl[0] br[0] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_3 
+ bl[1] br[1] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_4 
+ bl[2] br[2] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_5 
+ bl[3] br[3] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_6 
+ bl[4] br[4] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_7 
+ bl[5] br[5] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_8 
+ bl[6] br[6] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_9 
+ bl[7] br[7] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_10 
+ bl[8] br[8] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_11 
+ bl[9] br[9] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_12 
+ bl[10] br[10] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_13 
+ bl[11] br[11] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_14 
+ bl[12] br[12] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_15 
+ bl[13] br[13] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_16 
+ bl[14] br[14] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_17 
+ bl[15] br[15] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_18 
+ bl[16] br[16] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_19 
+ bl[17] br[17] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_20 
+ bl[18] br[18] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_21 
+ bl[19] br[19] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_22 
+ bl[20] br[20] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_23 
+ bl[21] br[21] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_24 
+ bl[22] br[22] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_25 
+ bl[23] br[23] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_26 
+ bl[24] br[24] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_27 
+ bl[25] br[25] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_28 
+ bl[26] br[26] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_29 
+ bl[27] br[27] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_30 
+ bl[28] br[28] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_31 
+ bl[29] br[29] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_32 
+ bl[30] br[30] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_33 
+ bl[31] br[31] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_34 
+ bl[32] br[32] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_35 
+ bl[33] br[33] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_36 
+ bl[34] br[34] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_37 
+ bl[35] br[35] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_38 
+ bl[36] br[36] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_39 
+ bl[37] br[37] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_40 
+ bl[38] br[38] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_41 
+ bl[39] br[39] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_42 
+ bl[40] br[40] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_43 
+ bl[41] br[41] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_44 
+ bl[42] br[42] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_45 
+ bl[43] br[43] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_46 
+ bl[44] br[44] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_47 
+ bl[45] br[45] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_48 
+ bl[46] br[46] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_49 
+ bl[47] br[47] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_50 
+ bl[48] br[48] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_51 
+ bl[49] br[49] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_52 
+ bl[50] br[50] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_53 
+ bl[51] br[51] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_54 
+ bl[52] br[52] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_55 
+ bl[53] br[53] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_56 
+ bl[54] br[54] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_57 
+ bl[55] br[55] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_58 
+ bl[56] br[56] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_59 
+ bl[57] br[57] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_60 
+ bl[58] br[58] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_61 
+ bl[59] br[59] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_62 
+ bl[60] br[60] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_63 
+ bl[61] br[61] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_64 
+ bl[62] br[62] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_65 
+ bl[63] br[63] vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_66 
+ vdd vdd vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_425_67 
+ vdd vdd vdd vss wl[423] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_0 
+ vdd vdd vss vdd vpb vnb wl[424] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_426_1 
+ rbl rbr vss vdd vpb vnb wl[424] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_426_2 
+ bl[0] br[0] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_3 
+ bl[1] br[1] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_4 
+ bl[2] br[2] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_5 
+ bl[3] br[3] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_6 
+ bl[4] br[4] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_7 
+ bl[5] br[5] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_8 
+ bl[6] br[6] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_9 
+ bl[7] br[7] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_10 
+ bl[8] br[8] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_11 
+ bl[9] br[9] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_12 
+ bl[10] br[10] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_13 
+ bl[11] br[11] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_14 
+ bl[12] br[12] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_15 
+ bl[13] br[13] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_16 
+ bl[14] br[14] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_17 
+ bl[15] br[15] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_18 
+ bl[16] br[16] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_19 
+ bl[17] br[17] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_20 
+ bl[18] br[18] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_21 
+ bl[19] br[19] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_22 
+ bl[20] br[20] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_23 
+ bl[21] br[21] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_24 
+ bl[22] br[22] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_25 
+ bl[23] br[23] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_26 
+ bl[24] br[24] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_27 
+ bl[25] br[25] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_28 
+ bl[26] br[26] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_29 
+ bl[27] br[27] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_30 
+ bl[28] br[28] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_31 
+ bl[29] br[29] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_32 
+ bl[30] br[30] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_33 
+ bl[31] br[31] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_34 
+ bl[32] br[32] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_35 
+ bl[33] br[33] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_36 
+ bl[34] br[34] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_37 
+ bl[35] br[35] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_38 
+ bl[36] br[36] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_39 
+ bl[37] br[37] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_40 
+ bl[38] br[38] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_41 
+ bl[39] br[39] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_42 
+ bl[40] br[40] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_43 
+ bl[41] br[41] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_44 
+ bl[42] br[42] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_45 
+ bl[43] br[43] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_46 
+ bl[44] br[44] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_47 
+ bl[45] br[45] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_48 
+ bl[46] br[46] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_49 
+ bl[47] br[47] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_50 
+ bl[48] br[48] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_51 
+ bl[49] br[49] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_52 
+ bl[50] br[50] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_53 
+ bl[51] br[51] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_54 
+ bl[52] br[52] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_55 
+ bl[53] br[53] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_56 
+ bl[54] br[54] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_57 
+ bl[55] br[55] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_58 
+ bl[56] br[56] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_59 
+ bl[57] br[57] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_60 
+ bl[58] br[58] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_61 
+ bl[59] br[59] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_62 
+ bl[60] br[60] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_63 
+ bl[61] br[61] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_64 
+ bl[62] br[62] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_65 
+ bl[63] br[63] vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_66 
+ vdd vdd vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_426_67 
+ vdd vdd vdd vss wl[424] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_0 
+ vdd vdd vss vdd vpb vnb wl[425] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_427_1 
+ rbl rbr vss vdd vpb vnb wl[425] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_427_2 
+ bl[0] br[0] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_3 
+ bl[1] br[1] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_4 
+ bl[2] br[2] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_5 
+ bl[3] br[3] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_6 
+ bl[4] br[4] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_7 
+ bl[5] br[5] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_8 
+ bl[6] br[6] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_9 
+ bl[7] br[7] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_10 
+ bl[8] br[8] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_11 
+ bl[9] br[9] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_12 
+ bl[10] br[10] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_13 
+ bl[11] br[11] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_14 
+ bl[12] br[12] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_15 
+ bl[13] br[13] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_16 
+ bl[14] br[14] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_17 
+ bl[15] br[15] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_18 
+ bl[16] br[16] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_19 
+ bl[17] br[17] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_20 
+ bl[18] br[18] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_21 
+ bl[19] br[19] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_22 
+ bl[20] br[20] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_23 
+ bl[21] br[21] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_24 
+ bl[22] br[22] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_25 
+ bl[23] br[23] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_26 
+ bl[24] br[24] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_27 
+ bl[25] br[25] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_28 
+ bl[26] br[26] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_29 
+ bl[27] br[27] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_30 
+ bl[28] br[28] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_31 
+ bl[29] br[29] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_32 
+ bl[30] br[30] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_33 
+ bl[31] br[31] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_34 
+ bl[32] br[32] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_35 
+ bl[33] br[33] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_36 
+ bl[34] br[34] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_37 
+ bl[35] br[35] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_38 
+ bl[36] br[36] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_39 
+ bl[37] br[37] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_40 
+ bl[38] br[38] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_41 
+ bl[39] br[39] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_42 
+ bl[40] br[40] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_43 
+ bl[41] br[41] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_44 
+ bl[42] br[42] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_45 
+ bl[43] br[43] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_46 
+ bl[44] br[44] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_47 
+ bl[45] br[45] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_48 
+ bl[46] br[46] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_49 
+ bl[47] br[47] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_50 
+ bl[48] br[48] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_51 
+ bl[49] br[49] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_52 
+ bl[50] br[50] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_53 
+ bl[51] br[51] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_54 
+ bl[52] br[52] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_55 
+ bl[53] br[53] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_56 
+ bl[54] br[54] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_57 
+ bl[55] br[55] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_58 
+ bl[56] br[56] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_59 
+ bl[57] br[57] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_60 
+ bl[58] br[58] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_61 
+ bl[59] br[59] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_62 
+ bl[60] br[60] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_63 
+ bl[61] br[61] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_64 
+ bl[62] br[62] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_65 
+ bl[63] br[63] vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_66 
+ vdd vdd vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_427_67 
+ vdd vdd vdd vss wl[425] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_0 
+ vdd vdd vss vdd vpb vnb wl[426] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_428_1 
+ rbl rbr vss vdd vpb vnb wl[426] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_428_2 
+ bl[0] br[0] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_3 
+ bl[1] br[1] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_4 
+ bl[2] br[2] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_5 
+ bl[3] br[3] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_6 
+ bl[4] br[4] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_7 
+ bl[5] br[5] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_8 
+ bl[6] br[6] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_9 
+ bl[7] br[7] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_10 
+ bl[8] br[8] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_11 
+ bl[9] br[9] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_12 
+ bl[10] br[10] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_13 
+ bl[11] br[11] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_14 
+ bl[12] br[12] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_15 
+ bl[13] br[13] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_16 
+ bl[14] br[14] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_17 
+ bl[15] br[15] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_18 
+ bl[16] br[16] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_19 
+ bl[17] br[17] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_20 
+ bl[18] br[18] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_21 
+ bl[19] br[19] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_22 
+ bl[20] br[20] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_23 
+ bl[21] br[21] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_24 
+ bl[22] br[22] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_25 
+ bl[23] br[23] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_26 
+ bl[24] br[24] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_27 
+ bl[25] br[25] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_28 
+ bl[26] br[26] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_29 
+ bl[27] br[27] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_30 
+ bl[28] br[28] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_31 
+ bl[29] br[29] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_32 
+ bl[30] br[30] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_33 
+ bl[31] br[31] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_34 
+ bl[32] br[32] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_35 
+ bl[33] br[33] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_36 
+ bl[34] br[34] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_37 
+ bl[35] br[35] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_38 
+ bl[36] br[36] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_39 
+ bl[37] br[37] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_40 
+ bl[38] br[38] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_41 
+ bl[39] br[39] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_42 
+ bl[40] br[40] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_43 
+ bl[41] br[41] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_44 
+ bl[42] br[42] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_45 
+ bl[43] br[43] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_46 
+ bl[44] br[44] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_47 
+ bl[45] br[45] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_48 
+ bl[46] br[46] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_49 
+ bl[47] br[47] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_50 
+ bl[48] br[48] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_51 
+ bl[49] br[49] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_52 
+ bl[50] br[50] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_53 
+ bl[51] br[51] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_54 
+ bl[52] br[52] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_55 
+ bl[53] br[53] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_56 
+ bl[54] br[54] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_57 
+ bl[55] br[55] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_58 
+ bl[56] br[56] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_59 
+ bl[57] br[57] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_60 
+ bl[58] br[58] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_61 
+ bl[59] br[59] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_62 
+ bl[60] br[60] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_63 
+ bl[61] br[61] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_64 
+ bl[62] br[62] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_65 
+ bl[63] br[63] vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_66 
+ vdd vdd vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_428_67 
+ vdd vdd vdd vss wl[426] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_0 
+ vdd vdd vss vdd vpb vnb wl[427] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_429_1 
+ rbl rbr vss vdd vpb vnb wl[427] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_429_2 
+ bl[0] br[0] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_3 
+ bl[1] br[1] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_4 
+ bl[2] br[2] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_5 
+ bl[3] br[3] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_6 
+ bl[4] br[4] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_7 
+ bl[5] br[5] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_8 
+ bl[6] br[6] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_9 
+ bl[7] br[7] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_10 
+ bl[8] br[8] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_11 
+ bl[9] br[9] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_12 
+ bl[10] br[10] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_13 
+ bl[11] br[11] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_14 
+ bl[12] br[12] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_15 
+ bl[13] br[13] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_16 
+ bl[14] br[14] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_17 
+ bl[15] br[15] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_18 
+ bl[16] br[16] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_19 
+ bl[17] br[17] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_20 
+ bl[18] br[18] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_21 
+ bl[19] br[19] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_22 
+ bl[20] br[20] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_23 
+ bl[21] br[21] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_24 
+ bl[22] br[22] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_25 
+ bl[23] br[23] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_26 
+ bl[24] br[24] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_27 
+ bl[25] br[25] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_28 
+ bl[26] br[26] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_29 
+ bl[27] br[27] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_30 
+ bl[28] br[28] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_31 
+ bl[29] br[29] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_32 
+ bl[30] br[30] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_33 
+ bl[31] br[31] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_34 
+ bl[32] br[32] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_35 
+ bl[33] br[33] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_36 
+ bl[34] br[34] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_37 
+ bl[35] br[35] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_38 
+ bl[36] br[36] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_39 
+ bl[37] br[37] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_40 
+ bl[38] br[38] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_41 
+ bl[39] br[39] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_42 
+ bl[40] br[40] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_43 
+ bl[41] br[41] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_44 
+ bl[42] br[42] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_45 
+ bl[43] br[43] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_46 
+ bl[44] br[44] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_47 
+ bl[45] br[45] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_48 
+ bl[46] br[46] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_49 
+ bl[47] br[47] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_50 
+ bl[48] br[48] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_51 
+ bl[49] br[49] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_52 
+ bl[50] br[50] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_53 
+ bl[51] br[51] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_54 
+ bl[52] br[52] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_55 
+ bl[53] br[53] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_56 
+ bl[54] br[54] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_57 
+ bl[55] br[55] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_58 
+ bl[56] br[56] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_59 
+ bl[57] br[57] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_60 
+ bl[58] br[58] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_61 
+ bl[59] br[59] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_62 
+ bl[60] br[60] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_63 
+ bl[61] br[61] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_64 
+ bl[62] br[62] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_65 
+ bl[63] br[63] vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_66 
+ vdd vdd vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_429_67 
+ vdd vdd vdd vss wl[427] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_0 
+ vdd vdd vss vdd vpb vnb wl[428] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_430_1 
+ rbl rbr vss vdd vpb vnb wl[428] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_430_2 
+ bl[0] br[0] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_3 
+ bl[1] br[1] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_4 
+ bl[2] br[2] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_5 
+ bl[3] br[3] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_6 
+ bl[4] br[4] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_7 
+ bl[5] br[5] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_8 
+ bl[6] br[6] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_9 
+ bl[7] br[7] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_10 
+ bl[8] br[8] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_11 
+ bl[9] br[9] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_12 
+ bl[10] br[10] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_13 
+ bl[11] br[11] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_14 
+ bl[12] br[12] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_15 
+ bl[13] br[13] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_16 
+ bl[14] br[14] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_17 
+ bl[15] br[15] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_18 
+ bl[16] br[16] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_19 
+ bl[17] br[17] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_20 
+ bl[18] br[18] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_21 
+ bl[19] br[19] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_22 
+ bl[20] br[20] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_23 
+ bl[21] br[21] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_24 
+ bl[22] br[22] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_25 
+ bl[23] br[23] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_26 
+ bl[24] br[24] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_27 
+ bl[25] br[25] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_28 
+ bl[26] br[26] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_29 
+ bl[27] br[27] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_30 
+ bl[28] br[28] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_31 
+ bl[29] br[29] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_32 
+ bl[30] br[30] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_33 
+ bl[31] br[31] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_34 
+ bl[32] br[32] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_35 
+ bl[33] br[33] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_36 
+ bl[34] br[34] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_37 
+ bl[35] br[35] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_38 
+ bl[36] br[36] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_39 
+ bl[37] br[37] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_40 
+ bl[38] br[38] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_41 
+ bl[39] br[39] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_42 
+ bl[40] br[40] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_43 
+ bl[41] br[41] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_44 
+ bl[42] br[42] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_45 
+ bl[43] br[43] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_46 
+ bl[44] br[44] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_47 
+ bl[45] br[45] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_48 
+ bl[46] br[46] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_49 
+ bl[47] br[47] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_50 
+ bl[48] br[48] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_51 
+ bl[49] br[49] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_52 
+ bl[50] br[50] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_53 
+ bl[51] br[51] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_54 
+ bl[52] br[52] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_55 
+ bl[53] br[53] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_56 
+ bl[54] br[54] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_57 
+ bl[55] br[55] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_58 
+ bl[56] br[56] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_59 
+ bl[57] br[57] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_60 
+ bl[58] br[58] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_61 
+ bl[59] br[59] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_62 
+ bl[60] br[60] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_63 
+ bl[61] br[61] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_64 
+ bl[62] br[62] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_65 
+ bl[63] br[63] vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_66 
+ vdd vdd vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_430_67 
+ vdd vdd vdd vss wl[428] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_0 
+ vdd vdd vss vdd vpb vnb wl[429] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_431_1 
+ rbl rbr vss vdd vpb vnb wl[429] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_431_2 
+ bl[0] br[0] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_3 
+ bl[1] br[1] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_4 
+ bl[2] br[2] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_5 
+ bl[3] br[3] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_6 
+ bl[4] br[4] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_7 
+ bl[5] br[5] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_8 
+ bl[6] br[6] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_9 
+ bl[7] br[7] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_10 
+ bl[8] br[8] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_11 
+ bl[9] br[9] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_12 
+ bl[10] br[10] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_13 
+ bl[11] br[11] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_14 
+ bl[12] br[12] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_15 
+ bl[13] br[13] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_16 
+ bl[14] br[14] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_17 
+ bl[15] br[15] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_18 
+ bl[16] br[16] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_19 
+ bl[17] br[17] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_20 
+ bl[18] br[18] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_21 
+ bl[19] br[19] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_22 
+ bl[20] br[20] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_23 
+ bl[21] br[21] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_24 
+ bl[22] br[22] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_25 
+ bl[23] br[23] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_26 
+ bl[24] br[24] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_27 
+ bl[25] br[25] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_28 
+ bl[26] br[26] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_29 
+ bl[27] br[27] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_30 
+ bl[28] br[28] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_31 
+ bl[29] br[29] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_32 
+ bl[30] br[30] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_33 
+ bl[31] br[31] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_34 
+ bl[32] br[32] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_35 
+ bl[33] br[33] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_36 
+ bl[34] br[34] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_37 
+ bl[35] br[35] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_38 
+ bl[36] br[36] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_39 
+ bl[37] br[37] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_40 
+ bl[38] br[38] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_41 
+ bl[39] br[39] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_42 
+ bl[40] br[40] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_43 
+ bl[41] br[41] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_44 
+ bl[42] br[42] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_45 
+ bl[43] br[43] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_46 
+ bl[44] br[44] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_47 
+ bl[45] br[45] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_48 
+ bl[46] br[46] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_49 
+ bl[47] br[47] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_50 
+ bl[48] br[48] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_51 
+ bl[49] br[49] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_52 
+ bl[50] br[50] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_53 
+ bl[51] br[51] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_54 
+ bl[52] br[52] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_55 
+ bl[53] br[53] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_56 
+ bl[54] br[54] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_57 
+ bl[55] br[55] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_58 
+ bl[56] br[56] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_59 
+ bl[57] br[57] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_60 
+ bl[58] br[58] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_61 
+ bl[59] br[59] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_62 
+ bl[60] br[60] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_63 
+ bl[61] br[61] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_64 
+ bl[62] br[62] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_65 
+ bl[63] br[63] vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_66 
+ vdd vdd vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_431_67 
+ vdd vdd vdd vss wl[429] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_0 
+ vdd vdd vss vdd vpb vnb wl[430] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_432_1 
+ rbl rbr vss vdd vpb vnb wl[430] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_432_2 
+ bl[0] br[0] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_3 
+ bl[1] br[1] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_4 
+ bl[2] br[2] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_5 
+ bl[3] br[3] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_6 
+ bl[4] br[4] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_7 
+ bl[5] br[5] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_8 
+ bl[6] br[6] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_9 
+ bl[7] br[7] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_10 
+ bl[8] br[8] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_11 
+ bl[9] br[9] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_12 
+ bl[10] br[10] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_13 
+ bl[11] br[11] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_14 
+ bl[12] br[12] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_15 
+ bl[13] br[13] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_16 
+ bl[14] br[14] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_17 
+ bl[15] br[15] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_18 
+ bl[16] br[16] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_19 
+ bl[17] br[17] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_20 
+ bl[18] br[18] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_21 
+ bl[19] br[19] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_22 
+ bl[20] br[20] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_23 
+ bl[21] br[21] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_24 
+ bl[22] br[22] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_25 
+ bl[23] br[23] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_26 
+ bl[24] br[24] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_27 
+ bl[25] br[25] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_28 
+ bl[26] br[26] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_29 
+ bl[27] br[27] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_30 
+ bl[28] br[28] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_31 
+ bl[29] br[29] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_32 
+ bl[30] br[30] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_33 
+ bl[31] br[31] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_34 
+ bl[32] br[32] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_35 
+ bl[33] br[33] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_36 
+ bl[34] br[34] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_37 
+ bl[35] br[35] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_38 
+ bl[36] br[36] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_39 
+ bl[37] br[37] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_40 
+ bl[38] br[38] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_41 
+ bl[39] br[39] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_42 
+ bl[40] br[40] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_43 
+ bl[41] br[41] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_44 
+ bl[42] br[42] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_45 
+ bl[43] br[43] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_46 
+ bl[44] br[44] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_47 
+ bl[45] br[45] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_48 
+ bl[46] br[46] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_49 
+ bl[47] br[47] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_50 
+ bl[48] br[48] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_51 
+ bl[49] br[49] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_52 
+ bl[50] br[50] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_53 
+ bl[51] br[51] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_54 
+ bl[52] br[52] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_55 
+ bl[53] br[53] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_56 
+ bl[54] br[54] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_57 
+ bl[55] br[55] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_58 
+ bl[56] br[56] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_59 
+ bl[57] br[57] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_60 
+ bl[58] br[58] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_61 
+ bl[59] br[59] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_62 
+ bl[60] br[60] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_63 
+ bl[61] br[61] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_64 
+ bl[62] br[62] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_65 
+ bl[63] br[63] vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_66 
+ vdd vdd vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_432_67 
+ vdd vdd vdd vss wl[430] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_0 
+ vdd vdd vss vdd vpb vnb wl[431] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_433_1 
+ rbl rbr vss vdd vpb vnb wl[431] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_433_2 
+ bl[0] br[0] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_3 
+ bl[1] br[1] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_4 
+ bl[2] br[2] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_5 
+ bl[3] br[3] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_6 
+ bl[4] br[4] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_7 
+ bl[5] br[5] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_8 
+ bl[6] br[6] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_9 
+ bl[7] br[7] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_10 
+ bl[8] br[8] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_11 
+ bl[9] br[9] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_12 
+ bl[10] br[10] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_13 
+ bl[11] br[11] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_14 
+ bl[12] br[12] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_15 
+ bl[13] br[13] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_16 
+ bl[14] br[14] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_17 
+ bl[15] br[15] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_18 
+ bl[16] br[16] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_19 
+ bl[17] br[17] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_20 
+ bl[18] br[18] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_21 
+ bl[19] br[19] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_22 
+ bl[20] br[20] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_23 
+ bl[21] br[21] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_24 
+ bl[22] br[22] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_25 
+ bl[23] br[23] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_26 
+ bl[24] br[24] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_27 
+ bl[25] br[25] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_28 
+ bl[26] br[26] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_29 
+ bl[27] br[27] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_30 
+ bl[28] br[28] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_31 
+ bl[29] br[29] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_32 
+ bl[30] br[30] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_33 
+ bl[31] br[31] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_34 
+ bl[32] br[32] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_35 
+ bl[33] br[33] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_36 
+ bl[34] br[34] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_37 
+ bl[35] br[35] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_38 
+ bl[36] br[36] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_39 
+ bl[37] br[37] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_40 
+ bl[38] br[38] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_41 
+ bl[39] br[39] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_42 
+ bl[40] br[40] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_43 
+ bl[41] br[41] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_44 
+ bl[42] br[42] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_45 
+ bl[43] br[43] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_46 
+ bl[44] br[44] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_47 
+ bl[45] br[45] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_48 
+ bl[46] br[46] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_49 
+ bl[47] br[47] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_50 
+ bl[48] br[48] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_51 
+ bl[49] br[49] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_52 
+ bl[50] br[50] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_53 
+ bl[51] br[51] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_54 
+ bl[52] br[52] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_55 
+ bl[53] br[53] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_56 
+ bl[54] br[54] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_57 
+ bl[55] br[55] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_58 
+ bl[56] br[56] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_59 
+ bl[57] br[57] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_60 
+ bl[58] br[58] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_61 
+ bl[59] br[59] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_62 
+ bl[60] br[60] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_63 
+ bl[61] br[61] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_64 
+ bl[62] br[62] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_65 
+ bl[63] br[63] vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_66 
+ vdd vdd vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_433_67 
+ vdd vdd vdd vss wl[431] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_0 
+ vdd vdd vss vdd vpb vnb wl[432] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_434_1 
+ rbl rbr vss vdd vpb vnb wl[432] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_434_2 
+ bl[0] br[0] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_3 
+ bl[1] br[1] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_4 
+ bl[2] br[2] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_5 
+ bl[3] br[3] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_6 
+ bl[4] br[4] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_7 
+ bl[5] br[5] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_8 
+ bl[6] br[6] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_9 
+ bl[7] br[7] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_10 
+ bl[8] br[8] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_11 
+ bl[9] br[9] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_12 
+ bl[10] br[10] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_13 
+ bl[11] br[11] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_14 
+ bl[12] br[12] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_15 
+ bl[13] br[13] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_16 
+ bl[14] br[14] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_17 
+ bl[15] br[15] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_18 
+ bl[16] br[16] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_19 
+ bl[17] br[17] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_20 
+ bl[18] br[18] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_21 
+ bl[19] br[19] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_22 
+ bl[20] br[20] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_23 
+ bl[21] br[21] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_24 
+ bl[22] br[22] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_25 
+ bl[23] br[23] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_26 
+ bl[24] br[24] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_27 
+ bl[25] br[25] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_28 
+ bl[26] br[26] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_29 
+ bl[27] br[27] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_30 
+ bl[28] br[28] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_31 
+ bl[29] br[29] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_32 
+ bl[30] br[30] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_33 
+ bl[31] br[31] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_34 
+ bl[32] br[32] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_35 
+ bl[33] br[33] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_36 
+ bl[34] br[34] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_37 
+ bl[35] br[35] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_38 
+ bl[36] br[36] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_39 
+ bl[37] br[37] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_40 
+ bl[38] br[38] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_41 
+ bl[39] br[39] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_42 
+ bl[40] br[40] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_43 
+ bl[41] br[41] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_44 
+ bl[42] br[42] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_45 
+ bl[43] br[43] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_46 
+ bl[44] br[44] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_47 
+ bl[45] br[45] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_48 
+ bl[46] br[46] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_49 
+ bl[47] br[47] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_50 
+ bl[48] br[48] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_51 
+ bl[49] br[49] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_52 
+ bl[50] br[50] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_53 
+ bl[51] br[51] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_54 
+ bl[52] br[52] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_55 
+ bl[53] br[53] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_56 
+ bl[54] br[54] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_57 
+ bl[55] br[55] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_58 
+ bl[56] br[56] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_59 
+ bl[57] br[57] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_60 
+ bl[58] br[58] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_61 
+ bl[59] br[59] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_62 
+ bl[60] br[60] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_63 
+ bl[61] br[61] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_64 
+ bl[62] br[62] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_65 
+ bl[63] br[63] vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_66 
+ vdd vdd vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_434_67 
+ vdd vdd vdd vss wl[432] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_0 
+ vdd vdd vss vdd vpb vnb wl[433] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_435_1 
+ rbl rbr vss vdd vpb vnb wl[433] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_435_2 
+ bl[0] br[0] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_3 
+ bl[1] br[1] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_4 
+ bl[2] br[2] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_5 
+ bl[3] br[3] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_6 
+ bl[4] br[4] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_7 
+ bl[5] br[5] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_8 
+ bl[6] br[6] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_9 
+ bl[7] br[7] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_10 
+ bl[8] br[8] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_11 
+ bl[9] br[9] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_12 
+ bl[10] br[10] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_13 
+ bl[11] br[11] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_14 
+ bl[12] br[12] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_15 
+ bl[13] br[13] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_16 
+ bl[14] br[14] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_17 
+ bl[15] br[15] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_18 
+ bl[16] br[16] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_19 
+ bl[17] br[17] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_20 
+ bl[18] br[18] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_21 
+ bl[19] br[19] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_22 
+ bl[20] br[20] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_23 
+ bl[21] br[21] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_24 
+ bl[22] br[22] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_25 
+ bl[23] br[23] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_26 
+ bl[24] br[24] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_27 
+ bl[25] br[25] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_28 
+ bl[26] br[26] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_29 
+ bl[27] br[27] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_30 
+ bl[28] br[28] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_31 
+ bl[29] br[29] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_32 
+ bl[30] br[30] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_33 
+ bl[31] br[31] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_34 
+ bl[32] br[32] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_35 
+ bl[33] br[33] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_36 
+ bl[34] br[34] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_37 
+ bl[35] br[35] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_38 
+ bl[36] br[36] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_39 
+ bl[37] br[37] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_40 
+ bl[38] br[38] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_41 
+ bl[39] br[39] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_42 
+ bl[40] br[40] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_43 
+ bl[41] br[41] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_44 
+ bl[42] br[42] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_45 
+ bl[43] br[43] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_46 
+ bl[44] br[44] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_47 
+ bl[45] br[45] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_48 
+ bl[46] br[46] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_49 
+ bl[47] br[47] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_50 
+ bl[48] br[48] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_51 
+ bl[49] br[49] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_52 
+ bl[50] br[50] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_53 
+ bl[51] br[51] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_54 
+ bl[52] br[52] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_55 
+ bl[53] br[53] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_56 
+ bl[54] br[54] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_57 
+ bl[55] br[55] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_58 
+ bl[56] br[56] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_59 
+ bl[57] br[57] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_60 
+ bl[58] br[58] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_61 
+ bl[59] br[59] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_62 
+ bl[60] br[60] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_63 
+ bl[61] br[61] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_64 
+ bl[62] br[62] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_65 
+ bl[63] br[63] vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_66 
+ vdd vdd vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_435_67 
+ vdd vdd vdd vss wl[433] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_0 
+ vdd vdd vss vdd vpb vnb wl[434] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_436_1 
+ rbl rbr vss vdd vpb vnb wl[434] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_436_2 
+ bl[0] br[0] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_3 
+ bl[1] br[1] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_4 
+ bl[2] br[2] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_5 
+ bl[3] br[3] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_6 
+ bl[4] br[4] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_7 
+ bl[5] br[5] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_8 
+ bl[6] br[6] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_9 
+ bl[7] br[7] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_10 
+ bl[8] br[8] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_11 
+ bl[9] br[9] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_12 
+ bl[10] br[10] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_13 
+ bl[11] br[11] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_14 
+ bl[12] br[12] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_15 
+ bl[13] br[13] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_16 
+ bl[14] br[14] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_17 
+ bl[15] br[15] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_18 
+ bl[16] br[16] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_19 
+ bl[17] br[17] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_20 
+ bl[18] br[18] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_21 
+ bl[19] br[19] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_22 
+ bl[20] br[20] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_23 
+ bl[21] br[21] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_24 
+ bl[22] br[22] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_25 
+ bl[23] br[23] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_26 
+ bl[24] br[24] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_27 
+ bl[25] br[25] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_28 
+ bl[26] br[26] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_29 
+ bl[27] br[27] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_30 
+ bl[28] br[28] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_31 
+ bl[29] br[29] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_32 
+ bl[30] br[30] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_33 
+ bl[31] br[31] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_34 
+ bl[32] br[32] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_35 
+ bl[33] br[33] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_36 
+ bl[34] br[34] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_37 
+ bl[35] br[35] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_38 
+ bl[36] br[36] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_39 
+ bl[37] br[37] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_40 
+ bl[38] br[38] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_41 
+ bl[39] br[39] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_42 
+ bl[40] br[40] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_43 
+ bl[41] br[41] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_44 
+ bl[42] br[42] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_45 
+ bl[43] br[43] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_46 
+ bl[44] br[44] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_47 
+ bl[45] br[45] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_48 
+ bl[46] br[46] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_49 
+ bl[47] br[47] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_50 
+ bl[48] br[48] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_51 
+ bl[49] br[49] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_52 
+ bl[50] br[50] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_53 
+ bl[51] br[51] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_54 
+ bl[52] br[52] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_55 
+ bl[53] br[53] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_56 
+ bl[54] br[54] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_57 
+ bl[55] br[55] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_58 
+ bl[56] br[56] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_59 
+ bl[57] br[57] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_60 
+ bl[58] br[58] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_61 
+ bl[59] br[59] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_62 
+ bl[60] br[60] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_63 
+ bl[61] br[61] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_64 
+ bl[62] br[62] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_65 
+ bl[63] br[63] vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_66 
+ vdd vdd vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_436_67 
+ vdd vdd vdd vss wl[434] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_0 
+ vdd vdd vss vdd vpb vnb wl[435] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_437_1 
+ rbl rbr vss vdd vpb vnb wl[435] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_437_2 
+ bl[0] br[0] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_3 
+ bl[1] br[1] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_4 
+ bl[2] br[2] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_5 
+ bl[3] br[3] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_6 
+ bl[4] br[4] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_7 
+ bl[5] br[5] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_8 
+ bl[6] br[6] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_9 
+ bl[7] br[7] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_10 
+ bl[8] br[8] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_11 
+ bl[9] br[9] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_12 
+ bl[10] br[10] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_13 
+ bl[11] br[11] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_14 
+ bl[12] br[12] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_15 
+ bl[13] br[13] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_16 
+ bl[14] br[14] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_17 
+ bl[15] br[15] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_18 
+ bl[16] br[16] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_19 
+ bl[17] br[17] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_20 
+ bl[18] br[18] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_21 
+ bl[19] br[19] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_22 
+ bl[20] br[20] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_23 
+ bl[21] br[21] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_24 
+ bl[22] br[22] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_25 
+ bl[23] br[23] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_26 
+ bl[24] br[24] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_27 
+ bl[25] br[25] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_28 
+ bl[26] br[26] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_29 
+ bl[27] br[27] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_30 
+ bl[28] br[28] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_31 
+ bl[29] br[29] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_32 
+ bl[30] br[30] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_33 
+ bl[31] br[31] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_34 
+ bl[32] br[32] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_35 
+ bl[33] br[33] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_36 
+ bl[34] br[34] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_37 
+ bl[35] br[35] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_38 
+ bl[36] br[36] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_39 
+ bl[37] br[37] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_40 
+ bl[38] br[38] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_41 
+ bl[39] br[39] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_42 
+ bl[40] br[40] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_43 
+ bl[41] br[41] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_44 
+ bl[42] br[42] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_45 
+ bl[43] br[43] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_46 
+ bl[44] br[44] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_47 
+ bl[45] br[45] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_48 
+ bl[46] br[46] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_49 
+ bl[47] br[47] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_50 
+ bl[48] br[48] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_51 
+ bl[49] br[49] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_52 
+ bl[50] br[50] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_53 
+ bl[51] br[51] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_54 
+ bl[52] br[52] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_55 
+ bl[53] br[53] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_56 
+ bl[54] br[54] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_57 
+ bl[55] br[55] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_58 
+ bl[56] br[56] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_59 
+ bl[57] br[57] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_60 
+ bl[58] br[58] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_61 
+ bl[59] br[59] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_62 
+ bl[60] br[60] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_63 
+ bl[61] br[61] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_64 
+ bl[62] br[62] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_65 
+ bl[63] br[63] vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_66 
+ vdd vdd vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_437_67 
+ vdd vdd vdd vss wl[435] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_0 
+ vdd vdd vss vdd vpb vnb wl[436] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_438_1 
+ rbl rbr vss vdd vpb vnb wl[436] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_438_2 
+ bl[0] br[0] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_3 
+ bl[1] br[1] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_4 
+ bl[2] br[2] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_5 
+ bl[3] br[3] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_6 
+ bl[4] br[4] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_7 
+ bl[5] br[5] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_8 
+ bl[6] br[6] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_9 
+ bl[7] br[7] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_10 
+ bl[8] br[8] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_11 
+ bl[9] br[9] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_12 
+ bl[10] br[10] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_13 
+ bl[11] br[11] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_14 
+ bl[12] br[12] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_15 
+ bl[13] br[13] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_16 
+ bl[14] br[14] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_17 
+ bl[15] br[15] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_18 
+ bl[16] br[16] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_19 
+ bl[17] br[17] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_20 
+ bl[18] br[18] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_21 
+ bl[19] br[19] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_22 
+ bl[20] br[20] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_23 
+ bl[21] br[21] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_24 
+ bl[22] br[22] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_25 
+ bl[23] br[23] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_26 
+ bl[24] br[24] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_27 
+ bl[25] br[25] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_28 
+ bl[26] br[26] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_29 
+ bl[27] br[27] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_30 
+ bl[28] br[28] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_31 
+ bl[29] br[29] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_32 
+ bl[30] br[30] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_33 
+ bl[31] br[31] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_34 
+ bl[32] br[32] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_35 
+ bl[33] br[33] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_36 
+ bl[34] br[34] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_37 
+ bl[35] br[35] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_38 
+ bl[36] br[36] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_39 
+ bl[37] br[37] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_40 
+ bl[38] br[38] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_41 
+ bl[39] br[39] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_42 
+ bl[40] br[40] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_43 
+ bl[41] br[41] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_44 
+ bl[42] br[42] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_45 
+ bl[43] br[43] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_46 
+ bl[44] br[44] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_47 
+ bl[45] br[45] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_48 
+ bl[46] br[46] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_49 
+ bl[47] br[47] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_50 
+ bl[48] br[48] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_51 
+ bl[49] br[49] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_52 
+ bl[50] br[50] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_53 
+ bl[51] br[51] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_54 
+ bl[52] br[52] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_55 
+ bl[53] br[53] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_56 
+ bl[54] br[54] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_57 
+ bl[55] br[55] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_58 
+ bl[56] br[56] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_59 
+ bl[57] br[57] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_60 
+ bl[58] br[58] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_61 
+ bl[59] br[59] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_62 
+ bl[60] br[60] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_63 
+ bl[61] br[61] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_64 
+ bl[62] br[62] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_65 
+ bl[63] br[63] vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_66 
+ vdd vdd vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_438_67 
+ vdd vdd vdd vss wl[436] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_0 
+ vdd vdd vss vdd vpb vnb wl[437] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_439_1 
+ rbl rbr vss vdd vpb vnb wl[437] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_439_2 
+ bl[0] br[0] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_3 
+ bl[1] br[1] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_4 
+ bl[2] br[2] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_5 
+ bl[3] br[3] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_6 
+ bl[4] br[4] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_7 
+ bl[5] br[5] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_8 
+ bl[6] br[6] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_9 
+ bl[7] br[7] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_10 
+ bl[8] br[8] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_11 
+ bl[9] br[9] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_12 
+ bl[10] br[10] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_13 
+ bl[11] br[11] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_14 
+ bl[12] br[12] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_15 
+ bl[13] br[13] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_16 
+ bl[14] br[14] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_17 
+ bl[15] br[15] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_18 
+ bl[16] br[16] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_19 
+ bl[17] br[17] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_20 
+ bl[18] br[18] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_21 
+ bl[19] br[19] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_22 
+ bl[20] br[20] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_23 
+ bl[21] br[21] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_24 
+ bl[22] br[22] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_25 
+ bl[23] br[23] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_26 
+ bl[24] br[24] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_27 
+ bl[25] br[25] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_28 
+ bl[26] br[26] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_29 
+ bl[27] br[27] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_30 
+ bl[28] br[28] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_31 
+ bl[29] br[29] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_32 
+ bl[30] br[30] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_33 
+ bl[31] br[31] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_34 
+ bl[32] br[32] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_35 
+ bl[33] br[33] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_36 
+ bl[34] br[34] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_37 
+ bl[35] br[35] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_38 
+ bl[36] br[36] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_39 
+ bl[37] br[37] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_40 
+ bl[38] br[38] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_41 
+ bl[39] br[39] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_42 
+ bl[40] br[40] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_43 
+ bl[41] br[41] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_44 
+ bl[42] br[42] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_45 
+ bl[43] br[43] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_46 
+ bl[44] br[44] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_47 
+ bl[45] br[45] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_48 
+ bl[46] br[46] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_49 
+ bl[47] br[47] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_50 
+ bl[48] br[48] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_51 
+ bl[49] br[49] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_52 
+ bl[50] br[50] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_53 
+ bl[51] br[51] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_54 
+ bl[52] br[52] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_55 
+ bl[53] br[53] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_56 
+ bl[54] br[54] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_57 
+ bl[55] br[55] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_58 
+ bl[56] br[56] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_59 
+ bl[57] br[57] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_60 
+ bl[58] br[58] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_61 
+ bl[59] br[59] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_62 
+ bl[60] br[60] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_63 
+ bl[61] br[61] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_64 
+ bl[62] br[62] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_65 
+ bl[63] br[63] vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_66 
+ vdd vdd vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_439_67 
+ vdd vdd vdd vss wl[437] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_0 
+ vdd vdd vss vdd vpb vnb wl[438] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_440_1 
+ rbl rbr vss vdd vpb vnb wl[438] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_440_2 
+ bl[0] br[0] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_3 
+ bl[1] br[1] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_4 
+ bl[2] br[2] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_5 
+ bl[3] br[3] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_6 
+ bl[4] br[4] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_7 
+ bl[5] br[5] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_8 
+ bl[6] br[6] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_9 
+ bl[7] br[7] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_10 
+ bl[8] br[8] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_11 
+ bl[9] br[9] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_12 
+ bl[10] br[10] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_13 
+ bl[11] br[11] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_14 
+ bl[12] br[12] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_15 
+ bl[13] br[13] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_16 
+ bl[14] br[14] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_17 
+ bl[15] br[15] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_18 
+ bl[16] br[16] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_19 
+ bl[17] br[17] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_20 
+ bl[18] br[18] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_21 
+ bl[19] br[19] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_22 
+ bl[20] br[20] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_23 
+ bl[21] br[21] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_24 
+ bl[22] br[22] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_25 
+ bl[23] br[23] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_26 
+ bl[24] br[24] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_27 
+ bl[25] br[25] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_28 
+ bl[26] br[26] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_29 
+ bl[27] br[27] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_30 
+ bl[28] br[28] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_31 
+ bl[29] br[29] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_32 
+ bl[30] br[30] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_33 
+ bl[31] br[31] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_34 
+ bl[32] br[32] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_35 
+ bl[33] br[33] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_36 
+ bl[34] br[34] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_37 
+ bl[35] br[35] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_38 
+ bl[36] br[36] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_39 
+ bl[37] br[37] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_40 
+ bl[38] br[38] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_41 
+ bl[39] br[39] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_42 
+ bl[40] br[40] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_43 
+ bl[41] br[41] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_44 
+ bl[42] br[42] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_45 
+ bl[43] br[43] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_46 
+ bl[44] br[44] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_47 
+ bl[45] br[45] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_48 
+ bl[46] br[46] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_49 
+ bl[47] br[47] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_50 
+ bl[48] br[48] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_51 
+ bl[49] br[49] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_52 
+ bl[50] br[50] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_53 
+ bl[51] br[51] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_54 
+ bl[52] br[52] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_55 
+ bl[53] br[53] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_56 
+ bl[54] br[54] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_57 
+ bl[55] br[55] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_58 
+ bl[56] br[56] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_59 
+ bl[57] br[57] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_60 
+ bl[58] br[58] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_61 
+ bl[59] br[59] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_62 
+ bl[60] br[60] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_63 
+ bl[61] br[61] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_64 
+ bl[62] br[62] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_65 
+ bl[63] br[63] vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_66 
+ vdd vdd vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_440_67 
+ vdd vdd vdd vss wl[438] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_0 
+ vdd vdd vss vdd vpb vnb wl[439] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_441_1 
+ rbl rbr vss vdd vpb vnb wl[439] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_441_2 
+ bl[0] br[0] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_3 
+ bl[1] br[1] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_4 
+ bl[2] br[2] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_5 
+ bl[3] br[3] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_6 
+ bl[4] br[4] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_7 
+ bl[5] br[5] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_8 
+ bl[6] br[6] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_9 
+ bl[7] br[7] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_10 
+ bl[8] br[8] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_11 
+ bl[9] br[9] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_12 
+ bl[10] br[10] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_13 
+ bl[11] br[11] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_14 
+ bl[12] br[12] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_15 
+ bl[13] br[13] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_16 
+ bl[14] br[14] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_17 
+ bl[15] br[15] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_18 
+ bl[16] br[16] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_19 
+ bl[17] br[17] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_20 
+ bl[18] br[18] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_21 
+ bl[19] br[19] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_22 
+ bl[20] br[20] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_23 
+ bl[21] br[21] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_24 
+ bl[22] br[22] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_25 
+ bl[23] br[23] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_26 
+ bl[24] br[24] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_27 
+ bl[25] br[25] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_28 
+ bl[26] br[26] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_29 
+ bl[27] br[27] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_30 
+ bl[28] br[28] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_31 
+ bl[29] br[29] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_32 
+ bl[30] br[30] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_33 
+ bl[31] br[31] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_34 
+ bl[32] br[32] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_35 
+ bl[33] br[33] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_36 
+ bl[34] br[34] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_37 
+ bl[35] br[35] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_38 
+ bl[36] br[36] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_39 
+ bl[37] br[37] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_40 
+ bl[38] br[38] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_41 
+ bl[39] br[39] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_42 
+ bl[40] br[40] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_43 
+ bl[41] br[41] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_44 
+ bl[42] br[42] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_45 
+ bl[43] br[43] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_46 
+ bl[44] br[44] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_47 
+ bl[45] br[45] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_48 
+ bl[46] br[46] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_49 
+ bl[47] br[47] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_50 
+ bl[48] br[48] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_51 
+ bl[49] br[49] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_52 
+ bl[50] br[50] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_53 
+ bl[51] br[51] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_54 
+ bl[52] br[52] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_55 
+ bl[53] br[53] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_56 
+ bl[54] br[54] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_57 
+ bl[55] br[55] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_58 
+ bl[56] br[56] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_59 
+ bl[57] br[57] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_60 
+ bl[58] br[58] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_61 
+ bl[59] br[59] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_62 
+ bl[60] br[60] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_63 
+ bl[61] br[61] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_64 
+ bl[62] br[62] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_65 
+ bl[63] br[63] vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_66 
+ vdd vdd vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_441_67 
+ vdd vdd vdd vss wl[439] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_0 
+ vdd vdd vss vdd vpb vnb wl[440] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_442_1 
+ rbl rbr vss vdd vpb vnb wl[440] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_442_2 
+ bl[0] br[0] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_3 
+ bl[1] br[1] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_4 
+ bl[2] br[2] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_5 
+ bl[3] br[3] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_6 
+ bl[4] br[4] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_7 
+ bl[5] br[5] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_8 
+ bl[6] br[6] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_9 
+ bl[7] br[7] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_10 
+ bl[8] br[8] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_11 
+ bl[9] br[9] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_12 
+ bl[10] br[10] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_13 
+ bl[11] br[11] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_14 
+ bl[12] br[12] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_15 
+ bl[13] br[13] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_16 
+ bl[14] br[14] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_17 
+ bl[15] br[15] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_18 
+ bl[16] br[16] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_19 
+ bl[17] br[17] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_20 
+ bl[18] br[18] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_21 
+ bl[19] br[19] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_22 
+ bl[20] br[20] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_23 
+ bl[21] br[21] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_24 
+ bl[22] br[22] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_25 
+ bl[23] br[23] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_26 
+ bl[24] br[24] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_27 
+ bl[25] br[25] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_28 
+ bl[26] br[26] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_29 
+ bl[27] br[27] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_30 
+ bl[28] br[28] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_31 
+ bl[29] br[29] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_32 
+ bl[30] br[30] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_33 
+ bl[31] br[31] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_34 
+ bl[32] br[32] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_35 
+ bl[33] br[33] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_36 
+ bl[34] br[34] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_37 
+ bl[35] br[35] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_38 
+ bl[36] br[36] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_39 
+ bl[37] br[37] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_40 
+ bl[38] br[38] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_41 
+ bl[39] br[39] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_42 
+ bl[40] br[40] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_43 
+ bl[41] br[41] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_44 
+ bl[42] br[42] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_45 
+ bl[43] br[43] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_46 
+ bl[44] br[44] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_47 
+ bl[45] br[45] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_48 
+ bl[46] br[46] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_49 
+ bl[47] br[47] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_50 
+ bl[48] br[48] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_51 
+ bl[49] br[49] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_52 
+ bl[50] br[50] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_53 
+ bl[51] br[51] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_54 
+ bl[52] br[52] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_55 
+ bl[53] br[53] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_56 
+ bl[54] br[54] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_57 
+ bl[55] br[55] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_58 
+ bl[56] br[56] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_59 
+ bl[57] br[57] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_60 
+ bl[58] br[58] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_61 
+ bl[59] br[59] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_62 
+ bl[60] br[60] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_63 
+ bl[61] br[61] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_64 
+ bl[62] br[62] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_65 
+ bl[63] br[63] vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_66 
+ vdd vdd vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_442_67 
+ vdd vdd vdd vss wl[440] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_0 
+ vdd vdd vss vdd vpb vnb wl[441] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_443_1 
+ rbl rbr vss vdd vpb vnb wl[441] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_443_2 
+ bl[0] br[0] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_3 
+ bl[1] br[1] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_4 
+ bl[2] br[2] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_5 
+ bl[3] br[3] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_6 
+ bl[4] br[4] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_7 
+ bl[5] br[5] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_8 
+ bl[6] br[6] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_9 
+ bl[7] br[7] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_10 
+ bl[8] br[8] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_11 
+ bl[9] br[9] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_12 
+ bl[10] br[10] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_13 
+ bl[11] br[11] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_14 
+ bl[12] br[12] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_15 
+ bl[13] br[13] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_16 
+ bl[14] br[14] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_17 
+ bl[15] br[15] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_18 
+ bl[16] br[16] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_19 
+ bl[17] br[17] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_20 
+ bl[18] br[18] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_21 
+ bl[19] br[19] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_22 
+ bl[20] br[20] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_23 
+ bl[21] br[21] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_24 
+ bl[22] br[22] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_25 
+ bl[23] br[23] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_26 
+ bl[24] br[24] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_27 
+ bl[25] br[25] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_28 
+ bl[26] br[26] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_29 
+ bl[27] br[27] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_30 
+ bl[28] br[28] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_31 
+ bl[29] br[29] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_32 
+ bl[30] br[30] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_33 
+ bl[31] br[31] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_34 
+ bl[32] br[32] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_35 
+ bl[33] br[33] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_36 
+ bl[34] br[34] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_37 
+ bl[35] br[35] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_38 
+ bl[36] br[36] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_39 
+ bl[37] br[37] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_40 
+ bl[38] br[38] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_41 
+ bl[39] br[39] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_42 
+ bl[40] br[40] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_43 
+ bl[41] br[41] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_44 
+ bl[42] br[42] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_45 
+ bl[43] br[43] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_46 
+ bl[44] br[44] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_47 
+ bl[45] br[45] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_48 
+ bl[46] br[46] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_49 
+ bl[47] br[47] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_50 
+ bl[48] br[48] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_51 
+ bl[49] br[49] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_52 
+ bl[50] br[50] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_53 
+ bl[51] br[51] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_54 
+ bl[52] br[52] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_55 
+ bl[53] br[53] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_56 
+ bl[54] br[54] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_57 
+ bl[55] br[55] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_58 
+ bl[56] br[56] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_59 
+ bl[57] br[57] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_60 
+ bl[58] br[58] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_61 
+ bl[59] br[59] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_62 
+ bl[60] br[60] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_63 
+ bl[61] br[61] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_64 
+ bl[62] br[62] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_65 
+ bl[63] br[63] vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_66 
+ vdd vdd vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_443_67 
+ vdd vdd vdd vss wl[441] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_0 
+ vdd vdd vss vdd vpb vnb wl[442] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_444_1 
+ rbl rbr vss vdd vpb vnb wl[442] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_444_2 
+ bl[0] br[0] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_3 
+ bl[1] br[1] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_4 
+ bl[2] br[2] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_5 
+ bl[3] br[3] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_6 
+ bl[4] br[4] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_7 
+ bl[5] br[5] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_8 
+ bl[6] br[6] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_9 
+ bl[7] br[7] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_10 
+ bl[8] br[8] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_11 
+ bl[9] br[9] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_12 
+ bl[10] br[10] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_13 
+ bl[11] br[11] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_14 
+ bl[12] br[12] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_15 
+ bl[13] br[13] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_16 
+ bl[14] br[14] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_17 
+ bl[15] br[15] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_18 
+ bl[16] br[16] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_19 
+ bl[17] br[17] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_20 
+ bl[18] br[18] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_21 
+ bl[19] br[19] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_22 
+ bl[20] br[20] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_23 
+ bl[21] br[21] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_24 
+ bl[22] br[22] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_25 
+ bl[23] br[23] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_26 
+ bl[24] br[24] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_27 
+ bl[25] br[25] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_28 
+ bl[26] br[26] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_29 
+ bl[27] br[27] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_30 
+ bl[28] br[28] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_31 
+ bl[29] br[29] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_32 
+ bl[30] br[30] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_33 
+ bl[31] br[31] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_34 
+ bl[32] br[32] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_35 
+ bl[33] br[33] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_36 
+ bl[34] br[34] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_37 
+ bl[35] br[35] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_38 
+ bl[36] br[36] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_39 
+ bl[37] br[37] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_40 
+ bl[38] br[38] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_41 
+ bl[39] br[39] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_42 
+ bl[40] br[40] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_43 
+ bl[41] br[41] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_44 
+ bl[42] br[42] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_45 
+ bl[43] br[43] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_46 
+ bl[44] br[44] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_47 
+ bl[45] br[45] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_48 
+ bl[46] br[46] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_49 
+ bl[47] br[47] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_50 
+ bl[48] br[48] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_51 
+ bl[49] br[49] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_52 
+ bl[50] br[50] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_53 
+ bl[51] br[51] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_54 
+ bl[52] br[52] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_55 
+ bl[53] br[53] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_56 
+ bl[54] br[54] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_57 
+ bl[55] br[55] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_58 
+ bl[56] br[56] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_59 
+ bl[57] br[57] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_60 
+ bl[58] br[58] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_61 
+ bl[59] br[59] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_62 
+ bl[60] br[60] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_63 
+ bl[61] br[61] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_64 
+ bl[62] br[62] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_65 
+ bl[63] br[63] vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_66 
+ vdd vdd vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_444_67 
+ vdd vdd vdd vss wl[442] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_0 
+ vdd vdd vss vdd vpb vnb wl[443] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_445_1 
+ rbl rbr vss vdd vpb vnb wl[443] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_445_2 
+ bl[0] br[0] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_3 
+ bl[1] br[1] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_4 
+ bl[2] br[2] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_5 
+ bl[3] br[3] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_6 
+ bl[4] br[4] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_7 
+ bl[5] br[5] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_8 
+ bl[6] br[6] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_9 
+ bl[7] br[7] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_10 
+ bl[8] br[8] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_11 
+ bl[9] br[9] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_12 
+ bl[10] br[10] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_13 
+ bl[11] br[11] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_14 
+ bl[12] br[12] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_15 
+ bl[13] br[13] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_16 
+ bl[14] br[14] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_17 
+ bl[15] br[15] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_18 
+ bl[16] br[16] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_19 
+ bl[17] br[17] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_20 
+ bl[18] br[18] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_21 
+ bl[19] br[19] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_22 
+ bl[20] br[20] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_23 
+ bl[21] br[21] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_24 
+ bl[22] br[22] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_25 
+ bl[23] br[23] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_26 
+ bl[24] br[24] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_27 
+ bl[25] br[25] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_28 
+ bl[26] br[26] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_29 
+ bl[27] br[27] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_30 
+ bl[28] br[28] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_31 
+ bl[29] br[29] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_32 
+ bl[30] br[30] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_33 
+ bl[31] br[31] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_34 
+ bl[32] br[32] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_35 
+ bl[33] br[33] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_36 
+ bl[34] br[34] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_37 
+ bl[35] br[35] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_38 
+ bl[36] br[36] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_39 
+ bl[37] br[37] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_40 
+ bl[38] br[38] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_41 
+ bl[39] br[39] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_42 
+ bl[40] br[40] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_43 
+ bl[41] br[41] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_44 
+ bl[42] br[42] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_45 
+ bl[43] br[43] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_46 
+ bl[44] br[44] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_47 
+ bl[45] br[45] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_48 
+ bl[46] br[46] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_49 
+ bl[47] br[47] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_50 
+ bl[48] br[48] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_51 
+ bl[49] br[49] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_52 
+ bl[50] br[50] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_53 
+ bl[51] br[51] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_54 
+ bl[52] br[52] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_55 
+ bl[53] br[53] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_56 
+ bl[54] br[54] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_57 
+ bl[55] br[55] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_58 
+ bl[56] br[56] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_59 
+ bl[57] br[57] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_60 
+ bl[58] br[58] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_61 
+ bl[59] br[59] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_62 
+ bl[60] br[60] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_63 
+ bl[61] br[61] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_64 
+ bl[62] br[62] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_65 
+ bl[63] br[63] vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_66 
+ vdd vdd vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_445_67 
+ vdd vdd vdd vss wl[443] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_0 
+ vdd vdd vss vdd vpb vnb wl[444] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_446_1 
+ rbl rbr vss vdd vpb vnb wl[444] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_446_2 
+ bl[0] br[0] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_3 
+ bl[1] br[1] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_4 
+ bl[2] br[2] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_5 
+ bl[3] br[3] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_6 
+ bl[4] br[4] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_7 
+ bl[5] br[5] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_8 
+ bl[6] br[6] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_9 
+ bl[7] br[7] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_10 
+ bl[8] br[8] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_11 
+ bl[9] br[9] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_12 
+ bl[10] br[10] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_13 
+ bl[11] br[11] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_14 
+ bl[12] br[12] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_15 
+ bl[13] br[13] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_16 
+ bl[14] br[14] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_17 
+ bl[15] br[15] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_18 
+ bl[16] br[16] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_19 
+ bl[17] br[17] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_20 
+ bl[18] br[18] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_21 
+ bl[19] br[19] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_22 
+ bl[20] br[20] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_23 
+ bl[21] br[21] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_24 
+ bl[22] br[22] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_25 
+ bl[23] br[23] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_26 
+ bl[24] br[24] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_27 
+ bl[25] br[25] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_28 
+ bl[26] br[26] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_29 
+ bl[27] br[27] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_30 
+ bl[28] br[28] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_31 
+ bl[29] br[29] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_32 
+ bl[30] br[30] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_33 
+ bl[31] br[31] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_34 
+ bl[32] br[32] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_35 
+ bl[33] br[33] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_36 
+ bl[34] br[34] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_37 
+ bl[35] br[35] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_38 
+ bl[36] br[36] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_39 
+ bl[37] br[37] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_40 
+ bl[38] br[38] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_41 
+ bl[39] br[39] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_42 
+ bl[40] br[40] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_43 
+ bl[41] br[41] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_44 
+ bl[42] br[42] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_45 
+ bl[43] br[43] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_46 
+ bl[44] br[44] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_47 
+ bl[45] br[45] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_48 
+ bl[46] br[46] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_49 
+ bl[47] br[47] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_50 
+ bl[48] br[48] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_51 
+ bl[49] br[49] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_52 
+ bl[50] br[50] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_53 
+ bl[51] br[51] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_54 
+ bl[52] br[52] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_55 
+ bl[53] br[53] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_56 
+ bl[54] br[54] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_57 
+ bl[55] br[55] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_58 
+ bl[56] br[56] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_59 
+ bl[57] br[57] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_60 
+ bl[58] br[58] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_61 
+ bl[59] br[59] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_62 
+ bl[60] br[60] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_63 
+ bl[61] br[61] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_64 
+ bl[62] br[62] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_65 
+ bl[63] br[63] vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_66 
+ vdd vdd vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_446_67 
+ vdd vdd vdd vss wl[444] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_0 
+ vdd vdd vss vdd vpb vnb wl[445] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_447_1 
+ rbl rbr vss vdd vpb vnb wl[445] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_447_2 
+ bl[0] br[0] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_3 
+ bl[1] br[1] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_4 
+ bl[2] br[2] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_5 
+ bl[3] br[3] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_6 
+ bl[4] br[4] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_7 
+ bl[5] br[5] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_8 
+ bl[6] br[6] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_9 
+ bl[7] br[7] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_10 
+ bl[8] br[8] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_11 
+ bl[9] br[9] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_12 
+ bl[10] br[10] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_13 
+ bl[11] br[11] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_14 
+ bl[12] br[12] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_15 
+ bl[13] br[13] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_16 
+ bl[14] br[14] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_17 
+ bl[15] br[15] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_18 
+ bl[16] br[16] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_19 
+ bl[17] br[17] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_20 
+ bl[18] br[18] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_21 
+ bl[19] br[19] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_22 
+ bl[20] br[20] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_23 
+ bl[21] br[21] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_24 
+ bl[22] br[22] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_25 
+ bl[23] br[23] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_26 
+ bl[24] br[24] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_27 
+ bl[25] br[25] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_28 
+ bl[26] br[26] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_29 
+ bl[27] br[27] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_30 
+ bl[28] br[28] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_31 
+ bl[29] br[29] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_32 
+ bl[30] br[30] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_33 
+ bl[31] br[31] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_34 
+ bl[32] br[32] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_35 
+ bl[33] br[33] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_36 
+ bl[34] br[34] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_37 
+ bl[35] br[35] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_38 
+ bl[36] br[36] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_39 
+ bl[37] br[37] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_40 
+ bl[38] br[38] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_41 
+ bl[39] br[39] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_42 
+ bl[40] br[40] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_43 
+ bl[41] br[41] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_44 
+ bl[42] br[42] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_45 
+ bl[43] br[43] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_46 
+ bl[44] br[44] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_47 
+ bl[45] br[45] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_48 
+ bl[46] br[46] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_49 
+ bl[47] br[47] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_50 
+ bl[48] br[48] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_51 
+ bl[49] br[49] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_52 
+ bl[50] br[50] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_53 
+ bl[51] br[51] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_54 
+ bl[52] br[52] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_55 
+ bl[53] br[53] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_56 
+ bl[54] br[54] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_57 
+ bl[55] br[55] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_58 
+ bl[56] br[56] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_59 
+ bl[57] br[57] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_60 
+ bl[58] br[58] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_61 
+ bl[59] br[59] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_62 
+ bl[60] br[60] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_63 
+ bl[61] br[61] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_64 
+ bl[62] br[62] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_65 
+ bl[63] br[63] vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_66 
+ vdd vdd vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_447_67 
+ vdd vdd vdd vss wl[445] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_0 
+ vdd vdd vss vdd vpb vnb wl[446] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_448_1 
+ rbl rbr vss vdd vpb vnb wl[446] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_448_2 
+ bl[0] br[0] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_3 
+ bl[1] br[1] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_4 
+ bl[2] br[2] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_5 
+ bl[3] br[3] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_6 
+ bl[4] br[4] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_7 
+ bl[5] br[5] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_8 
+ bl[6] br[6] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_9 
+ bl[7] br[7] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_10 
+ bl[8] br[8] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_11 
+ bl[9] br[9] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_12 
+ bl[10] br[10] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_13 
+ bl[11] br[11] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_14 
+ bl[12] br[12] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_15 
+ bl[13] br[13] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_16 
+ bl[14] br[14] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_17 
+ bl[15] br[15] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_18 
+ bl[16] br[16] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_19 
+ bl[17] br[17] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_20 
+ bl[18] br[18] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_21 
+ bl[19] br[19] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_22 
+ bl[20] br[20] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_23 
+ bl[21] br[21] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_24 
+ bl[22] br[22] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_25 
+ bl[23] br[23] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_26 
+ bl[24] br[24] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_27 
+ bl[25] br[25] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_28 
+ bl[26] br[26] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_29 
+ bl[27] br[27] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_30 
+ bl[28] br[28] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_31 
+ bl[29] br[29] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_32 
+ bl[30] br[30] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_33 
+ bl[31] br[31] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_34 
+ bl[32] br[32] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_35 
+ bl[33] br[33] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_36 
+ bl[34] br[34] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_37 
+ bl[35] br[35] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_38 
+ bl[36] br[36] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_39 
+ bl[37] br[37] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_40 
+ bl[38] br[38] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_41 
+ bl[39] br[39] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_42 
+ bl[40] br[40] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_43 
+ bl[41] br[41] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_44 
+ bl[42] br[42] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_45 
+ bl[43] br[43] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_46 
+ bl[44] br[44] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_47 
+ bl[45] br[45] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_48 
+ bl[46] br[46] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_49 
+ bl[47] br[47] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_50 
+ bl[48] br[48] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_51 
+ bl[49] br[49] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_52 
+ bl[50] br[50] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_53 
+ bl[51] br[51] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_54 
+ bl[52] br[52] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_55 
+ bl[53] br[53] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_56 
+ bl[54] br[54] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_57 
+ bl[55] br[55] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_58 
+ bl[56] br[56] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_59 
+ bl[57] br[57] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_60 
+ bl[58] br[58] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_61 
+ bl[59] br[59] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_62 
+ bl[60] br[60] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_63 
+ bl[61] br[61] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_64 
+ bl[62] br[62] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_65 
+ bl[63] br[63] vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_66 
+ vdd vdd vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_448_67 
+ vdd vdd vdd vss wl[446] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_0 
+ vdd vdd vss vdd vpb vnb wl[447] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_449_1 
+ rbl rbr vss vdd vpb vnb wl[447] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_449_2 
+ bl[0] br[0] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_3 
+ bl[1] br[1] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_4 
+ bl[2] br[2] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_5 
+ bl[3] br[3] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_6 
+ bl[4] br[4] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_7 
+ bl[5] br[5] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_8 
+ bl[6] br[6] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_9 
+ bl[7] br[7] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_10 
+ bl[8] br[8] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_11 
+ bl[9] br[9] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_12 
+ bl[10] br[10] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_13 
+ bl[11] br[11] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_14 
+ bl[12] br[12] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_15 
+ bl[13] br[13] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_16 
+ bl[14] br[14] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_17 
+ bl[15] br[15] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_18 
+ bl[16] br[16] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_19 
+ bl[17] br[17] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_20 
+ bl[18] br[18] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_21 
+ bl[19] br[19] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_22 
+ bl[20] br[20] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_23 
+ bl[21] br[21] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_24 
+ bl[22] br[22] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_25 
+ bl[23] br[23] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_26 
+ bl[24] br[24] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_27 
+ bl[25] br[25] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_28 
+ bl[26] br[26] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_29 
+ bl[27] br[27] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_30 
+ bl[28] br[28] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_31 
+ bl[29] br[29] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_32 
+ bl[30] br[30] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_33 
+ bl[31] br[31] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_34 
+ bl[32] br[32] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_35 
+ bl[33] br[33] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_36 
+ bl[34] br[34] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_37 
+ bl[35] br[35] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_38 
+ bl[36] br[36] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_39 
+ bl[37] br[37] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_40 
+ bl[38] br[38] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_41 
+ bl[39] br[39] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_42 
+ bl[40] br[40] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_43 
+ bl[41] br[41] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_44 
+ bl[42] br[42] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_45 
+ bl[43] br[43] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_46 
+ bl[44] br[44] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_47 
+ bl[45] br[45] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_48 
+ bl[46] br[46] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_49 
+ bl[47] br[47] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_50 
+ bl[48] br[48] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_51 
+ bl[49] br[49] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_52 
+ bl[50] br[50] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_53 
+ bl[51] br[51] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_54 
+ bl[52] br[52] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_55 
+ bl[53] br[53] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_56 
+ bl[54] br[54] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_57 
+ bl[55] br[55] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_58 
+ bl[56] br[56] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_59 
+ bl[57] br[57] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_60 
+ bl[58] br[58] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_61 
+ bl[59] br[59] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_62 
+ bl[60] br[60] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_63 
+ bl[61] br[61] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_64 
+ bl[62] br[62] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_65 
+ bl[63] br[63] vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_66 
+ vdd vdd vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_449_67 
+ vdd vdd vdd vss wl[447] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_0 
+ vdd vdd vss vdd vpb vnb wl[448] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_450_1 
+ rbl rbr vss vdd vpb vnb wl[448] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_450_2 
+ bl[0] br[0] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_3 
+ bl[1] br[1] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_4 
+ bl[2] br[2] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_5 
+ bl[3] br[3] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_6 
+ bl[4] br[4] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_7 
+ bl[5] br[5] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_8 
+ bl[6] br[6] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_9 
+ bl[7] br[7] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_10 
+ bl[8] br[8] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_11 
+ bl[9] br[9] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_12 
+ bl[10] br[10] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_13 
+ bl[11] br[11] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_14 
+ bl[12] br[12] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_15 
+ bl[13] br[13] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_16 
+ bl[14] br[14] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_17 
+ bl[15] br[15] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_18 
+ bl[16] br[16] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_19 
+ bl[17] br[17] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_20 
+ bl[18] br[18] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_21 
+ bl[19] br[19] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_22 
+ bl[20] br[20] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_23 
+ bl[21] br[21] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_24 
+ bl[22] br[22] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_25 
+ bl[23] br[23] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_26 
+ bl[24] br[24] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_27 
+ bl[25] br[25] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_28 
+ bl[26] br[26] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_29 
+ bl[27] br[27] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_30 
+ bl[28] br[28] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_31 
+ bl[29] br[29] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_32 
+ bl[30] br[30] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_33 
+ bl[31] br[31] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_34 
+ bl[32] br[32] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_35 
+ bl[33] br[33] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_36 
+ bl[34] br[34] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_37 
+ bl[35] br[35] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_38 
+ bl[36] br[36] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_39 
+ bl[37] br[37] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_40 
+ bl[38] br[38] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_41 
+ bl[39] br[39] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_42 
+ bl[40] br[40] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_43 
+ bl[41] br[41] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_44 
+ bl[42] br[42] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_45 
+ bl[43] br[43] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_46 
+ bl[44] br[44] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_47 
+ bl[45] br[45] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_48 
+ bl[46] br[46] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_49 
+ bl[47] br[47] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_50 
+ bl[48] br[48] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_51 
+ bl[49] br[49] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_52 
+ bl[50] br[50] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_53 
+ bl[51] br[51] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_54 
+ bl[52] br[52] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_55 
+ bl[53] br[53] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_56 
+ bl[54] br[54] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_57 
+ bl[55] br[55] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_58 
+ bl[56] br[56] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_59 
+ bl[57] br[57] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_60 
+ bl[58] br[58] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_61 
+ bl[59] br[59] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_62 
+ bl[60] br[60] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_63 
+ bl[61] br[61] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_64 
+ bl[62] br[62] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_65 
+ bl[63] br[63] vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_66 
+ vdd vdd vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_450_67 
+ vdd vdd vdd vss wl[448] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_0 
+ vdd vdd vss vdd vpb vnb wl[449] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_451_1 
+ rbl rbr vss vdd vpb vnb wl[449] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_451_2 
+ bl[0] br[0] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_3 
+ bl[1] br[1] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_4 
+ bl[2] br[2] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_5 
+ bl[3] br[3] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_6 
+ bl[4] br[4] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_7 
+ bl[5] br[5] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_8 
+ bl[6] br[6] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_9 
+ bl[7] br[7] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_10 
+ bl[8] br[8] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_11 
+ bl[9] br[9] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_12 
+ bl[10] br[10] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_13 
+ bl[11] br[11] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_14 
+ bl[12] br[12] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_15 
+ bl[13] br[13] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_16 
+ bl[14] br[14] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_17 
+ bl[15] br[15] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_18 
+ bl[16] br[16] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_19 
+ bl[17] br[17] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_20 
+ bl[18] br[18] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_21 
+ bl[19] br[19] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_22 
+ bl[20] br[20] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_23 
+ bl[21] br[21] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_24 
+ bl[22] br[22] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_25 
+ bl[23] br[23] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_26 
+ bl[24] br[24] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_27 
+ bl[25] br[25] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_28 
+ bl[26] br[26] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_29 
+ bl[27] br[27] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_30 
+ bl[28] br[28] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_31 
+ bl[29] br[29] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_32 
+ bl[30] br[30] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_33 
+ bl[31] br[31] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_34 
+ bl[32] br[32] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_35 
+ bl[33] br[33] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_36 
+ bl[34] br[34] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_37 
+ bl[35] br[35] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_38 
+ bl[36] br[36] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_39 
+ bl[37] br[37] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_40 
+ bl[38] br[38] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_41 
+ bl[39] br[39] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_42 
+ bl[40] br[40] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_43 
+ bl[41] br[41] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_44 
+ bl[42] br[42] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_45 
+ bl[43] br[43] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_46 
+ bl[44] br[44] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_47 
+ bl[45] br[45] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_48 
+ bl[46] br[46] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_49 
+ bl[47] br[47] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_50 
+ bl[48] br[48] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_51 
+ bl[49] br[49] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_52 
+ bl[50] br[50] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_53 
+ bl[51] br[51] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_54 
+ bl[52] br[52] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_55 
+ bl[53] br[53] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_56 
+ bl[54] br[54] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_57 
+ bl[55] br[55] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_58 
+ bl[56] br[56] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_59 
+ bl[57] br[57] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_60 
+ bl[58] br[58] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_61 
+ bl[59] br[59] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_62 
+ bl[60] br[60] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_63 
+ bl[61] br[61] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_64 
+ bl[62] br[62] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_65 
+ bl[63] br[63] vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_66 
+ vdd vdd vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_451_67 
+ vdd vdd vdd vss wl[449] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_0 
+ vdd vdd vss vdd vpb vnb wl[450] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_452_1 
+ rbl rbr vss vdd vpb vnb wl[450] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_452_2 
+ bl[0] br[0] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_3 
+ bl[1] br[1] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_4 
+ bl[2] br[2] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_5 
+ bl[3] br[3] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_6 
+ bl[4] br[4] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_7 
+ bl[5] br[5] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_8 
+ bl[6] br[6] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_9 
+ bl[7] br[7] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_10 
+ bl[8] br[8] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_11 
+ bl[9] br[9] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_12 
+ bl[10] br[10] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_13 
+ bl[11] br[11] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_14 
+ bl[12] br[12] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_15 
+ bl[13] br[13] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_16 
+ bl[14] br[14] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_17 
+ bl[15] br[15] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_18 
+ bl[16] br[16] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_19 
+ bl[17] br[17] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_20 
+ bl[18] br[18] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_21 
+ bl[19] br[19] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_22 
+ bl[20] br[20] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_23 
+ bl[21] br[21] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_24 
+ bl[22] br[22] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_25 
+ bl[23] br[23] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_26 
+ bl[24] br[24] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_27 
+ bl[25] br[25] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_28 
+ bl[26] br[26] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_29 
+ bl[27] br[27] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_30 
+ bl[28] br[28] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_31 
+ bl[29] br[29] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_32 
+ bl[30] br[30] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_33 
+ bl[31] br[31] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_34 
+ bl[32] br[32] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_35 
+ bl[33] br[33] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_36 
+ bl[34] br[34] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_37 
+ bl[35] br[35] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_38 
+ bl[36] br[36] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_39 
+ bl[37] br[37] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_40 
+ bl[38] br[38] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_41 
+ bl[39] br[39] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_42 
+ bl[40] br[40] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_43 
+ bl[41] br[41] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_44 
+ bl[42] br[42] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_45 
+ bl[43] br[43] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_46 
+ bl[44] br[44] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_47 
+ bl[45] br[45] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_48 
+ bl[46] br[46] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_49 
+ bl[47] br[47] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_50 
+ bl[48] br[48] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_51 
+ bl[49] br[49] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_52 
+ bl[50] br[50] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_53 
+ bl[51] br[51] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_54 
+ bl[52] br[52] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_55 
+ bl[53] br[53] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_56 
+ bl[54] br[54] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_57 
+ bl[55] br[55] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_58 
+ bl[56] br[56] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_59 
+ bl[57] br[57] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_60 
+ bl[58] br[58] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_61 
+ bl[59] br[59] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_62 
+ bl[60] br[60] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_63 
+ bl[61] br[61] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_64 
+ bl[62] br[62] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_65 
+ bl[63] br[63] vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_66 
+ vdd vdd vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_452_67 
+ vdd vdd vdd vss wl[450] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_0 
+ vdd vdd vss vdd vpb vnb wl[451] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_453_1 
+ rbl rbr vss vdd vpb vnb wl[451] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_453_2 
+ bl[0] br[0] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_3 
+ bl[1] br[1] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_4 
+ bl[2] br[2] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_5 
+ bl[3] br[3] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_6 
+ bl[4] br[4] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_7 
+ bl[5] br[5] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_8 
+ bl[6] br[6] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_9 
+ bl[7] br[7] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_10 
+ bl[8] br[8] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_11 
+ bl[9] br[9] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_12 
+ bl[10] br[10] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_13 
+ bl[11] br[11] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_14 
+ bl[12] br[12] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_15 
+ bl[13] br[13] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_16 
+ bl[14] br[14] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_17 
+ bl[15] br[15] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_18 
+ bl[16] br[16] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_19 
+ bl[17] br[17] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_20 
+ bl[18] br[18] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_21 
+ bl[19] br[19] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_22 
+ bl[20] br[20] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_23 
+ bl[21] br[21] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_24 
+ bl[22] br[22] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_25 
+ bl[23] br[23] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_26 
+ bl[24] br[24] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_27 
+ bl[25] br[25] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_28 
+ bl[26] br[26] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_29 
+ bl[27] br[27] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_30 
+ bl[28] br[28] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_31 
+ bl[29] br[29] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_32 
+ bl[30] br[30] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_33 
+ bl[31] br[31] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_34 
+ bl[32] br[32] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_35 
+ bl[33] br[33] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_36 
+ bl[34] br[34] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_37 
+ bl[35] br[35] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_38 
+ bl[36] br[36] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_39 
+ bl[37] br[37] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_40 
+ bl[38] br[38] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_41 
+ bl[39] br[39] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_42 
+ bl[40] br[40] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_43 
+ bl[41] br[41] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_44 
+ bl[42] br[42] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_45 
+ bl[43] br[43] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_46 
+ bl[44] br[44] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_47 
+ bl[45] br[45] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_48 
+ bl[46] br[46] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_49 
+ bl[47] br[47] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_50 
+ bl[48] br[48] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_51 
+ bl[49] br[49] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_52 
+ bl[50] br[50] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_53 
+ bl[51] br[51] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_54 
+ bl[52] br[52] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_55 
+ bl[53] br[53] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_56 
+ bl[54] br[54] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_57 
+ bl[55] br[55] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_58 
+ bl[56] br[56] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_59 
+ bl[57] br[57] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_60 
+ bl[58] br[58] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_61 
+ bl[59] br[59] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_62 
+ bl[60] br[60] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_63 
+ bl[61] br[61] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_64 
+ bl[62] br[62] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_65 
+ bl[63] br[63] vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_66 
+ vdd vdd vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_453_67 
+ vdd vdd vdd vss wl[451] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_0 
+ vdd vdd vss vdd vpb vnb wl[452] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_454_1 
+ rbl rbr vss vdd vpb vnb wl[452] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_454_2 
+ bl[0] br[0] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_3 
+ bl[1] br[1] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_4 
+ bl[2] br[2] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_5 
+ bl[3] br[3] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_6 
+ bl[4] br[4] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_7 
+ bl[5] br[5] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_8 
+ bl[6] br[6] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_9 
+ bl[7] br[7] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_10 
+ bl[8] br[8] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_11 
+ bl[9] br[9] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_12 
+ bl[10] br[10] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_13 
+ bl[11] br[11] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_14 
+ bl[12] br[12] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_15 
+ bl[13] br[13] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_16 
+ bl[14] br[14] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_17 
+ bl[15] br[15] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_18 
+ bl[16] br[16] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_19 
+ bl[17] br[17] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_20 
+ bl[18] br[18] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_21 
+ bl[19] br[19] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_22 
+ bl[20] br[20] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_23 
+ bl[21] br[21] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_24 
+ bl[22] br[22] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_25 
+ bl[23] br[23] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_26 
+ bl[24] br[24] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_27 
+ bl[25] br[25] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_28 
+ bl[26] br[26] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_29 
+ bl[27] br[27] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_30 
+ bl[28] br[28] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_31 
+ bl[29] br[29] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_32 
+ bl[30] br[30] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_33 
+ bl[31] br[31] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_34 
+ bl[32] br[32] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_35 
+ bl[33] br[33] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_36 
+ bl[34] br[34] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_37 
+ bl[35] br[35] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_38 
+ bl[36] br[36] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_39 
+ bl[37] br[37] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_40 
+ bl[38] br[38] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_41 
+ bl[39] br[39] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_42 
+ bl[40] br[40] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_43 
+ bl[41] br[41] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_44 
+ bl[42] br[42] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_45 
+ bl[43] br[43] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_46 
+ bl[44] br[44] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_47 
+ bl[45] br[45] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_48 
+ bl[46] br[46] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_49 
+ bl[47] br[47] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_50 
+ bl[48] br[48] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_51 
+ bl[49] br[49] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_52 
+ bl[50] br[50] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_53 
+ bl[51] br[51] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_54 
+ bl[52] br[52] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_55 
+ bl[53] br[53] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_56 
+ bl[54] br[54] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_57 
+ bl[55] br[55] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_58 
+ bl[56] br[56] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_59 
+ bl[57] br[57] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_60 
+ bl[58] br[58] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_61 
+ bl[59] br[59] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_62 
+ bl[60] br[60] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_63 
+ bl[61] br[61] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_64 
+ bl[62] br[62] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_65 
+ bl[63] br[63] vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_66 
+ vdd vdd vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_454_67 
+ vdd vdd vdd vss wl[452] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_0 
+ vdd vdd vss vdd vpb vnb wl[453] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_455_1 
+ rbl rbr vss vdd vpb vnb wl[453] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_455_2 
+ bl[0] br[0] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_3 
+ bl[1] br[1] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_4 
+ bl[2] br[2] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_5 
+ bl[3] br[3] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_6 
+ bl[4] br[4] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_7 
+ bl[5] br[5] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_8 
+ bl[6] br[6] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_9 
+ bl[7] br[7] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_10 
+ bl[8] br[8] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_11 
+ bl[9] br[9] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_12 
+ bl[10] br[10] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_13 
+ bl[11] br[11] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_14 
+ bl[12] br[12] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_15 
+ bl[13] br[13] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_16 
+ bl[14] br[14] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_17 
+ bl[15] br[15] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_18 
+ bl[16] br[16] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_19 
+ bl[17] br[17] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_20 
+ bl[18] br[18] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_21 
+ bl[19] br[19] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_22 
+ bl[20] br[20] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_23 
+ bl[21] br[21] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_24 
+ bl[22] br[22] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_25 
+ bl[23] br[23] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_26 
+ bl[24] br[24] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_27 
+ bl[25] br[25] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_28 
+ bl[26] br[26] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_29 
+ bl[27] br[27] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_30 
+ bl[28] br[28] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_31 
+ bl[29] br[29] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_32 
+ bl[30] br[30] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_33 
+ bl[31] br[31] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_34 
+ bl[32] br[32] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_35 
+ bl[33] br[33] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_36 
+ bl[34] br[34] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_37 
+ bl[35] br[35] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_38 
+ bl[36] br[36] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_39 
+ bl[37] br[37] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_40 
+ bl[38] br[38] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_41 
+ bl[39] br[39] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_42 
+ bl[40] br[40] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_43 
+ bl[41] br[41] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_44 
+ bl[42] br[42] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_45 
+ bl[43] br[43] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_46 
+ bl[44] br[44] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_47 
+ bl[45] br[45] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_48 
+ bl[46] br[46] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_49 
+ bl[47] br[47] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_50 
+ bl[48] br[48] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_51 
+ bl[49] br[49] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_52 
+ bl[50] br[50] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_53 
+ bl[51] br[51] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_54 
+ bl[52] br[52] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_55 
+ bl[53] br[53] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_56 
+ bl[54] br[54] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_57 
+ bl[55] br[55] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_58 
+ bl[56] br[56] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_59 
+ bl[57] br[57] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_60 
+ bl[58] br[58] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_61 
+ bl[59] br[59] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_62 
+ bl[60] br[60] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_63 
+ bl[61] br[61] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_64 
+ bl[62] br[62] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_65 
+ bl[63] br[63] vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_66 
+ vdd vdd vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_455_67 
+ vdd vdd vdd vss wl[453] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_0 
+ vdd vdd vss vdd vpb vnb wl[454] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_456_1 
+ rbl rbr vss vdd vpb vnb wl[454] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_456_2 
+ bl[0] br[0] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_3 
+ bl[1] br[1] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_4 
+ bl[2] br[2] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_5 
+ bl[3] br[3] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_6 
+ bl[4] br[4] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_7 
+ bl[5] br[5] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_8 
+ bl[6] br[6] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_9 
+ bl[7] br[7] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_10 
+ bl[8] br[8] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_11 
+ bl[9] br[9] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_12 
+ bl[10] br[10] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_13 
+ bl[11] br[11] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_14 
+ bl[12] br[12] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_15 
+ bl[13] br[13] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_16 
+ bl[14] br[14] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_17 
+ bl[15] br[15] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_18 
+ bl[16] br[16] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_19 
+ bl[17] br[17] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_20 
+ bl[18] br[18] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_21 
+ bl[19] br[19] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_22 
+ bl[20] br[20] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_23 
+ bl[21] br[21] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_24 
+ bl[22] br[22] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_25 
+ bl[23] br[23] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_26 
+ bl[24] br[24] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_27 
+ bl[25] br[25] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_28 
+ bl[26] br[26] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_29 
+ bl[27] br[27] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_30 
+ bl[28] br[28] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_31 
+ bl[29] br[29] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_32 
+ bl[30] br[30] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_33 
+ bl[31] br[31] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_34 
+ bl[32] br[32] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_35 
+ bl[33] br[33] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_36 
+ bl[34] br[34] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_37 
+ bl[35] br[35] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_38 
+ bl[36] br[36] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_39 
+ bl[37] br[37] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_40 
+ bl[38] br[38] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_41 
+ bl[39] br[39] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_42 
+ bl[40] br[40] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_43 
+ bl[41] br[41] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_44 
+ bl[42] br[42] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_45 
+ bl[43] br[43] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_46 
+ bl[44] br[44] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_47 
+ bl[45] br[45] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_48 
+ bl[46] br[46] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_49 
+ bl[47] br[47] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_50 
+ bl[48] br[48] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_51 
+ bl[49] br[49] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_52 
+ bl[50] br[50] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_53 
+ bl[51] br[51] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_54 
+ bl[52] br[52] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_55 
+ bl[53] br[53] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_56 
+ bl[54] br[54] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_57 
+ bl[55] br[55] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_58 
+ bl[56] br[56] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_59 
+ bl[57] br[57] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_60 
+ bl[58] br[58] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_61 
+ bl[59] br[59] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_62 
+ bl[60] br[60] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_63 
+ bl[61] br[61] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_64 
+ bl[62] br[62] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_65 
+ bl[63] br[63] vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_66 
+ vdd vdd vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_456_67 
+ vdd vdd vdd vss wl[454] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_0 
+ vdd vdd vss vdd vpb vnb wl[455] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_457_1 
+ rbl rbr vss vdd vpb vnb wl[455] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_457_2 
+ bl[0] br[0] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_3 
+ bl[1] br[1] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_4 
+ bl[2] br[2] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_5 
+ bl[3] br[3] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_6 
+ bl[4] br[4] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_7 
+ bl[5] br[5] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_8 
+ bl[6] br[6] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_9 
+ bl[7] br[7] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_10 
+ bl[8] br[8] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_11 
+ bl[9] br[9] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_12 
+ bl[10] br[10] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_13 
+ bl[11] br[11] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_14 
+ bl[12] br[12] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_15 
+ bl[13] br[13] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_16 
+ bl[14] br[14] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_17 
+ bl[15] br[15] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_18 
+ bl[16] br[16] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_19 
+ bl[17] br[17] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_20 
+ bl[18] br[18] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_21 
+ bl[19] br[19] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_22 
+ bl[20] br[20] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_23 
+ bl[21] br[21] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_24 
+ bl[22] br[22] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_25 
+ bl[23] br[23] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_26 
+ bl[24] br[24] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_27 
+ bl[25] br[25] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_28 
+ bl[26] br[26] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_29 
+ bl[27] br[27] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_30 
+ bl[28] br[28] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_31 
+ bl[29] br[29] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_32 
+ bl[30] br[30] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_33 
+ bl[31] br[31] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_34 
+ bl[32] br[32] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_35 
+ bl[33] br[33] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_36 
+ bl[34] br[34] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_37 
+ bl[35] br[35] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_38 
+ bl[36] br[36] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_39 
+ bl[37] br[37] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_40 
+ bl[38] br[38] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_41 
+ bl[39] br[39] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_42 
+ bl[40] br[40] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_43 
+ bl[41] br[41] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_44 
+ bl[42] br[42] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_45 
+ bl[43] br[43] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_46 
+ bl[44] br[44] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_47 
+ bl[45] br[45] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_48 
+ bl[46] br[46] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_49 
+ bl[47] br[47] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_50 
+ bl[48] br[48] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_51 
+ bl[49] br[49] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_52 
+ bl[50] br[50] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_53 
+ bl[51] br[51] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_54 
+ bl[52] br[52] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_55 
+ bl[53] br[53] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_56 
+ bl[54] br[54] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_57 
+ bl[55] br[55] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_58 
+ bl[56] br[56] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_59 
+ bl[57] br[57] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_60 
+ bl[58] br[58] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_61 
+ bl[59] br[59] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_62 
+ bl[60] br[60] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_63 
+ bl[61] br[61] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_64 
+ bl[62] br[62] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_65 
+ bl[63] br[63] vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_66 
+ vdd vdd vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_457_67 
+ vdd vdd vdd vss wl[455] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_0 
+ vdd vdd vss vdd vpb vnb wl[456] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_458_1 
+ rbl rbr vss vdd vpb vnb wl[456] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_458_2 
+ bl[0] br[0] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_3 
+ bl[1] br[1] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_4 
+ bl[2] br[2] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_5 
+ bl[3] br[3] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_6 
+ bl[4] br[4] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_7 
+ bl[5] br[5] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_8 
+ bl[6] br[6] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_9 
+ bl[7] br[7] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_10 
+ bl[8] br[8] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_11 
+ bl[9] br[9] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_12 
+ bl[10] br[10] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_13 
+ bl[11] br[11] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_14 
+ bl[12] br[12] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_15 
+ bl[13] br[13] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_16 
+ bl[14] br[14] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_17 
+ bl[15] br[15] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_18 
+ bl[16] br[16] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_19 
+ bl[17] br[17] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_20 
+ bl[18] br[18] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_21 
+ bl[19] br[19] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_22 
+ bl[20] br[20] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_23 
+ bl[21] br[21] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_24 
+ bl[22] br[22] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_25 
+ bl[23] br[23] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_26 
+ bl[24] br[24] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_27 
+ bl[25] br[25] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_28 
+ bl[26] br[26] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_29 
+ bl[27] br[27] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_30 
+ bl[28] br[28] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_31 
+ bl[29] br[29] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_32 
+ bl[30] br[30] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_33 
+ bl[31] br[31] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_34 
+ bl[32] br[32] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_35 
+ bl[33] br[33] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_36 
+ bl[34] br[34] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_37 
+ bl[35] br[35] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_38 
+ bl[36] br[36] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_39 
+ bl[37] br[37] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_40 
+ bl[38] br[38] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_41 
+ bl[39] br[39] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_42 
+ bl[40] br[40] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_43 
+ bl[41] br[41] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_44 
+ bl[42] br[42] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_45 
+ bl[43] br[43] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_46 
+ bl[44] br[44] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_47 
+ bl[45] br[45] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_48 
+ bl[46] br[46] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_49 
+ bl[47] br[47] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_50 
+ bl[48] br[48] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_51 
+ bl[49] br[49] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_52 
+ bl[50] br[50] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_53 
+ bl[51] br[51] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_54 
+ bl[52] br[52] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_55 
+ bl[53] br[53] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_56 
+ bl[54] br[54] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_57 
+ bl[55] br[55] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_58 
+ bl[56] br[56] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_59 
+ bl[57] br[57] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_60 
+ bl[58] br[58] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_61 
+ bl[59] br[59] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_62 
+ bl[60] br[60] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_63 
+ bl[61] br[61] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_64 
+ bl[62] br[62] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_65 
+ bl[63] br[63] vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_66 
+ vdd vdd vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_458_67 
+ vdd vdd vdd vss wl[456] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_0 
+ vdd vdd vss vdd vpb vnb wl[457] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_459_1 
+ rbl rbr vss vdd vpb vnb wl[457] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_459_2 
+ bl[0] br[0] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_3 
+ bl[1] br[1] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_4 
+ bl[2] br[2] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_5 
+ bl[3] br[3] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_6 
+ bl[4] br[4] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_7 
+ bl[5] br[5] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_8 
+ bl[6] br[6] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_9 
+ bl[7] br[7] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_10 
+ bl[8] br[8] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_11 
+ bl[9] br[9] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_12 
+ bl[10] br[10] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_13 
+ bl[11] br[11] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_14 
+ bl[12] br[12] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_15 
+ bl[13] br[13] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_16 
+ bl[14] br[14] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_17 
+ bl[15] br[15] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_18 
+ bl[16] br[16] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_19 
+ bl[17] br[17] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_20 
+ bl[18] br[18] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_21 
+ bl[19] br[19] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_22 
+ bl[20] br[20] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_23 
+ bl[21] br[21] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_24 
+ bl[22] br[22] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_25 
+ bl[23] br[23] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_26 
+ bl[24] br[24] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_27 
+ bl[25] br[25] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_28 
+ bl[26] br[26] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_29 
+ bl[27] br[27] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_30 
+ bl[28] br[28] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_31 
+ bl[29] br[29] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_32 
+ bl[30] br[30] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_33 
+ bl[31] br[31] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_34 
+ bl[32] br[32] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_35 
+ bl[33] br[33] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_36 
+ bl[34] br[34] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_37 
+ bl[35] br[35] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_38 
+ bl[36] br[36] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_39 
+ bl[37] br[37] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_40 
+ bl[38] br[38] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_41 
+ bl[39] br[39] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_42 
+ bl[40] br[40] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_43 
+ bl[41] br[41] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_44 
+ bl[42] br[42] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_45 
+ bl[43] br[43] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_46 
+ bl[44] br[44] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_47 
+ bl[45] br[45] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_48 
+ bl[46] br[46] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_49 
+ bl[47] br[47] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_50 
+ bl[48] br[48] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_51 
+ bl[49] br[49] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_52 
+ bl[50] br[50] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_53 
+ bl[51] br[51] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_54 
+ bl[52] br[52] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_55 
+ bl[53] br[53] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_56 
+ bl[54] br[54] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_57 
+ bl[55] br[55] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_58 
+ bl[56] br[56] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_59 
+ bl[57] br[57] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_60 
+ bl[58] br[58] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_61 
+ bl[59] br[59] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_62 
+ bl[60] br[60] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_63 
+ bl[61] br[61] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_64 
+ bl[62] br[62] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_65 
+ bl[63] br[63] vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_66 
+ vdd vdd vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_459_67 
+ vdd vdd vdd vss wl[457] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_0 
+ vdd vdd vss vdd vpb vnb wl[458] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_460_1 
+ rbl rbr vss vdd vpb vnb wl[458] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_460_2 
+ bl[0] br[0] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_3 
+ bl[1] br[1] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_4 
+ bl[2] br[2] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_5 
+ bl[3] br[3] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_6 
+ bl[4] br[4] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_7 
+ bl[5] br[5] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_8 
+ bl[6] br[6] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_9 
+ bl[7] br[7] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_10 
+ bl[8] br[8] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_11 
+ bl[9] br[9] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_12 
+ bl[10] br[10] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_13 
+ bl[11] br[11] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_14 
+ bl[12] br[12] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_15 
+ bl[13] br[13] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_16 
+ bl[14] br[14] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_17 
+ bl[15] br[15] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_18 
+ bl[16] br[16] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_19 
+ bl[17] br[17] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_20 
+ bl[18] br[18] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_21 
+ bl[19] br[19] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_22 
+ bl[20] br[20] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_23 
+ bl[21] br[21] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_24 
+ bl[22] br[22] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_25 
+ bl[23] br[23] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_26 
+ bl[24] br[24] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_27 
+ bl[25] br[25] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_28 
+ bl[26] br[26] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_29 
+ bl[27] br[27] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_30 
+ bl[28] br[28] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_31 
+ bl[29] br[29] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_32 
+ bl[30] br[30] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_33 
+ bl[31] br[31] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_34 
+ bl[32] br[32] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_35 
+ bl[33] br[33] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_36 
+ bl[34] br[34] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_37 
+ bl[35] br[35] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_38 
+ bl[36] br[36] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_39 
+ bl[37] br[37] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_40 
+ bl[38] br[38] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_41 
+ bl[39] br[39] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_42 
+ bl[40] br[40] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_43 
+ bl[41] br[41] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_44 
+ bl[42] br[42] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_45 
+ bl[43] br[43] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_46 
+ bl[44] br[44] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_47 
+ bl[45] br[45] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_48 
+ bl[46] br[46] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_49 
+ bl[47] br[47] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_50 
+ bl[48] br[48] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_51 
+ bl[49] br[49] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_52 
+ bl[50] br[50] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_53 
+ bl[51] br[51] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_54 
+ bl[52] br[52] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_55 
+ bl[53] br[53] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_56 
+ bl[54] br[54] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_57 
+ bl[55] br[55] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_58 
+ bl[56] br[56] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_59 
+ bl[57] br[57] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_60 
+ bl[58] br[58] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_61 
+ bl[59] br[59] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_62 
+ bl[60] br[60] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_63 
+ bl[61] br[61] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_64 
+ bl[62] br[62] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_65 
+ bl[63] br[63] vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_66 
+ vdd vdd vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_460_67 
+ vdd vdd vdd vss wl[458] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_0 
+ vdd vdd vss vdd vpb vnb wl[459] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_461_1 
+ rbl rbr vss vdd vpb vnb wl[459] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_461_2 
+ bl[0] br[0] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_3 
+ bl[1] br[1] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_4 
+ bl[2] br[2] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_5 
+ bl[3] br[3] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_6 
+ bl[4] br[4] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_7 
+ bl[5] br[5] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_8 
+ bl[6] br[6] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_9 
+ bl[7] br[7] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_10 
+ bl[8] br[8] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_11 
+ bl[9] br[9] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_12 
+ bl[10] br[10] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_13 
+ bl[11] br[11] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_14 
+ bl[12] br[12] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_15 
+ bl[13] br[13] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_16 
+ bl[14] br[14] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_17 
+ bl[15] br[15] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_18 
+ bl[16] br[16] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_19 
+ bl[17] br[17] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_20 
+ bl[18] br[18] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_21 
+ bl[19] br[19] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_22 
+ bl[20] br[20] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_23 
+ bl[21] br[21] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_24 
+ bl[22] br[22] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_25 
+ bl[23] br[23] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_26 
+ bl[24] br[24] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_27 
+ bl[25] br[25] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_28 
+ bl[26] br[26] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_29 
+ bl[27] br[27] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_30 
+ bl[28] br[28] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_31 
+ bl[29] br[29] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_32 
+ bl[30] br[30] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_33 
+ bl[31] br[31] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_34 
+ bl[32] br[32] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_35 
+ bl[33] br[33] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_36 
+ bl[34] br[34] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_37 
+ bl[35] br[35] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_38 
+ bl[36] br[36] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_39 
+ bl[37] br[37] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_40 
+ bl[38] br[38] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_41 
+ bl[39] br[39] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_42 
+ bl[40] br[40] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_43 
+ bl[41] br[41] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_44 
+ bl[42] br[42] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_45 
+ bl[43] br[43] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_46 
+ bl[44] br[44] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_47 
+ bl[45] br[45] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_48 
+ bl[46] br[46] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_49 
+ bl[47] br[47] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_50 
+ bl[48] br[48] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_51 
+ bl[49] br[49] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_52 
+ bl[50] br[50] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_53 
+ bl[51] br[51] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_54 
+ bl[52] br[52] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_55 
+ bl[53] br[53] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_56 
+ bl[54] br[54] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_57 
+ bl[55] br[55] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_58 
+ bl[56] br[56] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_59 
+ bl[57] br[57] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_60 
+ bl[58] br[58] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_61 
+ bl[59] br[59] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_62 
+ bl[60] br[60] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_63 
+ bl[61] br[61] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_64 
+ bl[62] br[62] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_65 
+ bl[63] br[63] vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_66 
+ vdd vdd vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_461_67 
+ vdd vdd vdd vss wl[459] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_0 
+ vdd vdd vss vdd vpb vnb wl[460] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_462_1 
+ rbl rbr vss vdd vpb vnb wl[460] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_462_2 
+ bl[0] br[0] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_3 
+ bl[1] br[1] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_4 
+ bl[2] br[2] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_5 
+ bl[3] br[3] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_6 
+ bl[4] br[4] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_7 
+ bl[5] br[5] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_8 
+ bl[6] br[6] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_9 
+ bl[7] br[7] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_10 
+ bl[8] br[8] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_11 
+ bl[9] br[9] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_12 
+ bl[10] br[10] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_13 
+ bl[11] br[11] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_14 
+ bl[12] br[12] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_15 
+ bl[13] br[13] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_16 
+ bl[14] br[14] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_17 
+ bl[15] br[15] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_18 
+ bl[16] br[16] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_19 
+ bl[17] br[17] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_20 
+ bl[18] br[18] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_21 
+ bl[19] br[19] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_22 
+ bl[20] br[20] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_23 
+ bl[21] br[21] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_24 
+ bl[22] br[22] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_25 
+ bl[23] br[23] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_26 
+ bl[24] br[24] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_27 
+ bl[25] br[25] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_28 
+ bl[26] br[26] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_29 
+ bl[27] br[27] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_30 
+ bl[28] br[28] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_31 
+ bl[29] br[29] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_32 
+ bl[30] br[30] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_33 
+ bl[31] br[31] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_34 
+ bl[32] br[32] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_35 
+ bl[33] br[33] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_36 
+ bl[34] br[34] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_37 
+ bl[35] br[35] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_38 
+ bl[36] br[36] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_39 
+ bl[37] br[37] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_40 
+ bl[38] br[38] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_41 
+ bl[39] br[39] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_42 
+ bl[40] br[40] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_43 
+ bl[41] br[41] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_44 
+ bl[42] br[42] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_45 
+ bl[43] br[43] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_46 
+ bl[44] br[44] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_47 
+ bl[45] br[45] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_48 
+ bl[46] br[46] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_49 
+ bl[47] br[47] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_50 
+ bl[48] br[48] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_51 
+ bl[49] br[49] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_52 
+ bl[50] br[50] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_53 
+ bl[51] br[51] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_54 
+ bl[52] br[52] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_55 
+ bl[53] br[53] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_56 
+ bl[54] br[54] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_57 
+ bl[55] br[55] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_58 
+ bl[56] br[56] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_59 
+ bl[57] br[57] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_60 
+ bl[58] br[58] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_61 
+ bl[59] br[59] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_62 
+ bl[60] br[60] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_63 
+ bl[61] br[61] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_64 
+ bl[62] br[62] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_65 
+ bl[63] br[63] vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_66 
+ vdd vdd vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_462_67 
+ vdd vdd vdd vss wl[460] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_0 
+ vdd vdd vss vdd vpb vnb wl[461] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_463_1 
+ rbl rbr vss vdd vpb vnb wl[461] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_463_2 
+ bl[0] br[0] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_3 
+ bl[1] br[1] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_4 
+ bl[2] br[2] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_5 
+ bl[3] br[3] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_6 
+ bl[4] br[4] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_7 
+ bl[5] br[5] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_8 
+ bl[6] br[6] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_9 
+ bl[7] br[7] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_10 
+ bl[8] br[8] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_11 
+ bl[9] br[9] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_12 
+ bl[10] br[10] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_13 
+ bl[11] br[11] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_14 
+ bl[12] br[12] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_15 
+ bl[13] br[13] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_16 
+ bl[14] br[14] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_17 
+ bl[15] br[15] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_18 
+ bl[16] br[16] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_19 
+ bl[17] br[17] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_20 
+ bl[18] br[18] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_21 
+ bl[19] br[19] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_22 
+ bl[20] br[20] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_23 
+ bl[21] br[21] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_24 
+ bl[22] br[22] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_25 
+ bl[23] br[23] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_26 
+ bl[24] br[24] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_27 
+ bl[25] br[25] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_28 
+ bl[26] br[26] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_29 
+ bl[27] br[27] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_30 
+ bl[28] br[28] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_31 
+ bl[29] br[29] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_32 
+ bl[30] br[30] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_33 
+ bl[31] br[31] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_34 
+ bl[32] br[32] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_35 
+ bl[33] br[33] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_36 
+ bl[34] br[34] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_37 
+ bl[35] br[35] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_38 
+ bl[36] br[36] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_39 
+ bl[37] br[37] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_40 
+ bl[38] br[38] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_41 
+ bl[39] br[39] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_42 
+ bl[40] br[40] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_43 
+ bl[41] br[41] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_44 
+ bl[42] br[42] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_45 
+ bl[43] br[43] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_46 
+ bl[44] br[44] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_47 
+ bl[45] br[45] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_48 
+ bl[46] br[46] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_49 
+ bl[47] br[47] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_50 
+ bl[48] br[48] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_51 
+ bl[49] br[49] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_52 
+ bl[50] br[50] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_53 
+ bl[51] br[51] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_54 
+ bl[52] br[52] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_55 
+ bl[53] br[53] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_56 
+ bl[54] br[54] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_57 
+ bl[55] br[55] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_58 
+ bl[56] br[56] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_59 
+ bl[57] br[57] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_60 
+ bl[58] br[58] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_61 
+ bl[59] br[59] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_62 
+ bl[60] br[60] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_63 
+ bl[61] br[61] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_64 
+ bl[62] br[62] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_65 
+ bl[63] br[63] vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_66 
+ vdd vdd vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_463_67 
+ vdd vdd vdd vss wl[461] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_0 
+ vdd vdd vss vdd vpb vnb wl[462] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_464_1 
+ rbl rbr vss vdd vpb vnb wl[462] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_464_2 
+ bl[0] br[0] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_3 
+ bl[1] br[1] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_4 
+ bl[2] br[2] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_5 
+ bl[3] br[3] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_6 
+ bl[4] br[4] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_7 
+ bl[5] br[5] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_8 
+ bl[6] br[6] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_9 
+ bl[7] br[7] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_10 
+ bl[8] br[8] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_11 
+ bl[9] br[9] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_12 
+ bl[10] br[10] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_13 
+ bl[11] br[11] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_14 
+ bl[12] br[12] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_15 
+ bl[13] br[13] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_16 
+ bl[14] br[14] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_17 
+ bl[15] br[15] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_18 
+ bl[16] br[16] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_19 
+ bl[17] br[17] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_20 
+ bl[18] br[18] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_21 
+ bl[19] br[19] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_22 
+ bl[20] br[20] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_23 
+ bl[21] br[21] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_24 
+ bl[22] br[22] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_25 
+ bl[23] br[23] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_26 
+ bl[24] br[24] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_27 
+ bl[25] br[25] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_28 
+ bl[26] br[26] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_29 
+ bl[27] br[27] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_30 
+ bl[28] br[28] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_31 
+ bl[29] br[29] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_32 
+ bl[30] br[30] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_33 
+ bl[31] br[31] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_34 
+ bl[32] br[32] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_35 
+ bl[33] br[33] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_36 
+ bl[34] br[34] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_37 
+ bl[35] br[35] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_38 
+ bl[36] br[36] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_39 
+ bl[37] br[37] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_40 
+ bl[38] br[38] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_41 
+ bl[39] br[39] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_42 
+ bl[40] br[40] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_43 
+ bl[41] br[41] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_44 
+ bl[42] br[42] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_45 
+ bl[43] br[43] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_46 
+ bl[44] br[44] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_47 
+ bl[45] br[45] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_48 
+ bl[46] br[46] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_49 
+ bl[47] br[47] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_50 
+ bl[48] br[48] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_51 
+ bl[49] br[49] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_52 
+ bl[50] br[50] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_53 
+ bl[51] br[51] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_54 
+ bl[52] br[52] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_55 
+ bl[53] br[53] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_56 
+ bl[54] br[54] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_57 
+ bl[55] br[55] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_58 
+ bl[56] br[56] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_59 
+ bl[57] br[57] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_60 
+ bl[58] br[58] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_61 
+ bl[59] br[59] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_62 
+ bl[60] br[60] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_63 
+ bl[61] br[61] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_64 
+ bl[62] br[62] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_65 
+ bl[63] br[63] vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_66 
+ vdd vdd vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_464_67 
+ vdd vdd vdd vss wl[462] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_0 
+ vdd vdd vss vdd vpb vnb wl[463] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_465_1 
+ rbl rbr vss vdd vpb vnb wl[463] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_465_2 
+ bl[0] br[0] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_3 
+ bl[1] br[1] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_4 
+ bl[2] br[2] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_5 
+ bl[3] br[3] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_6 
+ bl[4] br[4] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_7 
+ bl[5] br[5] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_8 
+ bl[6] br[6] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_9 
+ bl[7] br[7] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_10 
+ bl[8] br[8] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_11 
+ bl[9] br[9] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_12 
+ bl[10] br[10] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_13 
+ bl[11] br[11] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_14 
+ bl[12] br[12] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_15 
+ bl[13] br[13] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_16 
+ bl[14] br[14] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_17 
+ bl[15] br[15] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_18 
+ bl[16] br[16] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_19 
+ bl[17] br[17] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_20 
+ bl[18] br[18] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_21 
+ bl[19] br[19] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_22 
+ bl[20] br[20] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_23 
+ bl[21] br[21] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_24 
+ bl[22] br[22] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_25 
+ bl[23] br[23] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_26 
+ bl[24] br[24] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_27 
+ bl[25] br[25] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_28 
+ bl[26] br[26] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_29 
+ bl[27] br[27] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_30 
+ bl[28] br[28] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_31 
+ bl[29] br[29] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_32 
+ bl[30] br[30] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_33 
+ bl[31] br[31] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_34 
+ bl[32] br[32] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_35 
+ bl[33] br[33] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_36 
+ bl[34] br[34] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_37 
+ bl[35] br[35] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_38 
+ bl[36] br[36] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_39 
+ bl[37] br[37] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_40 
+ bl[38] br[38] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_41 
+ bl[39] br[39] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_42 
+ bl[40] br[40] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_43 
+ bl[41] br[41] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_44 
+ bl[42] br[42] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_45 
+ bl[43] br[43] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_46 
+ bl[44] br[44] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_47 
+ bl[45] br[45] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_48 
+ bl[46] br[46] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_49 
+ bl[47] br[47] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_50 
+ bl[48] br[48] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_51 
+ bl[49] br[49] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_52 
+ bl[50] br[50] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_53 
+ bl[51] br[51] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_54 
+ bl[52] br[52] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_55 
+ bl[53] br[53] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_56 
+ bl[54] br[54] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_57 
+ bl[55] br[55] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_58 
+ bl[56] br[56] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_59 
+ bl[57] br[57] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_60 
+ bl[58] br[58] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_61 
+ bl[59] br[59] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_62 
+ bl[60] br[60] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_63 
+ bl[61] br[61] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_64 
+ bl[62] br[62] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_65 
+ bl[63] br[63] vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_66 
+ vdd vdd vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_465_67 
+ vdd vdd vdd vss wl[463] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_0 
+ vdd vdd vss vdd vpb vnb wl[464] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_466_1 
+ rbl rbr vss vdd vpb vnb wl[464] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_466_2 
+ bl[0] br[0] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_3 
+ bl[1] br[1] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_4 
+ bl[2] br[2] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_5 
+ bl[3] br[3] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_6 
+ bl[4] br[4] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_7 
+ bl[5] br[5] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_8 
+ bl[6] br[6] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_9 
+ bl[7] br[7] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_10 
+ bl[8] br[8] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_11 
+ bl[9] br[9] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_12 
+ bl[10] br[10] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_13 
+ bl[11] br[11] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_14 
+ bl[12] br[12] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_15 
+ bl[13] br[13] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_16 
+ bl[14] br[14] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_17 
+ bl[15] br[15] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_18 
+ bl[16] br[16] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_19 
+ bl[17] br[17] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_20 
+ bl[18] br[18] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_21 
+ bl[19] br[19] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_22 
+ bl[20] br[20] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_23 
+ bl[21] br[21] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_24 
+ bl[22] br[22] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_25 
+ bl[23] br[23] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_26 
+ bl[24] br[24] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_27 
+ bl[25] br[25] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_28 
+ bl[26] br[26] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_29 
+ bl[27] br[27] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_30 
+ bl[28] br[28] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_31 
+ bl[29] br[29] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_32 
+ bl[30] br[30] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_33 
+ bl[31] br[31] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_34 
+ bl[32] br[32] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_35 
+ bl[33] br[33] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_36 
+ bl[34] br[34] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_37 
+ bl[35] br[35] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_38 
+ bl[36] br[36] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_39 
+ bl[37] br[37] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_40 
+ bl[38] br[38] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_41 
+ bl[39] br[39] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_42 
+ bl[40] br[40] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_43 
+ bl[41] br[41] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_44 
+ bl[42] br[42] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_45 
+ bl[43] br[43] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_46 
+ bl[44] br[44] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_47 
+ bl[45] br[45] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_48 
+ bl[46] br[46] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_49 
+ bl[47] br[47] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_50 
+ bl[48] br[48] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_51 
+ bl[49] br[49] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_52 
+ bl[50] br[50] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_53 
+ bl[51] br[51] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_54 
+ bl[52] br[52] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_55 
+ bl[53] br[53] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_56 
+ bl[54] br[54] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_57 
+ bl[55] br[55] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_58 
+ bl[56] br[56] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_59 
+ bl[57] br[57] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_60 
+ bl[58] br[58] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_61 
+ bl[59] br[59] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_62 
+ bl[60] br[60] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_63 
+ bl[61] br[61] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_64 
+ bl[62] br[62] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_65 
+ bl[63] br[63] vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_66 
+ vdd vdd vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_466_67 
+ vdd vdd vdd vss wl[464] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_0 
+ vdd vdd vss vdd vpb vnb wl[465] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_467_1 
+ rbl rbr vss vdd vpb vnb wl[465] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_467_2 
+ bl[0] br[0] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_3 
+ bl[1] br[1] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_4 
+ bl[2] br[2] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_5 
+ bl[3] br[3] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_6 
+ bl[4] br[4] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_7 
+ bl[5] br[5] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_8 
+ bl[6] br[6] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_9 
+ bl[7] br[7] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_10 
+ bl[8] br[8] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_11 
+ bl[9] br[9] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_12 
+ bl[10] br[10] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_13 
+ bl[11] br[11] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_14 
+ bl[12] br[12] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_15 
+ bl[13] br[13] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_16 
+ bl[14] br[14] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_17 
+ bl[15] br[15] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_18 
+ bl[16] br[16] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_19 
+ bl[17] br[17] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_20 
+ bl[18] br[18] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_21 
+ bl[19] br[19] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_22 
+ bl[20] br[20] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_23 
+ bl[21] br[21] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_24 
+ bl[22] br[22] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_25 
+ bl[23] br[23] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_26 
+ bl[24] br[24] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_27 
+ bl[25] br[25] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_28 
+ bl[26] br[26] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_29 
+ bl[27] br[27] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_30 
+ bl[28] br[28] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_31 
+ bl[29] br[29] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_32 
+ bl[30] br[30] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_33 
+ bl[31] br[31] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_34 
+ bl[32] br[32] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_35 
+ bl[33] br[33] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_36 
+ bl[34] br[34] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_37 
+ bl[35] br[35] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_38 
+ bl[36] br[36] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_39 
+ bl[37] br[37] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_40 
+ bl[38] br[38] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_41 
+ bl[39] br[39] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_42 
+ bl[40] br[40] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_43 
+ bl[41] br[41] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_44 
+ bl[42] br[42] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_45 
+ bl[43] br[43] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_46 
+ bl[44] br[44] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_47 
+ bl[45] br[45] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_48 
+ bl[46] br[46] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_49 
+ bl[47] br[47] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_50 
+ bl[48] br[48] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_51 
+ bl[49] br[49] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_52 
+ bl[50] br[50] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_53 
+ bl[51] br[51] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_54 
+ bl[52] br[52] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_55 
+ bl[53] br[53] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_56 
+ bl[54] br[54] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_57 
+ bl[55] br[55] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_58 
+ bl[56] br[56] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_59 
+ bl[57] br[57] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_60 
+ bl[58] br[58] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_61 
+ bl[59] br[59] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_62 
+ bl[60] br[60] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_63 
+ bl[61] br[61] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_64 
+ bl[62] br[62] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_65 
+ bl[63] br[63] vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_66 
+ vdd vdd vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_467_67 
+ vdd vdd vdd vss wl[465] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_0 
+ vdd vdd vss vdd vpb vnb wl[466] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_468_1 
+ rbl rbr vss vdd vpb vnb wl[466] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_468_2 
+ bl[0] br[0] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_3 
+ bl[1] br[1] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_4 
+ bl[2] br[2] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_5 
+ bl[3] br[3] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_6 
+ bl[4] br[4] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_7 
+ bl[5] br[5] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_8 
+ bl[6] br[6] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_9 
+ bl[7] br[7] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_10 
+ bl[8] br[8] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_11 
+ bl[9] br[9] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_12 
+ bl[10] br[10] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_13 
+ bl[11] br[11] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_14 
+ bl[12] br[12] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_15 
+ bl[13] br[13] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_16 
+ bl[14] br[14] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_17 
+ bl[15] br[15] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_18 
+ bl[16] br[16] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_19 
+ bl[17] br[17] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_20 
+ bl[18] br[18] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_21 
+ bl[19] br[19] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_22 
+ bl[20] br[20] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_23 
+ bl[21] br[21] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_24 
+ bl[22] br[22] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_25 
+ bl[23] br[23] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_26 
+ bl[24] br[24] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_27 
+ bl[25] br[25] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_28 
+ bl[26] br[26] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_29 
+ bl[27] br[27] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_30 
+ bl[28] br[28] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_31 
+ bl[29] br[29] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_32 
+ bl[30] br[30] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_33 
+ bl[31] br[31] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_34 
+ bl[32] br[32] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_35 
+ bl[33] br[33] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_36 
+ bl[34] br[34] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_37 
+ bl[35] br[35] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_38 
+ bl[36] br[36] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_39 
+ bl[37] br[37] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_40 
+ bl[38] br[38] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_41 
+ bl[39] br[39] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_42 
+ bl[40] br[40] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_43 
+ bl[41] br[41] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_44 
+ bl[42] br[42] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_45 
+ bl[43] br[43] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_46 
+ bl[44] br[44] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_47 
+ bl[45] br[45] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_48 
+ bl[46] br[46] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_49 
+ bl[47] br[47] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_50 
+ bl[48] br[48] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_51 
+ bl[49] br[49] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_52 
+ bl[50] br[50] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_53 
+ bl[51] br[51] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_54 
+ bl[52] br[52] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_55 
+ bl[53] br[53] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_56 
+ bl[54] br[54] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_57 
+ bl[55] br[55] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_58 
+ bl[56] br[56] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_59 
+ bl[57] br[57] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_60 
+ bl[58] br[58] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_61 
+ bl[59] br[59] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_62 
+ bl[60] br[60] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_63 
+ bl[61] br[61] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_64 
+ bl[62] br[62] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_65 
+ bl[63] br[63] vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_66 
+ vdd vdd vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_468_67 
+ vdd vdd vdd vss wl[466] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_0 
+ vdd vdd vss vdd vpb vnb wl[467] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_469_1 
+ rbl rbr vss vdd vpb vnb wl[467] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_469_2 
+ bl[0] br[0] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_3 
+ bl[1] br[1] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_4 
+ bl[2] br[2] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_5 
+ bl[3] br[3] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_6 
+ bl[4] br[4] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_7 
+ bl[5] br[5] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_8 
+ bl[6] br[6] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_9 
+ bl[7] br[7] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_10 
+ bl[8] br[8] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_11 
+ bl[9] br[9] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_12 
+ bl[10] br[10] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_13 
+ bl[11] br[11] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_14 
+ bl[12] br[12] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_15 
+ bl[13] br[13] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_16 
+ bl[14] br[14] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_17 
+ bl[15] br[15] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_18 
+ bl[16] br[16] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_19 
+ bl[17] br[17] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_20 
+ bl[18] br[18] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_21 
+ bl[19] br[19] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_22 
+ bl[20] br[20] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_23 
+ bl[21] br[21] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_24 
+ bl[22] br[22] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_25 
+ bl[23] br[23] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_26 
+ bl[24] br[24] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_27 
+ bl[25] br[25] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_28 
+ bl[26] br[26] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_29 
+ bl[27] br[27] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_30 
+ bl[28] br[28] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_31 
+ bl[29] br[29] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_32 
+ bl[30] br[30] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_33 
+ bl[31] br[31] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_34 
+ bl[32] br[32] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_35 
+ bl[33] br[33] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_36 
+ bl[34] br[34] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_37 
+ bl[35] br[35] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_38 
+ bl[36] br[36] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_39 
+ bl[37] br[37] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_40 
+ bl[38] br[38] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_41 
+ bl[39] br[39] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_42 
+ bl[40] br[40] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_43 
+ bl[41] br[41] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_44 
+ bl[42] br[42] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_45 
+ bl[43] br[43] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_46 
+ bl[44] br[44] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_47 
+ bl[45] br[45] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_48 
+ bl[46] br[46] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_49 
+ bl[47] br[47] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_50 
+ bl[48] br[48] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_51 
+ bl[49] br[49] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_52 
+ bl[50] br[50] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_53 
+ bl[51] br[51] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_54 
+ bl[52] br[52] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_55 
+ bl[53] br[53] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_56 
+ bl[54] br[54] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_57 
+ bl[55] br[55] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_58 
+ bl[56] br[56] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_59 
+ bl[57] br[57] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_60 
+ bl[58] br[58] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_61 
+ bl[59] br[59] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_62 
+ bl[60] br[60] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_63 
+ bl[61] br[61] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_64 
+ bl[62] br[62] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_65 
+ bl[63] br[63] vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_66 
+ vdd vdd vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_469_67 
+ vdd vdd vdd vss wl[467] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_0 
+ vdd vdd vss vdd vpb vnb wl[468] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_470_1 
+ rbl rbr vss vdd vpb vnb wl[468] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_470_2 
+ bl[0] br[0] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_3 
+ bl[1] br[1] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_4 
+ bl[2] br[2] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_5 
+ bl[3] br[3] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_6 
+ bl[4] br[4] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_7 
+ bl[5] br[5] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_8 
+ bl[6] br[6] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_9 
+ bl[7] br[7] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_10 
+ bl[8] br[8] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_11 
+ bl[9] br[9] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_12 
+ bl[10] br[10] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_13 
+ bl[11] br[11] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_14 
+ bl[12] br[12] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_15 
+ bl[13] br[13] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_16 
+ bl[14] br[14] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_17 
+ bl[15] br[15] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_18 
+ bl[16] br[16] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_19 
+ bl[17] br[17] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_20 
+ bl[18] br[18] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_21 
+ bl[19] br[19] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_22 
+ bl[20] br[20] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_23 
+ bl[21] br[21] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_24 
+ bl[22] br[22] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_25 
+ bl[23] br[23] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_26 
+ bl[24] br[24] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_27 
+ bl[25] br[25] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_28 
+ bl[26] br[26] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_29 
+ bl[27] br[27] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_30 
+ bl[28] br[28] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_31 
+ bl[29] br[29] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_32 
+ bl[30] br[30] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_33 
+ bl[31] br[31] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_34 
+ bl[32] br[32] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_35 
+ bl[33] br[33] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_36 
+ bl[34] br[34] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_37 
+ bl[35] br[35] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_38 
+ bl[36] br[36] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_39 
+ bl[37] br[37] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_40 
+ bl[38] br[38] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_41 
+ bl[39] br[39] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_42 
+ bl[40] br[40] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_43 
+ bl[41] br[41] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_44 
+ bl[42] br[42] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_45 
+ bl[43] br[43] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_46 
+ bl[44] br[44] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_47 
+ bl[45] br[45] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_48 
+ bl[46] br[46] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_49 
+ bl[47] br[47] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_50 
+ bl[48] br[48] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_51 
+ bl[49] br[49] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_52 
+ bl[50] br[50] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_53 
+ bl[51] br[51] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_54 
+ bl[52] br[52] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_55 
+ bl[53] br[53] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_56 
+ bl[54] br[54] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_57 
+ bl[55] br[55] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_58 
+ bl[56] br[56] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_59 
+ bl[57] br[57] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_60 
+ bl[58] br[58] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_61 
+ bl[59] br[59] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_62 
+ bl[60] br[60] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_63 
+ bl[61] br[61] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_64 
+ bl[62] br[62] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_65 
+ bl[63] br[63] vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_66 
+ vdd vdd vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_470_67 
+ vdd vdd vdd vss wl[468] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_0 
+ vdd vdd vss vdd vpb vnb wl[469] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_471_1 
+ rbl rbr vss vdd vpb vnb wl[469] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_471_2 
+ bl[0] br[0] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_3 
+ bl[1] br[1] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_4 
+ bl[2] br[2] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_5 
+ bl[3] br[3] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_6 
+ bl[4] br[4] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_7 
+ bl[5] br[5] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_8 
+ bl[6] br[6] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_9 
+ bl[7] br[7] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_10 
+ bl[8] br[8] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_11 
+ bl[9] br[9] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_12 
+ bl[10] br[10] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_13 
+ bl[11] br[11] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_14 
+ bl[12] br[12] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_15 
+ bl[13] br[13] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_16 
+ bl[14] br[14] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_17 
+ bl[15] br[15] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_18 
+ bl[16] br[16] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_19 
+ bl[17] br[17] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_20 
+ bl[18] br[18] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_21 
+ bl[19] br[19] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_22 
+ bl[20] br[20] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_23 
+ bl[21] br[21] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_24 
+ bl[22] br[22] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_25 
+ bl[23] br[23] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_26 
+ bl[24] br[24] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_27 
+ bl[25] br[25] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_28 
+ bl[26] br[26] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_29 
+ bl[27] br[27] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_30 
+ bl[28] br[28] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_31 
+ bl[29] br[29] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_32 
+ bl[30] br[30] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_33 
+ bl[31] br[31] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_34 
+ bl[32] br[32] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_35 
+ bl[33] br[33] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_36 
+ bl[34] br[34] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_37 
+ bl[35] br[35] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_38 
+ bl[36] br[36] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_39 
+ bl[37] br[37] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_40 
+ bl[38] br[38] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_41 
+ bl[39] br[39] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_42 
+ bl[40] br[40] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_43 
+ bl[41] br[41] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_44 
+ bl[42] br[42] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_45 
+ bl[43] br[43] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_46 
+ bl[44] br[44] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_47 
+ bl[45] br[45] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_48 
+ bl[46] br[46] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_49 
+ bl[47] br[47] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_50 
+ bl[48] br[48] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_51 
+ bl[49] br[49] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_52 
+ bl[50] br[50] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_53 
+ bl[51] br[51] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_54 
+ bl[52] br[52] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_55 
+ bl[53] br[53] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_56 
+ bl[54] br[54] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_57 
+ bl[55] br[55] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_58 
+ bl[56] br[56] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_59 
+ bl[57] br[57] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_60 
+ bl[58] br[58] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_61 
+ bl[59] br[59] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_62 
+ bl[60] br[60] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_63 
+ bl[61] br[61] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_64 
+ bl[62] br[62] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_65 
+ bl[63] br[63] vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_66 
+ vdd vdd vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_471_67 
+ vdd vdd vdd vss wl[469] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_0 
+ vdd vdd vss vdd vpb vnb wl[470] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_472_1 
+ rbl rbr vss vdd vpb vnb wl[470] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_472_2 
+ bl[0] br[0] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_3 
+ bl[1] br[1] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_4 
+ bl[2] br[2] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_5 
+ bl[3] br[3] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_6 
+ bl[4] br[4] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_7 
+ bl[5] br[5] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_8 
+ bl[6] br[6] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_9 
+ bl[7] br[7] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_10 
+ bl[8] br[8] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_11 
+ bl[9] br[9] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_12 
+ bl[10] br[10] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_13 
+ bl[11] br[11] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_14 
+ bl[12] br[12] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_15 
+ bl[13] br[13] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_16 
+ bl[14] br[14] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_17 
+ bl[15] br[15] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_18 
+ bl[16] br[16] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_19 
+ bl[17] br[17] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_20 
+ bl[18] br[18] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_21 
+ bl[19] br[19] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_22 
+ bl[20] br[20] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_23 
+ bl[21] br[21] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_24 
+ bl[22] br[22] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_25 
+ bl[23] br[23] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_26 
+ bl[24] br[24] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_27 
+ bl[25] br[25] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_28 
+ bl[26] br[26] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_29 
+ bl[27] br[27] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_30 
+ bl[28] br[28] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_31 
+ bl[29] br[29] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_32 
+ bl[30] br[30] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_33 
+ bl[31] br[31] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_34 
+ bl[32] br[32] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_35 
+ bl[33] br[33] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_36 
+ bl[34] br[34] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_37 
+ bl[35] br[35] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_38 
+ bl[36] br[36] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_39 
+ bl[37] br[37] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_40 
+ bl[38] br[38] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_41 
+ bl[39] br[39] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_42 
+ bl[40] br[40] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_43 
+ bl[41] br[41] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_44 
+ bl[42] br[42] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_45 
+ bl[43] br[43] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_46 
+ bl[44] br[44] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_47 
+ bl[45] br[45] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_48 
+ bl[46] br[46] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_49 
+ bl[47] br[47] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_50 
+ bl[48] br[48] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_51 
+ bl[49] br[49] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_52 
+ bl[50] br[50] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_53 
+ bl[51] br[51] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_54 
+ bl[52] br[52] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_55 
+ bl[53] br[53] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_56 
+ bl[54] br[54] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_57 
+ bl[55] br[55] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_58 
+ bl[56] br[56] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_59 
+ bl[57] br[57] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_60 
+ bl[58] br[58] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_61 
+ bl[59] br[59] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_62 
+ bl[60] br[60] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_63 
+ bl[61] br[61] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_64 
+ bl[62] br[62] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_65 
+ bl[63] br[63] vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_66 
+ vdd vdd vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_472_67 
+ vdd vdd vdd vss wl[470] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_0 
+ vdd vdd vss vdd vpb vnb wl[471] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_473_1 
+ rbl rbr vss vdd vpb vnb wl[471] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_473_2 
+ bl[0] br[0] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_3 
+ bl[1] br[1] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_4 
+ bl[2] br[2] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_5 
+ bl[3] br[3] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_6 
+ bl[4] br[4] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_7 
+ bl[5] br[5] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_8 
+ bl[6] br[6] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_9 
+ bl[7] br[7] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_10 
+ bl[8] br[8] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_11 
+ bl[9] br[9] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_12 
+ bl[10] br[10] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_13 
+ bl[11] br[11] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_14 
+ bl[12] br[12] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_15 
+ bl[13] br[13] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_16 
+ bl[14] br[14] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_17 
+ bl[15] br[15] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_18 
+ bl[16] br[16] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_19 
+ bl[17] br[17] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_20 
+ bl[18] br[18] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_21 
+ bl[19] br[19] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_22 
+ bl[20] br[20] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_23 
+ bl[21] br[21] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_24 
+ bl[22] br[22] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_25 
+ bl[23] br[23] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_26 
+ bl[24] br[24] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_27 
+ bl[25] br[25] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_28 
+ bl[26] br[26] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_29 
+ bl[27] br[27] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_30 
+ bl[28] br[28] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_31 
+ bl[29] br[29] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_32 
+ bl[30] br[30] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_33 
+ bl[31] br[31] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_34 
+ bl[32] br[32] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_35 
+ bl[33] br[33] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_36 
+ bl[34] br[34] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_37 
+ bl[35] br[35] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_38 
+ bl[36] br[36] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_39 
+ bl[37] br[37] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_40 
+ bl[38] br[38] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_41 
+ bl[39] br[39] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_42 
+ bl[40] br[40] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_43 
+ bl[41] br[41] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_44 
+ bl[42] br[42] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_45 
+ bl[43] br[43] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_46 
+ bl[44] br[44] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_47 
+ bl[45] br[45] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_48 
+ bl[46] br[46] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_49 
+ bl[47] br[47] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_50 
+ bl[48] br[48] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_51 
+ bl[49] br[49] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_52 
+ bl[50] br[50] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_53 
+ bl[51] br[51] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_54 
+ bl[52] br[52] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_55 
+ bl[53] br[53] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_56 
+ bl[54] br[54] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_57 
+ bl[55] br[55] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_58 
+ bl[56] br[56] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_59 
+ bl[57] br[57] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_60 
+ bl[58] br[58] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_61 
+ bl[59] br[59] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_62 
+ bl[60] br[60] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_63 
+ bl[61] br[61] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_64 
+ bl[62] br[62] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_65 
+ bl[63] br[63] vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_66 
+ vdd vdd vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_473_67 
+ vdd vdd vdd vss wl[471] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_0 
+ vdd vdd vss vdd vpb vnb wl[472] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_474_1 
+ rbl rbr vss vdd vpb vnb wl[472] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_474_2 
+ bl[0] br[0] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_3 
+ bl[1] br[1] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_4 
+ bl[2] br[2] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_5 
+ bl[3] br[3] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_6 
+ bl[4] br[4] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_7 
+ bl[5] br[5] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_8 
+ bl[6] br[6] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_9 
+ bl[7] br[7] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_10 
+ bl[8] br[8] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_11 
+ bl[9] br[9] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_12 
+ bl[10] br[10] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_13 
+ bl[11] br[11] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_14 
+ bl[12] br[12] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_15 
+ bl[13] br[13] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_16 
+ bl[14] br[14] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_17 
+ bl[15] br[15] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_18 
+ bl[16] br[16] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_19 
+ bl[17] br[17] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_20 
+ bl[18] br[18] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_21 
+ bl[19] br[19] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_22 
+ bl[20] br[20] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_23 
+ bl[21] br[21] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_24 
+ bl[22] br[22] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_25 
+ bl[23] br[23] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_26 
+ bl[24] br[24] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_27 
+ bl[25] br[25] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_28 
+ bl[26] br[26] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_29 
+ bl[27] br[27] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_30 
+ bl[28] br[28] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_31 
+ bl[29] br[29] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_32 
+ bl[30] br[30] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_33 
+ bl[31] br[31] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_34 
+ bl[32] br[32] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_35 
+ bl[33] br[33] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_36 
+ bl[34] br[34] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_37 
+ bl[35] br[35] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_38 
+ bl[36] br[36] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_39 
+ bl[37] br[37] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_40 
+ bl[38] br[38] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_41 
+ bl[39] br[39] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_42 
+ bl[40] br[40] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_43 
+ bl[41] br[41] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_44 
+ bl[42] br[42] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_45 
+ bl[43] br[43] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_46 
+ bl[44] br[44] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_47 
+ bl[45] br[45] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_48 
+ bl[46] br[46] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_49 
+ bl[47] br[47] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_50 
+ bl[48] br[48] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_51 
+ bl[49] br[49] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_52 
+ bl[50] br[50] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_53 
+ bl[51] br[51] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_54 
+ bl[52] br[52] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_55 
+ bl[53] br[53] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_56 
+ bl[54] br[54] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_57 
+ bl[55] br[55] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_58 
+ bl[56] br[56] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_59 
+ bl[57] br[57] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_60 
+ bl[58] br[58] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_61 
+ bl[59] br[59] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_62 
+ bl[60] br[60] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_63 
+ bl[61] br[61] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_64 
+ bl[62] br[62] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_65 
+ bl[63] br[63] vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_66 
+ vdd vdd vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_474_67 
+ vdd vdd vdd vss wl[472] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_0 
+ vdd vdd vss vdd vpb vnb wl[473] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_475_1 
+ rbl rbr vss vdd vpb vnb wl[473] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_475_2 
+ bl[0] br[0] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_3 
+ bl[1] br[1] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_4 
+ bl[2] br[2] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_5 
+ bl[3] br[3] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_6 
+ bl[4] br[4] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_7 
+ bl[5] br[5] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_8 
+ bl[6] br[6] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_9 
+ bl[7] br[7] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_10 
+ bl[8] br[8] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_11 
+ bl[9] br[9] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_12 
+ bl[10] br[10] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_13 
+ bl[11] br[11] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_14 
+ bl[12] br[12] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_15 
+ bl[13] br[13] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_16 
+ bl[14] br[14] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_17 
+ bl[15] br[15] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_18 
+ bl[16] br[16] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_19 
+ bl[17] br[17] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_20 
+ bl[18] br[18] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_21 
+ bl[19] br[19] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_22 
+ bl[20] br[20] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_23 
+ bl[21] br[21] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_24 
+ bl[22] br[22] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_25 
+ bl[23] br[23] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_26 
+ bl[24] br[24] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_27 
+ bl[25] br[25] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_28 
+ bl[26] br[26] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_29 
+ bl[27] br[27] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_30 
+ bl[28] br[28] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_31 
+ bl[29] br[29] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_32 
+ bl[30] br[30] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_33 
+ bl[31] br[31] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_34 
+ bl[32] br[32] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_35 
+ bl[33] br[33] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_36 
+ bl[34] br[34] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_37 
+ bl[35] br[35] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_38 
+ bl[36] br[36] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_39 
+ bl[37] br[37] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_40 
+ bl[38] br[38] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_41 
+ bl[39] br[39] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_42 
+ bl[40] br[40] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_43 
+ bl[41] br[41] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_44 
+ bl[42] br[42] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_45 
+ bl[43] br[43] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_46 
+ bl[44] br[44] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_47 
+ bl[45] br[45] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_48 
+ bl[46] br[46] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_49 
+ bl[47] br[47] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_50 
+ bl[48] br[48] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_51 
+ bl[49] br[49] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_52 
+ bl[50] br[50] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_53 
+ bl[51] br[51] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_54 
+ bl[52] br[52] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_55 
+ bl[53] br[53] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_56 
+ bl[54] br[54] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_57 
+ bl[55] br[55] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_58 
+ bl[56] br[56] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_59 
+ bl[57] br[57] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_60 
+ bl[58] br[58] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_61 
+ bl[59] br[59] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_62 
+ bl[60] br[60] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_63 
+ bl[61] br[61] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_64 
+ bl[62] br[62] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_65 
+ bl[63] br[63] vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_66 
+ vdd vdd vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_475_67 
+ vdd vdd vdd vss wl[473] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_0 
+ vdd vdd vss vdd vpb vnb wl[474] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_476_1 
+ rbl rbr vss vdd vpb vnb wl[474] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_476_2 
+ bl[0] br[0] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_3 
+ bl[1] br[1] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_4 
+ bl[2] br[2] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_5 
+ bl[3] br[3] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_6 
+ bl[4] br[4] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_7 
+ bl[5] br[5] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_8 
+ bl[6] br[6] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_9 
+ bl[7] br[7] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_10 
+ bl[8] br[8] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_11 
+ bl[9] br[9] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_12 
+ bl[10] br[10] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_13 
+ bl[11] br[11] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_14 
+ bl[12] br[12] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_15 
+ bl[13] br[13] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_16 
+ bl[14] br[14] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_17 
+ bl[15] br[15] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_18 
+ bl[16] br[16] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_19 
+ bl[17] br[17] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_20 
+ bl[18] br[18] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_21 
+ bl[19] br[19] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_22 
+ bl[20] br[20] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_23 
+ bl[21] br[21] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_24 
+ bl[22] br[22] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_25 
+ bl[23] br[23] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_26 
+ bl[24] br[24] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_27 
+ bl[25] br[25] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_28 
+ bl[26] br[26] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_29 
+ bl[27] br[27] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_30 
+ bl[28] br[28] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_31 
+ bl[29] br[29] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_32 
+ bl[30] br[30] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_33 
+ bl[31] br[31] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_34 
+ bl[32] br[32] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_35 
+ bl[33] br[33] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_36 
+ bl[34] br[34] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_37 
+ bl[35] br[35] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_38 
+ bl[36] br[36] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_39 
+ bl[37] br[37] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_40 
+ bl[38] br[38] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_41 
+ bl[39] br[39] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_42 
+ bl[40] br[40] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_43 
+ bl[41] br[41] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_44 
+ bl[42] br[42] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_45 
+ bl[43] br[43] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_46 
+ bl[44] br[44] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_47 
+ bl[45] br[45] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_48 
+ bl[46] br[46] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_49 
+ bl[47] br[47] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_50 
+ bl[48] br[48] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_51 
+ bl[49] br[49] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_52 
+ bl[50] br[50] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_53 
+ bl[51] br[51] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_54 
+ bl[52] br[52] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_55 
+ bl[53] br[53] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_56 
+ bl[54] br[54] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_57 
+ bl[55] br[55] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_58 
+ bl[56] br[56] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_59 
+ bl[57] br[57] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_60 
+ bl[58] br[58] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_61 
+ bl[59] br[59] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_62 
+ bl[60] br[60] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_63 
+ bl[61] br[61] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_64 
+ bl[62] br[62] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_65 
+ bl[63] br[63] vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_66 
+ vdd vdd vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_476_67 
+ vdd vdd vdd vss wl[474] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_0 
+ vdd vdd vss vdd vpb vnb wl[475] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_477_1 
+ rbl rbr vss vdd vpb vnb wl[475] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_477_2 
+ bl[0] br[0] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_3 
+ bl[1] br[1] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_4 
+ bl[2] br[2] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_5 
+ bl[3] br[3] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_6 
+ bl[4] br[4] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_7 
+ bl[5] br[5] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_8 
+ bl[6] br[6] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_9 
+ bl[7] br[7] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_10 
+ bl[8] br[8] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_11 
+ bl[9] br[9] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_12 
+ bl[10] br[10] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_13 
+ bl[11] br[11] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_14 
+ bl[12] br[12] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_15 
+ bl[13] br[13] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_16 
+ bl[14] br[14] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_17 
+ bl[15] br[15] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_18 
+ bl[16] br[16] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_19 
+ bl[17] br[17] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_20 
+ bl[18] br[18] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_21 
+ bl[19] br[19] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_22 
+ bl[20] br[20] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_23 
+ bl[21] br[21] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_24 
+ bl[22] br[22] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_25 
+ bl[23] br[23] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_26 
+ bl[24] br[24] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_27 
+ bl[25] br[25] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_28 
+ bl[26] br[26] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_29 
+ bl[27] br[27] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_30 
+ bl[28] br[28] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_31 
+ bl[29] br[29] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_32 
+ bl[30] br[30] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_33 
+ bl[31] br[31] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_34 
+ bl[32] br[32] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_35 
+ bl[33] br[33] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_36 
+ bl[34] br[34] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_37 
+ bl[35] br[35] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_38 
+ bl[36] br[36] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_39 
+ bl[37] br[37] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_40 
+ bl[38] br[38] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_41 
+ bl[39] br[39] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_42 
+ bl[40] br[40] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_43 
+ bl[41] br[41] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_44 
+ bl[42] br[42] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_45 
+ bl[43] br[43] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_46 
+ bl[44] br[44] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_47 
+ bl[45] br[45] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_48 
+ bl[46] br[46] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_49 
+ bl[47] br[47] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_50 
+ bl[48] br[48] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_51 
+ bl[49] br[49] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_52 
+ bl[50] br[50] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_53 
+ bl[51] br[51] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_54 
+ bl[52] br[52] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_55 
+ bl[53] br[53] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_56 
+ bl[54] br[54] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_57 
+ bl[55] br[55] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_58 
+ bl[56] br[56] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_59 
+ bl[57] br[57] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_60 
+ bl[58] br[58] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_61 
+ bl[59] br[59] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_62 
+ bl[60] br[60] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_63 
+ bl[61] br[61] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_64 
+ bl[62] br[62] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_65 
+ bl[63] br[63] vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_66 
+ vdd vdd vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_477_67 
+ vdd vdd vdd vss wl[475] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_0 
+ vdd vdd vss vdd vpb vnb wl[476] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_478_1 
+ rbl rbr vss vdd vpb vnb wl[476] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_478_2 
+ bl[0] br[0] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_3 
+ bl[1] br[1] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_4 
+ bl[2] br[2] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_5 
+ bl[3] br[3] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_6 
+ bl[4] br[4] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_7 
+ bl[5] br[5] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_8 
+ bl[6] br[6] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_9 
+ bl[7] br[7] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_10 
+ bl[8] br[8] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_11 
+ bl[9] br[9] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_12 
+ bl[10] br[10] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_13 
+ bl[11] br[11] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_14 
+ bl[12] br[12] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_15 
+ bl[13] br[13] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_16 
+ bl[14] br[14] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_17 
+ bl[15] br[15] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_18 
+ bl[16] br[16] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_19 
+ bl[17] br[17] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_20 
+ bl[18] br[18] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_21 
+ bl[19] br[19] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_22 
+ bl[20] br[20] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_23 
+ bl[21] br[21] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_24 
+ bl[22] br[22] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_25 
+ bl[23] br[23] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_26 
+ bl[24] br[24] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_27 
+ bl[25] br[25] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_28 
+ bl[26] br[26] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_29 
+ bl[27] br[27] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_30 
+ bl[28] br[28] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_31 
+ bl[29] br[29] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_32 
+ bl[30] br[30] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_33 
+ bl[31] br[31] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_34 
+ bl[32] br[32] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_35 
+ bl[33] br[33] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_36 
+ bl[34] br[34] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_37 
+ bl[35] br[35] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_38 
+ bl[36] br[36] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_39 
+ bl[37] br[37] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_40 
+ bl[38] br[38] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_41 
+ bl[39] br[39] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_42 
+ bl[40] br[40] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_43 
+ bl[41] br[41] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_44 
+ bl[42] br[42] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_45 
+ bl[43] br[43] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_46 
+ bl[44] br[44] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_47 
+ bl[45] br[45] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_48 
+ bl[46] br[46] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_49 
+ bl[47] br[47] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_50 
+ bl[48] br[48] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_51 
+ bl[49] br[49] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_52 
+ bl[50] br[50] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_53 
+ bl[51] br[51] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_54 
+ bl[52] br[52] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_55 
+ bl[53] br[53] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_56 
+ bl[54] br[54] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_57 
+ bl[55] br[55] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_58 
+ bl[56] br[56] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_59 
+ bl[57] br[57] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_60 
+ bl[58] br[58] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_61 
+ bl[59] br[59] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_62 
+ bl[60] br[60] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_63 
+ bl[61] br[61] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_64 
+ bl[62] br[62] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_65 
+ bl[63] br[63] vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_66 
+ vdd vdd vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_478_67 
+ vdd vdd vdd vss wl[476] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_0 
+ vdd vdd vss vdd vpb vnb wl[477] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_479_1 
+ rbl rbr vss vdd vpb vnb wl[477] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_479_2 
+ bl[0] br[0] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_3 
+ bl[1] br[1] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_4 
+ bl[2] br[2] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_5 
+ bl[3] br[3] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_6 
+ bl[4] br[4] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_7 
+ bl[5] br[5] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_8 
+ bl[6] br[6] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_9 
+ bl[7] br[7] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_10 
+ bl[8] br[8] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_11 
+ bl[9] br[9] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_12 
+ bl[10] br[10] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_13 
+ bl[11] br[11] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_14 
+ bl[12] br[12] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_15 
+ bl[13] br[13] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_16 
+ bl[14] br[14] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_17 
+ bl[15] br[15] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_18 
+ bl[16] br[16] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_19 
+ bl[17] br[17] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_20 
+ bl[18] br[18] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_21 
+ bl[19] br[19] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_22 
+ bl[20] br[20] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_23 
+ bl[21] br[21] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_24 
+ bl[22] br[22] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_25 
+ bl[23] br[23] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_26 
+ bl[24] br[24] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_27 
+ bl[25] br[25] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_28 
+ bl[26] br[26] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_29 
+ bl[27] br[27] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_30 
+ bl[28] br[28] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_31 
+ bl[29] br[29] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_32 
+ bl[30] br[30] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_33 
+ bl[31] br[31] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_34 
+ bl[32] br[32] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_35 
+ bl[33] br[33] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_36 
+ bl[34] br[34] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_37 
+ bl[35] br[35] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_38 
+ bl[36] br[36] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_39 
+ bl[37] br[37] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_40 
+ bl[38] br[38] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_41 
+ bl[39] br[39] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_42 
+ bl[40] br[40] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_43 
+ bl[41] br[41] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_44 
+ bl[42] br[42] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_45 
+ bl[43] br[43] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_46 
+ bl[44] br[44] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_47 
+ bl[45] br[45] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_48 
+ bl[46] br[46] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_49 
+ bl[47] br[47] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_50 
+ bl[48] br[48] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_51 
+ bl[49] br[49] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_52 
+ bl[50] br[50] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_53 
+ bl[51] br[51] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_54 
+ bl[52] br[52] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_55 
+ bl[53] br[53] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_56 
+ bl[54] br[54] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_57 
+ bl[55] br[55] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_58 
+ bl[56] br[56] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_59 
+ bl[57] br[57] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_60 
+ bl[58] br[58] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_61 
+ bl[59] br[59] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_62 
+ bl[60] br[60] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_63 
+ bl[61] br[61] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_64 
+ bl[62] br[62] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_65 
+ bl[63] br[63] vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_66 
+ vdd vdd vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_479_67 
+ vdd vdd vdd vss wl[477] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_0 
+ vdd vdd vss vdd vpb vnb wl[478] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_480_1 
+ rbl rbr vss vdd vpb vnb wl[478] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_480_2 
+ bl[0] br[0] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_3 
+ bl[1] br[1] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_4 
+ bl[2] br[2] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_5 
+ bl[3] br[3] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_6 
+ bl[4] br[4] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_7 
+ bl[5] br[5] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_8 
+ bl[6] br[6] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_9 
+ bl[7] br[7] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_10 
+ bl[8] br[8] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_11 
+ bl[9] br[9] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_12 
+ bl[10] br[10] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_13 
+ bl[11] br[11] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_14 
+ bl[12] br[12] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_15 
+ bl[13] br[13] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_16 
+ bl[14] br[14] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_17 
+ bl[15] br[15] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_18 
+ bl[16] br[16] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_19 
+ bl[17] br[17] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_20 
+ bl[18] br[18] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_21 
+ bl[19] br[19] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_22 
+ bl[20] br[20] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_23 
+ bl[21] br[21] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_24 
+ bl[22] br[22] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_25 
+ bl[23] br[23] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_26 
+ bl[24] br[24] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_27 
+ bl[25] br[25] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_28 
+ bl[26] br[26] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_29 
+ bl[27] br[27] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_30 
+ bl[28] br[28] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_31 
+ bl[29] br[29] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_32 
+ bl[30] br[30] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_33 
+ bl[31] br[31] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_34 
+ bl[32] br[32] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_35 
+ bl[33] br[33] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_36 
+ bl[34] br[34] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_37 
+ bl[35] br[35] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_38 
+ bl[36] br[36] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_39 
+ bl[37] br[37] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_40 
+ bl[38] br[38] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_41 
+ bl[39] br[39] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_42 
+ bl[40] br[40] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_43 
+ bl[41] br[41] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_44 
+ bl[42] br[42] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_45 
+ bl[43] br[43] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_46 
+ bl[44] br[44] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_47 
+ bl[45] br[45] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_48 
+ bl[46] br[46] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_49 
+ bl[47] br[47] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_50 
+ bl[48] br[48] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_51 
+ bl[49] br[49] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_52 
+ bl[50] br[50] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_53 
+ bl[51] br[51] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_54 
+ bl[52] br[52] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_55 
+ bl[53] br[53] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_56 
+ bl[54] br[54] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_57 
+ bl[55] br[55] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_58 
+ bl[56] br[56] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_59 
+ bl[57] br[57] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_60 
+ bl[58] br[58] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_61 
+ bl[59] br[59] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_62 
+ bl[60] br[60] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_63 
+ bl[61] br[61] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_64 
+ bl[62] br[62] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_65 
+ bl[63] br[63] vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_66 
+ vdd vdd vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_480_67 
+ vdd vdd vdd vss wl[478] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_0 
+ vdd vdd vss vdd vpb vnb wl[479] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_481_1 
+ rbl rbr vss vdd vpb vnb wl[479] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_481_2 
+ bl[0] br[0] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_3 
+ bl[1] br[1] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_4 
+ bl[2] br[2] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_5 
+ bl[3] br[3] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_6 
+ bl[4] br[4] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_7 
+ bl[5] br[5] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_8 
+ bl[6] br[6] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_9 
+ bl[7] br[7] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_10 
+ bl[8] br[8] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_11 
+ bl[9] br[9] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_12 
+ bl[10] br[10] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_13 
+ bl[11] br[11] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_14 
+ bl[12] br[12] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_15 
+ bl[13] br[13] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_16 
+ bl[14] br[14] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_17 
+ bl[15] br[15] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_18 
+ bl[16] br[16] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_19 
+ bl[17] br[17] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_20 
+ bl[18] br[18] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_21 
+ bl[19] br[19] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_22 
+ bl[20] br[20] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_23 
+ bl[21] br[21] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_24 
+ bl[22] br[22] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_25 
+ bl[23] br[23] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_26 
+ bl[24] br[24] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_27 
+ bl[25] br[25] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_28 
+ bl[26] br[26] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_29 
+ bl[27] br[27] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_30 
+ bl[28] br[28] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_31 
+ bl[29] br[29] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_32 
+ bl[30] br[30] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_33 
+ bl[31] br[31] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_34 
+ bl[32] br[32] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_35 
+ bl[33] br[33] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_36 
+ bl[34] br[34] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_37 
+ bl[35] br[35] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_38 
+ bl[36] br[36] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_39 
+ bl[37] br[37] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_40 
+ bl[38] br[38] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_41 
+ bl[39] br[39] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_42 
+ bl[40] br[40] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_43 
+ bl[41] br[41] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_44 
+ bl[42] br[42] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_45 
+ bl[43] br[43] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_46 
+ bl[44] br[44] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_47 
+ bl[45] br[45] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_48 
+ bl[46] br[46] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_49 
+ bl[47] br[47] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_50 
+ bl[48] br[48] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_51 
+ bl[49] br[49] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_52 
+ bl[50] br[50] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_53 
+ bl[51] br[51] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_54 
+ bl[52] br[52] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_55 
+ bl[53] br[53] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_56 
+ bl[54] br[54] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_57 
+ bl[55] br[55] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_58 
+ bl[56] br[56] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_59 
+ bl[57] br[57] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_60 
+ bl[58] br[58] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_61 
+ bl[59] br[59] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_62 
+ bl[60] br[60] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_63 
+ bl[61] br[61] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_64 
+ bl[62] br[62] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_65 
+ bl[63] br[63] vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_66 
+ vdd vdd vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_481_67 
+ vdd vdd vdd vss wl[479] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_0 
+ vdd vdd vss vdd vpb vnb wl[480] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_482_1 
+ rbl rbr vss vdd vpb vnb wl[480] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_482_2 
+ bl[0] br[0] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_3 
+ bl[1] br[1] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_4 
+ bl[2] br[2] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_5 
+ bl[3] br[3] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_6 
+ bl[4] br[4] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_7 
+ bl[5] br[5] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_8 
+ bl[6] br[6] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_9 
+ bl[7] br[7] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_10 
+ bl[8] br[8] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_11 
+ bl[9] br[9] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_12 
+ bl[10] br[10] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_13 
+ bl[11] br[11] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_14 
+ bl[12] br[12] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_15 
+ bl[13] br[13] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_16 
+ bl[14] br[14] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_17 
+ bl[15] br[15] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_18 
+ bl[16] br[16] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_19 
+ bl[17] br[17] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_20 
+ bl[18] br[18] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_21 
+ bl[19] br[19] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_22 
+ bl[20] br[20] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_23 
+ bl[21] br[21] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_24 
+ bl[22] br[22] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_25 
+ bl[23] br[23] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_26 
+ bl[24] br[24] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_27 
+ bl[25] br[25] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_28 
+ bl[26] br[26] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_29 
+ bl[27] br[27] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_30 
+ bl[28] br[28] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_31 
+ bl[29] br[29] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_32 
+ bl[30] br[30] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_33 
+ bl[31] br[31] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_34 
+ bl[32] br[32] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_35 
+ bl[33] br[33] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_36 
+ bl[34] br[34] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_37 
+ bl[35] br[35] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_38 
+ bl[36] br[36] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_39 
+ bl[37] br[37] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_40 
+ bl[38] br[38] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_41 
+ bl[39] br[39] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_42 
+ bl[40] br[40] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_43 
+ bl[41] br[41] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_44 
+ bl[42] br[42] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_45 
+ bl[43] br[43] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_46 
+ bl[44] br[44] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_47 
+ bl[45] br[45] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_48 
+ bl[46] br[46] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_49 
+ bl[47] br[47] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_50 
+ bl[48] br[48] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_51 
+ bl[49] br[49] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_52 
+ bl[50] br[50] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_53 
+ bl[51] br[51] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_54 
+ bl[52] br[52] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_55 
+ bl[53] br[53] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_56 
+ bl[54] br[54] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_57 
+ bl[55] br[55] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_58 
+ bl[56] br[56] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_59 
+ bl[57] br[57] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_60 
+ bl[58] br[58] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_61 
+ bl[59] br[59] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_62 
+ bl[60] br[60] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_63 
+ bl[61] br[61] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_64 
+ bl[62] br[62] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_65 
+ bl[63] br[63] vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_66 
+ vdd vdd vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_482_67 
+ vdd vdd vdd vss wl[480] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_0 
+ vdd vdd vss vdd vpb vnb wl[481] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_483_1 
+ rbl rbr vss vdd vpb vnb wl[481] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_483_2 
+ bl[0] br[0] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_3 
+ bl[1] br[1] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_4 
+ bl[2] br[2] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_5 
+ bl[3] br[3] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_6 
+ bl[4] br[4] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_7 
+ bl[5] br[5] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_8 
+ bl[6] br[6] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_9 
+ bl[7] br[7] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_10 
+ bl[8] br[8] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_11 
+ bl[9] br[9] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_12 
+ bl[10] br[10] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_13 
+ bl[11] br[11] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_14 
+ bl[12] br[12] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_15 
+ bl[13] br[13] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_16 
+ bl[14] br[14] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_17 
+ bl[15] br[15] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_18 
+ bl[16] br[16] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_19 
+ bl[17] br[17] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_20 
+ bl[18] br[18] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_21 
+ bl[19] br[19] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_22 
+ bl[20] br[20] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_23 
+ bl[21] br[21] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_24 
+ bl[22] br[22] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_25 
+ bl[23] br[23] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_26 
+ bl[24] br[24] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_27 
+ bl[25] br[25] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_28 
+ bl[26] br[26] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_29 
+ bl[27] br[27] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_30 
+ bl[28] br[28] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_31 
+ bl[29] br[29] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_32 
+ bl[30] br[30] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_33 
+ bl[31] br[31] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_34 
+ bl[32] br[32] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_35 
+ bl[33] br[33] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_36 
+ bl[34] br[34] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_37 
+ bl[35] br[35] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_38 
+ bl[36] br[36] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_39 
+ bl[37] br[37] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_40 
+ bl[38] br[38] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_41 
+ bl[39] br[39] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_42 
+ bl[40] br[40] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_43 
+ bl[41] br[41] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_44 
+ bl[42] br[42] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_45 
+ bl[43] br[43] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_46 
+ bl[44] br[44] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_47 
+ bl[45] br[45] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_48 
+ bl[46] br[46] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_49 
+ bl[47] br[47] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_50 
+ bl[48] br[48] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_51 
+ bl[49] br[49] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_52 
+ bl[50] br[50] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_53 
+ bl[51] br[51] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_54 
+ bl[52] br[52] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_55 
+ bl[53] br[53] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_56 
+ bl[54] br[54] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_57 
+ bl[55] br[55] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_58 
+ bl[56] br[56] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_59 
+ bl[57] br[57] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_60 
+ bl[58] br[58] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_61 
+ bl[59] br[59] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_62 
+ bl[60] br[60] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_63 
+ bl[61] br[61] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_64 
+ bl[62] br[62] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_65 
+ bl[63] br[63] vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_66 
+ vdd vdd vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_483_67 
+ vdd vdd vdd vss wl[481] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_0 
+ vdd vdd vss vdd vpb vnb wl[482] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_484_1 
+ rbl rbr vss vdd vpb vnb wl[482] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_484_2 
+ bl[0] br[0] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_3 
+ bl[1] br[1] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_4 
+ bl[2] br[2] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_5 
+ bl[3] br[3] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_6 
+ bl[4] br[4] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_7 
+ bl[5] br[5] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_8 
+ bl[6] br[6] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_9 
+ bl[7] br[7] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_10 
+ bl[8] br[8] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_11 
+ bl[9] br[9] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_12 
+ bl[10] br[10] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_13 
+ bl[11] br[11] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_14 
+ bl[12] br[12] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_15 
+ bl[13] br[13] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_16 
+ bl[14] br[14] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_17 
+ bl[15] br[15] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_18 
+ bl[16] br[16] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_19 
+ bl[17] br[17] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_20 
+ bl[18] br[18] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_21 
+ bl[19] br[19] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_22 
+ bl[20] br[20] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_23 
+ bl[21] br[21] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_24 
+ bl[22] br[22] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_25 
+ bl[23] br[23] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_26 
+ bl[24] br[24] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_27 
+ bl[25] br[25] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_28 
+ bl[26] br[26] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_29 
+ bl[27] br[27] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_30 
+ bl[28] br[28] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_31 
+ bl[29] br[29] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_32 
+ bl[30] br[30] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_33 
+ bl[31] br[31] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_34 
+ bl[32] br[32] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_35 
+ bl[33] br[33] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_36 
+ bl[34] br[34] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_37 
+ bl[35] br[35] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_38 
+ bl[36] br[36] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_39 
+ bl[37] br[37] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_40 
+ bl[38] br[38] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_41 
+ bl[39] br[39] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_42 
+ bl[40] br[40] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_43 
+ bl[41] br[41] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_44 
+ bl[42] br[42] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_45 
+ bl[43] br[43] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_46 
+ bl[44] br[44] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_47 
+ bl[45] br[45] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_48 
+ bl[46] br[46] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_49 
+ bl[47] br[47] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_50 
+ bl[48] br[48] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_51 
+ bl[49] br[49] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_52 
+ bl[50] br[50] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_53 
+ bl[51] br[51] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_54 
+ bl[52] br[52] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_55 
+ bl[53] br[53] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_56 
+ bl[54] br[54] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_57 
+ bl[55] br[55] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_58 
+ bl[56] br[56] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_59 
+ bl[57] br[57] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_60 
+ bl[58] br[58] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_61 
+ bl[59] br[59] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_62 
+ bl[60] br[60] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_63 
+ bl[61] br[61] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_64 
+ bl[62] br[62] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_65 
+ bl[63] br[63] vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_66 
+ vdd vdd vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_484_67 
+ vdd vdd vdd vss wl[482] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_0 
+ vdd vdd vss vdd vpb vnb wl[483] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_485_1 
+ rbl rbr vss vdd vpb vnb wl[483] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_485_2 
+ bl[0] br[0] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_3 
+ bl[1] br[1] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_4 
+ bl[2] br[2] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_5 
+ bl[3] br[3] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_6 
+ bl[4] br[4] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_7 
+ bl[5] br[5] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_8 
+ bl[6] br[6] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_9 
+ bl[7] br[7] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_10 
+ bl[8] br[8] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_11 
+ bl[9] br[9] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_12 
+ bl[10] br[10] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_13 
+ bl[11] br[11] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_14 
+ bl[12] br[12] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_15 
+ bl[13] br[13] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_16 
+ bl[14] br[14] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_17 
+ bl[15] br[15] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_18 
+ bl[16] br[16] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_19 
+ bl[17] br[17] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_20 
+ bl[18] br[18] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_21 
+ bl[19] br[19] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_22 
+ bl[20] br[20] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_23 
+ bl[21] br[21] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_24 
+ bl[22] br[22] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_25 
+ bl[23] br[23] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_26 
+ bl[24] br[24] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_27 
+ bl[25] br[25] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_28 
+ bl[26] br[26] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_29 
+ bl[27] br[27] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_30 
+ bl[28] br[28] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_31 
+ bl[29] br[29] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_32 
+ bl[30] br[30] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_33 
+ bl[31] br[31] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_34 
+ bl[32] br[32] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_35 
+ bl[33] br[33] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_36 
+ bl[34] br[34] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_37 
+ bl[35] br[35] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_38 
+ bl[36] br[36] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_39 
+ bl[37] br[37] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_40 
+ bl[38] br[38] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_41 
+ bl[39] br[39] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_42 
+ bl[40] br[40] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_43 
+ bl[41] br[41] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_44 
+ bl[42] br[42] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_45 
+ bl[43] br[43] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_46 
+ bl[44] br[44] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_47 
+ bl[45] br[45] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_48 
+ bl[46] br[46] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_49 
+ bl[47] br[47] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_50 
+ bl[48] br[48] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_51 
+ bl[49] br[49] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_52 
+ bl[50] br[50] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_53 
+ bl[51] br[51] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_54 
+ bl[52] br[52] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_55 
+ bl[53] br[53] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_56 
+ bl[54] br[54] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_57 
+ bl[55] br[55] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_58 
+ bl[56] br[56] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_59 
+ bl[57] br[57] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_60 
+ bl[58] br[58] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_61 
+ bl[59] br[59] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_62 
+ bl[60] br[60] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_63 
+ bl[61] br[61] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_64 
+ bl[62] br[62] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_65 
+ bl[63] br[63] vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_66 
+ vdd vdd vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_485_67 
+ vdd vdd vdd vss wl[483] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_0 
+ vdd vdd vss vdd vpb vnb wl[484] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_486_1 
+ rbl rbr vss vdd vpb vnb wl[484] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_486_2 
+ bl[0] br[0] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_3 
+ bl[1] br[1] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_4 
+ bl[2] br[2] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_5 
+ bl[3] br[3] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_6 
+ bl[4] br[4] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_7 
+ bl[5] br[5] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_8 
+ bl[6] br[6] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_9 
+ bl[7] br[7] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_10 
+ bl[8] br[8] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_11 
+ bl[9] br[9] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_12 
+ bl[10] br[10] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_13 
+ bl[11] br[11] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_14 
+ bl[12] br[12] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_15 
+ bl[13] br[13] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_16 
+ bl[14] br[14] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_17 
+ bl[15] br[15] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_18 
+ bl[16] br[16] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_19 
+ bl[17] br[17] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_20 
+ bl[18] br[18] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_21 
+ bl[19] br[19] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_22 
+ bl[20] br[20] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_23 
+ bl[21] br[21] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_24 
+ bl[22] br[22] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_25 
+ bl[23] br[23] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_26 
+ bl[24] br[24] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_27 
+ bl[25] br[25] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_28 
+ bl[26] br[26] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_29 
+ bl[27] br[27] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_30 
+ bl[28] br[28] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_31 
+ bl[29] br[29] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_32 
+ bl[30] br[30] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_33 
+ bl[31] br[31] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_34 
+ bl[32] br[32] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_35 
+ bl[33] br[33] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_36 
+ bl[34] br[34] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_37 
+ bl[35] br[35] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_38 
+ bl[36] br[36] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_39 
+ bl[37] br[37] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_40 
+ bl[38] br[38] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_41 
+ bl[39] br[39] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_42 
+ bl[40] br[40] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_43 
+ bl[41] br[41] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_44 
+ bl[42] br[42] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_45 
+ bl[43] br[43] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_46 
+ bl[44] br[44] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_47 
+ bl[45] br[45] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_48 
+ bl[46] br[46] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_49 
+ bl[47] br[47] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_50 
+ bl[48] br[48] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_51 
+ bl[49] br[49] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_52 
+ bl[50] br[50] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_53 
+ bl[51] br[51] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_54 
+ bl[52] br[52] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_55 
+ bl[53] br[53] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_56 
+ bl[54] br[54] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_57 
+ bl[55] br[55] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_58 
+ bl[56] br[56] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_59 
+ bl[57] br[57] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_60 
+ bl[58] br[58] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_61 
+ bl[59] br[59] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_62 
+ bl[60] br[60] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_63 
+ bl[61] br[61] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_64 
+ bl[62] br[62] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_65 
+ bl[63] br[63] vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_66 
+ vdd vdd vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_486_67 
+ vdd vdd vdd vss wl[484] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_0 
+ vdd vdd vss vdd vpb vnb wl[485] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_487_1 
+ rbl rbr vss vdd vpb vnb wl[485] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_487_2 
+ bl[0] br[0] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_3 
+ bl[1] br[1] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_4 
+ bl[2] br[2] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_5 
+ bl[3] br[3] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_6 
+ bl[4] br[4] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_7 
+ bl[5] br[5] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_8 
+ bl[6] br[6] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_9 
+ bl[7] br[7] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_10 
+ bl[8] br[8] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_11 
+ bl[9] br[9] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_12 
+ bl[10] br[10] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_13 
+ bl[11] br[11] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_14 
+ bl[12] br[12] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_15 
+ bl[13] br[13] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_16 
+ bl[14] br[14] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_17 
+ bl[15] br[15] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_18 
+ bl[16] br[16] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_19 
+ bl[17] br[17] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_20 
+ bl[18] br[18] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_21 
+ bl[19] br[19] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_22 
+ bl[20] br[20] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_23 
+ bl[21] br[21] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_24 
+ bl[22] br[22] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_25 
+ bl[23] br[23] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_26 
+ bl[24] br[24] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_27 
+ bl[25] br[25] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_28 
+ bl[26] br[26] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_29 
+ bl[27] br[27] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_30 
+ bl[28] br[28] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_31 
+ bl[29] br[29] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_32 
+ bl[30] br[30] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_33 
+ bl[31] br[31] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_34 
+ bl[32] br[32] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_35 
+ bl[33] br[33] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_36 
+ bl[34] br[34] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_37 
+ bl[35] br[35] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_38 
+ bl[36] br[36] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_39 
+ bl[37] br[37] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_40 
+ bl[38] br[38] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_41 
+ bl[39] br[39] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_42 
+ bl[40] br[40] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_43 
+ bl[41] br[41] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_44 
+ bl[42] br[42] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_45 
+ bl[43] br[43] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_46 
+ bl[44] br[44] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_47 
+ bl[45] br[45] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_48 
+ bl[46] br[46] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_49 
+ bl[47] br[47] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_50 
+ bl[48] br[48] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_51 
+ bl[49] br[49] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_52 
+ bl[50] br[50] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_53 
+ bl[51] br[51] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_54 
+ bl[52] br[52] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_55 
+ bl[53] br[53] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_56 
+ bl[54] br[54] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_57 
+ bl[55] br[55] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_58 
+ bl[56] br[56] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_59 
+ bl[57] br[57] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_60 
+ bl[58] br[58] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_61 
+ bl[59] br[59] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_62 
+ bl[60] br[60] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_63 
+ bl[61] br[61] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_64 
+ bl[62] br[62] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_65 
+ bl[63] br[63] vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_66 
+ vdd vdd vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_487_67 
+ vdd vdd vdd vss wl[485] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_0 
+ vdd vdd vss vdd vpb vnb wl[486] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_488_1 
+ rbl rbr vss vdd vpb vnb wl[486] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_488_2 
+ bl[0] br[0] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_3 
+ bl[1] br[1] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_4 
+ bl[2] br[2] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_5 
+ bl[3] br[3] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_6 
+ bl[4] br[4] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_7 
+ bl[5] br[5] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_8 
+ bl[6] br[6] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_9 
+ bl[7] br[7] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_10 
+ bl[8] br[8] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_11 
+ bl[9] br[9] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_12 
+ bl[10] br[10] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_13 
+ bl[11] br[11] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_14 
+ bl[12] br[12] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_15 
+ bl[13] br[13] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_16 
+ bl[14] br[14] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_17 
+ bl[15] br[15] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_18 
+ bl[16] br[16] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_19 
+ bl[17] br[17] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_20 
+ bl[18] br[18] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_21 
+ bl[19] br[19] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_22 
+ bl[20] br[20] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_23 
+ bl[21] br[21] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_24 
+ bl[22] br[22] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_25 
+ bl[23] br[23] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_26 
+ bl[24] br[24] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_27 
+ bl[25] br[25] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_28 
+ bl[26] br[26] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_29 
+ bl[27] br[27] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_30 
+ bl[28] br[28] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_31 
+ bl[29] br[29] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_32 
+ bl[30] br[30] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_33 
+ bl[31] br[31] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_34 
+ bl[32] br[32] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_35 
+ bl[33] br[33] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_36 
+ bl[34] br[34] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_37 
+ bl[35] br[35] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_38 
+ bl[36] br[36] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_39 
+ bl[37] br[37] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_40 
+ bl[38] br[38] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_41 
+ bl[39] br[39] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_42 
+ bl[40] br[40] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_43 
+ bl[41] br[41] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_44 
+ bl[42] br[42] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_45 
+ bl[43] br[43] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_46 
+ bl[44] br[44] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_47 
+ bl[45] br[45] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_48 
+ bl[46] br[46] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_49 
+ bl[47] br[47] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_50 
+ bl[48] br[48] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_51 
+ bl[49] br[49] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_52 
+ bl[50] br[50] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_53 
+ bl[51] br[51] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_54 
+ bl[52] br[52] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_55 
+ bl[53] br[53] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_56 
+ bl[54] br[54] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_57 
+ bl[55] br[55] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_58 
+ bl[56] br[56] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_59 
+ bl[57] br[57] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_60 
+ bl[58] br[58] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_61 
+ bl[59] br[59] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_62 
+ bl[60] br[60] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_63 
+ bl[61] br[61] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_64 
+ bl[62] br[62] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_65 
+ bl[63] br[63] vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_66 
+ vdd vdd vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_488_67 
+ vdd vdd vdd vss wl[486] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_0 
+ vdd vdd vss vdd vpb vnb wl[487] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_489_1 
+ rbl rbr vss vdd vpb vnb wl[487] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_489_2 
+ bl[0] br[0] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_3 
+ bl[1] br[1] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_4 
+ bl[2] br[2] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_5 
+ bl[3] br[3] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_6 
+ bl[4] br[4] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_7 
+ bl[5] br[5] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_8 
+ bl[6] br[6] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_9 
+ bl[7] br[7] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_10 
+ bl[8] br[8] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_11 
+ bl[9] br[9] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_12 
+ bl[10] br[10] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_13 
+ bl[11] br[11] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_14 
+ bl[12] br[12] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_15 
+ bl[13] br[13] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_16 
+ bl[14] br[14] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_17 
+ bl[15] br[15] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_18 
+ bl[16] br[16] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_19 
+ bl[17] br[17] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_20 
+ bl[18] br[18] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_21 
+ bl[19] br[19] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_22 
+ bl[20] br[20] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_23 
+ bl[21] br[21] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_24 
+ bl[22] br[22] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_25 
+ bl[23] br[23] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_26 
+ bl[24] br[24] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_27 
+ bl[25] br[25] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_28 
+ bl[26] br[26] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_29 
+ bl[27] br[27] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_30 
+ bl[28] br[28] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_31 
+ bl[29] br[29] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_32 
+ bl[30] br[30] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_33 
+ bl[31] br[31] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_34 
+ bl[32] br[32] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_35 
+ bl[33] br[33] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_36 
+ bl[34] br[34] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_37 
+ bl[35] br[35] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_38 
+ bl[36] br[36] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_39 
+ bl[37] br[37] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_40 
+ bl[38] br[38] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_41 
+ bl[39] br[39] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_42 
+ bl[40] br[40] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_43 
+ bl[41] br[41] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_44 
+ bl[42] br[42] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_45 
+ bl[43] br[43] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_46 
+ bl[44] br[44] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_47 
+ bl[45] br[45] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_48 
+ bl[46] br[46] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_49 
+ bl[47] br[47] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_50 
+ bl[48] br[48] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_51 
+ bl[49] br[49] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_52 
+ bl[50] br[50] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_53 
+ bl[51] br[51] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_54 
+ bl[52] br[52] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_55 
+ bl[53] br[53] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_56 
+ bl[54] br[54] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_57 
+ bl[55] br[55] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_58 
+ bl[56] br[56] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_59 
+ bl[57] br[57] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_60 
+ bl[58] br[58] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_61 
+ bl[59] br[59] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_62 
+ bl[60] br[60] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_63 
+ bl[61] br[61] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_64 
+ bl[62] br[62] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_65 
+ bl[63] br[63] vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_66 
+ vdd vdd vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_489_67 
+ vdd vdd vdd vss wl[487] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_0 
+ vdd vdd vss vdd vpb vnb wl[488] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_490_1 
+ rbl rbr vss vdd vpb vnb wl[488] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_490_2 
+ bl[0] br[0] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_3 
+ bl[1] br[1] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_4 
+ bl[2] br[2] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_5 
+ bl[3] br[3] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_6 
+ bl[4] br[4] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_7 
+ bl[5] br[5] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_8 
+ bl[6] br[6] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_9 
+ bl[7] br[7] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_10 
+ bl[8] br[8] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_11 
+ bl[9] br[9] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_12 
+ bl[10] br[10] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_13 
+ bl[11] br[11] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_14 
+ bl[12] br[12] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_15 
+ bl[13] br[13] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_16 
+ bl[14] br[14] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_17 
+ bl[15] br[15] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_18 
+ bl[16] br[16] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_19 
+ bl[17] br[17] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_20 
+ bl[18] br[18] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_21 
+ bl[19] br[19] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_22 
+ bl[20] br[20] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_23 
+ bl[21] br[21] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_24 
+ bl[22] br[22] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_25 
+ bl[23] br[23] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_26 
+ bl[24] br[24] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_27 
+ bl[25] br[25] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_28 
+ bl[26] br[26] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_29 
+ bl[27] br[27] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_30 
+ bl[28] br[28] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_31 
+ bl[29] br[29] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_32 
+ bl[30] br[30] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_33 
+ bl[31] br[31] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_34 
+ bl[32] br[32] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_35 
+ bl[33] br[33] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_36 
+ bl[34] br[34] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_37 
+ bl[35] br[35] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_38 
+ bl[36] br[36] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_39 
+ bl[37] br[37] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_40 
+ bl[38] br[38] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_41 
+ bl[39] br[39] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_42 
+ bl[40] br[40] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_43 
+ bl[41] br[41] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_44 
+ bl[42] br[42] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_45 
+ bl[43] br[43] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_46 
+ bl[44] br[44] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_47 
+ bl[45] br[45] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_48 
+ bl[46] br[46] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_49 
+ bl[47] br[47] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_50 
+ bl[48] br[48] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_51 
+ bl[49] br[49] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_52 
+ bl[50] br[50] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_53 
+ bl[51] br[51] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_54 
+ bl[52] br[52] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_55 
+ bl[53] br[53] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_56 
+ bl[54] br[54] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_57 
+ bl[55] br[55] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_58 
+ bl[56] br[56] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_59 
+ bl[57] br[57] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_60 
+ bl[58] br[58] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_61 
+ bl[59] br[59] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_62 
+ bl[60] br[60] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_63 
+ bl[61] br[61] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_64 
+ bl[62] br[62] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_65 
+ bl[63] br[63] vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_66 
+ vdd vdd vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_490_67 
+ vdd vdd vdd vss wl[488] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_0 
+ vdd vdd vss vdd vpb vnb wl[489] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_491_1 
+ rbl rbr vss vdd vpb vnb wl[489] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_491_2 
+ bl[0] br[0] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_3 
+ bl[1] br[1] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_4 
+ bl[2] br[2] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_5 
+ bl[3] br[3] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_6 
+ bl[4] br[4] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_7 
+ bl[5] br[5] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_8 
+ bl[6] br[6] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_9 
+ bl[7] br[7] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_10 
+ bl[8] br[8] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_11 
+ bl[9] br[9] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_12 
+ bl[10] br[10] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_13 
+ bl[11] br[11] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_14 
+ bl[12] br[12] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_15 
+ bl[13] br[13] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_16 
+ bl[14] br[14] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_17 
+ bl[15] br[15] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_18 
+ bl[16] br[16] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_19 
+ bl[17] br[17] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_20 
+ bl[18] br[18] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_21 
+ bl[19] br[19] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_22 
+ bl[20] br[20] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_23 
+ bl[21] br[21] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_24 
+ bl[22] br[22] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_25 
+ bl[23] br[23] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_26 
+ bl[24] br[24] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_27 
+ bl[25] br[25] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_28 
+ bl[26] br[26] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_29 
+ bl[27] br[27] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_30 
+ bl[28] br[28] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_31 
+ bl[29] br[29] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_32 
+ bl[30] br[30] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_33 
+ bl[31] br[31] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_34 
+ bl[32] br[32] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_35 
+ bl[33] br[33] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_36 
+ bl[34] br[34] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_37 
+ bl[35] br[35] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_38 
+ bl[36] br[36] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_39 
+ bl[37] br[37] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_40 
+ bl[38] br[38] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_41 
+ bl[39] br[39] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_42 
+ bl[40] br[40] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_43 
+ bl[41] br[41] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_44 
+ bl[42] br[42] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_45 
+ bl[43] br[43] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_46 
+ bl[44] br[44] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_47 
+ bl[45] br[45] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_48 
+ bl[46] br[46] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_49 
+ bl[47] br[47] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_50 
+ bl[48] br[48] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_51 
+ bl[49] br[49] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_52 
+ bl[50] br[50] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_53 
+ bl[51] br[51] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_54 
+ bl[52] br[52] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_55 
+ bl[53] br[53] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_56 
+ bl[54] br[54] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_57 
+ bl[55] br[55] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_58 
+ bl[56] br[56] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_59 
+ bl[57] br[57] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_60 
+ bl[58] br[58] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_61 
+ bl[59] br[59] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_62 
+ bl[60] br[60] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_63 
+ bl[61] br[61] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_64 
+ bl[62] br[62] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_65 
+ bl[63] br[63] vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_66 
+ vdd vdd vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_491_67 
+ vdd vdd vdd vss wl[489] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_0 
+ vdd vdd vss vdd vpb vnb wl[490] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_492_1 
+ rbl rbr vss vdd vpb vnb wl[490] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_492_2 
+ bl[0] br[0] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_3 
+ bl[1] br[1] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_4 
+ bl[2] br[2] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_5 
+ bl[3] br[3] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_6 
+ bl[4] br[4] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_7 
+ bl[5] br[5] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_8 
+ bl[6] br[6] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_9 
+ bl[7] br[7] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_10 
+ bl[8] br[8] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_11 
+ bl[9] br[9] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_12 
+ bl[10] br[10] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_13 
+ bl[11] br[11] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_14 
+ bl[12] br[12] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_15 
+ bl[13] br[13] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_16 
+ bl[14] br[14] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_17 
+ bl[15] br[15] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_18 
+ bl[16] br[16] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_19 
+ bl[17] br[17] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_20 
+ bl[18] br[18] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_21 
+ bl[19] br[19] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_22 
+ bl[20] br[20] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_23 
+ bl[21] br[21] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_24 
+ bl[22] br[22] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_25 
+ bl[23] br[23] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_26 
+ bl[24] br[24] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_27 
+ bl[25] br[25] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_28 
+ bl[26] br[26] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_29 
+ bl[27] br[27] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_30 
+ bl[28] br[28] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_31 
+ bl[29] br[29] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_32 
+ bl[30] br[30] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_33 
+ bl[31] br[31] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_34 
+ bl[32] br[32] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_35 
+ bl[33] br[33] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_36 
+ bl[34] br[34] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_37 
+ bl[35] br[35] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_38 
+ bl[36] br[36] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_39 
+ bl[37] br[37] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_40 
+ bl[38] br[38] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_41 
+ bl[39] br[39] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_42 
+ bl[40] br[40] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_43 
+ bl[41] br[41] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_44 
+ bl[42] br[42] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_45 
+ bl[43] br[43] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_46 
+ bl[44] br[44] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_47 
+ bl[45] br[45] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_48 
+ bl[46] br[46] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_49 
+ bl[47] br[47] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_50 
+ bl[48] br[48] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_51 
+ bl[49] br[49] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_52 
+ bl[50] br[50] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_53 
+ bl[51] br[51] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_54 
+ bl[52] br[52] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_55 
+ bl[53] br[53] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_56 
+ bl[54] br[54] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_57 
+ bl[55] br[55] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_58 
+ bl[56] br[56] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_59 
+ bl[57] br[57] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_60 
+ bl[58] br[58] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_61 
+ bl[59] br[59] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_62 
+ bl[60] br[60] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_63 
+ bl[61] br[61] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_64 
+ bl[62] br[62] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_65 
+ bl[63] br[63] vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_66 
+ vdd vdd vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_492_67 
+ vdd vdd vdd vss wl[490] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_0 
+ vdd vdd vss vdd vpb vnb wl[491] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_493_1 
+ rbl rbr vss vdd vpb vnb wl[491] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_493_2 
+ bl[0] br[0] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_3 
+ bl[1] br[1] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_4 
+ bl[2] br[2] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_5 
+ bl[3] br[3] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_6 
+ bl[4] br[4] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_7 
+ bl[5] br[5] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_8 
+ bl[6] br[6] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_9 
+ bl[7] br[7] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_10 
+ bl[8] br[8] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_11 
+ bl[9] br[9] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_12 
+ bl[10] br[10] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_13 
+ bl[11] br[11] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_14 
+ bl[12] br[12] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_15 
+ bl[13] br[13] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_16 
+ bl[14] br[14] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_17 
+ bl[15] br[15] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_18 
+ bl[16] br[16] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_19 
+ bl[17] br[17] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_20 
+ bl[18] br[18] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_21 
+ bl[19] br[19] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_22 
+ bl[20] br[20] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_23 
+ bl[21] br[21] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_24 
+ bl[22] br[22] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_25 
+ bl[23] br[23] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_26 
+ bl[24] br[24] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_27 
+ bl[25] br[25] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_28 
+ bl[26] br[26] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_29 
+ bl[27] br[27] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_30 
+ bl[28] br[28] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_31 
+ bl[29] br[29] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_32 
+ bl[30] br[30] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_33 
+ bl[31] br[31] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_34 
+ bl[32] br[32] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_35 
+ bl[33] br[33] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_36 
+ bl[34] br[34] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_37 
+ bl[35] br[35] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_38 
+ bl[36] br[36] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_39 
+ bl[37] br[37] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_40 
+ bl[38] br[38] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_41 
+ bl[39] br[39] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_42 
+ bl[40] br[40] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_43 
+ bl[41] br[41] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_44 
+ bl[42] br[42] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_45 
+ bl[43] br[43] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_46 
+ bl[44] br[44] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_47 
+ bl[45] br[45] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_48 
+ bl[46] br[46] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_49 
+ bl[47] br[47] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_50 
+ bl[48] br[48] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_51 
+ bl[49] br[49] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_52 
+ bl[50] br[50] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_53 
+ bl[51] br[51] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_54 
+ bl[52] br[52] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_55 
+ bl[53] br[53] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_56 
+ bl[54] br[54] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_57 
+ bl[55] br[55] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_58 
+ bl[56] br[56] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_59 
+ bl[57] br[57] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_60 
+ bl[58] br[58] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_61 
+ bl[59] br[59] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_62 
+ bl[60] br[60] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_63 
+ bl[61] br[61] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_64 
+ bl[62] br[62] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_65 
+ bl[63] br[63] vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_66 
+ vdd vdd vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_493_67 
+ vdd vdd vdd vss wl[491] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_0 
+ vdd vdd vss vdd vpb vnb wl[492] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_494_1 
+ rbl rbr vss vdd vpb vnb wl[492] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_494_2 
+ bl[0] br[0] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_3 
+ bl[1] br[1] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_4 
+ bl[2] br[2] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_5 
+ bl[3] br[3] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_6 
+ bl[4] br[4] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_7 
+ bl[5] br[5] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_8 
+ bl[6] br[6] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_9 
+ bl[7] br[7] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_10 
+ bl[8] br[8] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_11 
+ bl[9] br[9] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_12 
+ bl[10] br[10] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_13 
+ bl[11] br[11] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_14 
+ bl[12] br[12] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_15 
+ bl[13] br[13] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_16 
+ bl[14] br[14] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_17 
+ bl[15] br[15] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_18 
+ bl[16] br[16] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_19 
+ bl[17] br[17] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_20 
+ bl[18] br[18] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_21 
+ bl[19] br[19] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_22 
+ bl[20] br[20] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_23 
+ bl[21] br[21] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_24 
+ bl[22] br[22] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_25 
+ bl[23] br[23] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_26 
+ bl[24] br[24] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_27 
+ bl[25] br[25] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_28 
+ bl[26] br[26] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_29 
+ bl[27] br[27] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_30 
+ bl[28] br[28] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_31 
+ bl[29] br[29] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_32 
+ bl[30] br[30] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_33 
+ bl[31] br[31] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_34 
+ bl[32] br[32] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_35 
+ bl[33] br[33] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_36 
+ bl[34] br[34] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_37 
+ bl[35] br[35] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_38 
+ bl[36] br[36] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_39 
+ bl[37] br[37] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_40 
+ bl[38] br[38] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_41 
+ bl[39] br[39] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_42 
+ bl[40] br[40] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_43 
+ bl[41] br[41] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_44 
+ bl[42] br[42] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_45 
+ bl[43] br[43] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_46 
+ bl[44] br[44] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_47 
+ bl[45] br[45] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_48 
+ bl[46] br[46] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_49 
+ bl[47] br[47] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_50 
+ bl[48] br[48] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_51 
+ bl[49] br[49] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_52 
+ bl[50] br[50] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_53 
+ bl[51] br[51] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_54 
+ bl[52] br[52] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_55 
+ bl[53] br[53] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_56 
+ bl[54] br[54] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_57 
+ bl[55] br[55] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_58 
+ bl[56] br[56] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_59 
+ bl[57] br[57] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_60 
+ bl[58] br[58] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_61 
+ bl[59] br[59] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_62 
+ bl[60] br[60] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_63 
+ bl[61] br[61] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_64 
+ bl[62] br[62] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_65 
+ bl[63] br[63] vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_66 
+ vdd vdd vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_494_67 
+ vdd vdd vdd vss wl[492] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_0 
+ vdd vdd vss vdd vpb vnb wl[493] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_495_1 
+ rbl rbr vss vdd vpb vnb wl[493] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_495_2 
+ bl[0] br[0] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_3 
+ bl[1] br[1] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_4 
+ bl[2] br[2] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_5 
+ bl[3] br[3] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_6 
+ bl[4] br[4] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_7 
+ bl[5] br[5] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_8 
+ bl[6] br[6] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_9 
+ bl[7] br[7] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_10 
+ bl[8] br[8] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_11 
+ bl[9] br[9] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_12 
+ bl[10] br[10] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_13 
+ bl[11] br[11] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_14 
+ bl[12] br[12] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_15 
+ bl[13] br[13] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_16 
+ bl[14] br[14] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_17 
+ bl[15] br[15] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_18 
+ bl[16] br[16] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_19 
+ bl[17] br[17] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_20 
+ bl[18] br[18] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_21 
+ bl[19] br[19] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_22 
+ bl[20] br[20] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_23 
+ bl[21] br[21] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_24 
+ bl[22] br[22] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_25 
+ bl[23] br[23] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_26 
+ bl[24] br[24] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_27 
+ bl[25] br[25] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_28 
+ bl[26] br[26] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_29 
+ bl[27] br[27] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_30 
+ bl[28] br[28] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_31 
+ bl[29] br[29] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_32 
+ bl[30] br[30] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_33 
+ bl[31] br[31] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_34 
+ bl[32] br[32] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_35 
+ bl[33] br[33] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_36 
+ bl[34] br[34] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_37 
+ bl[35] br[35] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_38 
+ bl[36] br[36] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_39 
+ bl[37] br[37] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_40 
+ bl[38] br[38] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_41 
+ bl[39] br[39] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_42 
+ bl[40] br[40] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_43 
+ bl[41] br[41] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_44 
+ bl[42] br[42] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_45 
+ bl[43] br[43] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_46 
+ bl[44] br[44] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_47 
+ bl[45] br[45] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_48 
+ bl[46] br[46] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_49 
+ bl[47] br[47] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_50 
+ bl[48] br[48] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_51 
+ bl[49] br[49] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_52 
+ bl[50] br[50] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_53 
+ bl[51] br[51] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_54 
+ bl[52] br[52] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_55 
+ bl[53] br[53] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_56 
+ bl[54] br[54] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_57 
+ bl[55] br[55] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_58 
+ bl[56] br[56] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_59 
+ bl[57] br[57] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_60 
+ bl[58] br[58] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_61 
+ bl[59] br[59] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_62 
+ bl[60] br[60] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_63 
+ bl[61] br[61] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_64 
+ bl[62] br[62] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_65 
+ bl[63] br[63] vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_66 
+ vdd vdd vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_495_67 
+ vdd vdd vdd vss wl[493] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_0 
+ vdd vdd vss vdd vpb vnb wl[494] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_496_1 
+ rbl rbr vss vdd vpb vnb wl[494] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_496_2 
+ bl[0] br[0] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_3 
+ bl[1] br[1] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_4 
+ bl[2] br[2] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_5 
+ bl[3] br[3] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_6 
+ bl[4] br[4] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_7 
+ bl[5] br[5] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_8 
+ bl[6] br[6] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_9 
+ bl[7] br[7] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_10 
+ bl[8] br[8] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_11 
+ bl[9] br[9] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_12 
+ bl[10] br[10] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_13 
+ bl[11] br[11] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_14 
+ bl[12] br[12] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_15 
+ bl[13] br[13] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_16 
+ bl[14] br[14] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_17 
+ bl[15] br[15] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_18 
+ bl[16] br[16] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_19 
+ bl[17] br[17] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_20 
+ bl[18] br[18] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_21 
+ bl[19] br[19] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_22 
+ bl[20] br[20] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_23 
+ bl[21] br[21] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_24 
+ bl[22] br[22] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_25 
+ bl[23] br[23] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_26 
+ bl[24] br[24] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_27 
+ bl[25] br[25] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_28 
+ bl[26] br[26] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_29 
+ bl[27] br[27] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_30 
+ bl[28] br[28] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_31 
+ bl[29] br[29] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_32 
+ bl[30] br[30] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_33 
+ bl[31] br[31] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_34 
+ bl[32] br[32] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_35 
+ bl[33] br[33] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_36 
+ bl[34] br[34] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_37 
+ bl[35] br[35] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_38 
+ bl[36] br[36] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_39 
+ bl[37] br[37] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_40 
+ bl[38] br[38] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_41 
+ bl[39] br[39] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_42 
+ bl[40] br[40] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_43 
+ bl[41] br[41] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_44 
+ bl[42] br[42] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_45 
+ bl[43] br[43] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_46 
+ bl[44] br[44] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_47 
+ bl[45] br[45] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_48 
+ bl[46] br[46] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_49 
+ bl[47] br[47] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_50 
+ bl[48] br[48] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_51 
+ bl[49] br[49] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_52 
+ bl[50] br[50] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_53 
+ bl[51] br[51] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_54 
+ bl[52] br[52] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_55 
+ bl[53] br[53] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_56 
+ bl[54] br[54] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_57 
+ bl[55] br[55] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_58 
+ bl[56] br[56] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_59 
+ bl[57] br[57] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_60 
+ bl[58] br[58] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_61 
+ bl[59] br[59] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_62 
+ bl[60] br[60] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_63 
+ bl[61] br[61] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_64 
+ bl[62] br[62] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_65 
+ bl[63] br[63] vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_66 
+ vdd vdd vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_496_67 
+ vdd vdd vdd vss wl[494] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_0 
+ vdd vdd vss vdd vpb vnb wl[495] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_497_1 
+ rbl rbr vss vdd vpb vnb wl[495] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_497_2 
+ bl[0] br[0] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_3 
+ bl[1] br[1] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_4 
+ bl[2] br[2] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_5 
+ bl[3] br[3] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_6 
+ bl[4] br[4] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_7 
+ bl[5] br[5] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_8 
+ bl[6] br[6] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_9 
+ bl[7] br[7] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_10 
+ bl[8] br[8] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_11 
+ bl[9] br[9] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_12 
+ bl[10] br[10] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_13 
+ bl[11] br[11] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_14 
+ bl[12] br[12] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_15 
+ bl[13] br[13] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_16 
+ bl[14] br[14] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_17 
+ bl[15] br[15] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_18 
+ bl[16] br[16] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_19 
+ bl[17] br[17] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_20 
+ bl[18] br[18] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_21 
+ bl[19] br[19] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_22 
+ bl[20] br[20] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_23 
+ bl[21] br[21] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_24 
+ bl[22] br[22] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_25 
+ bl[23] br[23] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_26 
+ bl[24] br[24] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_27 
+ bl[25] br[25] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_28 
+ bl[26] br[26] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_29 
+ bl[27] br[27] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_30 
+ bl[28] br[28] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_31 
+ bl[29] br[29] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_32 
+ bl[30] br[30] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_33 
+ bl[31] br[31] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_34 
+ bl[32] br[32] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_35 
+ bl[33] br[33] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_36 
+ bl[34] br[34] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_37 
+ bl[35] br[35] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_38 
+ bl[36] br[36] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_39 
+ bl[37] br[37] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_40 
+ bl[38] br[38] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_41 
+ bl[39] br[39] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_42 
+ bl[40] br[40] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_43 
+ bl[41] br[41] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_44 
+ bl[42] br[42] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_45 
+ bl[43] br[43] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_46 
+ bl[44] br[44] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_47 
+ bl[45] br[45] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_48 
+ bl[46] br[46] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_49 
+ bl[47] br[47] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_50 
+ bl[48] br[48] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_51 
+ bl[49] br[49] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_52 
+ bl[50] br[50] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_53 
+ bl[51] br[51] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_54 
+ bl[52] br[52] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_55 
+ bl[53] br[53] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_56 
+ bl[54] br[54] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_57 
+ bl[55] br[55] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_58 
+ bl[56] br[56] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_59 
+ bl[57] br[57] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_60 
+ bl[58] br[58] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_61 
+ bl[59] br[59] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_62 
+ bl[60] br[60] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_63 
+ bl[61] br[61] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_64 
+ bl[62] br[62] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_65 
+ bl[63] br[63] vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_66 
+ vdd vdd vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_497_67 
+ vdd vdd vdd vss wl[495] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_0 
+ vdd vdd vss vdd vpb vnb wl[496] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_498_1 
+ rbl rbr vss vdd vpb vnb wl[496] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_498_2 
+ bl[0] br[0] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_3 
+ bl[1] br[1] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_4 
+ bl[2] br[2] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_5 
+ bl[3] br[3] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_6 
+ bl[4] br[4] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_7 
+ bl[5] br[5] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_8 
+ bl[6] br[6] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_9 
+ bl[7] br[7] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_10 
+ bl[8] br[8] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_11 
+ bl[9] br[9] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_12 
+ bl[10] br[10] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_13 
+ bl[11] br[11] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_14 
+ bl[12] br[12] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_15 
+ bl[13] br[13] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_16 
+ bl[14] br[14] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_17 
+ bl[15] br[15] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_18 
+ bl[16] br[16] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_19 
+ bl[17] br[17] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_20 
+ bl[18] br[18] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_21 
+ bl[19] br[19] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_22 
+ bl[20] br[20] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_23 
+ bl[21] br[21] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_24 
+ bl[22] br[22] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_25 
+ bl[23] br[23] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_26 
+ bl[24] br[24] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_27 
+ bl[25] br[25] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_28 
+ bl[26] br[26] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_29 
+ bl[27] br[27] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_30 
+ bl[28] br[28] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_31 
+ bl[29] br[29] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_32 
+ bl[30] br[30] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_33 
+ bl[31] br[31] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_34 
+ bl[32] br[32] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_35 
+ bl[33] br[33] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_36 
+ bl[34] br[34] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_37 
+ bl[35] br[35] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_38 
+ bl[36] br[36] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_39 
+ bl[37] br[37] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_40 
+ bl[38] br[38] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_41 
+ bl[39] br[39] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_42 
+ bl[40] br[40] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_43 
+ bl[41] br[41] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_44 
+ bl[42] br[42] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_45 
+ bl[43] br[43] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_46 
+ bl[44] br[44] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_47 
+ bl[45] br[45] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_48 
+ bl[46] br[46] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_49 
+ bl[47] br[47] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_50 
+ bl[48] br[48] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_51 
+ bl[49] br[49] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_52 
+ bl[50] br[50] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_53 
+ bl[51] br[51] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_54 
+ bl[52] br[52] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_55 
+ bl[53] br[53] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_56 
+ bl[54] br[54] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_57 
+ bl[55] br[55] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_58 
+ bl[56] br[56] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_59 
+ bl[57] br[57] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_60 
+ bl[58] br[58] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_61 
+ bl[59] br[59] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_62 
+ bl[60] br[60] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_63 
+ bl[61] br[61] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_64 
+ bl[62] br[62] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_65 
+ bl[63] br[63] vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_66 
+ vdd vdd vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_498_67 
+ vdd vdd vdd vss wl[496] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_0 
+ vdd vdd vss vdd vpb vnb wl[497] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_499_1 
+ rbl rbr vss vdd vpb vnb wl[497] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_499_2 
+ bl[0] br[0] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_3 
+ bl[1] br[1] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_4 
+ bl[2] br[2] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_5 
+ bl[3] br[3] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_6 
+ bl[4] br[4] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_7 
+ bl[5] br[5] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_8 
+ bl[6] br[6] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_9 
+ bl[7] br[7] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_10 
+ bl[8] br[8] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_11 
+ bl[9] br[9] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_12 
+ bl[10] br[10] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_13 
+ bl[11] br[11] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_14 
+ bl[12] br[12] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_15 
+ bl[13] br[13] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_16 
+ bl[14] br[14] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_17 
+ bl[15] br[15] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_18 
+ bl[16] br[16] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_19 
+ bl[17] br[17] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_20 
+ bl[18] br[18] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_21 
+ bl[19] br[19] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_22 
+ bl[20] br[20] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_23 
+ bl[21] br[21] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_24 
+ bl[22] br[22] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_25 
+ bl[23] br[23] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_26 
+ bl[24] br[24] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_27 
+ bl[25] br[25] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_28 
+ bl[26] br[26] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_29 
+ bl[27] br[27] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_30 
+ bl[28] br[28] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_31 
+ bl[29] br[29] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_32 
+ bl[30] br[30] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_33 
+ bl[31] br[31] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_34 
+ bl[32] br[32] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_35 
+ bl[33] br[33] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_36 
+ bl[34] br[34] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_37 
+ bl[35] br[35] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_38 
+ bl[36] br[36] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_39 
+ bl[37] br[37] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_40 
+ bl[38] br[38] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_41 
+ bl[39] br[39] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_42 
+ bl[40] br[40] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_43 
+ bl[41] br[41] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_44 
+ bl[42] br[42] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_45 
+ bl[43] br[43] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_46 
+ bl[44] br[44] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_47 
+ bl[45] br[45] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_48 
+ bl[46] br[46] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_49 
+ bl[47] br[47] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_50 
+ bl[48] br[48] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_51 
+ bl[49] br[49] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_52 
+ bl[50] br[50] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_53 
+ bl[51] br[51] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_54 
+ bl[52] br[52] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_55 
+ bl[53] br[53] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_56 
+ bl[54] br[54] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_57 
+ bl[55] br[55] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_58 
+ bl[56] br[56] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_59 
+ bl[57] br[57] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_60 
+ bl[58] br[58] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_61 
+ bl[59] br[59] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_62 
+ bl[60] br[60] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_63 
+ bl[61] br[61] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_64 
+ bl[62] br[62] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_65 
+ bl[63] br[63] vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_66 
+ vdd vdd vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_499_67 
+ vdd vdd vdd vss wl[497] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_0 
+ vdd vdd vss vdd vpb vnb wl[498] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_500_1 
+ rbl rbr vss vdd vpb vnb wl[498] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_500_2 
+ bl[0] br[0] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_3 
+ bl[1] br[1] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_4 
+ bl[2] br[2] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_5 
+ bl[3] br[3] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_6 
+ bl[4] br[4] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_7 
+ bl[5] br[5] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_8 
+ bl[6] br[6] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_9 
+ bl[7] br[7] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_10 
+ bl[8] br[8] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_11 
+ bl[9] br[9] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_12 
+ bl[10] br[10] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_13 
+ bl[11] br[11] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_14 
+ bl[12] br[12] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_15 
+ bl[13] br[13] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_16 
+ bl[14] br[14] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_17 
+ bl[15] br[15] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_18 
+ bl[16] br[16] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_19 
+ bl[17] br[17] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_20 
+ bl[18] br[18] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_21 
+ bl[19] br[19] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_22 
+ bl[20] br[20] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_23 
+ bl[21] br[21] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_24 
+ bl[22] br[22] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_25 
+ bl[23] br[23] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_26 
+ bl[24] br[24] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_27 
+ bl[25] br[25] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_28 
+ bl[26] br[26] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_29 
+ bl[27] br[27] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_30 
+ bl[28] br[28] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_31 
+ bl[29] br[29] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_32 
+ bl[30] br[30] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_33 
+ bl[31] br[31] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_34 
+ bl[32] br[32] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_35 
+ bl[33] br[33] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_36 
+ bl[34] br[34] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_37 
+ bl[35] br[35] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_38 
+ bl[36] br[36] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_39 
+ bl[37] br[37] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_40 
+ bl[38] br[38] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_41 
+ bl[39] br[39] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_42 
+ bl[40] br[40] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_43 
+ bl[41] br[41] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_44 
+ bl[42] br[42] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_45 
+ bl[43] br[43] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_46 
+ bl[44] br[44] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_47 
+ bl[45] br[45] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_48 
+ bl[46] br[46] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_49 
+ bl[47] br[47] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_50 
+ bl[48] br[48] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_51 
+ bl[49] br[49] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_52 
+ bl[50] br[50] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_53 
+ bl[51] br[51] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_54 
+ bl[52] br[52] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_55 
+ bl[53] br[53] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_56 
+ bl[54] br[54] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_57 
+ bl[55] br[55] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_58 
+ bl[56] br[56] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_59 
+ bl[57] br[57] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_60 
+ bl[58] br[58] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_61 
+ bl[59] br[59] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_62 
+ bl[60] br[60] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_63 
+ bl[61] br[61] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_64 
+ bl[62] br[62] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_65 
+ bl[63] br[63] vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_66 
+ vdd vdd vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_500_67 
+ vdd vdd vdd vss wl[498] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_0 
+ vdd vdd vss vdd vpb vnb wl[499] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_501_1 
+ rbl rbr vss vdd vpb vnb wl[499] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_501_2 
+ bl[0] br[0] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_3 
+ bl[1] br[1] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_4 
+ bl[2] br[2] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_5 
+ bl[3] br[3] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_6 
+ bl[4] br[4] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_7 
+ bl[5] br[5] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_8 
+ bl[6] br[6] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_9 
+ bl[7] br[7] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_10 
+ bl[8] br[8] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_11 
+ bl[9] br[9] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_12 
+ bl[10] br[10] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_13 
+ bl[11] br[11] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_14 
+ bl[12] br[12] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_15 
+ bl[13] br[13] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_16 
+ bl[14] br[14] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_17 
+ bl[15] br[15] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_18 
+ bl[16] br[16] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_19 
+ bl[17] br[17] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_20 
+ bl[18] br[18] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_21 
+ bl[19] br[19] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_22 
+ bl[20] br[20] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_23 
+ bl[21] br[21] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_24 
+ bl[22] br[22] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_25 
+ bl[23] br[23] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_26 
+ bl[24] br[24] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_27 
+ bl[25] br[25] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_28 
+ bl[26] br[26] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_29 
+ bl[27] br[27] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_30 
+ bl[28] br[28] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_31 
+ bl[29] br[29] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_32 
+ bl[30] br[30] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_33 
+ bl[31] br[31] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_34 
+ bl[32] br[32] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_35 
+ bl[33] br[33] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_36 
+ bl[34] br[34] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_37 
+ bl[35] br[35] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_38 
+ bl[36] br[36] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_39 
+ bl[37] br[37] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_40 
+ bl[38] br[38] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_41 
+ bl[39] br[39] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_42 
+ bl[40] br[40] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_43 
+ bl[41] br[41] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_44 
+ bl[42] br[42] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_45 
+ bl[43] br[43] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_46 
+ bl[44] br[44] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_47 
+ bl[45] br[45] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_48 
+ bl[46] br[46] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_49 
+ bl[47] br[47] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_50 
+ bl[48] br[48] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_51 
+ bl[49] br[49] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_52 
+ bl[50] br[50] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_53 
+ bl[51] br[51] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_54 
+ bl[52] br[52] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_55 
+ bl[53] br[53] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_56 
+ bl[54] br[54] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_57 
+ bl[55] br[55] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_58 
+ bl[56] br[56] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_59 
+ bl[57] br[57] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_60 
+ bl[58] br[58] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_61 
+ bl[59] br[59] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_62 
+ bl[60] br[60] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_63 
+ bl[61] br[61] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_64 
+ bl[62] br[62] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_65 
+ bl[63] br[63] vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_66 
+ vdd vdd vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_501_67 
+ vdd vdd vdd vss wl[499] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_0 
+ vdd vdd vss vdd vpb vnb wl[500] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_502_1 
+ rbl rbr vss vdd vpb vnb wl[500] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_502_2 
+ bl[0] br[0] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_3 
+ bl[1] br[1] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_4 
+ bl[2] br[2] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_5 
+ bl[3] br[3] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_6 
+ bl[4] br[4] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_7 
+ bl[5] br[5] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_8 
+ bl[6] br[6] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_9 
+ bl[7] br[7] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_10 
+ bl[8] br[8] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_11 
+ bl[9] br[9] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_12 
+ bl[10] br[10] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_13 
+ bl[11] br[11] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_14 
+ bl[12] br[12] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_15 
+ bl[13] br[13] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_16 
+ bl[14] br[14] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_17 
+ bl[15] br[15] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_18 
+ bl[16] br[16] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_19 
+ bl[17] br[17] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_20 
+ bl[18] br[18] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_21 
+ bl[19] br[19] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_22 
+ bl[20] br[20] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_23 
+ bl[21] br[21] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_24 
+ bl[22] br[22] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_25 
+ bl[23] br[23] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_26 
+ bl[24] br[24] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_27 
+ bl[25] br[25] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_28 
+ bl[26] br[26] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_29 
+ bl[27] br[27] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_30 
+ bl[28] br[28] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_31 
+ bl[29] br[29] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_32 
+ bl[30] br[30] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_33 
+ bl[31] br[31] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_34 
+ bl[32] br[32] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_35 
+ bl[33] br[33] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_36 
+ bl[34] br[34] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_37 
+ bl[35] br[35] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_38 
+ bl[36] br[36] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_39 
+ bl[37] br[37] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_40 
+ bl[38] br[38] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_41 
+ bl[39] br[39] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_42 
+ bl[40] br[40] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_43 
+ bl[41] br[41] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_44 
+ bl[42] br[42] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_45 
+ bl[43] br[43] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_46 
+ bl[44] br[44] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_47 
+ bl[45] br[45] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_48 
+ bl[46] br[46] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_49 
+ bl[47] br[47] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_50 
+ bl[48] br[48] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_51 
+ bl[49] br[49] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_52 
+ bl[50] br[50] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_53 
+ bl[51] br[51] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_54 
+ bl[52] br[52] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_55 
+ bl[53] br[53] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_56 
+ bl[54] br[54] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_57 
+ bl[55] br[55] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_58 
+ bl[56] br[56] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_59 
+ bl[57] br[57] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_60 
+ bl[58] br[58] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_61 
+ bl[59] br[59] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_62 
+ bl[60] br[60] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_63 
+ bl[61] br[61] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_64 
+ bl[62] br[62] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_65 
+ bl[63] br[63] vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_66 
+ vdd vdd vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_502_67 
+ vdd vdd vdd vss wl[500] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_0 
+ vdd vdd vss vdd vpb vnb wl[501] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_503_1 
+ rbl rbr vss vdd vpb vnb wl[501] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_503_2 
+ bl[0] br[0] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_3 
+ bl[1] br[1] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_4 
+ bl[2] br[2] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_5 
+ bl[3] br[3] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_6 
+ bl[4] br[4] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_7 
+ bl[5] br[5] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_8 
+ bl[6] br[6] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_9 
+ bl[7] br[7] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_10 
+ bl[8] br[8] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_11 
+ bl[9] br[9] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_12 
+ bl[10] br[10] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_13 
+ bl[11] br[11] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_14 
+ bl[12] br[12] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_15 
+ bl[13] br[13] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_16 
+ bl[14] br[14] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_17 
+ bl[15] br[15] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_18 
+ bl[16] br[16] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_19 
+ bl[17] br[17] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_20 
+ bl[18] br[18] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_21 
+ bl[19] br[19] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_22 
+ bl[20] br[20] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_23 
+ bl[21] br[21] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_24 
+ bl[22] br[22] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_25 
+ bl[23] br[23] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_26 
+ bl[24] br[24] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_27 
+ bl[25] br[25] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_28 
+ bl[26] br[26] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_29 
+ bl[27] br[27] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_30 
+ bl[28] br[28] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_31 
+ bl[29] br[29] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_32 
+ bl[30] br[30] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_33 
+ bl[31] br[31] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_34 
+ bl[32] br[32] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_35 
+ bl[33] br[33] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_36 
+ bl[34] br[34] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_37 
+ bl[35] br[35] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_38 
+ bl[36] br[36] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_39 
+ bl[37] br[37] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_40 
+ bl[38] br[38] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_41 
+ bl[39] br[39] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_42 
+ bl[40] br[40] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_43 
+ bl[41] br[41] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_44 
+ bl[42] br[42] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_45 
+ bl[43] br[43] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_46 
+ bl[44] br[44] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_47 
+ bl[45] br[45] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_48 
+ bl[46] br[46] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_49 
+ bl[47] br[47] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_50 
+ bl[48] br[48] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_51 
+ bl[49] br[49] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_52 
+ bl[50] br[50] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_53 
+ bl[51] br[51] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_54 
+ bl[52] br[52] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_55 
+ bl[53] br[53] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_56 
+ bl[54] br[54] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_57 
+ bl[55] br[55] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_58 
+ bl[56] br[56] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_59 
+ bl[57] br[57] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_60 
+ bl[58] br[58] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_61 
+ bl[59] br[59] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_62 
+ bl[60] br[60] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_63 
+ bl[61] br[61] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_64 
+ bl[62] br[62] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_65 
+ bl[63] br[63] vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_66 
+ vdd vdd vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_503_67 
+ vdd vdd vdd vss wl[501] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_0 
+ vdd vdd vss vdd vpb vnb wl[502] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_504_1 
+ rbl rbr vss vdd vpb vnb wl[502] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_504_2 
+ bl[0] br[0] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_3 
+ bl[1] br[1] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_4 
+ bl[2] br[2] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_5 
+ bl[3] br[3] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_6 
+ bl[4] br[4] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_7 
+ bl[5] br[5] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_8 
+ bl[6] br[6] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_9 
+ bl[7] br[7] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_10 
+ bl[8] br[8] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_11 
+ bl[9] br[9] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_12 
+ bl[10] br[10] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_13 
+ bl[11] br[11] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_14 
+ bl[12] br[12] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_15 
+ bl[13] br[13] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_16 
+ bl[14] br[14] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_17 
+ bl[15] br[15] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_18 
+ bl[16] br[16] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_19 
+ bl[17] br[17] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_20 
+ bl[18] br[18] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_21 
+ bl[19] br[19] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_22 
+ bl[20] br[20] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_23 
+ bl[21] br[21] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_24 
+ bl[22] br[22] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_25 
+ bl[23] br[23] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_26 
+ bl[24] br[24] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_27 
+ bl[25] br[25] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_28 
+ bl[26] br[26] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_29 
+ bl[27] br[27] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_30 
+ bl[28] br[28] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_31 
+ bl[29] br[29] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_32 
+ bl[30] br[30] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_33 
+ bl[31] br[31] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_34 
+ bl[32] br[32] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_35 
+ bl[33] br[33] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_36 
+ bl[34] br[34] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_37 
+ bl[35] br[35] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_38 
+ bl[36] br[36] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_39 
+ bl[37] br[37] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_40 
+ bl[38] br[38] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_41 
+ bl[39] br[39] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_42 
+ bl[40] br[40] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_43 
+ bl[41] br[41] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_44 
+ bl[42] br[42] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_45 
+ bl[43] br[43] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_46 
+ bl[44] br[44] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_47 
+ bl[45] br[45] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_48 
+ bl[46] br[46] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_49 
+ bl[47] br[47] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_50 
+ bl[48] br[48] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_51 
+ bl[49] br[49] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_52 
+ bl[50] br[50] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_53 
+ bl[51] br[51] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_54 
+ bl[52] br[52] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_55 
+ bl[53] br[53] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_56 
+ bl[54] br[54] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_57 
+ bl[55] br[55] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_58 
+ bl[56] br[56] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_59 
+ bl[57] br[57] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_60 
+ bl[58] br[58] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_61 
+ bl[59] br[59] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_62 
+ bl[60] br[60] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_63 
+ bl[61] br[61] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_64 
+ bl[62] br[62] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_65 
+ bl[63] br[63] vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_66 
+ vdd vdd vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_504_67 
+ vdd vdd vdd vss wl[502] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_0 
+ vdd vdd vss vdd vpb vnb wl[503] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_505_1 
+ rbl rbr vss vdd vpb vnb wl[503] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_505_2 
+ bl[0] br[0] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_3 
+ bl[1] br[1] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_4 
+ bl[2] br[2] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_5 
+ bl[3] br[3] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_6 
+ bl[4] br[4] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_7 
+ bl[5] br[5] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_8 
+ bl[6] br[6] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_9 
+ bl[7] br[7] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_10 
+ bl[8] br[8] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_11 
+ bl[9] br[9] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_12 
+ bl[10] br[10] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_13 
+ bl[11] br[11] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_14 
+ bl[12] br[12] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_15 
+ bl[13] br[13] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_16 
+ bl[14] br[14] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_17 
+ bl[15] br[15] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_18 
+ bl[16] br[16] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_19 
+ bl[17] br[17] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_20 
+ bl[18] br[18] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_21 
+ bl[19] br[19] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_22 
+ bl[20] br[20] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_23 
+ bl[21] br[21] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_24 
+ bl[22] br[22] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_25 
+ bl[23] br[23] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_26 
+ bl[24] br[24] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_27 
+ bl[25] br[25] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_28 
+ bl[26] br[26] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_29 
+ bl[27] br[27] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_30 
+ bl[28] br[28] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_31 
+ bl[29] br[29] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_32 
+ bl[30] br[30] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_33 
+ bl[31] br[31] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_34 
+ bl[32] br[32] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_35 
+ bl[33] br[33] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_36 
+ bl[34] br[34] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_37 
+ bl[35] br[35] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_38 
+ bl[36] br[36] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_39 
+ bl[37] br[37] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_40 
+ bl[38] br[38] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_41 
+ bl[39] br[39] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_42 
+ bl[40] br[40] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_43 
+ bl[41] br[41] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_44 
+ bl[42] br[42] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_45 
+ bl[43] br[43] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_46 
+ bl[44] br[44] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_47 
+ bl[45] br[45] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_48 
+ bl[46] br[46] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_49 
+ bl[47] br[47] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_50 
+ bl[48] br[48] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_51 
+ bl[49] br[49] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_52 
+ bl[50] br[50] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_53 
+ bl[51] br[51] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_54 
+ bl[52] br[52] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_55 
+ bl[53] br[53] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_56 
+ bl[54] br[54] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_57 
+ bl[55] br[55] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_58 
+ bl[56] br[56] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_59 
+ bl[57] br[57] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_60 
+ bl[58] br[58] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_61 
+ bl[59] br[59] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_62 
+ bl[60] br[60] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_63 
+ bl[61] br[61] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_64 
+ bl[62] br[62] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_65 
+ bl[63] br[63] vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_66 
+ vdd vdd vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_505_67 
+ vdd vdd vdd vss wl[503] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_0 
+ vdd vdd vss vdd vpb vnb wl[504] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_506_1 
+ rbl rbr vss vdd vpb vnb wl[504] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_506_2 
+ bl[0] br[0] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_3 
+ bl[1] br[1] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_4 
+ bl[2] br[2] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_5 
+ bl[3] br[3] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_6 
+ bl[4] br[4] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_7 
+ bl[5] br[5] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_8 
+ bl[6] br[6] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_9 
+ bl[7] br[7] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_10 
+ bl[8] br[8] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_11 
+ bl[9] br[9] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_12 
+ bl[10] br[10] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_13 
+ bl[11] br[11] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_14 
+ bl[12] br[12] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_15 
+ bl[13] br[13] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_16 
+ bl[14] br[14] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_17 
+ bl[15] br[15] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_18 
+ bl[16] br[16] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_19 
+ bl[17] br[17] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_20 
+ bl[18] br[18] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_21 
+ bl[19] br[19] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_22 
+ bl[20] br[20] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_23 
+ bl[21] br[21] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_24 
+ bl[22] br[22] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_25 
+ bl[23] br[23] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_26 
+ bl[24] br[24] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_27 
+ bl[25] br[25] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_28 
+ bl[26] br[26] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_29 
+ bl[27] br[27] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_30 
+ bl[28] br[28] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_31 
+ bl[29] br[29] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_32 
+ bl[30] br[30] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_33 
+ bl[31] br[31] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_34 
+ bl[32] br[32] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_35 
+ bl[33] br[33] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_36 
+ bl[34] br[34] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_37 
+ bl[35] br[35] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_38 
+ bl[36] br[36] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_39 
+ bl[37] br[37] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_40 
+ bl[38] br[38] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_41 
+ bl[39] br[39] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_42 
+ bl[40] br[40] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_43 
+ bl[41] br[41] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_44 
+ bl[42] br[42] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_45 
+ bl[43] br[43] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_46 
+ bl[44] br[44] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_47 
+ bl[45] br[45] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_48 
+ bl[46] br[46] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_49 
+ bl[47] br[47] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_50 
+ bl[48] br[48] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_51 
+ bl[49] br[49] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_52 
+ bl[50] br[50] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_53 
+ bl[51] br[51] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_54 
+ bl[52] br[52] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_55 
+ bl[53] br[53] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_56 
+ bl[54] br[54] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_57 
+ bl[55] br[55] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_58 
+ bl[56] br[56] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_59 
+ bl[57] br[57] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_60 
+ bl[58] br[58] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_61 
+ bl[59] br[59] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_62 
+ bl[60] br[60] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_63 
+ bl[61] br[61] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_64 
+ bl[62] br[62] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_65 
+ bl[63] br[63] vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_66 
+ vdd vdd vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_506_67 
+ vdd vdd vdd vss wl[504] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_0 
+ vdd vdd vss vdd vpb vnb wl[505] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_507_1 
+ rbl rbr vss vdd vpb vnb wl[505] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_507_2 
+ bl[0] br[0] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_3 
+ bl[1] br[1] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_4 
+ bl[2] br[2] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_5 
+ bl[3] br[3] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_6 
+ bl[4] br[4] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_7 
+ bl[5] br[5] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_8 
+ bl[6] br[6] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_9 
+ bl[7] br[7] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_10 
+ bl[8] br[8] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_11 
+ bl[9] br[9] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_12 
+ bl[10] br[10] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_13 
+ bl[11] br[11] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_14 
+ bl[12] br[12] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_15 
+ bl[13] br[13] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_16 
+ bl[14] br[14] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_17 
+ bl[15] br[15] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_18 
+ bl[16] br[16] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_19 
+ bl[17] br[17] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_20 
+ bl[18] br[18] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_21 
+ bl[19] br[19] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_22 
+ bl[20] br[20] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_23 
+ bl[21] br[21] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_24 
+ bl[22] br[22] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_25 
+ bl[23] br[23] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_26 
+ bl[24] br[24] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_27 
+ bl[25] br[25] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_28 
+ bl[26] br[26] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_29 
+ bl[27] br[27] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_30 
+ bl[28] br[28] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_31 
+ bl[29] br[29] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_32 
+ bl[30] br[30] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_33 
+ bl[31] br[31] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_34 
+ bl[32] br[32] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_35 
+ bl[33] br[33] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_36 
+ bl[34] br[34] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_37 
+ bl[35] br[35] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_38 
+ bl[36] br[36] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_39 
+ bl[37] br[37] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_40 
+ bl[38] br[38] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_41 
+ bl[39] br[39] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_42 
+ bl[40] br[40] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_43 
+ bl[41] br[41] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_44 
+ bl[42] br[42] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_45 
+ bl[43] br[43] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_46 
+ bl[44] br[44] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_47 
+ bl[45] br[45] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_48 
+ bl[46] br[46] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_49 
+ bl[47] br[47] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_50 
+ bl[48] br[48] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_51 
+ bl[49] br[49] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_52 
+ bl[50] br[50] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_53 
+ bl[51] br[51] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_54 
+ bl[52] br[52] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_55 
+ bl[53] br[53] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_56 
+ bl[54] br[54] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_57 
+ bl[55] br[55] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_58 
+ bl[56] br[56] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_59 
+ bl[57] br[57] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_60 
+ bl[58] br[58] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_61 
+ bl[59] br[59] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_62 
+ bl[60] br[60] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_63 
+ bl[61] br[61] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_64 
+ bl[62] br[62] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_65 
+ bl[63] br[63] vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_66 
+ vdd vdd vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_507_67 
+ vdd vdd vdd vss wl[505] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_0 
+ vdd vdd vss vdd vpb vnb wl[506] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_508_1 
+ rbl rbr vss vdd vpb vnb wl[506] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_508_2 
+ bl[0] br[0] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_3 
+ bl[1] br[1] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_4 
+ bl[2] br[2] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_5 
+ bl[3] br[3] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_6 
+ bl[4] br[4] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_7 
+ bl[5] br[5] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_8 
+ bl[6] br[6] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_9 
+ bl[7] br[7] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_10 
+ bl[8] br[8] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_11 
+ bl[9] br[9] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_12 
+ bl[10] br[10] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_13 
+ bl[11] br[11] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_14 
+ bl[12] br[12] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_15 
+ bl[13] br[13] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_16 
+ bl[14] br[14] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_17 
+ bl[15] br[15] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_18 
+ bl[16] br[16] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_19 
+ bl[17] br[17] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_20 
+ bl[18] br[18] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_21 
+ bl[19] br[19] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_22 
+ bl[20] br[20] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_23 
+ bl[21] br[21] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_24 
+ bl[22] br[22] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_25 
+ bl[23] br[23] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_26 
+ bl[24] br[24] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_27 
+ bl[25] br[25] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_28 
+ bl[26] br[26] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_29 
+ bl[27] br[27] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_30 
+ bl[28] br[28] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_31 
+ bl[29] br[29] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_32 
+ bl[30] br[30] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_33 
+ bl[31] br[31] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_34 
+ bl[32] br[32] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_35 
+ bl[33] br[33] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_36 
+ bl[34] br[34] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_37 
+ bl[35] br[35] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_38 
+ bl[36] br[36] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_39 
+ bl[37] br[37] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_40 
+ bl[38] br[38] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_41 
+ bl[39] br[39] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_42 
+ bl[40] br[40] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_43 
+ bl[41] br[41] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_44 
+ bl[42] br[42] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_45 
+ bl[43] br[43] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_46 
+ bl[44] br[44] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_47 
+ bl[45] br[45] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_48 
+ bl[46] br[46] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_49 
+ bl[47] br[47] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_50 
+ bl[48] br[48] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_51 
+ bl[49] br[49] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_52 
+ bl[50] br[50] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_53 
+ bl[51] br[51] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_54 
+ bl[52] br[52] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_55 
+ bl[53] br[53] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_56 
+ bl[54] br[54] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_57 
+ bl[55] br[55] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_58 
+ bl[56] br[56] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_59 
+ bl[57] br[57] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_60 
+ bl[58] br[58] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_61 
+ bl[59] br[59] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_62 
+ bl[60] br[60] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_63 
+ bl[61] br[61] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_64 
+ bl[62] br[62] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_65 
+ bl[63] br[63] vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_66 
+ vdd vdd vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_508_67 
+ vdd vdd vdd vss wl[506] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_0 
+ vdd vdd vss vdd vpb vnb wl[507] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_509_1 
+ rbl rbr vss vdd vpb vnb wl[507] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_509_2 
+ bl[0] br[0] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_3 
+ bl[1] br[1] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_4 
+ bl[2] br[2] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_5 
+ bl[3] br[3] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_6 
+ bl[4] br[4] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_7 
+ bl[5] br[5] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_8 
+ bl[6] br[6] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_9 
+ bl[7] br[7] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_10 
+ bl[8] br[8] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_11 
+ bl[9] br[9] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_12 
+ bl[10] br[10] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_13 
+ bl[11] br[11] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_14 
+ bl[12] br[12] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_15 
+ bl[13] br[13] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_16 
+ bl[14] br[14] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_17 
+ bl[15] br[15] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_18 
+ bl[16] br[16] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_19 
+ bl[17] br[17] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_20 
+ bl[18] br[18] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_21 
+ bl[19] br[19] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_22 
+ bl[20] br[20] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_23 
+ bl[21] br[21] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_24 
+ bl[22] br[22] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_25 
+ bl[23] br[23] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_26 
+ bl[24] br[24] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_27 
+ bl[25] br[25] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_28 
+ bl[26] br[26] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_29 
+ bl[27] br[27] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_30 
+ bl[28] br[28] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_31 
+ bl[29] br[29] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_32 
+ bl[30] br[30] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_33 
+ bl[31] br[31] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_34 
+ bl[32] br[32] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_35 
+ bl[33] br[33] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_36 
+ bl[34] br[34] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_37 
+ bl[35] br[35] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_38 
+ bl[36] br[36] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_39 
+ bl[37] br[37] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_40 
+ bl[38] br[38] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_41 
+ bl[39] br[39] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_42 
+ bl[40] br[40] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_43 
+ bl[41] br[41] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_44 
+ bl[42] br[42] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_45 
+ bl[43] br[43] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_46 
+ bl[44] br[44] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_47 
+ bl[45] br[45] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_48 
+ bl[46] br[46] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_49 
+ bl[47] br[47] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_50 
+ bl[48] br[48] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_51 
+ bl[49] br[49] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_52 
+ bl[50] br[50] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_53 
+ bl[51] br[51] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_54 
+ bl[52] br[52] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_55 
+ bl[53] br[53] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_56 
+ bl[54] br[54] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_57 
+ bl[55] br[55] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_58 
+ bl[56] br[56] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_59 
+ bl[57] br[57] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_60 
+ bl[58] br[58] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_61 
+ bl[59] br[59] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_62 
+ bl[60] br[60] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_63 
+ bl[61] br[61] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_64 
+ bl[62] br[62] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_65 
+ bl[63] br[63] vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_66 
+ vdd vdd vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_509_67 
+ vdd vdd vdd vss wl[507] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_0 
+ vdd vdd vss vdd vpb vnb wl[508] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_510_1 
+ rbl rbr vss vdd vpb vnb wl[508] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_510_2 
+ bl[0] br[0] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_3 
+ bl[1] br[1] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_4 
+ bl[2] br[2] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_5 
+ bl[3] br[3] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_6 
+ bl[4] br[4] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_7 
+ bl[5] br[5] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_8 
+ bl[6] br[6] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_9 
+ bl[7] br[7] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_10 
+ bl[8] br[8] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_11 
+ bl[9] br[9] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_12 
+ bl[10] br[10] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_13 
+ bl[11] br[11] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_14 
+ bl[12] br[12] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_15 
+ bl[13] br[13] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_16 
+ bl[14] br[14] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_17 
+ bl[15] br[15] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_18 
+ bl[16] br[16] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_19 
+ bl[17] br[17] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_20 
+ bl[18] br[18] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_21 
+ bl[19] br[19] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_22 
+ bl[20] br[20] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_23 
+ bl[21] br[21] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_24 
+ bl[22] br[22] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_25 
+ bl[23] br[23] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_26 
+ bl[24] br[24] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_27 
+ bl[25] br[25] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_28 
+ bl[26] br[26] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_29 
+ bl[27] br[27] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_30 
+ bl[28] br[28] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_31 
+ bl[29] br[29] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_32 
+ bl[30] br[30] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_33 
+ bl[31] br[31] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_34 
+ bl[32] br[32] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_35 
+ bl[33] br[33] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_36 
+ bl[34] br[34] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_37 
+ bl[35] br[35] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_38 
+ bl[36] br[36] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_39 
+ bl[37] br[37] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_40 
+ bl[38] br[38] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_41 
+ bl[39] br[39] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_42 
+ bl[40] br[40] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_43 
+ bl[41] br[41] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_44 
+ bl[42] br[42] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_45 
+ bl[43] br[43] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_46 
+ bl[44] br[44] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_47 
+ bl[45] br[45] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_48 
+ bl[46] br[46] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_49 
+ bl[47] br[47] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_50 
+ bl[48] br[48] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_51 
+ bl[49] br[49] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_52 
+ bl[50] br[50] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_53 
+ bl[51] br[51] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_54 
+ bl[52] br[52] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_55 
+ bl[53] br[53] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_56 
+ bl[54] br[54] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_57 
+ bl[55] br[55] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_58 
+ bl[56] br[56] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_59 
+ bl[57] br[57] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_60 
+ bl[58] br[58] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_61 
+ bl[59] br[59] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_62 
+ bl[60] br[60] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_63 
+ bl[61] br[61] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_64 
+ bl[62] br[62] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_65 
+ bl[63] br[63] vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_66 
+ vdd vdd vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_510_67 
+ vdd vdd vdd vss wl[508] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_0 
+ vdd vdd vss vdd vpb vnb wl[509] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_511_1 
+ rbl rbr vss vdd vpb vnb wl[509] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_511_2 
+ bl[0] br[0] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_3 
+ bl[1] br[1] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_4 
+ bl[2] br[2] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_5 
+ bl[3] br[3] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_6 
+ bl[4] br[4] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_7 
+ bl[5] br[5] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_8 
+ bl[6] br[6] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_9 
+ bl[7] br[7] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_10 
+ bl[8] br[8] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_11 
+ bl[9] br[9] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_12 
+ bl[10] br[10] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_13 
+ bl[11] br[11] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_14 
+ bl[12] br[12] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_15 
+ bl[13] br[13] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_16 
+ bl[14] br[14] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_17 
+ bl[15] br[15] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_18 
+ bl[16] br[16] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_19 
+ bl[17] br[17] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_20 
+ bl[18] br[18] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_21 
+ bl[19] br[19] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_22 
+ bl[20] br[20] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_23 
+ bl[21] br[21] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_24 
+ bl[22] br[22] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_25 
+ bl[23] br[23] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_26 
+ bl[24] br[24] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_27 
+ bl[25] br[25] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_28 
+ bl[26] br[26] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_29 
+ bl[27] br[27] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_30 
+ bl[28] br[28] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_31 
+ bl[29] br[29] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_32 
+ bl[30] br[30] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_33 
+ bl[31] br[31] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_34 
+ bl[32] br[32] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_35 
+ bl[33] br[33] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_36 
+ bl[34] br[34] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_37 
+ bl[35] br[35] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_38 
+ bl[36] br[36] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_39 
+ bl[37] br[37] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_40 
+ bl[38] br[38] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_41 
+ bl[39] br[39] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_42 
+ bl[40] br[40] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_43 
+ bl[41] br[41] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_44 
+ bl[42] br[42] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_45 
+ bl[43] br[43] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_46 
+ bl[44] br[44] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_47 
+ bl[45] br[45] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_48 
+ bl[46] br[46] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_49 
+ bl[47] br[47] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_50 
+ bl[48] br[48] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_51 
+ bl[49] br[49] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_52 
+ bl[50] br[50] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_53 
+ bl[51] br[51] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_54 
+ bl[52] br[52] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_55 
+ bl[53] br[53] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_56 
+ bl[54] br[54] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_57 
+ bl[55] br[55] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_58 
+ bl[56] br[56] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_59 
+ bl[57] br[57] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_60 
+ bl[58] br[58] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_61 
+ bl[59] br[59] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_62 
+ bl[60] br[60] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_63 
+ bl[61] br[61] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_64 
+ bl[62] br[62] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_65 
+ bl[63] br[63] vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_66 
+ vdd vdd vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_511_67 
+ vdd vdd vdd vss wl[509] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_0 
+ vdd vdd vss vdd vpb vnb wl[510] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_512_1 
+ rbl rbr vss vdd vpb vnb wl[510] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_512_2 
+ bl[0] br[0] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_3 
+ bl[1] br[1] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_4 
+ bl[2] br[2] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_5 
+ bl[3] br[3] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_6 
+ bl[4] br[4] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_7 
+ bl[5] br[5] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_8 
+ bl[6] br[6] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_9 
+ bl[7] br[7] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_10 
+ bl[8] br[8] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_11 
+ bl[9] br[9] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_12 
+ bl[10] br[10] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_13 
+ bl[11] br[11] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_14 
+ bl[12] br[12] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_15 
+ bl[13] br[13] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_16 
+ bl[14] br[14] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_17 
+ bl[15] br[15] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_18 
+ bl[16] br[16] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_19 
+ bl[17] br[17] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_20 
+ bl[18] br[18] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_21 
+ bl[19] br[19] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_22 
+ bl[20] br[20] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_23 
+ bl[21] br[21] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_24 
+ bl[22] br[22] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_25 
+ bl[23] br[23] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_26 
+ bl[24] br[24] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_27 
+ bl[25] br[25] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_28 
+ bl[26] br[26] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_29 
+ bl[27] br[27] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_30 
+ bl[28] br[28] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_31 
+ bl[29] br[29] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_32 
+ bl[30] br[30] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_33 
+ bl[31] br[31] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_34 
+ bl[32] br[32] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_35 
+ bl[33] br[33] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_36 
+ bl[34] br[34] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_37 
+ bl[35] br[35] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_38 
+ bl[36] br[36] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_39 
+ bl[37] br[37] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_40 
+ bl[38] br[38] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_41 
+ bl[39] br[39] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_42 
+ bl[40] br[40] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_43 
+ bl[41] br[41] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_44 
+ bl[42] br[42] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_45 
+ bl[43] br[43] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_46 
+ bl[44] br[44] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_47 
+ bl[45] br[45] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_48 
+ bl[46] br[46] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_49 
+ bl[47] br[47] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_50 
+ bl[48] br[48] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_51 
+ bl[49] br[49] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_52 
+ bl[50] br[50] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_53 
+ bl[51] br[51] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_54 
+ bl[52] br[52] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_55 
+ bl[53] br[53] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_56 
+ bl[54] br[54] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_57 
+ bl[55] br[55] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_58 
+ bl[56] br[56] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_59 
+ bl[57] br[57] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_60 
+ bl[58] br[58] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_61 
+ bl[59] br[59] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_62 
+ bl[60] br[60] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_63 
+ bl[61] br[61] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_64 
+ bl[62] br[62] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_65 
+ bl[63] br[63] vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_66 
+ vdd vdd vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_512_67 
+ vdd vdd vdd vss wl[510] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_0 
+ vdd vdd vss vdd vpb vnb wl[511] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_513_1 
+ rbl rbr vss vdd vpb vnb wl[511] 
+ sram_sp_cell_replica 
* No parameters

xbitcell_513_2 
+ bl[0] br[0] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_3 
+ bl[1] br[1] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_4 
+ bl[2] br[2] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_5 
+ bl[3] br[3] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_6 
+ bl[4] br[4] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_7 
+ bl[5] br[5] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_8 
+ bl[6] br[6] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_9 
+ bl[7] br[7] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_10 
+ bl[8] br[8] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_11 
+ bl[9] br[9] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_12 
+ bl[10] br[10] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_13 
+ bl[11] br[11] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_14 
+ bl[12] br[12] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_15 
+ bl[13] br[13] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_16 
+ bl[14] br[14] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_17 
+ bl[15] br[15] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_18 
+ bl[16] br[16] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_19 
+ bl[17] br[17] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_20 
+ bl[18] br[18] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_21 
+ bl[19] br[19] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_22 
+ bl[20] br[20] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_23 
+ bl[21] br[21] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_24 
+ bl[22] br[22] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_25 
+ bl[23] br[23] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_26 
+ bl[24] br[24] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_27 
+ bl[25] br[25] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_28 
+ bl[26] br[26] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_29 
+ bl[27] br[27] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_30 
+ bl[28] br[28] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_31 
+ bl[29] br[29] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_32 
+ bl[30] br[30] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_33 
+ bl[31] br[31] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_34 
+ bl[32] br[32] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_35 
+ bl[33] br[33] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_36 
+ bl[34] br[34] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_37 
+ bl[35] br[35] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_38 
+ bl[36] br[36] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_39 
+ bl[37] br[37] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_40 
+ bl[38] br[38] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_41 
+ bl[39] br[39] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_42 
+ bl[40] br[40] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_43 
+ bl[41] br[41] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_44 
+ bl[42] br[42] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_45 
+ bl[43] br[43] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_46 
+ bl[44] br[44] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_47 
+ bl[45] br[45] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_48 
+ bl[46] br[46] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_49 
+ bl[47] br[47] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_50 
+ bl[48] br[48] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_51 
+ bl[49] br[49] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_52 
+ bl[50] br[50] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_53 
+ bl[51] br[51] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_54 
+ bl[52] br[52] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_55 
+ bl[53] br[53] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_56 
+ bl[54] br[54] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_57 
+ bl[55] br[55] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_58 
+ bl[56] br[56] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_59 
+ bl[57] br[57] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_60 
+ bl[58] br[58] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_61 
+ bl[59] br[59] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_62 
+ bl[60] br[60] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_63 
+ bl[61] br[61] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_64 
+ bl[62] br[62] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_65 
+ bl[63] br[63] vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_66 
+ vdd vdd vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_513_67 
+ vdd vdd vdd vss wl[511] vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_66 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_514_67 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_0 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_1 
+ rbl rbr vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_2 
+ bl[0] br[0] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_3 
+ bl[1] br[1] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_4 
+ bl[2] br[2] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_5 
+ bl[3] br[3] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_6 
+ bl[4] br[4] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_7 
+ bl[5] br[5] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_8 
+ bl[6] br[6] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_9 
+ bl[7] br[7] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_10 
+ bl[8] br[8] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_11 
+ bl[9] br[9] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_12 
+ bl[10] br[10] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_13 
+ bl[11] br[11] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_14 
+ bl[12] br[12] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_15 
+ bl[13] br[13] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_16 
+ bl[14] br[14] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_17 
+ bl[15] br[15] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_18 
+ bl[16] br[16] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_19 
+ bl[17] br[17] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_20 
+ bl[18] br[18] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_21 
+ bl[19] br[19] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_22 
+ bl[20] br[20] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_23 
+ bl[21] br[21] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_24 
+ bl[22] br[22] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_25 
+ bl[23] br[23] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_26 
+ bl[24] br[24] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_27 
+ bl[25] br[25] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_28 
+ bl[26] br[26] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_29 
+ bl[27] br[27] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_30 
+ bl[28] br[28] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_31 
+ bl[29] br[29] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_32 
+ bl[30] br[30] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_33 
+ bl[31] br[31] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_34 
+ bl[32] br[32] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_35 
+ bl[33] br[33] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_36 
+ bl[34] br[34] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_37 
+ bl[35] br[35] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_38 
+ bl[36] br[36] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_39 
+ bl[37] br[37] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_40 
+ bl[38] br[38] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_41 
+ bl[39] br[39] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_42 
+ bl[40] br[40] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_43 
+ bl[41] br[41] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_44 
+ bl[42] br[42] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_45 
+ bl[43] br[43] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_46 
+ bl[44] br[44] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_47 
+ bl[45] br[45] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_48 
+ bl[46] br[46] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_49 
+ bl[47] br[47] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_50 
+ bl[48] br[48] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_51 
+ bl[49] br[49] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_52 
+ bl[50] br[50] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_53 
+ bl[51] br[51] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_54 
+ bl[52] br[52] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_55 
+ bl[53] br[53] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_56 
+ bl[54] br[54] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_57 
+ bl[55] br[55] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_58 
+ bl[56] br[56] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_59 
+ bl[57] br[57] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_60 
+ bl[58] br[58] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_61 
+ bl[59] br[59] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_62 
+ bl[60] br[60] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_63 
+ bl[61] br[61] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_64 
+ bl[62] br[62] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_65 
+ bl[63] br[63] vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_66 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xbitcell_515_67 
+ vdd vdd vdd vss vss vnb vpb 
+ sram_sp_cell 
* No parameters

xcolend_0_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_0_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_1_bot 
+ rbr vdd vss rbl vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_1_top 
+ rbr vdd vss rbl vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_2_bot 
+ br[0] vdd vss bl[0] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_2_top 
+ br[0] vdd vss bl[0] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_3_bot 
+ br[1] vdd vss bl[1] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_3_top 
+ br[1] vdd vss bl[1] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_4_bot 
+ br[2] vdd vss bl[2] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_4_top 
+ br[2] vdd vss bl[2] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_5_bot 
+ br[3] vdd vss bl[3] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_5_top 
+ br[3] vdd vss bl[3] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_6_bot 
+ br[4] vdd vss bl[4] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_6_top 
+ br[4] vdd vss bl[4] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_7_bot 
+ br[5] vdd vss bl[5] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_7_top 
+ br[5] vdd vss bl[5] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_8_bot 
+ br[6] vdd vss bl[6] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_8_top 
+ br[6] vdd vss bl[6] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_9_bot 
+ br[7] vdd vss bl[7] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_9_top 
+ br[7] vdd vss bl[7] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_10_bot 
+ br[8] vdd vss bl[8] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_10_top 
+ br[8] vdd vss bl[8] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_11_bot 
+ br[9] vdd vss bl[9] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_11_top 
+ br[9] vdd vss bl[9] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_12_bot 
+ br[10] vdd vss bl[10] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_12_top 
+ br[10] vdd vss bl[10] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_13_bot 
+ br[11] vdd vss bl[11] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_13_top 
+ br[11] vdd vss bl[11] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_14_bot 
+ br[12] vdd vss bl[12] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_14_top 
+ br[12] vdd vss bl[12] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_15_bot 
+ br[13] vdd vss bl[13] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_15_top 
+ br[13] vdd vss bl[13] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_16_bot 
+ br[14] vdd vss bl[14] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_16_top 
+ br[14] vdd vss bl[14] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_17_bot 
+ br[15] vdd vss bl[15] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_17_top 
+ br[15] vdd vss bl[15] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_18_bot 
+ br[16] vdd vss bl[16] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_18_top 
+ br[16] vdd vss bl[16] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_19_bot 
+ br[17] vdd vss bl[17] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_19_top 
+ br[17] vdd vss bl[17] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_20_bot 
+ br[18] vdd vss bl[18] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_20_top 
+ br[18] vdd vss bl[18] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_21_bot 
+ br[19] vdd vss bl[19] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_21_top 
+ br[19] vdd vss bl[19] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_22_bot 
+ br[20] vdd vss bl[20] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_22_top 
+ br[20] vdd vss bl[20] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_23_bot 
+ br[21] vdd vss bl[21] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_23_top 
+ br[21] vdd vss bl[21] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_24_bot 
+ br[22] vdd vss bl[22] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_24_top 
+ br[22] vdd vss bl[22] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_25_bot 
+ br[23] vdd vss bl[23] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_25_top 
+ br[23] vdd vss bl[23] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_26_bot 
+ br[24] vdd vss bl[24] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_26_top 
+ br[24] vdd vss bl[24] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_27_bot 
+ br[25] vdd vss bl[25] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_27_top 
+ br[25] vdd vss bl[25] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_28_bot 
+ br[26] vdd vss bl[26] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_28_top 
+ br[26] vdd vss bl[26] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_29_bot 
+ br[27] vdd vss bl[27] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_29_top 
+ br[27] vdd vss bl[27] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_30_bot 
+ br[28] vdd vss bl[28] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_30_top 
+ br[28] vdd vss bl[28] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_31_bot 
+ br[29] vdd vss bl[29] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_31_top 
+ br[29] vdd vss bl[29] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_32_bot 
+ br[30] vdd vss bl[30] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_32_top 
+ br[30] vdd vss bl[30] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_33_bot 
+ br[31] vdd vss bl[31] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_33_top 
+ br[31] vdd vss bl[31] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_34_bot 
+ br[32] vdd vss bl[32] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_34_top 
+ br[32] vdd vss bl[32] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_35_bot 
+ br[33] vdd vss bl[33] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_35_top 
+ br[33] vdd vss bl[33] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_36_bot 
+ br[34] vdd vss bl[34] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_36_top 
+ br[34] vdd vss bl[34] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_37_bot 
+ br[35] vdd vss bl[35] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_37_top 
+ br[35] vdd vss bl[35] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_38_bot 
+ br[36] vdd vss bl[36] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_38_top 
+ br[36] vdd vss bl[36] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_39_bot 
+ br[37] vdd vss bl[37] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_39_top 
+ br[37] vdd vss bl[37] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_40_bot 
+ br[38] vdd vss bl[38] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_40_top 
+ br[38] vdd vss bl[38] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_41_bot 
+ br[39] vdd vss bl[39] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_41_top 
+ br[39] vdd vss bl[39] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_42_bot 
+ br[40] vdd vss bl[40] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_42_top 
+ br[40] vdd vss bl[40] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_43_bot 
+ br[41] vdd vss bl[41] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_43_top 
+ br[41] vdd vss bl[41] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_44_bot 
+ br[42] vdd vss bl[42] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_44_top 
+ br[42] vdd vss bl[42] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_45_bot 
+ br[43] vdd vss bl[43] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_45_top 
+ br[43] vdd vss bl[43] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_46_bot 
+ br[44] vdd vss bl[44] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_46_top 
+ br[44] vdd vss bl[44] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_47_bot 
+ br[45] vdd vss bl[45] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_47_top 
+ br[45] vdd vss bl[45] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_48_bot 
+ br[46] vdd vss bl[46] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_48_top 
+ br[46] vdd vss bl[46] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_49_bot 
+ br[47] vdd vss bl[47] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_49_top 
+ br[47] vdd vss bl[47] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_50_bot 
+ br[48] vdd vss bl[48] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_50_top 
+ br[48] vdd vss bl[48] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_51_bot 
+ br[49] vdd vss bl[49] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_51_top 
+ br[49] vdd vss bl[49] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_52_bot 
+ br[50] vdd vss bl[50] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_52_top 
+ br[50] vdd vss bl[50] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_53_bot 
+ br[51] vdd vss bl[51] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_53_top 
+ br[51] vdd vss bl[51] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_54_bot 
+ br[52] vdd vss bl[52] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_54_top 
+ br[52] vdd vss bl[52] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_55_bot 
+ br[53] vdd vss bl[53] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_55_top 
+ br[53] vdd vss bl[53] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_56_bot 
+ br[54] vdd vss bl[54] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_56_top 
+ br[54] vdd vss bl[54] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_57_bot 
+ br[55] vdd vss bl[55] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_57_top 
+ br[55] vdd vss bl[55] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_58_bot 
+ br[56] vdd vss bl[56] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_58_top 
+ br[56] vdd vss bl[56] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_59_bot 
+ br[57] vdd vss bl[57] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_59_top 
+ br[57] vdd vss bl[57] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_60_bot 
+ br[58] vdd vss bl[58] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_60_top 
+ br[58] vdd vss bl[58] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_61_bot 
+ br[59] vdd vss bl[59] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_61_top 
+ br[59] vdd vss bl[59] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_62_bot 
+ br[60] vdd vss bl[60] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_62_top 
+ br[60] vdd vss bl[60] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_63_bot 
+ br[61] vdd vss bl[61] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_63_top 
+ br[61] vdd vss bl[61] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_64_bot 
+ br[62] vdd vss bl[62] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_64_top 
+ br[62] vdd vss bl[62] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_65_bot 
+ br[63] vdd vss bl[63] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_65_top 
+ br[63] vdd vss bl[63] vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_66_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_66_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_67_bot 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

xcolend_67_top 
+ vdd vdd vss vdd vnb vpb 
+ sky130_fd_bd_sram__sram_sp_colend 
* No parameters

.ENDS

.SUBCKT precharge 
+ vdd bl br en_b 

xbl_pull_up 
+ bl en_b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

xbr_pull_up 
+ br en_b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

xequalizer 
+ bl en_b br vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.0' l='0.15' 

.ENDS

.SUBCKT precharge_array 
+ vdd en_b bl[64] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[64] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] 

xprecharge_0 
+ vdd bl[0] br[0] en_b 
+ precharge 
* No parameters

xprecharge_1 
+ vdd bl[1] br[1] en_b 
+ precharge 
* No parameters

xprecharge_2 
+ vdd bl[2] br[2] en_b 
+ precharge 
* No parameters

xprecharge_3 
+ vdd bl[3] br[3] en_b 
+ precharge 
* No parameters

xprecharge_4 
+ vdd bl[4] br[4] en_b 
+ precharge 
* No parameters

xprecharge_5 
+ vdd bl[5] br[5] en_b 
+ precharge 
* No parameters

xprecharge_6 
+ vdd bl[6] br[6] en_b 
+ precharge 
* No parameters

xprecharge_7 
+ vdd bl[7] br[7] en_b 
+ precharge 
* No parameters

xprecharge_8 
+ vdd bl[8] br[8] en_b 
+ precharge 
* No parameters

xprecharge_9 
+ vdd bl[9] br[9] en_b 
+ precharge 
* No parameters

xprecharge_10 
+ vdd bl[10] br[10] en_b 
+ precharge 
* No parameters

xprecharge_11 
+ vdd bl[11] br[11] en_b 
+ precharge 
* No parameters

xprecharge_12 
+ vdd bl[12] br[12] en_b 
+ precharge 
* No parameters

xprecharge_13 
+ vdd bl[13] br[13] en_b 
+ precharge 
* No parameters

xprecharge_14 
+ vdd bl[14] br[14] en_b 
+ precharge 
* No parameters

xprecharge_15 
+ vdd bl[15] br[15] en_b 
+ precharge 
* No parameters

xprecharge_16 
+ vdd bl[16] br[16] en_b 
+ precharge 
* No parameters

xprecharge_17 
+ vdd bl[17] br[17] en_b 
+ precharge 
* No parameters

xprecharge_18 
+ vdd bl[18] br[18] en_b 
+ precharge 
* No parameters

xprecharge_19 
+ vdd bl[19] br[19] en_b 
+ precharge 
* No parameters

xprecharge_20 
+ vdd bl[20] br[20] en_b 
+ precharge 
* No parameters

xprecharge_21 
+ vdd bl[21] br[21] en_b 
+ precharge 
* No parameters

xprecharge_22 
+ vdd bl[22] br[22] en_b 
+ precharge 
* No parameters

xprecharge_23 
+ vdd bl[23] br[23] en_b 
+ precharge 
* No parameters

xprecharge_24 
+ vdd bl[24] br[24] en_b 
+ precharge 
* No parameters

xprecharge_25 
+ vdd bl[25] br[25] en_b 
+ precharge 
* No parameters

xprecharge_26 
+ vdd bl[26] br[26] en_b 
+ precharge 
* No parameters

xprecharge_27 
+ vdd bl[27] br[27] en_b 
+ precharge 
* No parameters

xprecharge_28 
+ vdd bl[28] br[28] en_b 
+ precharge 
* No parameters

xprecharge_29 
+ vdd bl[29] br[29] en_b 
+ precharge 
* No parameters

xprecharge_30 
+ vdd bl[30] br[30] en_b 
+ precharge 
* No parameters

xprecharge_31 
+ vdd bl[31] br[31] en_b 
+ precharge 
* No parameters

xprecharge_32 
+ vdd bl[32] br[32] en_b 
+ precharge 
* No parameters

xprecharge_33 
+ vdd bl[33] br[33] en_b 
+ precharge 
* No parameters

xprecharge_34 
+ vdd bl[34] br[34] en_b 
+ precharge 
* No parameters

xprecharge_35 
+ vdd bl[35] br[35] en_b 
+ precharge 
* No parameters

xprecharge_36 
+ vdd bl[36] br[36] en_b 
+ precharge 
* No parameters

xprecharge_37 
+ vdd bl[37] br[37] en_b 
+ precharge 
* No parameters

xprecharge_38 
+ vdd bl[38] br[38] en_b 
+ precharge 
* No parameters

xprecharge_39 
+ vdd bl[39] br[39] en_b 
+ precharge 
* No parameters

xprecharge_40 
+ vdd bl[40] br[40] en_b 
+ precharge 
* No parameters

xprecharge_41 
+ vdd bl[41] br[41] en_b 
+ precharge 
* No parameters

xprecharge_42 
+ vdd bl[42] br[42] en_b 
+ precharge 
* No parameters

xprecharge_43 
+ vdd bl[43] br[43] en_b 
+ precharge 
* No parameters

xprecharge_44 
+ vdd bl[44] br[44] en_b 
+ precharge 
* No parameters

xprecharge_45 
+ vdd bl[45] br[45] en_b 
+ precharge 
* No parameters

xprecharge_46 
+ vdd bl[46] br[46] en_b 
+ precharge 
* No parameters

xprecharge_47 
+ vdd bl[47] br[47] en_b 
+ precharge 
* No parameters

xprecharge_48 
+ vdd bl[48] br[48] en_b 
+ precharge 
* No parameters

xprecharge_49 
+ vdd bl[49] br[49] en_b 
+ precharge 
* No parameters

xprecharge_50 
+ vdd bl[50] br[50] en_b 
+ precharge 
* No parameters

xprecharge_51 
+ vdd bl[51] br[51] en_b 
+ precharge 
* No parameters

xprecharge_52 
+ vdd bl[52] br[52] en_b 
+ precharge 
* No parameters

xprecharge_53 
+ vdd bl[53] br[53] en_b 
+ precharge 
* No parameters

xprecharge_54 
+ vdd bl[54] br[54] en_b 
+ precharge 
* No parameters

xprecharge_55 
+ vdd bl[55] br[55] en_b 
+ precharge 
* No parameters

xprecharge_56 
+ vdd bl[56] br[56] en_b 
+ precharge 
* No parameters

xprecharge_57 
+ vdd bl[57] br[57] en_b 
+ precharge 
* No parameters

xprecharge_58 
+ vdd bl[58] br[58] en_b 
+ precharge 
* No parameters

xprecharge_59 
+ vdd bl[59] br[59] en_b 
+ precharge 
* No parameters

xprecharge_60 
+ vdd bl[60] br[60] en_b 
+ precharge 
* No parameters

xprecharge_61 
+ vdd bl[61] br[61] en_b 
+ precharge 
* No parameters

xprecharge_62 
+ vdd bl[62] br[62] en_b 
+ precharge 
* No parameters

xprecharge_63 
+ vdd bl[63] br[63] en_b 
+ precharge 
* No parameters

xprecharge_64 
+ vdd bl[64] br[64] en_b 
+ precharge 
* No parameters

.ENDS

.SUBCKT read_mux 
+ sel_b bl br bl_out br_out vdd 

xMBL 
+ bl_out sel_b bl vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.2' l='0.15' 

xMBR 
+ br_out sel_b br vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.2' l='0.15' 

.ENDS

.SUBCKT read_mux_array 
+ sel_b[7] sel_b[6] sel_b[5] sel_b[4] sel_b[3] sel_b[2] sel_b[1] sel_b[0] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] bl_out[7] bl_out[6] bl_out[5] bl_out[4] bl_out[3] bl_out[2] bl_out[1] bl_out[0] br_out[7] br_out[6] br_out[5] br_out[4] br_out[3] br_out[2] br_out[1] br_out[0] vdd 

xmux_0 
+ sel_b[0] bl[0] br[0] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_1 
+ sel_b[1] bl[1] br[1] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_2 
+ sel_b[2] bl[2] br[2] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_3 
+ sel_b[3] bl[3] br[3] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_4 
+ sel_b[4] bl[4] br[4] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_5 
+ sel_b[5] bl[5] br[5] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_6 
+ sel_b[6] bl[6] br[6] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_7 
+ sel_b[7] bl[7] br[7] bl_out[0] br_out[0] vdd 
+ read_mux 
* No parameters

xmux_8 
+ sel_b[0] bl[8] br[8] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_9 
+ sel_b[1] bl[9] br[9] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_10 
+ sel_b[2] bl[10] br[10] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_11 
+ sel_b[3] bl[11] br[11] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_12 
+ sel_b[4] bl[12] br[12] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_13 
+ sel_b[5] bl[13] br[13] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_14 
+ sel_b[6] bl[14] br[14] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_15 
+ sel_b[7] bl[15] br[15] bl_out[1] br_out[1] vdd 
+ read_mux 
* No parameters

xmux_16 
+ sel_b[0] bl[16] br[16] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_17 
+ sel_b[1] bl[17] br[17] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_18 
+ sel_b[2] bl[18] br[18] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_19 
+ sel_b[3] bl[19] br[19] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_20 
+ sel_b[4] bl[20] br[20] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_21 
+ sel_b[5] bl[21] br[21] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_22 
+ sel_b[6] bl[22] br[22] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_23 
+ sel_b[7] bl[23] br[23] bl_out[2] br_out[2] vdd 
+ read_mux 
* No parameters

xmux_24 
+ sel_b[0] bl[24] br[24] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_25 
+ sel_b[1] bl[25] br[25] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_26 
+ sel_b[2] bl[26] br[26] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_27 
+ sel_b[3] bl[27] br[27] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_28 
+ sel_b[4] bl[28] br[28] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_29 
+ sel_b[5] bl[29] br[29] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_30 
+ sel_b[6] bl[30] br[30] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_31 
+ sel_b[7] bl[31] br[31] bl_out[3] br_out[3] vdd 
+ read_mux 
* No parameters

xmux_32 
+ sel_b[0] bl[32] br[32] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_33 
+ sel_b[1] bl[33] br[33] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_34 
+ sel_b[2] bl[34] br[34] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_35 
+ sel_b[3] bl[35] br[35] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_36 
+ sel_b[4] bl[36] br[36] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_37 
+ sel_b[5] bl[37] br[37] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_38 
+ sel_b[6] bl[38] br[38] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_39 
+ sel_b[7] bl[39] br[39] bl_out[4] br_out[4] vdd 
+ read_mux 
* No parameters

xmux_40 
+ sel_b[0] bl[40] br[40] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_41 
+ sel_b[1] bl[41] br[41] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_42 
+ sel_b[2] bl[42] br[42] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_43 
+ sel_b[3] bl[43] br[43] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_44 
+ sel_b[4] bl[44] br[44] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_45 
+ sel_b[5] bl[45] br[45] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_46 
+ sel_b[6] bl[46] br[46] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_47 
+ sel_b[7] bl[47] br[47] bl_out[5] br_out[5] vdd 
+ read_mux 
* No parameters

xmux_48 
+ sel_b[0] bl[48] br[48] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_49 
+ sel_b[1] bl[49] br[49] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_50 
+ sel_b[2] bl[50] br[50] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_51 
+ sel_b[3] bl[51] br[51] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_52 
+ sel_b[4] bl[52] br[52] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_53 
+ sel_b[5] bl[53] br[53] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_54 
+ sel_b[6] bl[54] br[54] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_55 
+ sel_b[7] bl[55] br[55] bl_out[6] br_out[6] vdd 
+ read_mux 
* No parameters

xmux_56 
+ sel_b[0] bl[56] br[56] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_57 
+ sel_b[1] bl[57] br[57] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_58 
+ sel_b[2] bl[58] br[58] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_59 
+ sel_b[3] bl[59] br[59] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_60 
+ sel_b[4] bl[60] br[60] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_61 
+ sel_b[5] bl[61] br[61] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_62 
+ sel_b[6] bl[62] br[62] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

xmux_63 
+ sel_b[7] bl[63] br[63] bl_out[7] br_out[7] vdd 
+ read_mux 
* No parameters

.ENDS

.SUBCKT write_mux 
+ we data data_b bl br vss 

xMMUXBR 
+ br data x vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMMUXBL 
+ bl data_b x vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMPD 
+ x we vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

.ENDS

.SUBCKT write_mux_array 
+ we[7] we[6] we[5] we[4] we[3] we[2] we[1] we[0] data[7] data[6] data[5] data[4] data[3] data[2] data[1] data[0] data_b[7] data_b[6] data_b[5] data_b[4] data_b[3] data_b[2] data_b[1] data_b[0] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] vss 

xmux_0 
+ we[0] data[0] data_b[0] bl[0] br[0] vss 
+ write_mux 
* No parameters

xmux_1 
+ we[1] data[0] data_b[0] bl[1] br[1] vss 
+ write_mux 
* No parameters

xmux_2 
+ we[2] data[0] data_b[0] bl[2] br[2] vss 
+ write_mux 
* No parameters

xmux_3 
+ we[3] data[0] data_b[0] bl[3] br[3] vss 
+ write_mux 
* No parameters

xmux_4 
+ we[4] data[0] data_b[0] bl[4] br[4] vss 
+ write_mux 
* No parameters

xmux_5 
+ we[5] data[0] data_b[0] bl[5] br[5] vss 
+ write_mux 
* No parameters

xmux_6 
+ we[6] data[0] data_b[0] bl[6] br[6] vss 
+ write_mux 
* No parameters

xmux_7 
+ we[7] data[0] data_b[0] bl[7] br[7] vss 
+ write_mux 
* No parameters

xmux_8 
+ we[0] data[1] data_b[1] bl[8] br[8] vss 
+ write_mux 
* No parameters

xmux_9 
+ we[1] data[1] data_b[1] bl[9] br[9] vss 
+ write_mux 
* No parameters

xmux_10 
+ we[2] data[1] data_b[1] bl[10] br[10] vss 
+ write_mux 
* No parameters

xmux_11 
+ we[3] data[1] data_b[1] bl[11] br[11] vss 
+ write_mux 
* No parameters

xmux_12 
+ we[4] data[1] data_b[1] bl[12] br[12] vss 
+ write_mux 
* No parameters

xmux_13 
+ we[5] data[1] data_b[1] bl[13] br[13] vss 
+ write_mux 
* No parameters

xmux_14 
+ we[6] data[1] data_b[1] bl[14] br[14] vss 
+ write_mux 
* No parameters

xmux_15 
+ we[7] data[1] data_b[1] bl[15] br[15] vss 
+ write_mux 
* No parameters

xmux_16 
+ we[0] data[2] data_b[2] bl[16] br[16] vss 
+ write_mux 
* No parameters

xmux_17 
+ we[1] data[2] data_b[2] bl[17] br[17] vss 
+ write_mux 
* No parameters

xmux_18 
+ we[2] data[2] data_b[2] bl[18] br[18] vss 
+ write_mux 
* No parameters

xmux_19 
+ we[3] data[2] data_b[2] bl[19] br[19] vss 
+ write_mux 
* No parameters

xmux_20 
+ we[4] data[2] data_b[2] bl[20] br[20] vss 
+ write_mux 
* No parameters

xmux_21 
+ we[5] data[2] data_b[2] bl[21] br[21] vss 
+ write_mux 
* No parameters

xmux_22 
+ we[6] data[2] data_b[2] bl[22] br[22] vss 
+ write_mux 
* No parameters

xmux_23 
+ we[7] data[2] data_b[2] bl[23] br[23] vss 
+ write_mux 
* No parameters

xmux_24 
+ we[0] data[3] data_b[3] bl[24] br[24] vss 
+ write_mux 
* No parameters

xmux_25 
+ we[1] data[3] data_b[3] bl[25] br[25] vss 
+ write_mux 
* No parameters

xmux_26 
+ we[2] data[3] data_b[3] bl[26] br[26] vss 
+ write_mux 
* No parameters

xmux_27 
+ we[3] data[3] data_b[3] bl[27] br[27] vss 
+ write_mux 
* No parameters

xmux_28 
+ we[4] data[3] data_b[3] bl[28] br[28] vss 
+ write_mux 
* No parameters

xmux_29 
+ we[5] data[3] data_b[3] bl[29] br[29] vss 
+ write_mux 
* No parameters

xmux_30 
+ we[6] data[3] data_b[3] bl[30] br[30] vss 
+ write_mux 
* No parameters

xmux_31 
+ we[7] data[3] data_b[3] bl[31] br[31] vss 
+ write_mux 
* No parameters

xmux_32 
+ we[0] data[4] data_b[4] bl[32] br[32] vss 
+ write_mux 
* No parameters

xmux_33 
+ we[1] data[4] data_b[4] bl[33] br[33] vss 
+ write_mux 
* No parameters

xmux_34 
+ we[2] data[4] data_b[4] bl[34] br[34] vss 
+ write_mux 
* No parameters

xmux_35 
+ we[3] data[4] data_b[4] bl[35] br[35] vss 
+ write_mux 
* No parameters

xmux_36 
+ we[4] data[4] data_b[4] bl[36] br[36] vss 
+ write_mux 
* No parameters

xmux_37 
+ we[5] data[4] data_b[4] bl[37] br[37] vss 
+ write_mux 
* No parameters

xmux_38 
+ we[6] data[4] data_b[4] bl[38] br[38] vss 
+ write_mux 
* No parameters

xmux_39 
+ we[7] data[4] data_b[4] bl[39] br[39] vss 
+ write_mux 
* No parameters

xmux_40 
+ we[0] data[5] data_b[5] bl[40] br[40] vss 
+ write_mux 
* No parameters

xmux_41 
+ we[1] data[5] data_b[5] bl[41] br[41] vss 
+ write_mux 
* No parameters

xmux_42 
+ we[2] data[5] data_b[5] bl[42] br[42] vss 
+ write_mux 
* No parameters

xmux_43 
+ we[3] data[5] data_b[5] bl[43] br[43] vss 
+ write_mux 
* No parameters

xmux_44 
+ we[4] data[5] data_b[5] bl[44] br[44] vss 
+ write_mux 
* No parameters

xmux_45 
+ we[5] data[5] data_b[5] bl[45] br[45] vss 
+ write_mux 
* No parameters

xmux_46 
+ we[6] data[5] data_b[5] bl[46] br[46] vss 
+ write_mux 
* No parameters

xmux_47 
+ we[7] data[5] data_b[5] bl[47] br[47] vss 
+ write_mux 
* No parameters

xmux_48 
+ we[0] data[6] data_b[6] bl[48] br[48] vss 
+ write_mux 
* No parameters

xmux_49 
+ we[1] data[6] data_b[6] bl[49] br[49] vss 
+ write_mux 
* No parameters

xmux_50 
+ we[2] data[6] data_b[6] bl[50] br[50] vss 
+ write_mux 
* No parameters

xmux_51 
+ we[3] data[6] data_b[6] bl[51] br[51] vss 
+ write_mux 
* No parameters

xmux_52 
+ we[4] data[6] data_b[6] bl[52] br[52] vss 
+ write_mux 
* No parameters

xmux_53 
+ we[5] data[6] data_b[6] bl[53] br[53] vss 
+ write_mux 
* No parameters

xmux_54 
+ we[6] data[6] data_b[6] bl[54] br[54] vss 
+ write_mux 
* No parameters

xmux_55 
+ we[7] data[6] data_b[6] bl[55] br[55] vss 
+ write_mux 
* No parameters

xmux_56 
+ we[0] data[7] data_b[7] bl[56] br[56] vss 
+ write_mux 
* No parameters

xmux_57 
+ we[1] data[7] data_b[7] bl[57] br[57] vss 
+ write_mux 
* No parameters

xmux_58 
+ we[2] data[7] data_b[7] bl[58] br[58] vss 
+ write_mux 
* No parameters

xmux_59 
+ we[3] data[7] data_b[7] bl[59] br[59] vss 
+ write_mux 
* No parameters

xmux_60 
+ we[4] data[7] data_b[7] bl[60] br[60] vss 
+ write_mux 
* No parameters

xmux_61 
+ we[5] data[7] data_b[7] bl[61] br[61] vss 
+ write_mux 
* No parameters

xmux_62 
+ we[6] data[7] data_b[7] bl[62] br[62] vss 
+ write_mux 
* No parameters

xmux_63 
+ we[7] data[7] data_b[7] bl[63] br[63] vss 
+ write_mux 
* No parameters

.ENDS

.SUBCKT data_dff_array 
+ vdd vss clk d[7] d[6] d[5] d[4] d[3] d[2] d[1] d[0] q[7] q[6] q[5] q[4] q[3] q[2] q[1] q[0] q_b[7] q_b[6] q_b[5] q_b[4] q_b[3] q_b[2] q_b[1] q_b[0] 

xdff_0 
+ vdd vss clk d[0] q[0] q_b[0] 
+ openram_dff 
* No parameters

xdff_1 
+ vdd vss clk d[1] q[1] q_b[1] 
+ openram_dff 
* No parameters

xdff_2 
+ vdd vss clk d[2] q[2] q_b[2] 
+ openram_dff 
* No parameters

xdff_3 
+ vdd vss clk d[3] q[3] q_b[3] 
+ openram_dff 
* No parameters

xdff_4 
+ vdd vss clk d[4] q[4] q_b[4] 
+ openram_dff 
* No parameters

xdff_5 
+ vdd vss clk d[5] q[5] q_b[5] 
+ openram_dff 
* No parameters

xdff_6 
+ vdd vss clk d[6] q[6] q_b[6] 
+ openram_dff 
* No parameters

xdff_7 
+ vdd vss clk d[7] q[7] q_b[7] 
+ openram_dff 
* No parameters

.ENDS

.SUBCKT addr_dff_array 
+ vdd vss clk d[11] d[10] d[9] d[8] d[7] d[6] d[5] d[4] d[3] d[2] d[1] d[0] q[11] q[10] q[9] q[8] q[7] q[6] q[5] q[4] q[3] q[2] q[1] q[0] q_b[11] q_b[10] q_b[9] q_b[8] q_b[7] q_b[6] q_b[5] q_b[4] q_b[3] q_b[2] q_b[1] q_b[0] 

xdff_0 
+ vdd vss clk d[0] q[0] q_b[0] 
+ openram_dff 
* No parameters

xdff_1 
+ vdd vss clk d[1] q[1] q_b[1] 
+ openram_dff 
* No parameters

xdff_2 
+ vdd vss clk d[2] q[2] q_b[2] 
+ openram_dff 
* No parameters

xdff_3 
+ vdd vss clk d[3] q[3] q_b[3] 
+ openram_dff 
* No parameters

xdff_4 
+ vdd vss clk d[4] q[4] q_b[4] 
+ openram_dff 
* No parameters

xdff_5 
+ vdd vss clk d[5] q[5] q_b[5] 
+ openram_dff 
* No parameters

xdff_6 
+ vdd vss clk d[6] q[6] q_b[6] 
+ openram_dff 
* No parameters

xdff_7 
+ vdd vss clk d[7] q[7] q_b[7] 
+ openram_dff 
* No parameters

xdff_8 
+ vdd vss clk d[8] q[8] q_b[8] 
+ openram_dff 
* No parameters

xdff_9 
+ vdd vss clk d[9] q[9] q_b[9] 
+ openram_dff 
* No parameters

xdff_10 
+ vdd vss clk d[10] q[10] q_b[10] 
+ openram_dff 
* No parameters

xdff_11 
+ vdd vss clk d[11] q[11] q_b[11] 
+ openram_dff 
* No parameters

.ENDS

.SUBCKT col_data_inv 
+ din din_b vdd vss 

xMP0 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='2.6' l='0.15' 

xMN0 
+ din_b din vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.4' l='0.15' 

.ENDS

.SUBCKT col_inv_array 
+ din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] din_b[7] din_b[6] din_b[5] din_b[4] din_b[3] din_b[2] din_b[1] din_b[0] vdd vss 

xinv_0 
+ din[0] din_b[0] vdd vss 
+ col_data_inv 
* No parameters

xinv_1 
+ din[1] din_b[1] vdd vss 
+ col_data_inv 
* No parameters

xinv_2 
+ din[2] din_b[2] vdd vss 
+ col_data_inv 
* No parameters

xinv_3 
+ din[3] din_b[3] vdd vss 
+ col_data_inv 
* No parameters

xinv_4 
+ din[4] din_b[4] vdd vss 
+ col_data_inv 
* No parameters

xinv_5 
+ din[5] din_b[5] vdd vss 
+ col_data_inv 
* No parameters

xinv_6 
+ din[6] din_b[6] vdd vss 
+ col_data_inv 
* No parameters

xinv_7 
+ din[7] din_b[7] vdd vss 
+ col_data_inv 
* No parameters

.ENDS

.SUBCKT sense_amp_array 
+ vdd vss clk bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] data[7] data[6] data[5] data[4] data[3] data[2] data[1] data[0] data_b[7] data_b[6] data_b[5] data_b[4] data_b[3] data_b[2] data_b[1] data_b[0] 

xsense_amp_0 
+ clk br[0] bl[0] data_b[0] data[0] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_1 
+ clk br[1] bl[1] data_b[1] data[1] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_2 
+ clk br[2] bl[2] data_b[2] data[2] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_3 
+ clk br[3] bl[3] data_b[3] data[3] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_4 
+ clk br[4] bl[4] data_b[4] data[4] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_5 
+ clk br[5] bl[5] data_b[5] data[5] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_6 
+ clk br[6] bl[6] data_b[6] data[6] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

xsense_amp_7 
+ clk br[7] bl[7] data_b[7] data[7] vdd vss 
+ sramgen_sp_sense_amp 
* No parameters

.ENDS

.SUBCKT dout_buf 
+ din1 din2 dout1 dout2 vdd vss 

xMP11 
+ x1 din1 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.6' l='0.15' 

xMN11 
+ x1 din1 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.0' l='0.15' 

xMP21 
+ dout1 x1 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='3.2' l='0.15' 

xMN21 
+ dout1 x1 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

xMP12 
+ x2 din2 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='1.6' l='0.15' 

xMN12 
+ x2 din2 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='1.0' l='0.15' 

xMP22 
+ dout2 x2 vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='3.2' l='0.15' 

xMN22 
+ dout2 x2 vss vss 
+ sky130_fd_pr__nfet_01v8 
+ w='2.0' l='0.15' 

.ENDS

.SUBCKT dout_buf_array 
+ din1[7] din1[6] din1[5] din1[4] din1[3] din1[2] din1[1] din1[0] din2[7] din2[6] din2[5] din2[4] din2[3] din2[2] din2[1] din2[0] dout1[7] dout1[6] dout1[5] dout1[4] dout1[3] dout1[2] dout1[1] dout1[0] dout2[7] dout2[6] dout2[5] dout2[4] dout2[3] dout2[2] dout2[1] dout2[0] vdd vss 

xbuf_0 
+ din1[0] din2[0] dout1[0] dout2[0] vdd vss 
+ dout_buf 
* No parameters

xbuf_1 
+ din1[1] din2[1] dout1[1] dout2[1] vdd vss 
+ dout_buf 
* No parameters

xbuf_2 
+ din1[2] din2[2] dout1[2] dout2[2] vdd vss 
+ dout_buf 
* No parameters

xbuf_3 
+ din1[3] din2[3] dout1[3] dout2[3] vdd vss 
+ dout_buf 
* No parameters

xbuf_4 
+ din1[4] din2[4] dout1[4] dout2[4] vdd vss 
+ dout_buf 
* No parameters

xbuf_5 
+ din1[5] din2[5] dout1[5] dout2[5] vdd vss 
+ dout_buf 
* No parameters

xbuf_6 
+ din1[6] din2[6] dout1[6] dout2[6] vdd vss 
+ dout_buf 
* No parameters

xbuf_7 
+ din1[7] din2[7] dout1[7] dout2[7] vdd vss 
+ dout_buf 
* No parameters

.ENDS

.SUBCKT we_control_and2_nand 
+ gnd vdd a b y 

xn1 
+ x a gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.0' l='0.15' 

xn2 
+ y b x gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='3.0' l='0.15' 

xp1 
+ y a vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='4.0' l='0.15' 

xp2 
+ y b vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='4.0' l='0.15' 

.ENDS

.SUBCKT we_control_and2_inv 
+ gnd vdd din din_b 

xn 
+ din_b din gnd gnd 
+ sky130_fd_pr__nfet_01v8 
+ w='8.0' l='0.15' 

xp 
+ din_b din vdd vdd 
+ sky130_fd_pr__pfet_01v8 
+ w='12.0' l='0.15' 

.ENDS

.SUBCKT we_control_and2 
+ a b y vdd vss 

xnand 
+ vss vdd a b tmp 
+ we_control_and2_nand 
* No parameters

xinv 
+ vss vdd tmp y 
+ we_control_and2_inv 
* No parameters

.ENDS

.SUBCKT we_control 
+ wr_en sel[7] sel[6] sel[5] sel[4] sel[3] sel[2] sel[1] sel[0] write_driver_en[7] write_driver_en[6] write_driver_en[5] write_driver_en[4] write_driver_en[3] write_driver_en[2] write_driver_en[1] write_driver_en[0] vdd vss 

xand2_0 
+ sel[0] wr_en write_driver_en[0] vdd vss 
+ we_control_and2 
* No parameters

xand2_1 
+ sel[1] wr_en write_driver_en[1] vdd vss 
+ we_control_and2 
* No parameters

xand2_2 
+ sel[2] wr_en write_driver_en[2] vdd vss 
+ we_control_and2 
* No parameters

xand2_3 
+ sel[3] wr_en write_driver_en[3] vdd vss 
+ we_control_and2 
* No parameters

xand2_4 
+ sel[4] wr_en write_driver_en[4] vdd vss 
+ we_control_and2 
* No parameters

xand2_5 
+ sel[5] wr_en write_driver_en[5] vdd vss 
+ we_control_and2 
* No parameters

xand2_6 
+ sel[6] wr_en write_driver_en[6] vdd vss 
+ we_control_and2 
* No parameters

xand2_7 
+ sel[7] wr_en write_driver_en[7] vdd vss 
+ we_control_and2 
* No parameters

.ENDS

.SUBCKT control_logic_delay_chain 
+ din dout vdd vss 

xinv_0 
+ din int[0] vdd vss 
+ control_logic_inv 
* No parameters

xinv_1 
+ int[0] int[1] vdd vss 
+ control_logic_inv 
* No parameters

xinv_2 
+ int[1] int[2] vdd vss 
+ control_logic_inv 
* No parameters

xinv_3 
+ int[2] int[3] vdd vss 
+ control_logic_inv 
* No parameters

xinv_4 
+ int[3] int[4] vdd vss 
+ control_logic_inv 
* No parameters

xinv_5 
+ int[4] int[5] vdd vss 
+ control_logic_inv 
* No parameters

xinv_6 
+ int[5] int[6] vdd vss 
+ control_logic_inv 
* No parameters

xinv_7 
+ int[6] int[7] vdd vss 
+ control_logic_inv 
* No parameters

xinv_8 
+ int[7] int[8] vdd vss 
+ control_logic_inv 
* No parameters

xinv_9 
+ int[8] int[9] vdd vss 
+ control_logic_inv 
* No parameters

xinv_10 
+ int[9] int[10] vdd vss 
+ control_logic_inv 
* No parameters

xinv_11 
+ int[10] int[11] vdd vss 
+ control_logic_inv 
* No parameters

xinv_12 
+ int[11] int[12] vdd vss 
+ control_logic_inv 
* No parameters

xinv_13 
+ int[12] int[13] vdd vss 
+ control_logic_inv 
* No parameters

xinv_14 
+ int[13] int[14] vdd vss 
+ control_logic_inv 
* No parameters

xinv_15 
+ int[14] int[15] vdd vss 
+ control_logic_inv 
* No parameters

xinv_16 
+ int[15] int[16] vdd vss 
+ control_logic_inv 
* No parameters

xinv_17 
+ int[16] int[17] vdd vss 
+ control_logic_inv 
* No parameters

xinv_18 
+ int[17] int[18] vdd vss 
+ control_logic_inv 
* No parameters

xinv_19 
+ int[18] int[19] vdd vss 
+ control_logic_inv 
* No parameters

xinv_20 
+ int[19] int[20] vdd vss 
+ control_logic_inv 
* No parameters

xinv_21 
+ int[20] int[21] vdd vss 
+ control_logic_inv 
* No parameters

xinv_22 
+ int[21] int[22] vdd vss 
+ control_logic_inv 
* No parameters

xinv_23 
+ int[22] int[23] vdd vss 
+ control_logic_inv 
* No parameters

xinv_24 
+ int[23] int[24] vdd vss 
+ control_logic_inv 
* No parameters

xinv_25 
+ int[24] int[25] vdd vss 
+ control_logic_inv 
* No parameters

xinv_26 
+ int[25] int[26] vdd vss 
+ control_logic_inv 
* No parameters

xinv_27 
+ int[26] int[27] vdd vss 
+ control_logic_inv 
* No parameters

xinv_28 
+ int[27] int[28] vdd vss 
+ control_logic_inv 
* No parameters

xinv_29 
+ int[28] int[29] vdd vss 
+ control_logic_inv 
* No parameters

xinv_30 
+ int[29] int[30] vdd vss 
+ control_logic_inv 
* No parameters

xinv_31 
+ int[30] int[31] vdd vss 
+ control_logic_inv 
* No parameters

xinv_32 
+ int[31] int[32] vdd vss 
+ control_logic_inv 
* No parameters

xinv_33 
+ int[32] int[33] vdd vss 
+ control_logic_inv 
* No parameters

xinv_34 
+ int[33] int[34] vdd vss 
+ control_logic_inv 
* No parameters

xinv_35 
+ int[34] int[35] vdd vss 
+ control_logic_inv 
* No parameters

xinv_36 
+ int[35] int[36] vdd vss 
+ control_logic_inv 
* No parameters

xinv_37 
+ int[36] int[37] vdd vss 
+ control_logic_inv 
* No parameters

xinv_38 
+ int[37] int[38] vdd vss 
+ control_logic_inv 
* No parameters

xinv_39 
+ int[38] int[39] vdd vss 
+ control_logic_inv 
* No parameters

xinv_40 
+ int[39] int[40] vdd vss 
+ control_logic_inv 
* No parameters

xinv_41 
+ int[40] int[41] vdd vss 
+ control_logic_inv 
* No parameters

xinv_42 
+ int[41] int[42] vdd vss 
+ control_logic_inv 
* No parameters

xinv_43 
+ int[42] int[43] vdd vss 
+ control_logic_inv 
* No parameters

xinv_44 
+ int[43] dout vdd vss 
+ control_logic_inv 
* No parameters

.ENDS

.SUBCKT sramgen_sram_4096x8m8w8_replica_v1 
+ vdd vss clk din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] dout[7] dout[6] dout[5] dout[4] dout[3] dout[2] dout[1] dout[0] we addr[11] addr[10] addr[9] addr[8] addr[7] addr[6] addr[5] addr[4] addr[3] addr[2] addr[1] addr[0] 

xdin_dffs 
+ vdd vss clk din[7] din[6] din[5] din[4] din[3] din[2] din[1] din[0] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] dff_din_b[7] dff_din_b[6] dff_din_b[5] dff_din_b[4] dff_din_b[3] dff_din_b[2] dff_din_b[1] dff_din_b[0] 
+ data_dff_array 
* No parameters

xaddr_dffs 
+ vdd vss clk addr[11] addr[10] addr[9] addr[8] addr[7] addr[6] addr[5] addr[4] addr[3] addr[2] addr[1] addr[0] bank_addr[11] bank_addr[10] bank_addr[9] bank_addr[8] bank_addr[7] bank_addr[6] bank_addr[5] bank_addr[4] bank_addr[3] bank_addr[2] bank_addr[1] bank_addr[0] bank_addr_b[11] bank_addr_b[10] bank_addr_b[9] bank_addr_b[8] bank_addr_b[7] bank_addr_b[6] bank_addr_b[5] bank_addr_b[4] bank_addr_b[3] bank_addr_b[2] bank_addr_b[1] bank_addr_b[0] 
+ addr_dff_array 
* No parameters

xwe_dff 
+ vdd vss clk we bank_we bank_we_b 
+ openram_dff 
* No parameters

xdecoder 
+ vdd vss bank_addr[11] bank_addr[10] bank_addr[9] bank_addr[8] bank_addr[7] bank_addr[6] bank_addr[5] bank_addr[4] bank_addr[3] bank_addr_b[11] bank_addr_b[10] bank_addr_b[9] bank_addr_b[8] bank_addr_b[7] bank_addr_b[6] bank_addr_b[5] bank_addr_b[4] bank_addr_b[3] wl_data[511] wl_data[510] wl_data[509] wl_data[508] wl_data[507] wl_data[506] wl_data[505] wl_data[504] wl_data[503] wl_data[502] wl_data[501] wl_data[500] wl_data[499] wl_data[498] wl_data[497] wl_data[496] wl_data[495] wl_data[494] wl_data[493] wl_data[492] wl_data[491] wl_data[490] wl_data[489] wl_data[488] wl_data[487] wl_data[486] wl_data[485] wl_data[484] wl_data[483] wl_data[482] wl_data[481] wl_data[480] wl_data[479] wl_data[478] wl_data[477] wl_data[476] wl_data[475] wl_data[474] wl_data[473] wl_data[472] wl_data[471] wl_data[470] wl_data[469] wl_data[468] wl_data[467] wl_data[466] wl_data[465] wl_data[464] wl_data[463] wl_data[462] wl_data[461] wl_data[460] wl_data[459] wl_data[458] wl_data[457] wl_data[456] wl_data[455] wl_data[454] wl_data[453] wl_data[452] wl_data[451] wl_data[450] wl_data[449] wl_data[448] wl_data[447] wl_data[446] wl_data[445] wl_data[444] wl_data[443] wl_data[442] wl_data[441] wl_data[440] wl_data[439] wl_data[438] wl_data[437] wl_data[436] wl_data[435] wl_data[434] wl_data[433] wl_data[432] wl_data[431] wl_data[430] wl_data[429] wl_data[428] wl_data[427] wl_data[426] wl_data[425] wl_data[424] wl_data[423] wl_data[422] wl_data[421] wl_data[420] wl_data[419] wl_data[418] wl_data[417] wl_data[416] wl_data[415] wl_data[414] wl_data[413] wl_data[412] wl_data[411] wl_data[410] wl_data[409] wl_data[408] wl_data[407] wl_data[406] wl_data[405] wl_data[404] wl_data[403] wl_data[402] wl_data[401] wl_data[400] wl_data[399] wl_data[398] wl_data[397] wl_data[396] wl_data[395] wl_data[394] wl_data[393] wl_data[392] wl_data[391] wl_data[390] wl_data[389] wl_data[388] wl_data[387] wl_data[386] wl_data[385] wl_data[384] wl_data[383] wl_data[382] wl_data[381] wl_data[380] wl_data[379] wl_data[378] wl_data[377] wl_data[376] wl_data[375] wl_data[374] wl_data[373] wl_data[372] wl_data[371] wl_data[370] wl_data[369] wl_data[368] wl_data[367] wl_data[366] wl_data[365] wl_data[364] wl_data[363] wl_data[362] wl_data[361] wl_data[360] wl_data[359] wl_data[358] wl_data[357] wl_data[356] wl_data[355] wl_data[354] wl_data[353] wl_data[352] wl_data[351] wl_data[350] wl_data[349] wl_data[348] wl_data[347] wl_data[346] wl_data[345] wl_data[344] wl_data[343] wl_data[342] wl_data[341] wl_data[340] wl_data[339] wl_data[338] wl_data[337] wl_data[336] wl_data[335] wl_data[334] wl_data[333] wl_data[332] wl_data[331] wl_data[330] wl_data[329] wl_data[328] wl_data[327] wl_data[326] wl_data[325] wl_data[324] wl_data[323] wl_data[322] wl_data[321] wl_data[320] wl_data[319] wl_data[318] wl_data[317] wl_data[316] wl_data[315] wl_data[314] wl_data[313] wl_data[312] wl_data[311] wl_data[310] wl_data[309] wl_data[308] wl_data[307] wl_data[306] wl_data[305] wl_data[304] wl_data[303] wl_data[302] wl_data[301] wl_data[300] wl_data[299] wl_data[298] wl_data[297] wl_data[296] wl_data[295] wl_data[294] wl_data[293] wl_data[292] wl_data[291] wl_data[290] wl_data[289] wl_data[288] wl_data[287] wl_data[286] wl_data[285] wl_data[284] wl_data[283] wl_data[282] wl_data[281] wl_data[280] wl_data[279] wl_data[278] wl_data[277] wl_data[276] wl_data[275] wl_data[274] wl_data[273] wl_data[272] wl_data[271] wl_data[270] wl_data[269] wl_data[268] wl_data[267] wl_data[266] wl_data[265] wl_data[264] wl_data[263] wl_data[262] wl_data[261] wl_data[260] wl_data[259] wl_data[258] wl_data[257] wl_data[256] wl_data[255] wl_data[254] wl_data[253] wl_data[252] wl_data[251] wl_data[250] wl_data[249] wl_data[248] wl_data[247] wl_data[246] wl_data[245] wl_data[244] wl_data[243] wl_data[242] wl_data[241] wl_data[240] wl_data[239] wl_data[238] wl_data[237] wl_data[236] wl_data[235] wl_data[234] wl_data[233] wl_data[232] wl_data[231] wl_data[230] wl_data[229] wl_data[228] wl_data[227] wl_data[226] wl_data[225] wl_data[224] wl_data[223] wl_data[222] wl_data[221] wl_data[220] wl_data[219] wl_data[218] wl_data[217] wl_data[216] wl_data[215] wl_data[214] wl_data[213] wl_data[212] wl_data[211] wl_data[210] wl_data[209] wl_data[208] wl_data[207] wl_data[206] wl_data[205] wl_data[204] wl_data[203] wl_data[202] wl_data[201] wl_data[200] wl_data[199] wl_data[198] wl_data[197] wl_data[196] wl_data[195] wl_data[194] wl_data[193] wl_data[192] wl_data[191] wl_data[190] wl_data[189] wl_data[188] wl_data[187] wl_data[186] wl_data[185] wl_data[184] wl_data[183] wl_data[182] wl_data[181] wl_data[180] wl_data[179] wl_data[178] wl_data[177] wl_data[176] wl_data[175] wl_data[174] wl_data[173] wl_data[172] wl_data[171] wl_data[170] wl_data[169] wl_data[168] wl_data[167] wl_data[166] wl_data[165] wl_data[164] wl_data[163] wl_data[162] wl_data[161] wl_data[160] wl_data[159] wl_data[158] wl_data[157] wl_data[156] wl_data[155] wl_data[154] wl_data[153] wl_data[152] wl_data[151] wl_data[150] wl_data[149] wl_data[148] wl_data[147] wl_data[146] wl_data[145] wl_data[144] wl_data[143] wl_data[142] wl_data[141] wl_data[140] wl_data[139] wl_data[138] wl_data[137] wl_data[136] wl_data[135] wl_data[134] wl_data[133] wl_data[132] wl_data[131] wl_data[130] wl_data[129] wl_data[128] wl_data[127] wl_data[126] wl_data[125] wl_data[124] wl_data[123] wl_data[122] wl_data[121] wl_data[120] wl_data[119] wl_data[118] wl_data[117] wl_data[116] wl_data[115] wl_data[114] wl_data[113] wl_data[112] wl_data[111] wl_data[110] wl_data[109] wl_data[108] wl_data[107] wl_data[106] wl_data[105] wl_data[104] wl_data[103] wl_data[102] wl_data[101] wl_data[100] wl_data[99] wl_data[98] wl_data[97] wl_data[96] wl_data[95] wl_data[94] wl_data[93] wl_data[92] wl_data[91] wl_data[90] wl_data[89] wl_data[88] wl_data[87] wl_data[86] wl_data[85] wl_data[84] wl_data[83] wl_data[82] wl_data[81] wl_data[80] wl_data[79] wl_data[78] wl_data[77] wl_data[76] wl_data[75] wl_data[74] wl_data[73] wl_data[72] wl_data[71] wl_data[70] wl_data[69] wl_data[68] wl_data[67] wl_data[66] wl_data[65] wl_data[64] wl_data[63] wl_data[62] wl_data[61] wl_data[60] wl_data[59] wl_data[58] wl_data[57] wl_data[56] wl_data[55] wl_data[54] wl_data[53] wl_data[52] wl_data[51] wl_data[50] wl_data[49] wl_data[48] wl_data[47] wl_data[46] wl_data[45] wl_data[44] wl_data[43] wl_data[42] wl_data[41] wl_data[40] wl_data[39] wl_data[38] wl_data[37] wl_data[36] wl_data[35] wl_data[34] wl_data[33] wl_data[32] wl_data[31] wl_data[30] wl_data[29] wl_data[28] wl_data[27] wl_data[26] wl_data[25] wl_data[24] wl_data[23] wl_data[22] wl_data[21] wl_data[20] wl_data[19] wl_data[18] wl_data[17] wl_data[16] wl_data[15] wl_data[14] wl_data[13] wl_data[12] wl_data[11] wl_data[10] wl_data[9] wl_data[8] wl_data[7] wl_data[6] wl_data[5] wl_data[4] wl_data[3] wl_data[2] wl_data[1] wl_data[0] wl_data_b[511] wl_data_b[510] wl_data_b[509] wl_data_b[508] wl_data_b[507] wl_data_b[506] wl_data_b[505] wl_data_b[504] wl_data_b[503] wl_data_b[502] wl_data_b[501] wl_data_b[500] wl_data_b[499] wl_data_b[498] wl_data_b[497] wl_data_b[496] wl_data_b[495] wl_data_b[494] wl_data_b[493] wl_data_b[492] wl_data_b[491] wl_data_b[490] wl_data_b[489] wl_data_b[488] wl_data_b[487] wl_data_b[486] wl_data_b[485] wl_data_b[484] wl_data_b[483] wl_data_b[482] wl_data_b[481] wl_data_b[480] wl_data_b[479] wl_data_b[478] wl_data_b[477] wl_data_b[476] wl_data_b[475] wl_data_b[474] wl_data_b[473] wl_data_b[472] wl_data_b[471] wl_data_b[470] wl_data_b[469] wl_data_b[468] wl_data_b[467] wl_data_b[466] wl_data_b[465] wl_data_b[464] wl_data_b[463] wl_data_b[462] wl_data_b[461] wl_data_b[460] wl_data_b[459] wl_data_b[458] wl_data_b[457] wl_data_b[456] wl_data_b[455] wl_data_b[454] wl_data_b[453] wl_data_b[452] wl_data_b[451] wl_data_b[450] wl_data_b[449] wl_data_b[448] wl_data_b[447] wl_data_b[446] wl_data_b[445] wl_data_b[444] wl_data_b[443] wl_data_b[442] wl_data_b[441] wl_data_b[440] wl_data_b[439] wl_data_b[438] wl_data_b[437] wl_data_b[436] wl_data_b[435] wl_data_b[434] wl_data_b[433] wl_data_b[432] wl_data_b[431] wl_data_b[430] wl_data_b[429] wl_data_b[428] wl_data_b[427] wl_data_b[426] wl_data_b[425] wl_data_b[424] wl_data_b[423] wl_data_b[422] wl_data_b[421] wl_data_b[420] wl_data_b[419] wl_data_b[418] wl_data_b[417] wl_data_b[416] wl_data_b[415] wl_data_b[414] wl_data_b[413] wl_data_b[412] wl_data_b[411] wl_data_b[410] wl_data_b[409] wl_data_b[408] wl_data_b[407] wl_data_b[406] wl_data_b[405] wl_data_b[404] wl_data_b[403] wl_data_b[402] wl_data_b[401] wl_data_b[400] wl_data_b[399] wl_data_b[398] wl_data_b[397] wl_data_b[396] wl_data_b[395] wl_data_b[394] wl_data_b[393] wl_data_b[392] wl_data_b[391] wl_data_b[390] wl_data_b[389] wl_data_b[388] wl_data_b[387] wl_data_b[386] wl_data_b[385] wl_data_b[384] wl_data_b[383] wl_data_b[382] wl_data_b[381] wl_data_b[380] wl_data_b[379] wl_data_b[378] wl_data_b[377] wl_data_b[376] wl_data_b[375] wl_data_b[374] wl_data_b[373] wl_data_b[372] wl_data_b[371] wl_data_b[370] wl_data_b[369] wl_data_b[368] wl_data_b[367] wl_data_b[366] wl_data_b[365] wl_data_b[364] wl_data_b[363] wl_data_b[362] wl_data_b[361] wl_data_b[360] wl_data_b[359] wl_data_b[358] wl_data_b[357] wl_data_b[356] wl_data_b[355] wl_data_b[354] wl_data_b[353] wl_data_b[352] wl_data_b[351] wl_data_b[350] wl_data_b[349] wl_data_b[348] wl_data_b[347] wl_data_b[346] wl_data_b[345] wl_data_b[344] wl_data_b[343] wl_data_b[342] wl_data_b[341] wl_data_b[340] wl_data_b[339] wl_data_b[338] wl_data_b[337] wl_data_b[336] wl_data_b[335] wl_data_b[334] wl_data_b[333] wl_data_b[332] wl_data_b[331] wl_data_b[330] wl_data_b[329] wl_data_b[328] wl_data_b[327] wl_data_b[326] wl_data_b[325] wl_data_b[324] wl_data_b[323] wl_data_b[322] wl_data_b[321] wl_data_b[320] wl_data_b[319] wl_data_b[318] wl_data_b[317] wl_data_b[316] wl_data_b[315] wl_data_b[314] wl_data_b[313] wl_data_b[312] wl_data_b[311] wl_data_b[310] wl_data_b[309] wl_data_b[308] wl_data_b[307] wl_data_b[306] wl_data_b[305] wl_data_b[304] wl_data_b[303] wl_data_b[302] wl_data_b[301] wl_data_b[300] wl_data_b[299] wl_data_b[298] wl_data_b[297] wl_data_b[296] wl_data_b[295] wl_data_b[294] wl_data_b[293] wl_data_b[292] wl_data_b[291] wl_data_b[290] wl_data_b[289] wl_data_b[288] wl_data_b[287] wl_data_b[286] wl_data_b[285] wl_data_b[284] wl_data_b[283] wl_data_b[282] wl_data_b[281] wl_data_b[280] wl_data_b[279] wl_data_b[278] wl_data_b[277] wl_data_b[276] wl_data_b[275] wl_data_b[274] wl_data_b[273] wl_data_b[272] wl_data_b[271] wl_data_b[270] wl_data_b[269] wl_data_b[268] wl_data_b[267] wl_data_b[266] wl_data_b[265] wl_data_b[264] wl_data_b[263] wl_data_b[262] wl_data_b[261] wl_data_b[260] wl_data_b[259] wl_data_b[258] wl_data_b[257] wl_data_b[256] wl_data_b[255] wl_data_b[254] wl_data_b[253] wl_data_b[252] wl_data_b[251] wl_data_b[250] wl_data_b[249] wl_data_b[248] wl_data_b[247] wl_data_b[246] wl_data_b[245] wl_data_b[244] wl_data_b[243] wl_data_b[242] wl_data_b[241] wl_data_b[240] wl_data_b[239] wl_data_b[238] wl_data_b[237] wl_data_b[236] wl_data_b[235] wl_data_b[234] wl_data_b[233] wl_data_b[232] wl_data_b[231] wl_data_b[230] wl_data_b[229] wl_data_b[228] wl_data_b[227] wl_data_b[226] wl_data_b[225] wl_data_b[224] wl_data_b[223] wl_data_b[222] wl_data_b[221] wl_data_b[220] wl_data_b[219] wl_data_b[218] wl_data_b[217] wl_data_b[216] wl_data_b[215] wl_data_b[214] wl_data_b[213] wl_data_b[212] wl_data_b[211] wl_data_b[210] wl_data_b[209] wl_data_b[208] wl_data_b[207] wl_data_b[206] wl_data_b[205] wl_data_b[204] wl_data_b[203] wl_data_b[202] wl_data_b[201] wl_data_b[200] wl_data_b[199] wl_data_b[198] wl_data_b[197] wl_data_b[196] wl_data_b[195] wl_data_b[194] wl_data_b[193] wl_data_b[192] wl_data_b[191] wl_data_b[190] wl_data_b[189] wl_data_b[188] wl_data_b[187] wl_data_b[186] wl_data_b[185] wl_data_b[184] wl_data_b[183] wl_data_b[182] wl_data_b[181] wl_data_b[180] wl_data_b[179] wl_data_b[178] wl_data_b[177] wl_data_b[176] wl_data_b[175] wl_data_b[174] wl_data_b[173] wl_data_b[172] wl_data_b[171] wl_data_b[170] wl_data_b[169] wl_data_b[168] wl_data_b[167] wl_data_b[166] wl_data_b[165] wl_data_b[164] wl_data_b[163] wl_data_b[162] wl_data_b[161] wl_data_b[160] wl_data_b[159] wl_data_b[158] wl_data_b[157] wl_data_b[156] wl_data_b[155] wl_data_b[154] wl_data_b[153] wl_data_b[152] wl_data_b[151] wl_data_b[150] wl_data_b[149] wl_data_b[148] wl_data_b[147] wl_data_b[146] wl_data_b[145] wl_data_b[144] wl_data_b[143] wl_data_b[142] wl_data_b[141] wl_data_b[140] wl_data_b[139] wl_data_b[138] wl_data_b[137] wl_data_b[136] wl_data_b[135] wl_data_b[134] wl_data_b[133] wl_data_b[132] wl_data_b[131] wl_data_b[130] wl_data_b[129] wl_data_b[128] wl_data_b[127] wl_data_b[126] wl_data_b[125] wl_data_b[124] wl_data_b[123] wl_data_b[122] wl_data_b[121] wl_data_b[120] wl_data_b[119] wl_data_b[118] wl_data_b[117] wl_data_b[116] wl_data_b[115] wl_data_b[114] wl_data_b[113] wl_data_b[112] wl_data_b[111] wl_data_b[110] wl_data_b[109] wl_data_b[108] wl_data_b[107] wl_data_b[106] wl_data_b[105] wl_data_b[104] wl_data_b[103] wl_data_b[102] wl_data_b[101] wl_data_b[100] wl_data_b[99] wl_data_b[98] wl_data_b[97] wl_data_b[96] wl_data_b[95] wl_data_b[94] wl_data_b[93] wl_data_b[92] wl_data_b[91] wl_data_b[90] wl_data_b[89] wl_data_b[88] wl_data_b[87] wl_data_b[86] wl_data_b[85] wl_data_b[84] wl_data_b[83] wl_data_b[82] wl_data_b[81] wl_data_b[80] wl_data_b[79] wl_data_b[78] wl_data_b[77] wl_data_b[76] wl_data_b[75] wl_data_b[74] wl_data_b[73] wl_data_b[72] wl_data_b[71] wl_data_b[70] wl_data_b[69] wl_data_b[68] wl_data_b[67] wl_data_b[66] wl_data_b[65] wl_data_b[64] wl_data_b[63] wl_data_b[62] wl_data_b[61] wl_data_b[60] wl_data_b[59] wl_data_b[58] wl_data_b[57] wl_data_b[56] wl_data_b[55] wl_data_b[54] wl_data_b[53] wl_data_b[52] wl_data_b[51] wl_data_b[50] wl_data_b[49] wl_data_b[48] wl_data_b[47] wl_data_b[46] wl_data_b[45] wl_data_b[44] wl_data_b[43] wl_data_b[42] wl_data_b[41] wl_data_b[40] wl_data_b[39] wl_data_b[38] wl_data_b[37] wl_data_b[36] wl_data_b[35] wl_data_b[34] wl_data_b[33] wl_data_b[32] wl_data_b[31] wl_data_b[30] wl_data_b[29] wl_data_b[28] wl_data_b[27] wl_data_b[26] wl_data_b[25] wl_data_b[24] wl_data_b[23] wl_data_b[22] wl_data_b[21] wl_data_b[20] wl_data_b[19] wl_data_b[18] wl_data_b[17] wl_data_b[16] wl_data_b[15] wl_data_b[14] wl_data_b[13] wl_data_b[12] wl_data_b[11] wl_data_b[10] wl_data_b[9] wl_data_b[8] wl_data_b[7] wl_data_b[6] wl_data_b[5] wl_data_b[4] wl_data_b[3] wl_data_b[2] wl_data_b[1] wl_data_b[0] 
+ hierarchical_decoder 
* No parameters

xwl_driver_array 
+ vdd vss wl_data[511] wl_data[510] wl_data[509] wl_data[508] wl_data[507] wl_data[506] wl_data[505] wl_data[504] wl_data[503] wl_data[502] wl_data[501] wl_data[500] wl_data[499] wl_data[498] wl_data[497] wl_data[496] wl_data[495] wl_data[494] wl_data[493] wl_data[492] wl_data[491] wl_data[490] wl_data[489] wl_data[488] wl_data[487] wl_data[486] wl_data[485] wl_data[484] wl_data[483] wl_data[482] wl_data[481] wl_data[480] wl_data[479] wl_data[478] wl_data[477] wl_data[476] wl_data[475] wl_data[474] wl_data[473] wl_data[472] wl_data[471] wl_data[470] wl_data[469] wl_data[468] wl_data[467] wl_data[466] wl_data[465] wl_data[464] wl_data[463] wl_data[462] wl_data[461] wl_data[460] wl_data[459] wl_data[458] wl_data[457] wl_data[456] wl_data[455] wl_data[454] wl_data[453] wl_data[452] wl_data[451] wl_data[450] wl_data[449] wl_data[448] wl_data[447] wl_data[446] wl_data[445] wl_data[444] wl_data[443] wl_data[442] wl_data[441] wl_data[440] wl_data[439] wl_data[438] wl_data[437] wl_data[436] wl_data[435] wl_data[434] wl_data[433] wl_data[432] wl_data[431] wl_data[430] wl_data[429] wl_data[428] wl_data[427] wl_data[426] wl_data[425] wl_data[424] wl_data[423] wl_data[422] wl_data[421] wl_data[420] wl_data[419] wl_data[418] wl_data[417] wl_data[416] wl_data[415] wl_data[414] wl_data[413] wl_data[412] wl_data[411] wl_data[410] wl_data[409] wl_data[408] wl_data[407] wl_data[406] wl_data[405] wl_data[404] wl_data[403] wl_data[402] wl_data[401] wl_data[400] wl_data[399] wl_data[398] wl_data[397] wl_data[396] wl_data[395] wl_data[394] wl_data[393] wl_data[392] wl_data[391] wl_data[390] wl_data[389] wl_data[388] wl_data[387] wl_data[386] wl_data[385] wl_data[384] wl_data[383] wl_data[382] wl_data[381] wl_data[380] wl_data[379] wl_data[378] wl_data[377] wl_data[376] wl_data[375] wl_data[374] wl_data[373] wl_data[372] wl_data[371] wl_data[370] wl_data[369] wl_data[368] wl_data[367] wl_data[366] wl_data[365] wl_data[364] wl_data[363] wl_data[362] wl_data[361] wl_data[360] wl_data[359] wl_data[358] wl_data[357] wl_data[356] wl_data[355] wl_data[354] wl_data[353] wl_data[352] wl_data[351] wl_data[350] wl_data[349] wl_data[348] wl_data[347] wl_data[346] wl_data[345] wl_data[344] wl_data[343] wl_data[342] wl_data[341] wl_data[340] wl_data[339] wl_data[338] wl_data[337] wl_data[336] wl_data[335] wl_data[334] wl_data[333] wl_data[332] wl_data[331] wl_data[330] wl_data[329] wl_data[328] wl_data[327] wl_data[326] wl_data[325] wl_data[324] wl_data[323] wl_data[322] wl_data[321] wl_data[320] wl_data[319] wl_data[318] wl_data[317] wl_data[316] wl_data[315] wl_data[314] wl_data[313] wl_data[312] wl_data[311] wl_data[310] wl_data[309] wl_data[308] wl_data[307] wl_data[306] wl_data[305] wl_data[304] wl_data[303] wl_data[302] wl_data[301] wl_data[300] wl_data[299] wl_data[298] wl_data[297] wl_data[296] wl_data[295] wl_data[294] wl_data[293] wl_data[292] wl_data[291] wl_data[290] wl_data[289] wl_data[288] wl_data[287] wl_data[286] wl_data[285] wl_data[284] wl_data[283] wl_data[282] wl_data[281] wl_data[280] wl_data[279] wl_data[278] wl_data[277] wl_data[276] wl_data[275] wl_data[274] wl_data[273] wl_data[272] wl_data[271] wl_data[270] wl_data[269] wl_data[268] wl_data[267] wl_data[266] wl_data[265] wl_data[264] wl_data[263] wl_data[262] wl_data[261] wl_data[260] wl_data[259] wl_data[258] wl_data[257] wl_data[256] wl_data[255] wl_data[254] wl_data[253] wl_data[252] wl_data[251] wl_data[250] wl_data[249] wl_data[248] wl_data[247] wl_data[246] wl_data[245] wl_data[244] wl_data[243] wl_data[242] wl_data[241] wl_data[240] wl_data[239] wl_data[238] wl_data[237] wl_data[236] wl_data[235] wl_data[234] wl_data[233] wl_data[232] wl_data[231] wl_data[230] wl_data[229] wl_data[228] wl_data[227] wl_data[226] wl_data[225] wl_data[224] wl_data[223] wl_data[222] wl_data[221] wl_data[220] wl_data[219] wl_data[218] wl_data[217] wl_data[216] wl_data[215] wl_data[214] wl_data[213] wl_data[212] wl_data[211] wl_data[210] wl_data[209] wl_data[208] wl_data[207] wl_data[206] wl_data[205] wl_data[204] wl_data[203] wl_data[202] wl_data[201] wl_data[200] wl_data[199] wl_data[198] wl_data[197] wl_data[196] wl_data[195] wl_data[194] wl_data[193] wl_data[192] wl_data[191] wl_data[190] wl_data[189] wl_data[188] wl_data[187] wl_data[186] wl_data[185] wl_data[184] wl_data[183] wl_data[182] wl_data[181] wl_data[180] wl_data[179] wl_data[178] wl_data[177] wl_data[176] wl_data[175] wl_data[174] wl_data[173] wl_data[172] wl_data[171] wl_data[170] wl_data[169] wl_data[168] wl_data[167] wl_data[166] wl_data[165] wl_data[164] wl_data[163] wl_data[162] wl_data[161] wl_data[160] wl_data[159] wl_data[158] wl_data[157] wl_data[156] wl_data[155] wl_data[154] wl_data[153] wl_data[152] wl_data[151] wl_data[150] wl_data[149] wl_data[148] wl_data[147] wl_data[146] wl_data[145] wl_data[144] wl_data[143] wl_data[142] wl_data[141] wl_data[140] wl_data[139] wl_data[138] wl_data[137] wl_data[136] wl_data[135] wl_data[134] wl_data[133] wl_data[132] wl_data[131] wl_data[130] wl_data[129] wl_data[128] wl_data[127] wl_data[126] wl_data[125] wl_data[124] wl_data[123] wl_data[122] wl_data[121] wl_data[120] wl_data[119] wl_data[118] wl_data[117] wl_data[116] wl_data[115] wl_data[114] wl_data[113] wl_data[112] wl_data[111] wl_data[110] wl_data[109] wl_data[108] wl_data[107] wl_data[106] wl_data[105] wl_data[104] wl_data[103] wl_data[102] wl_data[101] wl_data[100] wl_data[99] wl_data[98] wl_data[97] wl_data[96] wl_data[95] wl_data[94] wl_data[93] wl_data[92] wl_data[91] wl_data[90] wl_data[89] wl_data[88] wl_data[87] wl_data[86] wl_data[85] wl_data[84] wl_data[83] wl_data[82] wl_data[81] wl_data[80] wl_data[79] wl_data[78] wl_data[77] wl_data[76] wl_data[75] wl_data[74] wl_data[73] wl_data[72] wl_data[71] wl_data[70] wl_data[69] wl_data[68] wl_data[67] wl_data[66] wl_data[65] wl_data[64] wl_data[63] wl_data[62] wl_data[61] wl_data[60] wl_data[59] wl_data[58] wl_data[57] wl_data[56] wl_data[55] wl_data[54] wl_data[53] wl_data[52] wl_data[51] wl_data[50] wl_data[49] wl_data[48] wl_data[47] wl_data[46] wl_data[45] wl_data[44] wl_data[43] wl_data[42] wl_data[41] wl_data[40] wl_data[39] wl_data[38] wl_data[37] wl_data[36] wl_data[35] wl_data[34] wl_data[33] wl_data[32] wl_data[31] wl_data[30] wl_data[29] wl_data[28] wl_data[27] wl_data[26] wl_data[25] wl_data[24] wl_data[23] wl_data[22] wl_data[21] wl_data[20] wl_data[19] wl_data[18] wl_data[17] wl_data[16] wl_data[15] wl_data[14] wl_data[13] wl_data[12] wl_data[11] wl_data[10] wl_data[9] wl_data[8] wl_data[7] wl_data[6] wl_data[5] wl_data[4] wl_data[3] wl_data[2] wl_data[1] wl_data[0] wl_en wl[511] wl[510] wl[509] wl[508] wl[507] wl[506] wl[505] wl[504] wl[503] wl[502] wl[501] wl[500] wl[499] wl[498] wl[497] wl[496] wl[495] wl[494] wl[493] wl[492] wl[491] wl[490] wl[489] wl[488] wl[487] wl[486] wl[485] wl[484] wl[483] wl[482] wl[481] wl[480] wl[479] wl[478] wl[477] wl[476] wl[475] wl[474] wl[473] wl[472] wl[471] wl[470] wl[469] wl[468] wl[467] wl[466] wl[465] wl[464] wl[463] wl[462] wl[461] wl[460] wl[459] wl[458] wl[457] wl[456] wl[455] wl[454] wl[453] wl[452] wl[451] wl[450] wl[449] wl[448] wl[447] wl[446] wl[445] wl[444] wl[443] wl[442] wl[441] wl[440] wl[439] wl[438] wl[437] wl[436] wl[435] wl[434] wl[433] wl[432] wl[431] wl[430] wl[429] wl[428] wl[427] wl[426] wl[425] wl[424] wl[423] wl[422] wl[421] wl[420] wl[419] wl[418] wl[417] wl[416] wl[415] wl[414] wl[413] wl[412] wl[411] wl[410] wl[409] wl[408] wl[407] wl[406] wl[405] wl[404] wl[403] wl[402] wl[401] wl[400] wl[399] wl[398] wl[397] wl[396] wl[395] wl[394] wl[393] wl[392] wl[391] wl[390] wl[389] wl[388] wl[387] wl[386] wl[385] wl[384] wl[383] wl[382] wl[381] wl[380] wl[379] wl[378] wl[377] wl[376] wl[375] wl[374] wl[373] wl[372] wl[371] wl[370] wl[369] wl[368] wl[367] wl[366] wl[365] wl[364] wl[363] wl[362] wl[361] wl[360] wl[359] wl[358] wl[357] wl[356] wl[355] wl[354] wl[353] wl[352] wl[351] wl[350] wl[349] wl[348] wl[347] wl[346] wl[345] wl[344] wl[343] wl[342] wl[341] wl[340] wl[339] wl[338] wl[337] wl[336] wl[335] wl[334] wl[333] wl[332] wl[331] wl[330] wl[329] wl[328] wl[327] wl[326] wl[325] wl[324] wl[323] wl[322] wl[321] wl[320] wl[319] wl[318] wl[317] wl[316] wl[315] wl[314] wl[313] wl[312] wl[311] wl[310] wl[309] wl[308] wl[307] wl[306] wl[305] wl[304] wl[303] wl[302] wl[301] wl[300] wl[299] wl[298] wl[297] wl[296] wl[295] wl[294] wl[293] wl[292] wl[291] wl[290] wl[289] wl[288] wl[287] wl[286] wl[285] wl[284] wl[283] wl[282] wl[281] wl[280] wl[279] wl[278] wl[277] wl[276] wl[275] wl[274] wl[273] wl[272] wl[271] wl[270] wl[269] wl[268] wl[267] wl[266] wl[265] wl[264] wl[263] wl[262] wl[261] wl[260] wl[259] wl[258] wl[257] wl[256] wl[255] wl[254] wl[253] wl[252] wl[251] wl[250] wl[249] wl[248] wl[247] wl[246] wl[245] wl[244] wl[243] wl[242] wl[241] wl[240] wl[239] wl[238] wl[237] wl[236] wl[235] wl[234] wl[233] wl[232] wl[231] wl[230] wl[229] wl[228] wl[227] wl[226] wl[225] wl[224] wl[223] wl[222] wl[221] wl[220] wl[219] wl[218] wl[217] wl[216] wl[215] wl[214] wl[213] wl[212] wl[211] wl[210] wl[209] wl[208] wl[207] wl[206] wl[205] wl[204] wl[203] wl[202] wl[201] wl[200] wl[199] wl[198] wl[197] wl[196] wl[195] wl[194] wl[193] wl[192] wl[191] wl[190] wl[189] wl[188] wl[187] wl[186] wl[185] wl[184] wl[183] wl[182] wl[181] wl[180] wl[179] wl[178] wl[177] wl[176] wl[175] wl[174] wl[173] wl[172] wl[171] wl[170] wl[169] wl[168] wl[167] wl[166] wl[165] wl[164] wl[163] wl[162] wl[161] wl[160] wl[159] wl[158] wl[157] wl[156] wl[155] wl[154] wl[153] wl[152] wl[151] wl[150] wl[149] wl[148] wl[147] wl[146] wl[145] wl[144] wl[143] wl[142] wl[141] wl[140] wl[139] wl[138] wl[137] wl[136] wl[135] wl[134] wl[133] wl[132] wl[131] wl[130] wl[129] wl[128] wl[127] wl[126] wl[125] wl[124] wl[123] wl[122] wl[121] wl[120] wl[119] wl[118] wl[117] wl[116] wl[115] wl[114] wl[113] wl[112] wl[111] wl[110] wl[109] wl[108] wl[107] wl[106] wl[105] wl[104] wl[103] wl[102] wl[101] wl[100] wl[99] wl[98] wl[97] wl[96] wl[95] wl[94] wl[93] wl[92] wl[91] wl[90] wl[89] wl[88] wl[87] wl[86] wl[85] wl[84] wl[83] wl[82] wl[81] wl[80] wl[79] wl[78] wl[77] wl[76] wl[75] wl[74] wl[73] wl[72] wl[71] wl[70] wl[69] wl[68] wl[67] wl[66] wl[65] wl[64] wl[63] wl[62] wl[61] wl[60] wl[59] wl[58] wl[57] wl[56] wl[55] wl[54] wl[53] wl[52] wl[51] wl[50] wl[49] wl[48] wl[47] wl[46] wl[45] wl[44] wl[43] wl[42] wl[41] wl[40] wl[39] wl[38] wl[37] wl[36] wl[35] wl[34] wl[33] wl[32] wl[31] wl[30] wl[29] wl[28] wl[27] wl[26] wl[25] wl[24] wl[23] wl[22] wl[21] wl[20] wl[19] wl[18] wl[17] wl[16] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] 
+ wordline_driver_array 
* No parameters

xbitcells 
+ vdd vss bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] wl[511] wl[510] wl[509] wl[508] wl[507] wl[506] wl[505] wl[504] wl[503] wl[502] wl[501] wl[500] wl[499] wl[498] wl[497] wl[496] wl[495] wl[494] wl[493] wl[492] wl[491] wl[490] wl[489] wl[488] wl[487] wl[486] wl[485] wl[484] wl[483] wl[482] wl[481] wl[480] wl[479] wl[478] wl[477] wl[476] wl[475] wl[474] wl[473] wl[472] wl[471] wl[470] wl[469] wl[468] wl[467] wl[466] wl[465] wl[464] wl[463] wl[462] wl[461] wl[460] wl[459] wl[458] wl[457] wl[456] wl[455] wl[454] wl[453] wl[452] wl[451] wl[450] wl[449] wl[448] wl[447] wl[446] wl[445] wl[444] wl[443] wl[442] wl[441] wl[440] wl[439] wl[438] wl[437] wl[436] wl[435] wl[434] wl[433] wl[432] wl[431] wl[430] wl[429] wl[428] wl[427] wl[426] wl[425] wl[424] wl[423] wl[422] wl[421] wl[420] wl[419] wl[418] wl[417] wl[416] wl[415] wl[414] wl[413] wl[412] wl[411] wl[410] wl[409] wl[408] wl[407] wl[406] wl[405] wl[404] wl[403] wl[402] wl[401] wl[400] wl[399] wl[398] wl[397] wl[396] wl[395] wl[394] wl[393] wl[392] wl[391] wl[390] wl[389] wl[388] wl[387] wl[386] wl[385] wl[384] wl[383] wl[382] wl[381] wl[380] wl[379] wl[378] wl[377] wl[376] wl[375] wl[374] wl[373] wl[372] wl[371] wl[370] wl[369] wl[368] wl[367] wl[366] wl[365] wl[364] wl[363] wl[362] wl[361] wl[360] wl[359] wl[358] wl[357] wl[356] wl[355] wl[354] wl[353] wl[352] wl[351] wl[350] wl[349] wl[348] wl[347] wl[346] wl[345] wl[344] wl[343] wl[342] wl[341] wl[340] wl[339] wl[338] wl[337] wl[336] wl[335] wl[334] wl[333] wl[332] wl[331] wl[330] wl[329] wl[328] wl[327] wl[326] wl[325] wl[324] wl[323] wl[322] wl[321] wl[320] wl[319] wl[318] wl[317] wl[316] wl[315] wl[314] wl[313] wl[312] wl[311] wl[310] wl[309] wl[308] wl[307] wl[306] wl[305] wl[304] wl[303] wl[302] wl[301] wl[300] wl[299] wl[298] wl[297] wl[296] wl[295] wl[294] wl[293] wl[292] wl[291] wl[290] wl[289] wl[288] wl[287] wl[286] wl[285] wl[284] wl[283] wl[282] wl[281] wl[280] wl[279] wl[278] wl[277] wl[276] wl[275] wl[274] wl[273] wl[272] wl[271] wl[270] wl[269] wl[268] wl[267] wl[266] wl[265] wl[264] wl[263] wl[262] wl[261] wl[260] wl[259] wl[258] wl[257] wl[256] wl[255] wl[254] wl[253] wl[252] wl[251] wl[250] wl[249] wl[248] wl[247] wl[246] wl[245] wl[244] wl[243] wl[242] wl[241] wl[240] wl[239] wl[238] wl[237] wl[236] wl[235] wl[234] wl[233] wl[232] wl[231] wl[230] wl[229] wl[228] wl[227] wl[226] wl[225] wl[224] wl[223] wl[222] wl[221] wl[220] wl[219] wl[218] wl[217] wl[216] wl[215] wl[214] wl[213] wl[212] wl[211] wl[210] wl[209] wl[208] wl[207] wl[206] wl[205] wl[204] wl[203] wl[202] wl[201] wl[200] wl[199] wl[198] wl[197] wl[196] wl[195] wl[194] wl[193] wl[192] wl[191] wl[190] wl[189] wl[188] wl[187] wl[186] wl[185] wl[184] wl[183] wl[182] wl[181] wl[180] wl[179] wl[178] wl[177] wl[176] wl[175] wl[174] wl[173] wl[172] wl[171] wl[170] wl[169] wl[168] wl[167] wl[166] wl[165] wl[164] wl[163] wl[162] wl[161] wl[160] wl[159] wl[158] wl[157] wl[156] wl[155] wl[154] wl[153] wl[152] wl[151] wl[150] wl[149] wl[148] wl[147] wl[146] wl[145] wl[144] wl[143] wl[142] wl[141] wl[140] wl[139] wl[138] wl[137] wl[136] wl[135] wl[134] wl[133] wl[132] wl[131] wl[130] wl[129] wl[128] wl[127] wl[126] wl[125] wl[124] wl[123] wl[122] wl[121] wl[120] wl[119] wl[118] wl[117] wl[116] wl[115] wl[114] wl[113] wl[112] wl[111] wl[110] wl[109] wl[108] wl[107] wl[106] wl[105] wl[104] wl[103] wl[102] wl[101] wl[100] wl[99] wl[98] wl[97] wl[96] wl[95] wl[94] wl[93] wl[92] wl[91] wl[90] wl[89] wl[88] wl[87] wl[86] wl[85] wl[84] wl[83] wl[82] wl[81] wl[80] wl[79] wl[78] wl[77] wl[76] wl[75] wl[74] wl[73] wl[72] wl[71] wl[70] wl[69] wl[68] wl[67] wl[66] wl[65] wl[64] wl[63] wl[62] wl[61] wl[60] wl[59] wl[58] wl[57] wl[56] wl[55] wl[54] wl[53] wl[52] wl[51] wl[50] wl[49] wl[48] wl[47] wl[46] wl[45] wl[44] wl[43] wl[42] wl[41] wl[40] wl[39] wl[38] wl[37] wl[36] wl[35] wl[34] wl[33] wl[32] wl[31] wl[30] wl[29] wl[28] wl[27] wl[26] wl[25] wl[24] wl[23] wl[22] wl[21] wl[20] wl[19] wl[18] wl[17] wl[16] wl[15] wl[14] wl[13] wl[12] wl[11] wl[10] wl[9] wl[8] wl[7] wl[6] wl[5] wl[4] wl[3] wl[2] wl[1] wl[0] vss vdd rbl rbr 
+ bitcell_array 
* No parameters

xprecharge_array 
+ vdd pc_b rbl bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0]  rbr br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0]  
+ precharge_array 
* No parameters

xwrite_mux_array 
+ write_driver_en[7] write_driver_en[6] write_driver_en[5] write_driver_en[4] write_driver_en[3] write_driver_en[2] write_driver_en[1] write_driver_en[0] bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] bank_din_b[7] bank_din_b[6] bank_din_b[5] bank_din_b[4] bank_din_b[3] bank_din_b[2] bank_din_b[1] bank_din_b[0] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] vss 
+ write_mux_array 
* No parameters

xread_mux_array 
+ col_sel_b[7] col_sel_b[6] col_sel_b[5] col_sel_b[4] col_sel_b[3] col_sel_b[2] col_sel_b[1] col_sel_b[0] bl[63] bl[62] bl[61] bl[60] bl[59] bl[58] bl[57] bl[56] bl[55] bl[54] bl[53] bl[52] bl[51] bl[50] bl[49] bl[48] bl[47] bl[46] bl[45] bl[44] bl[43] bl[42] bl[41] bl[40] bl[39] bl[38] bl[37] bl[36] bl[35] bl[34] bl[33] bl[32] bl[31] bl[30] bl[29] bl[28] bl[27] bl[26] bl[25] bl[24] bl[23] bl[22] bl[21] bl[20] bl[19] bl[18] bl[17] bl[16] bl[15] bl[14] bl[13] bl[12] bl[11] bl[10] bl[9] bl[8] bl[7] bl[6] bl[5] bl[4] bl[3] bl[2] bl[1] bl[0] br[63] br[62] br[61] br[60] br[59] br[58] br[57] br[56] br[55] br[54] br[53] br[52] br[51] br[50] br[49] br[48] br[47] br[46] br[45] br[44] br[43] br[42] br[41] br[40] br[39] br[38] br[37] br[36] br[35] br[34] br[33] br[32] br[31] br[30] br[29] br[28] br[27] br[26] br[25] br[24] br[23] br[22] br[21] br[20] br[19] br[18] br[17] br[16] br[15] br[14] br[13] br[12] br[11] br[10] br[9] br[8] br[7] br[6] br[5] br[4] br[3] br[2] br[1] br[0] bl_read[7] bl_read[6] bl_read[5] bl_read[4] bl_read[3] bl_read[2] bl_read[1] bl_read[0] br_read[7] br_read[6] br_read[5] br_read[4] br_read[3] br_read[2] br_read[1] br_read[0] vdd 
+ read_mux_array 
* No parameters

xcol_inv_array 
+ bank_din[7] bank_din[6] bank_din[5] bank_din[4] bank_din[3] bank_din[2] bank_din[1] bank_din[0] bank_din_b[7] bank_din_b[6] bank_din_b[5] bank_din_b[4] bank_din_b[3] bank_din_b[2] bank_din_b[1] bank_din_b[0] vdd vss 
+ col_inv_array 
* No parameters

xsense_amp_array 
+ vdd vss sense_amp_en bl_read[7] bl_read[6] bl_read[5] bl_read[4] bl_read[3] bl_read[2] bl_read[1] bl_read[0] br_read[7] br_read[6] br_read[5] br_read[4] br_read[3] br_read[2] br_read[1] br_read[0] sa_outp[7] sa_outp[6] sa_outp[5] sa_outp[4] sa_outp[3] sa_outp[2] sa_outp[1] sa_outp[0] sa_outn[7] sa_outn[6] sa_outn[5] sa_outn[4] sa_outn[3] sa_outn[2] sa_outn[1] sa_outn[0] 
+ sense_amp_array 
* No parameters

xdout_buf_array 
+ sa_outp[7] sa_outp[6] sa_outp[5] sa_outp[4] sa_outp[3] sa_outp[2] sa_outp[1] sa_outp[0] sa_outn[7] sa_outn[6] sa_outn[5] sa_outn[4] sa_outn[3] sa_outn[2] sa_outn[1] sa_outn[0] dout[7] dout[6] dout[5] dout[4] dout[3] dout[2] dout[1] dout[0] dout_b[7] dout_b[6] dout_b[5] dout_b[4] dout_b[3] dout_b[2] dout_b[1] dout_b[0] vdd vss 
+ dout_buf_array 
* No parameters

xcontrol_logic 
+ clk bank_we rbl pc_b wl_en wr_en sense_amp_en vdd vss 
+ sramgen_control_replica_v1 
* No parameters

xcolumn_decoder 
+ vdd vss bank_addr[2] bank_addr[1] bank_addr[0] bank_addr_b[2] bank_addr_b[1] bank_addr_b[0] col_sel[7] col_sel[6] col_sel[5] col_sel[4] col_sel[3] col_sel[2] col_sel[1] col_sel[0] col_sel_b[7] col_sel_b[6] col_sel_b[5] col_sel_b[4] col_sel_b[3] col_sel_b[2] col_sel_b[1] col_sel_b[0] 
+ column_decoder 
* No parameters

xwe_control 
+ wr_en col_sel[7] col_sel[6] col_sel[5] col_sel[4] col_sel[3] col_sel[2] col_sel[1] col_sel[0] write_driver_en[7] write_driver_en[6] write_driver_en[5] write_driver_en[4] write_driver_en[3] write_driver_en[2] write_driver_en[1] write_driver_en[0] vdd vss 
+ we_control 
* No parameters

.ENDS

